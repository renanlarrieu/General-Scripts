-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of MultiPartiteAdder object for LNS arithmetic in base 2.0 with 8-bit integer part and 9-bit fractional part
-- wI = 13 bits
-- wO = 10 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnsadd_mpt_9 is
  component LNSAdd_MPT_T1_9 is
    port( x : in  std_logic_vector(12 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9 is
    port( x : in  std_logic_vector(11 downto 0);
          r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9_Clk is
    port( x   : in  std_logic_vector(11 downto 0);
          r   : out std_logic_vector(9 downto 0);
          clk : in  std_logic );
  end component;
end package;


-- SimpleTable: LNS addition function: [-16.0 0.0[ -> [0.0 2.0[
-- (bounded to [-16.0; -8.0[)
-- wI = 13 bits
-- wO = 3 bits

library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T1_9 is
  port( x : in  std_logic_vector(12 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T1_9 is
begin
  with x select
    r <=
      "000" when "0000000000000", -- t[0] = 0
      "000" when "0000000000001", -- t[1] = 0
      "000" when "0000000000010", -- t[2] = 0
      "000" when "0000000000011", -- t[3] = 0
      "000" when "0000000000100", -- t[4] = 0
      "000" when "0000000000101", -- t[5] = 0
      "000" when "0000000000110", -- t[6] = 0
      "000" when "0000000000111", -- t[7] = 0
      "000" when "0000000001000", -- t[8] = 0
      "000" when "0000000001001", -- t[9] = 0
      "000" when "0000000001010", -- t[10] = 0
      "000" when "0000000001011", -- t[11] = 0
      "000" when "0000000001100", -- t[12] = 0
      "000" when "0000000001101", -- t[13] = 0
      "000" when "0000000001110", -- t[14] = 0
      "000" when "0000000001111", -- t[15] = 0
      "000" when "0000000010000", -- t[16] = 0
      "000" when "0000000010001", -- t[17] = 0
      "000" when "0000000010010", -- t[18] = 0
      "000" when "0000000010011", -- t[19] = 0
      "000" when "0000000010100", -- t[20] = 0
      "000" when "0000000010101", -- t[21] = 0
      "000" when "0000000010110", -- t[22] = 0
      "000" when "0000000010111", -- t[23] = 0
      "000" when "0000000011000", -- t[24] = 0
      "000" when "0000000011001", -- t[25] = 0
      "000" when "0000000011010", -- t[26] = 0
      "000" when "0000000011011", -- t[27] = 0
      "000" when "0000000011100", -- t[28] = 0
      "000" when "0000000011101", -- t[29] = 0
      "000" when "0000000011110", -- t[30] = 0
      "000" when "0000000011111", -- t[31] = 0
      "000" when "0000000100000", -- t[32] = 0
      "000" when "0000000100001", -- t[33] = 0
      "000" when "0000000100010", -- t[34] = 0
      "000" when "0000000100011", -- t[35] = 0
      "000" when "0000000100100", -- t[36] = 0
      "000" when "0000000100101", -- t[37] = 0
      "000" when "0000000100110", -- t[38] = 0
      "000" when "0000000100111", -- t[39] = 0
      "000" when "0000000101000", -- t[40] = 0
      "000" when "0000000101001", -- t[41] = 0
      "000" when "0000000101010", -- t[42] = 0
      "000" when "0000000101011", -- t[43] = 0
      "000" when "0000000101100", -- t[44] = 0
      "000" when "0000000101101", -- t[45] = 0
      "000" when "0000000101110", -- t[46] = 0
      "000" when "0000000101111", -- t[47] = 0
      "000" when "0000000110000", -- t[48] = 0
      "000" when "0000000110001", -- t[49] = 0
      "000" when "0000000110010", -- t[50] = 0
      "000" when "0000000110011", -- t[51] = 0
      "000" when "0000000110100", -- t[52] = 0
      "000" when "0000000110101", -- t[53] = 0
      "000" when "0000000110110", -- t[54] = 0
      "000" when "0000000110111", -- t[55] = 0
      "000" when "0000000111000", -- t[56] = 0
      "000" when "0000000111001", -- t[57] = 0
      "000" when "0000000111010", -- t[58] = 0
      "000" when "0000000111011", -- t[59] = 0
      "000" when "0000000111100", -- t[60] = 0
      "000" when "0000000111101", -- t[61] = 0
      "000" when "0000000111110", -- t[62] = 0
      "000" when "0000000111111", -- t[63] = 0
      "000" when "0000001000000", -- t[64] = 0
      "000" when "0000001000001", -- t[65] = 0
      "000" when "0000001000010", -- t[66] = 0
      "000" when "0000001000011", -- t[67] = 0
      "000" when "0000001000100", -- t[68] = 0
      "000" when "0000001000101", -- t[69] = 0
      "000" when "0000001000110", -- t[70] = 0
      "000" when "0000001000111", -- t[71] = 0
      "000" when "0000001001000", -- t[72] = 0
      "000" when "0000001001001", -- t[73] = 0
      "000" when "0000001001010", -- t[74] = 0
      "000" when "0000001001011", -- t[75] = 0
      "000" when "0000001001100", -- t[76] = 0
      "000" when "0000001001101", -- t[77] = 0
      "000" when "0000001001110", -- t[78] = 0
      "000" when "0000001001111", -- t[79] = 0
      "000" when "0000001010000", -- t[80] = 0
      "000" when "0000001010001", -- t[81] = 0
      "000" when "0000001010010", -- t[82] = 0
      "000" when "0000001010011", -- t[83] = 0
      "000" when "0000001010100", -- t[84] = 0
      "000" when "0000001010101", -- t[85] = 0
      "000" when "0000001010110", -- t[86] = 0
      "000" when "0000001010111", -- t[87] = 0
      "000" when "0000001011000", -- t[88] = 0
      "000" when "0000001011001", -- t[89] = 0
      "000" when "0000001011010", -- t[90] = 0
      "000" when "0000001011011", -- t[91] = 0
      "000" when "0000001011100", -- t[92] = 0
      "000" when "0000001011101", -- t[93] = 0
      "000" when "0000001011110", -- t[94] = 0
      "000" when "0000001011111", -- t[95] = 0
      "000" when "0000001100000", -- t[96] = 0
      "000" when "0000001100001", -- t[97] = 0
      "000" when "0000001100010", -- t[98] = 0
      "000" when "0000001100011", -- t[99] = 0
      "000" when "0000001100100", -- t[100] = 0
      "000" when "0000001100101", -- t[101] = 0
      "000" when "0000001100110", -- t[102] = 0
      "000" when "0000001100111", -- t[103] = 0
      "000" when "0000001101000", -- t[104] = 0
      "000" when "0000001101001", -- t[105] = 0
      "000" when "0000001101010", -- t[106] = 0
      "000" when "0000001101011", -- t[107] = 0
      "000" when "0000001101100", -- t[108] = 0
      "000" when "0000001101101", -- t[109] = 0
      "000" when "0000001101110", -- t[110] = 0
      "000" when "0000001101111", -- t[111] = 0
      "000" when "0000001110000", -- t[112] = 0
      "000" when "0000001110001", -- t[113] = 0
      "000" when "0000001110010", -- t[114] = 0
      "000" when "0000001110011", -- t[115] = 0
      "000" when "0000001110100", -- t[116] = 0
      "000" when "0000001110101", -- t[117] = 0
      "000" when "0000001110110", -- t[118] = 0
      "000" when "0000001110111", -- t[119] = 0
      "000" when "0000001111000", -- t[120] = 0
      "000" when "0000001111001", -- t[121] = 0
      "000" when "0000001111010", -- t[122] = 0
      "000" when "0000001111011", -- t[123] = 0
      "000" when "0000001111100", -- t[124] = 0
      "000" when "0000001111101", -- t[125] = 0
      "000" when "0000001111110", -- t[126] = 0
      "000" when "0000001111111", -- t[127] = 0
      "000" when "0000010000000", -- t[128] = 0
      "000" when "0000010000001", -- t[129] = 0
      "000" when "0000010000010", -- t[130] = 0
      "000" when "0000010000011", -- t[131] = 0
      "000" when "0000010000100", -- t[132] = 0
      "000" when "0000010000101", -- t[133] = 0
      "000" when "0000010000110", -- t[134] = 0
      "000" when "0000010000111", -- t[135] = 0
      "000" when "0000010001000", -- t[136] = 0
      "000" when "0000010001001", -- t[137] = 0
      "000" when "0000010001010", -- t[138] = 0
      "000" when "0000010001011", -- t[139] = 0
      "000" when "0000010001100", -- t[140] = 0
      "000" when "0000010001101", -- t[141] = 0
      "000" when "0000010001110", -- t[142] = 0
      "000" when "0000010001111", -- t[143] = 0
      "000" when "0000010010000", -- t[144] = 0
      "000" when "0000010010001", -- t[145] = 0
      "000" when "0000010010010", -- t[146] = 0
      "000" when "0000010010011", -- t[147] = 0
      "000" when "0000010010100", -- t[148] = 0
      "000" when "0000010010101", -- t[149] = 0
      "000" when "0000010010110", -- t[150] = 0
      "000" when "0000010010111", -- t[151] = 0
      "000" when "0000010011000", -- t[152] = 0
      "000" when "0000010011001", -- t[153] = 0
      "000" when "0000010011010", -- t[154] = 0
      "000" when "0000010011011", -- t[155] = 0
      "000" when "0000010011100", -- t[156] = 0
      "000" when "0000010011101", -- t[157] = 0
      "000" when "0000010011110", -- t[158] = 0
      "000" when "0000010011111", -- t[159] = 0
      "000" when "0000010100000", -- t[160] = 0
      "000" when "0000010100001", -- t[161] = 0
      "000" when "0000010100010", -- t[162] = 0
      "000" when "0000010100011", -- t[163] = 0
      "000" when "0000010100100", -- t[164] = 0
      "000" when "0000010100101", -- t[165] = 0
      "000" when "0000010100110", -- t[166] = 0
      "000" when "0000010100111", -- t[167] = 0
      "000" when "0000010101000", -- t[168] = 0
      "000" when "0000010101001", -- t[169] = 0
      "000" when "0000010101010", -- t[170] = 0
      "000" when "0000010101011", -- t[171] = 0
      "000" when "0000010101100", -- t[172] = 0
      "000" when "0000010101101", -- t[173] = 0
      "000" when "0000010101110", -- t[174] = 0
      "000" when "0000010101111", -- t[175] = 0
      "000" when "0000010110000", -- t[176] = 0
      "000" when "0000010110001", -- t[177] = 0
      "000" when "0000010110010", -- t[178] = 0
      "000" when "0000010110011", -- t[179] = 0
      "000" when "0000010110100", -- t[180] = 0
      "000" when "0000010110101", -- t[181] = 0
      "000" when "0000010110110", -- t[182] = 0
      "000" when "0000010110111", -- t[183] = 0
      "000" when "0000010111000", -- t[184] = 0
      "000" when "0000010111001", -- t[185] = 0
      "000" when "0000010111010", -- t[186] = 0
      "000" when "0000010111011", -- t[187] = 0
      "000" when "0000010111100", -- t[188] = 0
      "000" when "0000010111101", -- t[189] = 0
      "000" when "0000010111110", -- t[190] = 0
      "000" when "0000010111111", -- t[191] = 0
      "000" when "0000011000000", -- t[192] = 0
      "000" when "0000011000001", -- t[193] = 0
      "000" when "0000011000010", -- t[194] = 0
      "000" when "0000011000011", -- t[195] = 0
      "000" when "0000011000100", -- t[196] = 0
      "000" when "0000011000101", -- t[197] = 0
      "000" when "0000011000110", -- t[198] = 0
      "000" when "0000011000111", -- t[199] = 0
      "000" when "0000011001000", -- t[200] = 0
      "000" when "0000011001001", -- t[201] = 0
      "000" when "0000011001010", -- t[202] = 0
      "000" when "0000011001011", -- t[203] = 0
      "000" when "0000011001100", -- t[204] = 0
      "000" when "0000011001101", -- t[205] = 0
      "000" when "0000011001110", -- t[206] = 0
      "000" when "0000011001111", -- t[207] = 0
      "000" when "0000011010000", -- t[208] = 0
      "000" when "0000011010001", -- t[209] = 0
      "000" when "0000011010010", -- t[210] = 0
      "000" when "0000011010011", -- t[211] = 0
      "000" when "0000011010100", -- t[212] = 0
      "000" when "0000011010101", -- t[213] = 0
      "000" when "0000011010110", -- t[214] = 0
      "000" when "0000011010111", -- t[215] = 0
      "000" when "0000011011000", -- t[216] = 0
      "000" when "0000011011001", -- t[217] = 0
      "000" when "0000011011010", -- t[218] = 0
      "000" when "0000011011011", -- t[219] = 0
      "000" when "0000011011100", -- t[220] = 0
      "000" when "0000011011101", -- t[221] = 0
      "000" when "0000011011110", -- t[222] = 0
      "000" when "0000011011111", -- t[223] = 0
      "000" when "0000011100000", -- t[224] = 0
      "000" when "0000011100001", -- t[225] = 0
      "000" when "0000011100010", -- t[226] = 0
      "000" when "0000011100011", -- t[227] = 0
      "000" when "0000011100100", -- t[228] = 0
      "000" when "0000011100101", -- t[229] = 0
      "000" when "0000011100110", -- t[230] = 0
      "000" when "0000011100111", -- t[231] = 0
      "000" when "0000011101000", -- t[232] = 0
      "000" when "0000011101001", -- t[233] = 0
      "000" when "0000011101010", -- t[234] = 0
      "000" when "0000011101011", -- t[235] = 0
      "000" when "0000011101100", -- t[236] = 0
      "000" when "0000011101101", -- t[237] = 0
      "000" when "0000011101110", -- t[238] = 0
      "000" when "0000011101111", -- t[239] = 0
      "000" when "0000011110000", -- t[240] = 0
      "000" when "0000011110001", -- t[241] = 0
      "000" when "0000011110010", -- t[242] = 0
      "000" when "0000011110011", -- t[243] = 0
      "000" when "0000011110100", -- t[244] = 0
      "000" when "0000011110101", -- t[245] = 0
      "000" when "0000011110110", -- t[246] = 0
      "000" when "0000011110111", -- t[247] = 0
      "000" when "0000011111000", -- t[248] = 0
      "000" when "0000011111001", -- t[249] = 0
      "000" when "0000011111010", -- t[250] = 0
      "000" when "0000011111011", -- t[251] = 0
      "000" when "0000011111100", -- t[252] = 0
      "000" when "0000011111101", -- t[253] = 0
      "000" when "0000011111110", -- t[254] = 0
      "000" when "0000011111111", -- t[255] = 0
      "000" when "0000100000000", -- t[256] = 0
      "000" when "0000100000001", -- t[257] = 0
      "000" when "0000100000010", -- t[258] = 0
      "000" when "0000100000011", -- t[259] = 0
      "000" when "0000100000100", -- t[260] = 0
      "000" when "0000100000101", -- t[261] = 0
      "000" when "0000100000110", -- t[262] = 0
      "000" when "0000100000111", -- t[263] = 0
      "000" when "0000100001000", -- t[264] = 0
      "000" when "0000100001001", -- t[265] = 0
      "000" when "0000100001010", -- t[266] = 0
      "000" when "0000100001011", -- t[267] = 0
      "000" when "0000100001100", -- t[268] = 0
      "000" when "0000100001101", -- t[269] = 0
      "000" when "0000100001110", -- t[270] = 0
      "000" when "0000100001111", -- t[271] = 0
      "000" when "0000100010000", -- t[272] = 0
      "000" when "0000100010001", -- t[273] = 0
      "000" when "0000100010010", -- t[274] = 0
      "000" when "0000100010011", -- t[275] = 0
      "000" when "0000100010100", -- t[276] = 0
      "000" when "0000100010101", -- t[277] = 0
      "000" when "0000100010110", -- t[278] = 0
      "000" when "0000100010111", -- t[279] = 0
      "000" when "0000100011000", -- t[280] = 0
      "000" when "0000100011001", -- t[281] = 0
      "000" when "0000100011010", -- t[282] = 0
      "000" when "0000100011011", -- t[283] = 0
      "000" when "0000100011100", -- t[284] = 0
      "000" when "0000100011101", -- t[285] = 0
      "000" when "0000100011110", -- t[286] = 0
      "000" when "0000100011111", -- t[287] = 0
      "000" when "0000100100000", -- t[288] = 0
      "000" when "0000100100001", -- t[289] = 0
      "000" when "0000100100010", -- t[290] = 0
      "000" when "0000100100011", -- t[291] = 0
      "000" when "0000100100100", -- t[292] = 0
      "000" when "0000100100101", -- t[293] = 0
      "000" when "0000100100110", -- t[294] = 0
      "000" when "0000100100111", -- t[295] = 0
      "000" when "0000100101000", -- t[296] = 0
      "000" when "0000100101001", -- t[297] = 0
      "000" when "0000100101010", -- t[298] = 0
      "000" when "0000100101011", -- t[299] = 0
      "000" when "0000100101100", -- t[300] = 0
      "000" when "0000100101101", -- t[301] = 0
      "000" when "0000100101110", -- t[302] = 0
      "000" when "0000100101111", -- t[303] = 0
      "000" when "0000100110000", -- t[304] = 0
      "000" when "0000100110001", -- t[305] = 0
      "000" when "0000100110010", -- t[306] = 0
      "000" when "0000100110011", -- t[307] = 0
      "000" when "0000100110100", -- t[308] = 0
      "000" when "0000100110101", -- t[309] = 0
      "000" when "0000100110110", -- t[310] = 0
      "000" when "0000100110111", -- t[311] = 0
      "000" when "0000100111000", -- t[312] = 0
      "000" when "0000100111001", -- t[313] = 0
      "000" when "0000100111010", -- t[314] = 0
      "000" when "0000100111011", -- t[315] = 0
      "000" when "0000100111100", -- t[316] = 0
      "000" when "0000100111101", -- t[317] = 0
      "000" when "0000100111110", -- t[318] = 0
      "000" when "0000100111111", -- t[319] = 0
      "000" when "0000101000000", -- t[320] = 0
      "000" when "0000101000001", -- t[321] = 0
      "000" when "0000101000010", -- t[322] = 0
      "000" when "0000101000011", -- t[323] = 0
      "000" when "0000101000100", -- t[324] = 0
      "000" when "0000101000101", -- t[325] = 0
      "000" when "0000101000110", -- t[326] = 0
      "000" when "0000101000111", -- t[327] = 0
      "000" when "0000101001000", -- t[328] = 0
      "000" when "0000101001001", -- t[329] = 0
      "000" when "0000101001010", -- t[330] = 0
      "000" when "0000101001011", -- t[331] = 0
      "000" when "0000101001100", -- t[332] = 0
      "000" when "0000101001101", -- t[333] = 0
      "000" when "0000101001110", -- t[334] = 0
      "000" when "0000101001111", -- t[335] = 0
      "000" when "0000101010000", -- t[336] = 0
      "000" when "0000101010001", -- t[337] = 0
      "000" when "0000101010010", -- t[338] = 0
      "000" when "0000101010011", -- t[339] = 0
      "000" when "0000101010100", -- t[340] = 0
      "000" when "0000101010101", -- t[341] = 0
      "000" when "0000101010110", -- t[342] = 0
      "000" when "0000101010111", -- t[343] = 0
      "000" when "0000101011000", -- t[344] = 0
      "000" when "0000101011001", -- t[345] = 0
      "000" when "0000101011010", -- t[346] = 0
      "000" when "0000101011011", -- t[347] = 0
      "000" when "0000101011100", -- t[348] = 0
      "000" when "0000101011101", -- t[349] = 0
      "000" when "0000101011110", -- t[350] = 0
      "000" when "0000101011111", -- t[351] = 0
      "000" when "0000101100000", -- t[352] = 0
      "000" when "0000101100001", -- t[353] = 0
      "000" when "0000101100010", -- t[354] = 0
      "000" when "0000101100011", -- t[355] = 0
      "000" when "0000101100100", -- t[356] = 0
      "000" when "0000101100101", -- t[357] = 0
      "000" when "0000101100110", -- t[358] = 0
      "000" when "0000101100111", -- t[359] = 0
      "000" when "0000101101000", -- t[360] = 0
      "000" when "0000101101001", -- t[361] = 0
      "000" when "0000101101010", -- t[362] = 0
      "000" when "0000101101011", -- t[363] = 0
      "000" when "0000101101100", -- t[364] = 0
      "000" when "0000101101101", -- t[365] = 0
      "000" when "0000101101110", -- t[366] = 0
      "000" when "0000101101111", -- t[367] = 0
      "000" when "0000101110000", -- t[368] = 0
      "000" when "0000101110001", -- t[369] = 0
      "000" when "0000101110010", -- t[370] = 0
      "000" when "0000101110011", -- t[371] = 0
      "000" when "0000101110100", -- t[372] = 0
      "000" when "0000101110101", -- t[373] = 0
      "000" when "0000101110110", -- t[374] = 0
      "000" when "0000101110111", -- t[375] = 0
      "000" when "0000101111000", -- t[376] = 0
      "000" when "0000101111001", -- t[377] = 0
      "000" when "0000101111010", -- t[378] = 0
      "000" when "0000101111011", -- t[379] = 0
      "000" when "0000101111100", -- t[380] = 0
      "000" when "0000101111101", -- t[381] = 0
      "000" when "0000101111110", -- t[382] = 0
      "000" when "0000101111111", -- t[383] = 0
      "000" when "0000110000000", -- t[384] = 0
      "000" when "0000110000001", -- t[385] = 0
      "000" when "0000110000010", -- t[386] = 0
      "000" when "0000110000011", -- t[387] = 0
      "000" when "0000110000100", -- t[388] = 0
      "000" when "0000110000101", -- t[389] = 0
      "000" when "0000110000110", -- t[390] = 0
      "000" when "0000110000111", -- t[391] = 0
      "000" when "0000110001000", -- t[392] = 0
      "000" when "0000110001001", -- t[393] = 0
      "000" when "0000110001010", -- t[394] = 0
      "000" when "0000110001011", -- t[395] = 0
      "000" when "0000110001100", -- t[396] = 0
      "000" when "0000110001101", -- t[397] = 0
      "000" when "0000110001110", -- t[398] = 0
      "000" when "0000110001111", -- t[399] = 0
      "000" when "0000110010000", -- t[400] = 0
      "000" when "0000110010001", -- t[401] = 0
      "000" when "0000110010010", -- t[402] = 0
      "000" when "0000110010011", -- t[403] = 0
      "000" when "0000110010100", -- t[404] = 0
      "000" when "0000110010101", -- t[405] = 0
      "000" when "0000110010110", -- t[406] = 0
      "000" when "0000110010111", -- t[407] = 0
      "000" when "0000110011000", -- t[408] = 0
      "000" when "0000110011001", -- t[409] = 0
      "000" when "0000110011010", -- t[410] = 0
      "000" when "0000110011011", -- t[411] = 0
      "000" when "0000110011100", -- t[412] = 0
      "000" when "0000110011101", -- t[413] = 0
      "000" when "0000110011110", -- t[414] = 0
      "000" when "0000110011111", -- t[415] = 0
      "000" when "0000110100000", -- t[416] = 0
      "000" when "0000110100001", -- t[417] = 0
      "000" when "0000110100010", -- t[418] = 0
      "000" when "0000110100011", -- t[419] = 0
      "000" when "0000110100100", -- t[420] = 0
      "000" when "0000110100101", -- t[421] = 0
      "000" when "0000110100110", -- t[422] = 0
      "000" when "0000110100111", -- t[423] = 0
      "000" when "0000110101000", -- t[424] = 0
      "000" when "0000110101001", -- t[425] = 0
      "000" when "0000110101010", -- t[426] = 0
      "000" when "0000110101011", -- t[427] = 0
      "000" when "0000110101100", -- t[428] = 0
      "000" when "0000110101101", -- t[429] = 0
      "000" when "0000110101110", -- t[430] = 0
      "000" when "0000110101111", -- t[431] = 0
      "000" when "0000110110000", -- t[432] = 0
      "000" when "0000110110001", -- t[433] = 0
      "000" when "0000110110010", -- t[434] = 0
      "000" when "0000110110011", -- t[435] = 0
      "000" when "0000110110100", -- t[436] = 0
      "000" when "0000110110101", -- t[437] = 0
      "000" when "0000110110110", -- t[438] = 0
      "000" when "0000110110111", -- t[439] = 0
      "000" when "0000110111000", -- t[440] = 0
      "000" when "0000110111001", -- t[441] = 0
      "000" when "0000110111010", -- t[442] = 0
      "000" when "0000110111011", -- t[443] = 0
      "000" when "0000110111100", -- t[444] = 0
      "000" when "0000110111101", -- t[445] = 0
      "000" when "0000110111110", -- t[446] = 0
      "000" when "0000110111111", -- t[447] = 0
      "000" when "0000111000000", -- t[448] = 0
      "000" when "0000111000001", -- t[449] = 0
      "000" when "0000111000010", -- t[450] = 0
      "000" when "0000111000011", -- t[451] = 0
      "000" when "0000111000100", -- t[452] = 0
      "000" when "0000111000101", -- t[453] = 0
      "000" when "0000111000110", -- t[454] = 0
      "000" when "0000111000111", -- t[455] = 0
      "000" when "0000111001000", -- t[456] = 0
      "000" when "0000111001001", -- t[457] = 0
      "000" when "0000111001010", -- t[458] = 0
      "000" when "0000111001011", -- t[459] = 0
      "000" when "0000111001100", -- t[460] = 0
      "000" when "0000111001101", -- t[461] = 0
      "000" when "0000111001110", -- t[462] = 0
      "000" when "0000111001111", -- t[463] = 0
      "000" when "0000111010000", -- t[464] = 0
      "000" when "0000111010001", -- t[465] = 0
      "000" when "0000111010010", -- t[466] = 0
      "000" when "0000111010011", -- t[467] = 0
      "000" when "0000111010100", -- t[468] = 0
      "000" when "0000111010101", -- t[469] = 0
      "000" when "0000111010110", -- t[470] = 0
      "000" when "0000111010111", -- t[471] = 0
      "000" when "0000111011000", -- t[472] = 0
      "000" when "0000111011001", -- t[473] = 0
      "000" when "0000111011010", -- t[474] = 0
      "000" when "0000111011011", -- t[475] = 0
      "000" when "0000111011100", -- t[476] = 0
      "000" when "0000111011101", -- t[477] = 0
      "000" when "0000111011110", -- t[478] = 0
      "000" when "0000111011111", -- t[479] = 0
      "000" when "0000111100000", -- t[480] = 0
      "000" when "0000111100001", -- t[481] = 0
      "000" when "0000111100010", -- t[482] = 0
      "000" when "0000111100011", -- t[483] = 0
      "000" when "0000111100100", -- t[484] = 0
      "000" when "0000111100101", -- t[485] = 0
      "000" when "0000111100110", -- t[486] = 0
      "000" when "0000111100111", -- t[487] = 0
      "000" when "0000111101000", -- t[488] = 0
      "000" when "0000111101001", -- t[489] = 0
      "000" when "0000111101010", -- t[490] = 0
      "000" when "0000111101011", -- t[491] = 0
      "000" when "0000111101100", -- t[492] = 0
      "000" when "0000111101101", -- t[493] = 0
      "000" when "0000111101110", -- t[494] = 0
      "000" when "0000111101111", -- t[495] = 0
      "000" when "0000111110000", -- t[496] = 0
      "000" when "0000111110001", -- t[497] = 0
      "000" when "0000111110010", -- t[498] = 0
      "000" when "0000111110011", -- t[499] = 0
      "000" when "0000111110100", -- t[500] = 0
      "000" when "0000111110101", -- t[501] = 0
      "000" when "0000111110110", -- t[502] = 0
      "000" when "0000111110111", -- t[503] = 0
      "000" when "0000111111000", -- t[504] = 0
      "000" when "0000111111001", -- t[505] = 0
      "000" when "0000111111010", -- t[506] = 0
      "000" when "0000111111011", -- t[507] = 0
      "000" when "0000111111100", -- t[508] = 0
      "000" when "0000111111101", -- t[509] = 0
      "000" when "0000111111110", -- t[510] = 0
      "000" when "0000111111111", -- t[511] = 0
      "000" when "0001000000000", -- t[512] = 0
      "000" when "0001000000001", -- t[513] = 0
      "000" when "0001000000010", -- t[514] = 0
      "000" when "0001000000011", -- t[515] = 0
      "000" when "0001000000100", -- t[516] = 0
      "000" when "0001000000101", -- t[517] = 0
      "000" when "0001000000110", -- t[518] = 0
      "000" when "0001000000111", -- t[519] = 0
      "000" when "0001000001000", -- t[520] = 0
      "000" when "0001000001001", -- t[521] = 0
      "000" when "0001000001010", -- t[522] = 0
      "000" when "0001000001011", -- t[523] = 0
      "000" when "0001000001100", -- t[524] = 0
      "000" when "0001000001101", -- t[525] = 0
      "000" when "0001000001110", -- t[526] = 0
      "000" when "0001000001111", -- t[527] = 0
      "000" when "0001000010000", -- t[528] = 0
      "000" when "0001000010001", -- t[529] = 0
      "000" when "0001000010010", -- t[530] = 0
      "000" when "0001000010011", -- t[531] = 0
      "000" when "0001000010100", -- t[532] = 0
      "000" when "0001000010101", -- t[533] = 0
      "000" when "0001000010110", -- t[534] = 0
      "000" when "0001000010111", -- t[535] = 0
      "000" when "0001000011000", -- t[536] = 0
      "000" when "0001000011001", -- t[537] = 0
      "000" when "0001000011010", -- t[538] = 0
      "000" when "0001000011011", -- t[539] = 0
      "000" when "0001000011100", -- t[540] = 0
      "000" when "0001000011101", -- t[541] = 0
      "000" when "0001000011110", -- t[542] = 0
      "000" when "0001000011111", -- t[543] = 0
      "000" when "0001000100000", -- t[544] = 0
      "000" when "0001000100001", -- t[545] = 0
      "000" when "0001000100010", -- t[546] = 0
      "000" when "0001000100011", -- t[547] = 0
      "000" when "0001000100100", -- t[548] = 0
      "000" when "0001000100101", -- t[549] = 0
      "000" when "0001000100110", -- t[550] = 0
      "000" when "0001000100111", -- t[551] = 0
      "000" when "0001000101000", -- t[552] = 0
      "000" when "0001000101001", -- t[553] = 0
      "000" when "0001000101010", -- t[554] = 0
      "000" when "0001000101011", -- t[555] = 0
      "000" when "0001000101100", -- t[556] = 0
      "000" when "0001000101101", -- t[557] = 0
      "000" when "0001000101110", -- t[558] = 0
      "000" when "0001000101111", -- t[559] = 0
      "000" when "0001000110000", -- t[560] = 0
      "000" when "0001000110001", -- t[561] = 0
      "000" when "0001000110010", -- t[562] = 0
      "000" when "0001000110011", -- t[563] = 0
      "000" when "0001000110100", -- t[564] = 0
      "000" when "0001000110101", -- t[565] = 0
      "000" when "0001000110110", -- t[566] = 0
      "000" when "0001000110111", -- t[567] = 0
      "000" when "0001000111000", -- t[568] = 0
      "000" when "0001000111001", -- t[569] = 0
      "000" when "0001000111010", -- t[570] = 0
      "000" when "0001000111011", -- t[571] = 0
      "000" when "0001000111100", -- t[572] = 0
      "000" when "0001000111101", -- t[573] = 0
      "000" when "0001000111110", -- t[574] = 0
      "000" when "0001000111111", -- t[575] = 0
      "000" when "0001001000000", -- t[576] = 0
      "000" when "0001001000001", -- t[577] = 0
      "000" when "0001001000010", -- t[578] = 0
      "000" when "0001001000011", -- t[579] = 0
      "000" when "0001001000100", -- t[580] = 0
      "000" when "0001001000101", -- t[581] = 0
      "000" when "0001001000110", -- t[582] = 0
      "000" when "0001001000111", -- t[583] = 0
      "000" when "0001001001000", -- t[584] = 0
      "000" when "0001001001001", -- t[585] = 0
      "000" when "0001001001010", -- t[586] = 0
      "000" when "0001001001011", -- t[587] = 0
      "000" when "0001001001100", -- t[588] = 0
      "000" when "0001001001101", -- t[589] = 0
      "000" when "0001001001110", -- t[590] = 0
      "000" when "0001001001111", -- t[591] = 0
      "000" when "0001001010000", -- t[592] = 0
      "000" when "0001001010001", -- t[593] = 0
      "000" when "0001001010010", -- t[594] = 0
      "000" when "0001001010011", -- t[595] = 0
      "000" when "0001001010100", -- t[596] = 0
      "000" when "0001001010101", -- t[597] = 0
      "000" when "0001001010110", -- t[598] = 0
      "000" when "0001001010111", -- t[599] = 0
      "000" when "0001001011000", -- t[600] = 0
      "000" when "0001001011001", -- t[601] = 0
      "000" when "0001001011010", -- t[602] = 0
      "000" when "0001001011011", -- t[603] = 0
      "000" when "0001001011100", -- t[604] = 0
      "000" when "0001001011101", -- t[605] = 0
      "000" when "0001001011110", -- t[606] = 0
      "000" when "0001001011111", -- t[607] = 0
      "000" when "0001001100000", -- t[608] = 0
      "000" when "0001001100001", -- t[609] = 0
      "000" when "0001001100010", -- t[610] = 0
      "000" when "0001001100011", -- t[611] = 0
      "000" when "0001001100100", -- t[612] = 0
      "000" when "0001001100101", -- t[613] = 0
      "000" when "0001001100110", -- t[614] = 0
      "000" when "0001001100111", -- t[615] = 0
      "000" when "0001001101000", -- t[616] = 0
      "000" when "0001001101001", -- t[617] = 0
      "000" when "0001001101010", -- t[618] = 0
      "000" when "0001001101011", -- t[619] = 0
      "000" when "0001001101100", -- t[620] = 0
      "000" when "0001001101101", -- t[621] = 0
      "000" when "0001001101110", -- t[622] = 0
      "000" when "0001001101111", -- t[623] = 0
      "000" when "0001001110000", -- t[624] = 0
      "000" when "0001001110001", -- t[625] = 0
      "000" when "0001001110010", -- t[626] = 0
      "000" when "0001001110011", -- t[627] = 0
      "000" when "0001001110100", -- t[628] = 0
      "000" when "0001001110101", -- t[629] = 0
      "000" when "0001001110110", -- t[630] = 0
      "000" when "0001001110111", -- t[631] = 0
      "000" when "0001001111000", -- t[632] = 0
      "000" when "0001001111001", -- t[633] = 0
      "000" when "0001001111010", -- t[634] = 0
      "000" when "0001001111011", -- t[635] = 0
      "000" when "0001001111100", -- t[636] = 0
      "000" when "0001001111101", -- t[637] = 0
      "000" when "0001001111110", -- t[638] = 0
      "000" when "0001001111111", -- t[639] = 0
      "000" when "0001010000000", -- t[640] = 0
      "000" when "0001010000001", -- t[641] = 0
      "000" when "0001010000010", -- t[642] = 0
      "000" when "0001010000011", -- t[643] = 0
      "000" when "0001010000100", -- t[644] = 0
      "000" when "0001010000101", -- t[645] = 0
      "000" when "0001010000110", -- t[646] = 0
      "000" when "0001010000111", -- t[647] = 0
      "000" when "0001010001000", -- t[648] = 0
      "000" when "0001010001001", -- t[649] = 0
      "000" when "0001010001010", -- t[650] = 0
      "000" when "0001010001011", -- t[651] = 0
      "000" when "0001010001100", -- t[652] = 0
      "000" when "0001010001101", -- t[653] = 0
      "000" when "0001010001110", -- t[654] = 0
      "000" when "0001010001111", -- t[655] = 0
      "000" when "0001010010000", -- t[656] = 0
      "000" when "0001010010001", -- t[657] = 0
      "000" when "0001010010010", -- t[658] = 0
      "000" when "0001010010011", -- t[659] = 0
      "000" when "0001010010100", -- t[660] = 0
      "000" when "0001010010101", -- t[661] = 0
      "000" when "0001010010110", -- t[662] = 0
      "000" when "0001010010111", -- t[663] = 0
      "000" when "0001010011000", -- t[664] = 0
      "000" when "0001010011001", -- t[665] = 0
      "000" when "0001010011010", -- t[666] = 0
      "000" when "0001010011011", -- t[667] = 0
      "000" when "0001010011100", -- t[668] = 0
      "000" when "0001010011101", -- t[669] = 0
      "000" when "0001010011110", -- t[670] = 0
      "000" when "0001010011111", -- t[671] = 0
      "000" when "0001010100000", -- t[672] = 0
      "000" when "0001010100001", -- t[673] = 0
      "000" when "0001010100010", -- t[674] = 0
      "000" when "0001010100011", -- t[675] = 0
      "000" when "0001010100100", -- t[676] = 0
      "000" when "0001010100101", -- t[677] = 0
      "000" when "0001010100110", -- t[678] = 0
      "000" when "0001010100111", -- t[679] = 0
      "000" when "0001010101000", -- t[680] = 0
      "000" when "0001010101001", -- t[681] = 0
      "000" when "0001010101010", -- t[682] = 0
      "000" when "0001010101011", -- t[683] = 0
      "000" when "0001010101100", -- t[684] = 0
      "000" when "0001010101101", -- t[685] = 0
      "000" when "0001010101110", -- t[686] = 0
      "000" when "0001010101111", -- t[687] = 0
      "000" when "0001010110000", -- t[688] = 0
      "000" when "0001010110001", -- t[689] = 0
      "000" when "0001010110010", -- t[690] = 0
      "000" when "0001010110011", -- t[691] = 0
      "000" when "0001010110100", -- t[692] = 0
      "000" when "0001010110101", -- t[693] = 0
      "000" when "0001010110110", -- t[694] = 0
      "000" when "0001010110111", -- t[695] = 0
      "000" when "0001010111000", -- t[696] = 0
      "000" when "0001010111001", -- t[697] = 0
      "000" when "0001010111010", -- t[698] = 0
      "000" when "0001010111011", -- t[699] = 0
      "000" when "0001010111100", -- t[700] = 0
      "000" when "0001010111101", -- t[701] = 0
      "000" when "0001010111110", -- t[702] = 0
      "000" when "0001010111111", -- t[703] = 0
      "000" when "0001011000000", -- t[704] = 0
      "000" when "0001011000001", -- t[705] = 0
      "000" when "0001011000010", -- t[706] = 0
      "000" when "0001011000011", -- t[707] = 0
      "000" when "0001011000100", -- t[708] = 0
      "000" when "0001011000101", -- t[709] = 0
      "000" when "0001011000110", -- t[710] = 0
      "000" when "0001011000111", -- t[711] = 0
      "000" when "0001011001000", -- t[712] = 0
      "000" when "0001011001001", -- t[713] = 0
      "000" when "0001011001010", -- t[714] = 0
      "000" when "0001011001011", -- t[715] = 0
      "000" when "0001011001100", -- t[716] = 0
      "000" when "0001011001101", -- t[717] = 0
      "000" when "0001011001110", -- t[718] = 0
      "000" when "0001011001111", -- t[719] = 0
      "000" when "0001011010000", -- t[720] = 0
      "000" when "0001011010001", -- t[721] = 0
      "000" when "0001011010010", -- t[722] = 0
      "000" when "0001011010011", -- t[723] = 0
      "000" when "0001011010100", -- t[724] = 0
      "000" when "0001011010101", -- t[725] = 0
      "000" when "0001011010110", -- t[726] = 0
      "000" when "0001011010111", -- t[727] = 0
      "000" when "0001011011000", -- t[728] = 0
      "000" when "0001011011001", -- t[729] = 0
      "000" when "0001011011010", -- t[730] = 0
      "000" when "0001011011011", -- t[731] = 0
      "000" when "0001011011100", -- t[732] = 0
      "000" when "0001011011101", -- t[733] = 0
      "000" when "0001011011110", -- t[734] = 0
      "000" when "0001011011111", -- t[735] = 0
      "000" when "0001011100000", -- t[736] = 0
      "000" when "0001011100001", -- t[737] = 0
      "000" when "0001011100010", -- t[738] = 0
      "000" when "0001011100011", -- t[739] = 0
      "000" when "0001011100100", -- t[740] = 0
      "000" when "0001011100101", -- t[741] = 0
      "000" when "0001011100110", -- t[742] = 0
      "000" when "0001011100111", -- t[743] = 0
      "000" when "0001011101000", -- t[744] = 0
      "000" when "0001011101001", -- t[745] = 0
      "000" when "0001011101010", -- t[746] = 0
      "000" when "0001011101011", -- t[747] = 0
      "000" when "0001011101100", -- t[748] = 0
      "000" when "0001011101101", -- t[749] = 0
      "000" when "0001011101110", -- t[750] = 0
      "000" when "0001011101111", -- t[751] = 0
      "000" when "0001011110000", -- t[752] = 0
      "000" when "0001011110001", -- t[753] = 0
      "000" when "0001011110010", -- t[754] = 0
      "000" when "0001011110011", -- t[755] = 0
      "000" when "0001011110100", -- t[756] = 0
      "000" when "0001011110101", -- t[757] = 0
      "000" when "0001011110110", -- t[758] = 0
      "000" when "0001011110111", -- t[759] = 0
      "000" when "0001011111000", -- t[760] = 0
      "000" when "0001011111001", -- t[761] = 0
      "000" when "0001011111010", -- t[762] = 0
      "000" when "0001011111011", -- t[763] = 0
      "000" when "0001011111100", -- t[764] = 0
      "000" when "0001011111101", -- t[765] = 0
      "000" when "0001011111110", -- t[766] = 0
      "000" when "0001011111111", -- t[767] = 0
      "000" when "0001100000000", -- t[768] = 0
      "000" when "0001100000001", -- t[769] = 0
      "000" when "0001100000010", -- t[770] = 0
      "000" when "0001100000011", -- t[771] = 0
      "000" when "0001100000100", -- t[772] = 0
      "000" when "0001100000101", -- t[773] = 0
      "000" when "0001100000110", -- t[774] = 0
      "000" when "0001100000111", -- t[775] = 0
      "000" when "0001100001000", -- t[776] = 0
      "000" when "0001100001001", -- t[777] = 0
      "000" when "0001100001010", -- t[778] = 0
      "000" when "0001100001011", -- t[779] = 0
      "000" when "0001100001100", -- t[780] = 0
      "000" when "0001100001101", -- t[781] = 0
      "000" when "0001100001110", -- t[782] = 0
      "000" when "0001100001111", -- t[783] = 0
      "000" when "0001100010000", -- t[784] = 0
      "000" when "0001100010001", -- t[785] = 0
      "000" when "0001100010010", -- t[786] = 0
      "000" when "0001100010011", -- t[787] = 0
      "000" when "0001100010100", -- t[788] = 0
      "000" when "0001100010101", -- t[789] = 0
      "000" when "0001100010110", -- t[790] = 0
      "000" when "0001100010111", -- t[791] = 0
      "000" when "0001100011000", -- t[792] = 0
      "000" when "0001100011001", -- t[793] = 0
      "000" when "0001100011010", -- t[794] = 0
      "000" when "0001100011011", -- t[795] = 0
      "000" when "0001100011100", -- t[796] = 0
      "000" when "0001100011101", -- t[797] = 0
      "000" when "0001100011110", -- t[798] = 0
      "000" when "0001100011111", -- t[799] = 0
      "000" when "0001100100000", -- t[800] = 0
      "000" when "0001100100001", -- t[801] = 0
      "000" when "0001100100010", -- t[802] = 0
      "000" when "0001100100011", -- t[803] = 0
      "000" when "0001100100100", -- t[804] = 0
      "000" when "0001100100101", -- t[805] = 0
      "000" when "0001100100110", -- t[806] = 0
      "000" when "0001100100111", -- t[807] = 0
      "000" when "0001100101000", -- t[808] = 0
      "000" when "0001100101001", -- t[809] = 0
      "000" when "0001100101010", -- t[810] = 0
      "000" when "0001100101011", -- t[811] = 0
      "000" when "0001100101100", -- t[812] = 0
      "000" when "0001100101101", -- t[813] = 0
      "000" when "0001100101110", -- t[814] = 0
      "000" when "0001100101111", -- t[815] = 0
      "000" when "0001100110000", -- t[816] = 0
      "000" when "0001100110001", -- t[817] = 0
      "000" when "0001100110010", -- t[818] = 0
      "000" when "0001100110011", -- t[819] = 0
      "000" when "0001100110100", -- t[820] = 0
      "000" when "0001100110101", -- t[821] = 0
      "000" when "0001100110110", -- t[822] = 0
      "000" when "0001100110111", -- t[823] = 0
      "000" when "0001100111000", -- t[824] = 0
      "000" when "0001100111001", -- t[825] = 0
      "000" when "0001100111010", -- t[826] = 0
      "000" when "0001100111011", -- t[827] = 0
      "000" when "0001100111100", -- t[828] = 0
      "000" when "0001100111101", -- t[829] = 0
      "000" when "0001100111110", -- t[830] = 0
      "000" when "0001100111111", -- t[831] = 0
      "000" when "0001101000000", -- t[832] = 0
      "000" when "0001101000001", -- t[833] = 0
      "000" when "0001101000010", -- t[834] = 0
      "000" when "0001101000011", -- t[835] = 0
      "000" when "0001101000100", -- t[836] = 0
      "000" when "0001101000101", -- t[837] = 0
      "000" when "0001101000110", -- t[838] = 0
      "000" when "0001101000111", -- t[839] = 0
      "000" when "0001101001000", -- t[840] = 0
      "000" when "0001101001001", -- t[841] = 0
      "000" when "0001101001010", -- t[842] = 0
      "000" when "0001101001011", -- t[843] = 0
      "000" when "0001101001100", -- t[844] = 0
      "000" when "0001101001101", -- t[845] = 0
      "000" when "0001101001110", -- t[846] = 0
      "000" when "0001101001111", -- t[847] = 0
      "000" when "0001101010000", -- t[848] = 0
      "000" when "0001101010001", -- t[849] = 0
      "000" when "0001101010010", -- t[850] = 0
      "000" when "0001101010011", -- t[851] = 0
      "000" when "0001101010100", -- t[852] = 0
      "000" when "0001101010101", -- t[853] = 0
      "000" when "0001101010110", -- t[854] = 0
      "000" when "0001101010111", -- t[855] = 0
      "000" when "0001101011000", -- t[856] = 0
      "000" when "0001101011001", -- t[857] = 0
      "000" when "0001101011010", -- t[858] = 0
      "000" when "0001101011011", -- t[859] = 0
      "000" when "0001101011100", -- t[860] = 0
      "000" when "0001101011101", -- t[861] = 0
      "000" when "0001101011110", -- t[862] = 0
      "000" when "0001101011111", -- t[863] = 0
      "000" when "0001101100000", -- t[864] = 0
      "000" when "0001101100001", -- t[865] = 0
      "000" when "0001101100010", -- t[866] = 0
      "000" when "0001101100011", -- t[867] = 0
      "000" when "0001101100100", -- t[868] = 0
      "000" when "0001101100101", -- t[869] = 0
      "000" when "0001101100110", -- t[870] = 0
      "000" when "0001101100111", -- t[871] = 0
      "000" when "0001101101000", -- t[872] = 0
      "000" when "0001101101001", -- t[873] = 0
      "000" when "0001101101010", -- t[874] = 0
      "000" when "0001101101011", -- t[875] = 0
      "000" when "0001101101100", -- t[876] = 0
      "000" when "0001101101101", -- t[877] = 0
      "000" when "0001101101110", -- t[878] = 0
      "000" when "0001101101111", -- t[879] = 0
      "000" when "0001101110000", -- t[880] = 0
      "000" when "0001101110001", -- t[881] = 0
      "000" when "0001101110010", -- t[882] = 0
      "000" when "0001101110011", -- t[883] = 0
      "000" when "0001101110100", -- t[884] = 0
      "000" when "0001101110101", -- t[885] = 0
      "000" when "0001101110110", -- t[886] = 0
      "000" when "0001101110111", -- t[887] = 0
      "000" when "0001101111000", -- t[888] = 0
      "000" when "0001101111001", -- t[889] = 0
      "000" when "0001101111010", -- t[890] = 0
      "000" when "0001101111011", -- t[891] = 0
      "000" when "0001101111100", -- t[892] = 0
      "000" when "0001101111101", -- t[893] = 0
      "000" when "0001101111110", -- t[894] = 0
      "000" when "0001101111111", -- t[895] = 0
      "000" when "0001110000000", -- t[896] = 0
      "000" when "0001110000001", -- t[897] = 0
      "000" when "0001110000010", -- t[898] = 0
      "000" when "0001110000011", -- t[899] = 0
      "000" when "0001110000100", -- t[900] = 0
      "000" when "0001110000101", -- t[901] = 0
      "000" when "0001110000110", -- t[902] = 0
      "000" when "0001110000111", -- t[903] = 0
      "000" when "0001110001000", -- t[904] = 0
      "000" when "0001110001001", -- t[905] = 0
      "000" when "0001110001010", -- t[906] = 0
      "000" when "0001110001011", -- t[907] = 0
      "000" when "0001110001100", -- t[908] = 0
      "000" when "0001110001101", -- t[909] = 0
      "000" when "0001110001110", -- t[910] = 0
      "000" when "0001110001111", -- t[911] = 0
      "000" when "0001110010000", -- t[912] = 0
      "000" when "0001110010001", -- t[913] = 0
      "000" when "0001110010010", -- t[914] = 0
      "000" when "0001110010011", -- t[915] = 0
      "000" when "0001110010100", -- t[916] = 0
      "000" when "0001110010101", -- t[917] = 0
      "000" when "0001110010110", -- t[918] = 0
      "000" when "0001110010111", -- t[919] = 0
      "000" when "0001110011000", -- t[920] = 0
      "000" when "0001110011001", -- t[921] = 0
      "000" when "0001110011010", -- t[922] = 0
      "000" when "0001110011011", -- t[923] = 0
      "000" when "0001110011100", -- t[924] = 0
      "000" when "0001110011101", -- t[925] = 0
      "000" when "0001110011110", -- t[926] = 0
      "000" when "0001110011111", -- t[927] = 0
      "000" when "0001110100000", -- t[928] = 0
      "000" when "0001110100001", -- t[929] = 0
      "000" when "0001110100010", -- t[930] = 0
      "000" when "0001110100011", -- t[931] = 0
      "000" when "0001110100100", -- t[932] = 0
      "000" when "0001110100101", -- t[933] = 0
      "000" when "0001110100110", -- t[934] = 0
      "000" when "0001110100111", -- t[935] = 0
      "000" when "0001110101000", -- t[936] = 0
      "000" when "0001110101001", -- t[937] = 0
      "000" when "0001110101010", -- t[938] = 0
      "000" when "0001110101011", -- t[939] = 0
      "000" when "0001110101100", -- t[940] = 0
      "000" when "0001110101101", -- t[941] = 0
      "000" when "0001110101110", -- t[942] = 0
      "000" when "0001110101111", -- t[943] = 0
      "000" when "0001110110000", -- t[944] = 0
      "000" when "0001110110001", -- t[945] = 0
      "000" when "0001110110010", -- t[946] = 0
      "000" when "0001110110011", -- t[947] = 0
      "000" when "0001110110100", -- t[948] = 0
      "000" when "0001110110101", -- t[949] = 0
      "000" when "0001110110110", -- t[950] = 0
      "000" when "0001110110111", -- t[951] = 0
      "000" when "0001110111000", -- t[952] = 0
      "000" when "0001110111001", -- t[953] = 0
      "000" when "0001110111010", -- t[954] = 0
      "000" when "0001110111011", -- t[955] = 0
      "000" when "0001110111100", -- t[956] = 0
      "000" when "0001110111101", -- t[957] = 0
      "000" when "0001110111110", -- t[958] = 0
      "000" when "0001110111111", -- t[959] = 0
      "000" when "0001111000000", -- t[960] = 0
      "000" when "0001111000001", -- t[961] = 0
      "000" when "0001111000010", -- t[962] = 0
      "000" when "0001111000011", -- t[963] = 0
      "000" when "0001111000100", -- t[964] = 0
      "000" when "0001111000101", -- t[965] = 0
      "000" when "0001111000110", -- t[966] = 0
      "000" when "0001111000111", -- t[967] = 0
      "000" when "0001111001000", -- t[968] = 0
      "000" when "0001111001001", -- t[969] = 0
      "000" when "0001111001010", -- t[970] = 0
      "000" when "0001111001011", -- t[971] = 0
      "000" when "0001111001100", -- t[972] = 0
      "000" when "0001111001101", -- t[973] = 0
      "000" when "0001111001110", -- t[974] = 0
      "000" when "0001111001111", -- t[975] = 0
      "000" when "0001111010000", -- t[976] = 0
      "000" when "0001111010001", -- t[977] = 0
      "000" when "0001111010010", -- t[978] = 0
      "000" when "0001111010011", -- t[979] = 0
      "000" when "0001111010100", -- t[980] = 0
      "000" when "0001111010101", -- t[981] = 0
      "000" when "0001111010110", -- t[982] = 0
      "000" when "0001111010111", -- t[983] = 0
      "000" when "0001111011000", -- t[984] = 0
      "000" when "0001111011001", -- t[985] = 0
      "000" when "0001111011010", -- t[986] = 0
      "000" when "0001111011011", -- t[987] = 0
      "000" when "0001111011100", -- t[988] = 0
      "000" when "0001111011101", -- t[989] = 0
      "000" when "0001111011110", -- t[990] = 0
      "000" when "0001111011111", -- t[991] = 0
      "000" when "0001111100000", -- t[992] = 0
      "000" when "0001111100001", -- t[993] = 0
      "000" when "0001111100010", -- t[994] = 0
      "000" when "0001111100011", -- t[995] = 0
      "000" when "0001111100100", -- t[996] = 0
      "000" when "0001111100101", -- t[997] = 0
      "000" when "0001111100110", -- t[998] = 0
      "000" when "0001111100111", -- t[999] = 0
      "000" when "0001111101000", -- t[1000] = 0
      "000" when "0001111101001", -- t[1001] = 0
      "000" when "0001111101010", -- t[1002] = 0
      "000" when "0001111101011", -- t[1003] = 0
      "000" when "0001111101100", -- t[1004] = 0
      "000" when "0001111101101", -- t[1005] = 0
      "000" when "0001111101110", -- t[1006] = 0
      "000" when "0001111101111", -- t[1007] = 0
      "000" when "0001111110000", -- t[1008] = 0
      "000" when "0001111110001", -- t[1009] = 0
      "000" when "0001111110010", -- t[1010] = 0
      "000" when "0001111110011", -- t[1011] = 0
      "000" when "0001111110100", -- t[1012] = 0
      "000" when "0001111110101", -- t[1013] = 0
      "000" when "0001111110110", -- t[1014] = 0
      "000" when "0001111110111", -- t[1015] = 0
      "000" when "0001111111000", -- t[1016] = 0
      "000" when "0001111111001", -- t[1017] = 0
      "000" when "0001111111010", -- t[1018] = 0
      "000" when "0001111111011", -- t[1019] = 0
      "000" when "0001111111100", -- t[1020] = 0
      "000" when "0001111111101", -- t[1021] = 0
      "000" when "0001111111110", -- t[1022] = 0
      "000" when "0001111111111", -- t[1023] = 0
      "000" when "0010000000000", -- t[1024] = 0
      "000" when "0010000000001", -- t[1025] = 0
      "000" when "0010000000010", -- t[1026] = 0
      "000" when "0010000000011", -- t[1027] = 0
      "000" when "0010000000100", -- t[1028] = 0
      "000" when "0010000000101", -- t[1029] = 0
      "000" when "0010000000110", -- t[1030] = 0
      "000" when "0010000000111", -- t[1031] = 0
      "000" when "0010000001000", -- t[1032] = 0
      "000" when "0010000001001", -- t[1033] = 0
      "000" when "0010000001010", -- t[1034] = 0
      "000" when "0010000001011", -- t[1035] = 0
      "000" when "0010000001100", -- t[1036] = 0
      "000" when "0010000001101", -- t[1037] = 0
      "000" when "0010000001110", -- t[1038] = 0
      "000" when "0010000001111", -- t[1039] = 0
      "000" when "0010000010000", -- t[1040] = 0
      "000" when "0010000010001", -- t[1041] = 0
      "000" when "0010000010010", -- t[1042] = 0
      "000" when "0010000010011", -- t[1043] = 0
      "000" when "0010000010100", -- t[1044] = 0
      "000" when "0010000010101", -- t[1045] = 0
      "000" when "0010000010110", -- t[1046] = 0
      "000" when "0010000010111", -- t[1047] = 0
      "000" when "0010000011000", -- t[1048] = 0
      "000" when "0010000011001", -- t[1049] = 0
      "000" when "0010000011010", -- t[1050] = 0
      "000" when "0010000011011", -- t[1051] = 0
      "000" when "0010000011100", -- t[1052] = 0
      "000" when "0010000011101", -- t[1053] = 0
      "000" when "0010000011110", -- t[1054] = 0
      "000" when "0010000011111", -- t[1055] = 0
      "000" when "0010000100000", -- t[1056] = 0
      "000" when "0010000100001", -- t[1057] = 0
      "000" when "0010000100010", -- t[1058] = 0
      "000" when "0010000100011", -- t[1059] = 0
      "000" when "0010000100100", -- t[1060] = 0
      "000" when "0010000100101", -- t[1061] = 0
      "000" when "0010000100110", -- t[1062] = 0
      "000" when "0010000100111", -- t[1063] = 0
      "000" when "0010000101000", -- t[1064] = 0
      "000" when "0010000101001", -- t[1065] = 0
      "000" when "0010000101010", -- t[1066] = 0
      "000" when "0010000101011", -- t[1067] = 0
      "000" when "0010000101100", -- t[1068] = 0
      "000" when "0010000101101", -- t[1069] = 0
      "000" when "0010000101110", -- t[1070] = 0
      "000" when "0010000101111", -- t[1071] = 0
      "000" when "0010000110000", -- t[1072] = 0
      "000" when "0010000110001", -- t[1073] = 0
      "000" when "0010000110010", -- t[1074] = 0
      "000" when "0010000110011", -- t[1075] = 0
      "000" when "0010000110100", -- t[1076] = 0
      "000" when "0010000110101", -- t[1077] = 0
      "000" when "0010000110110", -- t[1078] = 0
      "000" when "0010000110111", -- t[1079] = 0
      "000" when "0010000111000", -- t[1080] = 0
      "000" when "0010000111001", -- t[1081] = 0
      "000" when "0010000111010", -- t[1082] = 0
      "000" when "0010000111011", -- t[1083] = 0
      "000" when "0010000111100", -- t[1084] = 0
      "000" when "0010000111101", -- t[1085] = 0
      "000" when "0010000111110", -- t[1086] = 0
      "000" when "0010000111111", -- t[1087] = 0
      "000" when "0010001000000", -- t[1088] = 0
      "000" when "0010001000001", -- t[1089] = 0
      "000" when "0010001000010", -- t[1090] = 0
      "000" when "0010001000011", -- t[1091] = 0
      "000" when "0010001000100", -- t[1092] = 0
      "000" when "0010001000101", -- t[1093] = 0
      "000" when "0010001000110", -- t[1094] = 0
      "000" when "0010001000111", -- t[1095] = 0
      "000" when "0010001001000", -- t[1096] = 0
      "000" when "0010001001001", -- t[1097] = 0
      "000" when "0010001001010", -- t[1098] = 0
      "000" when "0010001001011", -- t[1099] = 0
      "000" when "0010001001100", -- t[1100] = 0
      "000" when "0010001001101", -- t[1101] = 0
      "000" when "0010001001110", -- t[1102] = 0
      "000" when "0010001001111", -- t[1103] = 0
      "000" when "0010001010000", -- t[1104] = 0
      "000" when "0010001010001", -- t[1105] = 0
      "000" when "0010001010010", -- t[1106] = 0
      "000" when "0010001010011", -- t[1107] = 0
      "000" when "0010001010100", -- t[1108] = 0
      "000" when "0010001010101", -- t[1109] = 0
      "000" when "0010001010110", -- t[1110] = 0
      "000" when "0010001010111", -- t[1111] = 0
      "000" when "0010001011000", -- t[1112] = 0
      "000" when "0010001011001", -- t[1113] = 0
      "000" when "0010001011010", -- t[1114] = 0
      "000" when "0010001011011", -- t[1115] = 0
      "000" when "0010001011100", -- t[1116] = 0
      "000" when "0010001011101", -- t[1117] = 0
      "000" when "0010001011110", -- t[1118] = 0
      "000" when "0010001011111", -- t[1119] = 0
      "000" when "0010001100000", -- t[1120] = 0
      "000" when "0010001100001", -- t[1121] = 0
      "000" when "0010001100010", -- t[1122] = 0
      "000" when "0010001100011", -- t[1123] = 0
      "000" when "0010001100100", -- t[1124] = 0
      "000" when "0010001100101", -- t[1125] = 0
      "000" when "0010001100110", -- t[1126] = 0
      "000" when "0010001100111", -- t[1127] = 0
      "000" when "0010001101000", -- t[1128] = 0
      "000" when "0010001101001", -- t[1129] = 0
      "000" when "0010001101010", -- t[1130] = 0
      "000" when "0010001101011", -- t[1131] = 0
      "000" when "0010001101100", -- t[1132] = 0
      "000" when "0010001101101", -- t[1133] = 0
      "000" when "0010001101110", -- t[1134] = 0
      "000" when "0010001101111", -- t[1135] = 0
      "000" when "0010001110000", -- t[1136] = 0
      "000" when "0010001110001", -- t[1137] = 0
      "000" when "0010001110010", -- t[1138] = 0
      "000" when "0010001110011", -- t[1139] = 0
      "000" when "0010001110100", -- t[1140] = 0
      "000" when "0010001110101", -- t[1141] = 0
      "000" when "0010001110110", -- t[1142] = 0
      "000" when "0010001110111", -- t[1143] = 0
      "000" when "0010001111000", -- t[1144] = 0
      "000" when "0010001111001", -- t[1145] = 0
      "000" when "0010001111010", -- t[1146] = 0
      "000" when "0010001111011", -- t[1147] = 0
      "000" when "0010001111100", -- t[1148] = 0
      "000" when "0010001111101", -- t[1149] = 0
      "000" when "0010001111110", -- t[1150] = 0
      "000" when "0010001111111", -- t[1151] = 0
      "000" when "0010010000000", -- t[1152] = 0
      "000" when "0010010000001", -- t[1153] = 0
      "000" when "0010010000010", -- t[1154] = 0
      "000" when "0010010000011", -- t[1155] = 0
      "000" when "0010010000100", -- t[1156] = 0
      "000" when "0010010000101", -- t[1157] = 0
      "000" when "0010010000110", -- t[1158] = 0
      "000" when "0010010000111", -- t[1159] = 0
      "000" when "0010010001000", -- t[1160] = 0
      "000" when "0010010001001", -- t[1161] = 0
      "000" when "0010010001010", -- t[1162] = 0
      "000" when "0010010001011", -- t[1163] = 0
      "000" when "0010010001100", -- t[1164] = 0
      "000" when "0010010001101", -- t[1165] = 0
      "000" when "0010010001110", -- t[1166] = 0
      "000" when "0010010001111", -- t[1167] = 0
      "000" when "0010010010000", -- t[1168] = 0
      "000" when "0010010010001", -- t[1169] = 0
      "000" when "0010010010010", -- t[1170] = 0
      "000" when "0010010010011", -- t[1171] = 0
      "000" when "0010010010100", -- t[1172] = 0
      "000" when "0010010010101", -- t[1173] = 0
      "000" when "0010010010110", -- t[1174] = 0
      "000" when "0010010010111", -- t[1175] = 0
      "000" when "0010010011000", -- t[1176] = 0
      "000" when "0010010011001", -- t[1177] = 0
      "000" when "0010010011010", -- t[1178] = 0
      "000" when "0010010011011", -- t[1179] = 0
      "000" when "0010010011100", -- t[1180] = 0
      "000" when "0010010011101", -- t[1181] = 0
      "000" when "0010010011110", -- t[1182] = 0
      "000" when "0010010011111", -- t[1183] = 0
      "000" when "0010010100000", -- t[1184] = 0
      "000" when "0010010100001", -- t[1185] = 0
      "000" when "0010010100010", -- t[1186] = 0
      "000" when "0010010100011", -- t[1187] = 0
      "000" when "0010010100100", -- t[1188] = 0
      "000" when "0010010100101", -- t[1189] = 0
      "000" when "0010010100110", -- t[1190] = 0
      "000" when "0010010100111", -- t[1191] = 0
      "000" when "0010010101000", -- t[1192] = 0
      "000" when "0010010101001", -- t[1193] = 0
      "000" when "0010010101010", -- t[1194] = 0
      "000" when "0010010101011", -- t[1195] = 0
      "000" when "0010010101100", -- t[1196] = 0
      "000" when "0010010101101", -- t[1197] = 0
      "000" when "0010010101110", -- t[1198] = 0
      "000" when "0010010101111", -- t[1199] = 0
      "000" when "0010010110000", -- t[1200] = 0
      "000" when "0010010110001", -- t[1201] = 0
      "000" when "0010010110010", -- t[1202] = 0
      "000" when "0010010110011", -- t[1203] = 0
      "000" when "0010010110100", -- t[1204] = 0
      "000" when "0010010110101", -- t[1205] = 0
      "000" when "0010010110110", -- t[1206] = 0
      "000" when "0010010110111", -- t[1207] = 0
      "000" when "0010010111000", -- t[1208] = 0
      "000" when "0010010111001", -- t[1209] = 0
      "000" when "0010010111010", -- t[1210] = 0
      "000" when "0010010111011", -- t[1211] = 0
      "000" when "0010010111100", -- t[1212] = 0
      "000" when "0010010111101", -- t[1213] = 0
      "000" when "0010010111110", -- t[1214] = 0
      "000" when "0010010111111", -- t[1215] = 0
      "000" when "0010011000000", -- t[1216] = 0
      "000" when "0010011000001", -- t[1217] = 0
      "000" when "0010011000010", -- t[1218] = 0
      "000" when "0010011000011", -- t[1219] = 0
      "000" when "0010011000100", -- t[1220] = 0
      "000" when "0010011000101", -- t[1221] = 0
      "000" when "0010011000110", -- t[1222] = 0
      "000" when "0010011000111", -- t[1223] = 0
      "000" when "0010011001000", -- t[1224] = 0
      "000" when "0010011001001", -- t[1225] = 0
      "000" when "0010011001010", -- t[1226] = 0
      "000" when "0010011001011", -- t[1227] = 0
      "000" when "0010011001100", -- t[1228] = 0
      "000" when "0010011001101", -- t[1229] = 0
      "000" when "0010011001110", -- t[1230] = 0
      "000" when "0010011001111", -- t[1231] = 0
      "000" when "0010011010000", -- t[1232] = 0
      "000" when "0010011010001", -- t[1233] = 0
      "000" when "0010011010010", -- t[1234] = 0
      "000" when "0010011010011", -- t[1235] = 0
      "000" when "0010011010100", -- t[1236] = 0
      "000" when "0010011010101", -- t[1237] = 0
      "000" when "0010011010110", -- t[1238] = 0
      "000" when "0010011010111", -- t[1239] = 0
      "000" when "0010011011000", -- t[1240] = 0
      "000" when "0010011011001", -- t[1241] = 0
      "000" when "0010011011010", -- t[1242] = 0
      "000" when "0010011011011", -- t[1243] = 0
      "000" when "0010011011100", -- t[1244] = 0
      "000" when "0010011011101", -- t[1245] = 0
      "000" when "0010011011110", -- t[1246] = 0
      "000" when "0010011011111", -- t[1247] = 0
      "000" when "0010011100000", -- t[1248] = 0
      "000" when "0010011100001", -- t[1249] = 0
      "000" when "0010011100010", -- t[1250] = 0
      "000" when "0010011100011", -- t[1251] = 0
      "000" when "0010011100100", -- t[1252] = 0
      "000" when "0010011100101", -- t[1253] = 0
      "000" when "0010011100110", -- t[1254] = 0
      "000" when "0010011100111", -- t[1255] = 0
      "000" when "0010011101000", -- t[1256] = 0
      "000" when "0010011101001", -- t[1257] = 0
      "000" when "0010011101010", -- t[1258] = 0
      "000" when "0010011101011", -- t[1259] = 0
      "000" when "0010011101100", -- t[1260] = 0
      "000" when "0010011101101", -- t[1261] = 0
      "000" when "0010011101110", -- t[1262] = 0
      "000" when "0010011101111", -- t[1263] = 0
      "000" when "0010011110000", -- t[1264] = 0
      "000" when "0010011110001", -- t[1265] = 0
      "000" when "0010011110010", -- t[1266] = 0
      "000" when "0010011110011", -- t[1267] = 0
      "000" when "0010011110100", -- t[1268] = 0
      "000" when "0010011110101", -- t[1269] = 0
      "000" when "0010011110110", -- t[1270] = 0
      "000" when "0010011110111", -- t[1271] = 0
      "000" when "0010011111000", -- t[1272] = 0
      "000" when "0010011111001", -- t[1273] = 0
      "000" when "0010011111010", -- t[1274] = 0
      "000" when "0010011111011", -- t[1275] = 0
      "000" when "0010011111100", -- t[1276] = 0
      "000" when "0010011111101", -- t[1277] = 0
      "000" when "0010011111110", -- t[1278] = 0
      "000" when "0010011111111", -- t[1279] = 0
      "000" when "0010100000000", -- t[1280] = 0
      "000" when "0010100000001", -- t[1281] = 0
      "000" when "0010100000010", -- t[1282] = 0
      "000" when "0010100000011", -- t[1283] = 0
      "000" when "0010100000100", -- t[1284] = 0
      "000" when "0010100000101", -- t[1285] = 0
      "000" when "0010100000110", -- t[1286] = 0
      "000" when "0010100000111", -- t[1287] = 0
      "000" when "0010100001000", -- t[1288] = 0
      "000" when "0010100001001", -- t[1289] = 0
      "000" when "0010100001010", -- t[1290] = 0
      "000" when "0010100001011", -- t[1291] = 0
      "000" when "0010100001100", -- t[1292] = 0
      "000" when "0010100001101", -- t[1293] = 0
      "000" when "0010100001110", -- t[1294] = 0
      "000" when "0010100001111", -- t[1295] = 0
      "000" when "0010100010000", -- t[1296] = 0
      "000" when "0010100010001", -- t[1297] = 0
      "000" when "0010100010010", -- t[1298] = 0
      "000" when "0010100010011", -- t[1299] = 0
      "000" when "0010100010100", -- t[1300] = 0
      "000" when "0010100010101", -- t[1301] = 0
      "000" when "0010100010110", -- t[1302] = 0
      "000" when "0010100010111", -- t[1303] = 0
      "000" when "0010100011000", -- t[1304] = 0
      "000" when "0010100011001", -- t[1305] = 0
      "000" when "0010100011010", -- t[1306] = 0
      "000" when "0010100011011", -- t[1307] = 0
      "000" when "0010100011100", -- t[1308] = 0
      "000" when "0010100011101", -- t[1309] = 0
      "000" when "0010100011110", -- t[1310] = 0
      "000" when "0010100011111", -- t[1311] = 0
      "000" when "0010100100000", -- t[1312] = 0
      "000" when "0010100100001", -- t[1313] = 0
      "000" when "0010100100010", -- t[1314] = 0
      "000" when "0010100100011", -- t[1315] = 0
      "000" when "0010100100100", -- t[1316] = 0
      "000" when "0010100100101", -- t[1317] = 0
      "000" when "0010100100110", -- t[1318] = 0
      "000" when "0010100100111", -- t[1319] = 0
      "000" when "0010100101000", -- t[1320] = 0
      "000" when "0010100101001", -- t[1321] = 0
      "000" when "0010100101010", -- t[1322] = 0
      "000" when "0010100101011", -- t[1323] = 0
      "000" when "0010100101100", -- t[1324] = 0
      "000" when "0010100101101", -- t[1325] = 0
      "000" when "0010100101110", -- t[1326] = 0
      "000" when "0010100101111", -- t[1327] = 0
      "000" when "0010100110000", -- t[1328] = 0
      "000" when "0010100110001", -- t[1329] = 0
      "000" when "0010100110010", -- t[1330] = 0
      "000" when "0010100110011", -- t[1331] = 0
      "000" when "0010100110100", -- t[1332] = 0
      "000" when "0010100110101", -- t[1333] = 0
      "000" when "0010100110110", -- t[1334] = 0
      "000" when "0010100110111", -- t[1335] = 0
      "000" when "0010100111000", -- t[1336] = 0
      "000" when "0010100111001", -- t[1337] = 0
      "000" when "0010100111010", -- t[1338] = 0
      "000" when "0010100111011", -- t[1339] = 0
      "000" when "0010100111100", -- t[1340] = 0
      "000" when "0010100111101", -- t[1341] = 0
      "000" when "0010100111110", -- t[1342] = 0
      "000" when "0010100111111", -- t[1343] = 0
      "000" when "0010101000000", -- t[1344] = 0
      "000" when "0010101000001", -- t[1345] = 0
      "000" when "0010101000010", -- t[1346] = 0
      "000" when "0010101000011", -- t[1347] = 0
      "000" when "0010101000100", -- t[1348] = 0
      "000" when "0010101000101", -- t[1349] = 0
      "000" when "0010101000110", -- t[1350] = 0
      "000" when "0010101000111", -- t[1351] = 0
      "000" when "0010101001000", -- t[1352] = 0
      "000" when "0010101001001", -- t[1353] = 0
      "000" when "0010101001010", -- t[1354] = 0
      "000" when "0010101001011", -- t[1355] = 0
      "000" when "0010101001100", -- t[1356] = 0
      "000" when "0010101001101", -- t[1357] = 0
      "000" when "0010101001110", -- t[1358] = 0
      "000" when "0010101001111", -- t[1359] = 0
      "000" when "0010101010000", -- t[1360] = 0
      "000" when "0010101010001", -- t[1361] = 0
      "000" when "0010101010010", -- t[1362] = 0
      "000" when "0010101010011", -- t[1363] = 0
      "000" when "0010101010100", -- t[1364] = 0
      "000" when "0010101010101", -- t[1365] = 0
      "000" when "0010101010110", -- t[1366] = 0
      "000" when "0010101010111", -- t[1367] = 0
      "000" when "0010101011000", -- t[1368] = 0
      "000" when "0010101011001", -- t[1369] = 0
      "000" when "0010101011010", -- t[1370] = 0
      "000" when "0010101011011", -- t[1371] = 0
      "000" when "0010101011100", -- t[1372] = 0
      "000" when "0010101011101", -- t[1373] = 0
      "000" when "0010101011110", -- t[1374] = 0
      "000" when "0010101011111", -- t[1375] = 0
      "000" when "0010101100000", -- t[1376] = 0
      "000" when "0010101100001", -- t[1377] = 0
      "000" when "0010101100010", -- t[1378] = 0
      "000" when "0010101100011", -- t[1379] = 0
      "000" when "0010101100100", -- t[1380] = 0
      "000" when "0010101100101", -- t[1381] = 0
      "000" when "0010101100110", -- t[1382] = 0
      "000" when "0010101100111", -- t[1383] = 0
      "000" when "0010101101000", -- t[1384] = 0
      "000" when "0010101101001", -- t[1385] = 0
      "000" when "0010101101010", -- t[1386] = 0
      "000" when "0010101101011", -- t[1387] = 0
      "000" when "0010101101100", -- t[1388] = 0
      "000" when "0010101101101", -- t[1389] = 0
      "000" when "0010101101110", -- t[1390] = 0
      "000" when "0010101101111", -- t[1391] = 0
      "000" when "0010101110000", -- t[1392] = 0
      "000" when "0010101110001", -- t[1393] = 0
      "000" when "0010101110010", -- t[1394] = 0
      "000" when "0010101110011", -- t[1395] = 0
      "000" when "0010101110100", -- t[1396] = 0
      "000" when "0010101110101", -- t[1397] = 0
      "000" when "0010101110110", -- t[1398] = 0
      "000" when "0010101110111", -- t[1399] = 0
      "000" when "0010101111000", -- t[1400] = 0
      "000" when "0010101111001", -- t[1401] = 0
      "000" when "0010101111010", -- t[1402] = 0
      "000" when "0010101111011", -- t[1403] = 0
      "000" when "0010101111100", -- t[1404] = 0
      "000" when "0010101111101", -- t[1405] = 0
      "000" when "0010101111110", -- t[1406] = 0
      "000" when "0010101111111", -- t[1407] = 0
      "000" when "0010110000000", -- t[1408] = 0
      "000" when "0010110000001", -- t[1409] = 0
      "000" when "0010110000010", -- t[1410] = 0
      "000" when "0010110000011", -- t[1411] = 0
      "000" when "0010110000100", -- t[1412] = 0
      "000" when "0010110000101", -- t[1413] = 0
      "000" when "0010110000110", -- t[1414] = 0
      "000" when "0010110000111", -- t[1415] = 0
      "000" when "0010110001000", -- t[1416] = 0
      "000" when "0010110001001", -- t[1417] = 0
      "000" when "0010110001010", -- t[1418] = 0
      "000" when "0010110001011", -- t[1419] = 0
      "000" when "0010110001100", -- t[1420] = 0
      "000" when "0010110001101", -- t[1421] = 0
      "000" when "0010110001110", -- t[1422] = 0
      "000" when "0010110001111", -- t[1423] = 0
      "000" when "0010110010000", -- t[1424] = 0
      "000" when "0010110010001", -- t[1425] = 0
      "000" when "0010110010010", -- t[1426] = 0
      "000" when "0010110010011", -- t[1427] = 0
      "000" when "0010110010100", -- t[1428] = 0
      "000" when "0010110010101", -- t[1429] = 0
      "000" when "0010110010110", -- t[1430] = 0
      "000" when "0010110010111", -- t[1431] = 0
      "000" when "0010110011000", -- t[1432] = 0
      "000" when "0010110011001", -- t[1433] = 0
      "000" when "0010110011010", -- t[1434] = 0
      "000" when "0010110011011", -- t[1435] = 0
      "000" when "0010110011100", -- t[1436] = 0
      "000" when "0010110011101", -- t[1437] = 0
      "000" when "0010110011110", -- t[1438] = 0
      "000" when "0010110011111", -- t[1439] = 0
      "000" when "0010110100000", -- t[1440] = 0
      "000" when "0010110100001", -- t[1441] = 0
      "000" when "0010110100010", -- t[1442] = 0
      "000" when "0010110100011", -- t[1443] = 0
      "000" when "0010110100100", -- t[1444] = 0
      "000" when "0010110100101", -- t[1445] = 0
      "000" when "0010110100110", -- t[1446] = 0
      "000" when "0010110100111", -- t[1447] = 0
      "000" when "0010110101000", -- t[1448] = 0
      "000" when "0010110101001", -- t[1449] = 0
      "000" when "0010110101010", -- t[1450] = 0
      "000" when "0010110101011", -- t[1451] = 0
      "000" when "0010110101100", -- t[1452] = 0
      "000" when "0010110101101", -- t[1453] = 0
      "000" when "0010110101110", -- t[1454] = 0
      "000" when "0010110101111", -- t[1455] = 0
      "000" when "0010110110000", -- t[1456] = 0
      "000" when "0010110110001", -- t[1457] = 0
      "000" when "0010110110010", -- t[1458] = 0
      "000" when "0010110110011", -- t[1459] = 0
      "000" when "0010110110100", -- t[1460] = 0
      "000" when "0010110110101", -- t[1461] = 0
      "000" when "0010110110110", -- t[1462] = 0
      "000" when "0010110110111", -- t[1463] = 0
      "000" when "0010110111000", -- t[1464] = 0
      "000" when "0010110111001", -- t[1465] = 0
      "000" when "0010110111010", -- t[1466] = 0
      "000" when "0010110111011", -- t[1467] = 0
      "000" when "0010110111100", -- t[1468] = 0
      "000" when "0010110111101", -- t[1469] = 0
      "000" when "0010110111110", -- t[1470] = 0
      "000" when "0010110111111", -- t[1471] = 0
      "000" when "0010111000000", -- t[1472] = 0
      "000" when "0010111000001", -- t[1473] = 0
      "000" when "0010111000010", -- t[1474] = 0
      "000" when "0010111000011", -- t[1475] = 0
      "000" when "0010111000100", -- t[1476] = 0
      "000" when "0010111000101", -- t[1477] = 0
      "000" when "0010111000110", -- t[1478] = 0
      "000" when "0010111000111", -- t[1479] = 0
      "000" when "0010111001000", -- t[1480] = 0
      "000" when "0010111001001", -- t[1481] = 0
      "000" when "0010111001010", -- t[1482] = 0
      "000" when "0010111001011", -- t[1483] = 0
      "000" when "0010111001100", -- t[1484] = 0
      "000" when "0010111001101", -- t[1485] = 0
      "000" when "0010111001110", -- t[1486] = 0
      "000" when "0010111001111", -- t[1487] = 0
      "000" when "0010111010000", -- t[1488] = 0
      "000" when "0010111010001", -- t[1489] = 0
      "000" when "0010111010010", -- t[1490] = 0
      "000" when "0010111010011", -- t[1491] = 0
      "000" when "0010111010100", -- t[1492] = 0
      "000" when "0010111010101", -- t[1493] = 0
      "000" when "0010111010110", -- t[1494] = 0
      "000" when "0010111010111", -- t[1495] = 0
      "000" when "0010111011000", -- t[1496] = 0
      "000" when "0010111011001", -- t[1497] = 0
      "000" when "0010111011010", -- t[1498] = 0
      "000" when "0010111011011", -- t[1499] = 0
      "000" when "0010111011100", -- t[1500] = 0
      "000" when "0010111011101", -- t[1501] = 0
      "000" when "0010111011110", -- t[1502] = 0
      "000" when "0010111011111", -- t[1503] = 0
      "000" when "0010111100000", -- t[1504] = 0
      "000" when "0010111100001", -- t[1505] = 0
      "000" when "0010111100010", -- t[1506] = 0
      "000" when "0010111100011", -- t[1507] = 0
      "000" when "0010111100100", -- t[1508] = 0
      "000" when "0010111100101", -- t[1509] = 0
      "000" when "0010111100110", -- t[1510] = 0
      "000" when "0010111100111", -- t[1511] = 0
      "000" when "0010111101000", -- t[1512] = 0
      "000" when "0010111101001", -- t[1513] = 0
      "000" when "0010111101010", -- t[1514] = 0
      "000" when "0010111101011", -- t[1515] = 0
      "000" when "0010111101100", -- t[1516] = 0
      "000" when "0010111101101", -- t[1517] = 0
      "000" when "0010111101110", -- t[1518] = 0
      "000" when "0010111101111", -- t[1519] = 0
      "000" when "0010111110000", -- t[1520] = 0
      "000" when "0010111110001", -- t[1521] = 0
      "000" when "0010111110010", -- t[1522] = 0
      "000" when "0010111110011", -- t[1523] = 0
      "000" when "0010111110100", -- t[1524] = 0
      "000" when "0010111110101", -- t[1525] = 0
      "000" when "0010111110110", -- t[1526] = 0
      "000" when "0010111110111", -- t[1527] = 0
      "000" when "0010111111000", -- t[1528] = 0
      "000" when "0010111111001", -- t[1529] = 0
      "000" when "0010111111010", -- t[1530] = 0
      "000" when "0010111111011", -- t[1531] = 0
      "000" when "0010111111100", -- t[1532] = 0
      "000" when "0010111111101", -- t[1533] = 0
      "000" when "0010111111110", -- t[1534] = 0
      "000" when "0010111111111", -- t[1535] = 0
      "000" when "0011000000000", -- t[1536] = 0
      "000" when "0011000000001", -- t[1537] = 0
      "000" when "0011000000010", -- t[1538] = 0
      "000" when "0011000000011", -- t[1539] = 0
      "000" when "0011000000100", -- t[1540] = 0
      "000" when "0011000000101", -- t[1541] = 0
      "000" when "0011000000110", -- t[1542] = 0
      "000" when "0011000000111", -- t[1543] = 0
      "000" when "0011000001000", -- t[1544] = 0
      "000" when "0011000001001", -- t[1545] = 0
      "000" when "0011000001010", -- t[1546] = 0
      "000" when "0011000001011", -- t[1547] = 0
      "000" when "0011000001100", -- t[1548] = 0
      "000" when "0011000001101", -- t[1549] = 0
      "000" when "0011000001110", -- t[1550] = 0
      "000" when "0011000001111", -- t[1551] = 0
      "000" when "0011000010000", -- t[1552] = 0
      "000" when "0011000010001", -- t[1553] = 0
      "000" when "0011000010010", -- t[1554] = 0
      "000" when "0011000010011", -- t[1555] = 0
      "000" when "0011000010100", -- t[1556] = 0
      "000" when "0011000010101", -- t[1557] = 0
      "000" when "0011000010110", -- t[1558] = 0
      "000" when "0011000010111", -- t[1559] = 0
      "000" when "0011000011000", -- t[1560] = 0
      "000" when "0011000011001", -- t[1561] = 0
      "000" when "0011000011010", -- t[1562] = 0
      "000" when "0011000011011", -- t[1563] = 0
      "000" when "0011000011100", -- t[1564] = 0
      "000" when "0011000011101", -- t[1565] = 0
      "000" when "0011000011110", -- t[1566] = 0
      "000" when "0011000011111", -- t[1567] = 0
      "000" when "0011000100000", -- t[1568] = 0
      "000" when "0011000100001", -- t[1569] = 0
      "000" when "0011000100010", -- t[1570] = 0
      "000" when "0011000100011", -- t[1571] = 0
      "000" when "0011000100100", -- t[1572] = 0
      "000" when "0011000100101", -- t[1573] = 0
      "000" when "0011000100110", -- t[1574] = 0
      "000" when "0011000100111", -- t[1575] = 0
      "000" when "0011000101000", -- t[1576] = 0
      "000" when "0011000101001", -- t[1577] = 0
      "000" when "0011000101010", -- t[1578] = 0
      "000" when "0011000101011", -- t[1579] = 0
      "000" when "0011000101100", -- t[1580] = 0
      "000" when "0011000101101", -- t[1581] = 0
      "000" when "0011000101110", -- t[1582] = 0
      "000" when "0011000101111", -- t[1583] = 0
      "000" when "0011000110000", -- t[1584] = 0
      "000" when "0011000110001", -- t[1585] = 0
      "000" when "0011000110010", -- t[1586] = 0
      "000" when "0011000110011", -- t[1587] = 0
      "000" when "0011000110100", -- t[1588] = 0
      "000" when "0011000110101", -- t[1589] = 0
      "000" when "0011000110110", -- t[1590] = 0
      "000" when "0011000110111", -- t[1591] = 0
      "000" when "0011000111000", -- t[1592] = 0
      "000" when "0011000111001", -- t[1593] = 0
      "000" when "0011000111010", -- t[1594] = 0
      "000" when "0011000111011", -- t[1595] = 0
      "000" when "0011000111100", -- t[1596] = 0
      "000" when "0011000111101", -- t[1597] = 0
      "000" when "0011000111110", -- t[1598] = 0
      "000" when "0011000111111", -- t[1599] = 0
      "000" when "0011001000000", -- t[1600] = 0
      "000" when "0011001000001", -- t[1601] = 0
      "000" when "0011001000010", -- t[1602] = 0
      "000" when "0011001000011", -- t[1603] = 0
      "000" when "0011001000100", -- t[1604] = 0
      "000" when "0011001000101", -- t[1605] = 0
      "000" when "0011001000110", -- t[1606] = 0
      "000" when "0011001000111", -- t[1607] = 0
      "000" when "0011001001000", -- t[1608] = 0
      "000" when "0011001001001", -- t[1609] = 0
      "000" when "0011001001010", -- t[1610] = 0
      "000" when "0011001001011", -- t[1611] = 0
      "000" when "0011001001100", -- t[1612] = 0
      "000" when "0011001001101", -- t[1613] = 0
      "000" when "0011001001110", -- t[1614] = 0
      "000" when "0011001001111", -- t[1615] = 0
      "000" when "0011001010000", -- t[1616] = 0
      "000" when "0011001010001", -- t[1617] = 0
      "000" when "0011001010010", -- t[1618] = 0
      "000" when "0011001010011", -- t[1619] = 0
      "000" when "0011001010100", -- t[1620] = 0
      "000" when "0011001010101", -- t[1621] = 0
      "000" when "0011001010110", -- t[1622] = 0
      "000" when "0011001010111", -- t[1623] = 0
      "000" when "0011001011000", -- t[1624] = 0
      "000" when "0011001011001", -- t[1625] = 0
      "000" when "0011001011010", -- t[1626] = 0
      "000" when "0011001011011", -- t[1627] = 0
      "000" when "0011001011100", -- t[1628] = 0
      "000" when "0011001011101", -- t[1629] = 0
      "000" when "0011001011110", -- t[1630] = 0
      "000" when "0011001011111", -- t[1631] = 0
      "000" when "0011001100000", -- t[1632] = 0
      "000" when "0011001100001", -- t[1633] = 0
      "000" when "0011001100010", -- t[1634] = 0
      "000" when "0011001100011", -- t[1635] = 0
      "000" when "0011001100100", -- t[1636] = 0
      "000" when "0011001100101", -- t[1637] = 0
      "000" when "0011001100110", -- t[1638] = 0
      "000" when "0011001100111", -- t[1639] = 0
      "000" when "0011001101000", -- t[1640] = 0
      "000" when "0011001101001", -- t[1641] = 0
      "000" when "0011001101010", -- t[1642] = 0
      "000" when "0011001101011", -- t[1643] = 0
      "000" when "0011001101100", -- t[1644] = 0
      "000" when "0011001101101", -- t[1645] = 0
      "000" when "0011001101110", -- t[1646] = 0
      "000" when "0011001101111", -- t[1647] = 0
      "000" when "0011001110000", -- t[1648] = 0
      "000" when "0011001110001", -- t[1649] = 0
      "000" when "0011001110010", -- t[1650] = 0
      "000" when "0011001110011", -- t[1651] = 0
      "000" when "0011001110100", -- t[1652] = 0
      "000" when "0011001110101", -- t[1653] = 0
      "000" when "0011001110110", -- t[1654] = 0
      "000" when "0011001110111", -- t[1655] = 0
      "000" when "0011001111000", -- t[1656] = 0
      "000" when "0011001111001", -- t[1657] = 0
      "000" when "0011001111010", -- t[1658] = 0
      "000" when "0011001111011", -- t[1659] = 0
      "000" when "0011001111100", -- t[1660] = 0
      "000" when "0011001111101", -- t[1661] = 0
      "000" when "0011001111110", -- t[1662] = 0
      "000" when "0011001111111", -- t[1663] = 0
      "000" when "0011010000000", -- t[1664] = 0
      "000" when "0011010000001", -- t[1665] = 0
      "000" when "0011010000010", -- t[1666] = 0
      "000" when "0011010000011", -- t[1667] = 0
      "000" when "0011010000100", -- t[1668] = 0
      "000" when "0011010000101", -- t[1669] = 0
      "000" when "0011010000110", -- t[1670] = 0
      "000" when "0011010000111", -- t[1671] = 0
      "000" when "0011010001000", -- t[1672] = 0
      "000" when "0011010001001", -- t[1673] = 0
      "000" when "0011010001010", -- t[1674] = 0
      "000" when "0011010001011", -- t[1675] = 0
      "000" when "0011010001100", -- t[1676] = 0
      "000" when "0011010001101", -- t[1677] = 0
      "000" when "0011010001110", -- t[1678] = 0
      "000" when "0011010001111", -- t[1679] = 0
      "000" when "0011010010000", -- t[1680] = 0
      "000" when "0011010010001", -- t[1681] = 0
      "000" when "0011010010010", -- t[1682] = 0
      "000" when "0011010010011", -- t[1683] = 0
      "000" when "0011010010100", -- t[1684] = 0
      "000" when "0011010010101", -- t[1685] = 0
      "000" when "0011010010110", -- t[1686] = 0
      "000" when "0011010010111", -- t[1687] = 0
      "000" when "0011010011000", -- t[1688] = 0
      "000" when "0011010011001", -- t[1689] = 0
      "000" when "0011010011010", -- t[1690] = 0
      "000" when "0011010011011", -- t[1691] = 0
      "000" when "0011010011100", -- t[1692] = 0
      "000" when "0011010011101", -- t[1693] = 0
      "000" when "0011010011110", -- t[1694] = 0
      "000" when "0011010011111", -- t[1695] = 0
      "000" when "0011010100000", -- t[1696] = 0
      "000" when "0011010100001", -- t[1697] = 0
      "000" when "0011010100010", -- t[1698] = 0
      "000" when "0011010100011", -- t[1699] = 0
      "000" when "0011010100100", -- t[1700] = 0
      "000" when "0011010100101", -- t[1701] = 0
      "000" when "0011010100110", -- t[1702] = 0
      "000" when "0011010100111", -- t[1703] = 0
      "000" when "0011010101000", -- t[1704] = 0
      "000" when "0011010101001", -- t[1705] = 0
      "000" when "0011010101010", -- t[1706] = 0
      "000" when "0011010101011", -- t[1707] = 0
      "000" when "0011010101100", -- t[1708] = 0
      "000" when "0011010101101", -- t[1709] = 0
      "000" when "0011010101110", -- t[1710] = 0
      "000" when "0011010101111", -- t[1711] = 0
      "000" when "0011010110000", -- t[1712] = 0
      "000" when "0011010110001", -- t[1713] = 0
      "000" when "0011010110010", -- t[1714] = 0
      "000" when "0011010110011", -- t[1715] = 0
      "000" when "0011010110100", -- t[1716] = 0
      "000" when "0011010110101", -- t[1717] = 0
      "000" when "0011010110110", -- t[1718] = 0
      "000" when "0011010110111", -- t[1719] = 0
      "000" when "0011010111000", -- t[1720] = 0
      "000" when "0011010111001", -- t[1721] = 0
      "000" when "0011010111010", -- t[1722] = 0
      "000" when "0011010111011", -- t[1723] = 0
      "000" when "0011010111100", -- t[1724] = 0
      "000" when "0011010111101", -- t[1725] = 0
      "000" when "0011010111110", -- t[1726] = 0
      "000" when "0011010111111", -- t[1727] = 0
      "000" when "0011011000000", -- t[1728] = 0
      "000" when "0011011000001", -- t[1729] = 0
      "000" when "0011011000010", -- t[1730] = 0
      "000" when "0011011000011", -- t[1731] = 0
      "000" when "0011011000100", -- t[1732] = 0
      "000" when "0011011000101", -- t[1733] = 0
      "000" when "0011011000110", -- t[1734] = 0
      "000" when "0011011000111", -- t[1735] = 0
      "000" when "0011011001000", -- t[1736] = 0
      "000" when "0011011001001", -- t[1737] = 0
      "000" when "0011011001010", -- t[1738] = 0
      "000" when "0011011001011", -- t[1739] = 0
      "000" when "0011011001100", -- t[1740] = 0
      "000" when "0011011001101", -- t[1741] = 0
      "000" when "0011011001110", -- t[1742] = 0
      "000" when "0011011001111", -- t[1743] = 0
      "000" when "0011011010000", -- t[1744] = 0
      "000" when "0011011010001", -- t[1745] = 0
      "000" when "0011011010010", -- t[1746] = 0
      "000" when "0011011010011", -- t[1747] = 0
      "000" when "0011011010100", -- t[1748] = 0
      "000" when "0011011010101", -- t[1749] = 0
      "000" when "0011011010110", -- t[1750] = 0
      "000" when "0011011010111", -- t[1751] = 0
      "000" when "0011011011000", -- t[1752] = 0
      "000" when "0011011011001", -- t[1753] = 0
      "000" when "0011011011010", -- t[1754] = 0
      "000" when "0011011011011", -- t[1755] = 0
      "000" when "0011011011100", -- t[1756] = 0
      "000" when "0011011011101", -- t[1757] = 0
      "000" when "0011011011110", -- t[1758] = 0
      "000" when "0011011011111", -- t[1759] = 0
      "000" when "0011011100000", -- t[1760] = 0
      "000" when "0011011100001", -- t[1761] = 0
      "000" when "0011011100010", -- t[1762] = 0
      "000" when "0011011100011", -- t[1763] = 0
      "000" when "0011011100100", -- t[1764] = 0
      "000" when "0011011100101", -- t[1765] = 0
      "000" when "0011011100110", -- t[1766] = 0
      "000" when "0011011100111", -- t[1767] = 0
      "000" when "0011011101000", -- t[1768] = 0
      "000" when "0011011101001", -- t[1769] = 0
      "000" when "0011011101010", -- t[1770] = 0
      "000" when "0011011101011", -- t[1771] = 0
      "000" when "0011011101100", -- t[1772] = 0
      "000" when "0011011101101", -- t[1773] = 0
      "000" when "0011011101110", -- t[1774] = 0
      "000" when "0011011101111", -- t[1775] = 0
      "000" when "0011011110000", -- t[1776] = 0
      "000" when "0011011110001", -- t[1777] = 0
      "000" when "0011011110010", -- t[1778] = 0
      "000" when "0011011110011", -- t[1779] = 0
      "000" when "0011011110100", -- t[1780] = 0
      "000" when "0011011110101", -- t[1781] = 0
      "000" when "0011011110110", -- t[1782] = 0
      "000" when "0011011110111", -- t[1783] = 0
      "000" when "0011011111000", -- t[1784] = 0
      "000" when "0011011111001", -- t[1785] = 0
      "000" when "0011011111010", -- t[1786] = 0
      "000" when "0011011111011", -- t[1787] = 0
      "000" when "0011011111100", -- t[1788] = 0
      "000" when "0011011111101", -- t[1789] = 0
      "000" when "0011011111110", -- t[1790] = 0
      "000" when "0011011111111", -- t[1791] = 0
      "000" when "0011100000000", -- t[1792] = 0
      "000" when "0011100000001", -- t[1793] = 0
      "000" when "0011100000010", -- t[1794] = 0
      "000" when "0011100000011", -- t[1795] = 0
      "000" when "0011100000100", -- t[1796] = 0
      "000" when "0011100000101", -- t[1797] = 0
      "000" when "0011100000110", -- t[1798] = 0
      "000" when "0011100000111", -- t[1799] = 0
      "000" when "0011100001000", -- t[1800] = 0
      "000" when "0011100001001", -- t[1801] = 0
      "000" when "0011100001010", -- t[1802] = 0
      "000" when "0011100001011", -- t[1803] = 0
      "000" when "0011100001100", -- t[1804] = 0
      "000" when "0011100001101", -- t[1805] = 0
      "000" when "0011100001110", -- t[1806] = 0
      "000" when "0011100001111", -- t[1807] = 0
      "000" when "0011100010000", -- t[1808] = 0
      "000" when "0011100010001", -- t[1809] = 0
      "000" when "0011100010010", -- t[1810] = 0
      "000" when "0011100010011", -- t[1811] = 0
      "000" when "0011100010100", -- t[1812] = 0
      "000" when "0011100010101", -- t[1813] = 0
      "000" when "0011100010110", -- t[1814] = 0
      "000" when "0011100010111", -- t[1815] = 0
      "000" when "0011100011000", -- t[1816] = 0
      "000" when "0011100011001", -- t[1817] = 0
      "000" when "0011100011010", -- t[1818] = 0
      "000" when "0011100011011", -- t[1819] = 0
      "000" when "0011100011100", -- t[1820] = 0
      "000" when "0011100011101", -- t[1821] = 0
      "000" when "0011100011110", -- t[1822] = 0
      "000" when "0011100011111", -- t[1823] = 0
      "000" when "0011100100000", -- t[1824] = 0
      "000" when "0011100100001", -- t[1825] = 0
      "000" when "0011100100010", -- t[1826] = 0
      "000" when "0011100100011", -- t[1827] = 0
      "000" when "0011100100100", -- t[1828] = 0
      "000" when "0011100100101", -- t[1829] = 0
      "000" when "0011100100110", -- t[1830] = 0
      "000" when "0011100100111", -- t[1831] = 0
      "000" when "0011100101000", -- t[1832] = 0
      "000" when "0011100101001", -- t[1833] = 0
      "000" when "0011100101010", -- t[1834] = 0
      "000" when "0011100101011", -- t[1835] = 0
      "000" when "0011100101100", -- t[1836] = 0
      "000" when "0011100101101", -- t[1837] = 0
      "000" when "0011100101110", -- t[1838] = 0
      "000" when "0011100101111", -- t[1839] = 0
      "000" when "0011100110000", -- t[1840] = 0
      "000" when "0011100110001", -- t[1841] = 0
      "000" when "0011100110010", -- t[1842] = 0
      "000" when "0011100110011", -- t[1843] = 0
      "000" when "0011100110100", -- t[1844] = 0
      "000" when "0011100110101", -- t[1845] = 0
      "000" when "0011100110110", -- t[1846] = 0
      "000" when "0011100110111", -- t[1847] = 0
      "000" when "0011100111000", -- t[1848] = 0
      "000" when "0011100111001", -- t[1849] = 0
      "000" when "0011100111010", -- t[1850] = 0
      "000" when "0011100111011", -- t[1851] = 0
      "000" when "0011100111100", -- t[1852] = 0
      "000" when "0011100111101", -- t[1853] = 0
      "000" when "0011100111110", -- t[1854] = 0
      "000" when "0011100111111", -- t[1855] = 0
      "000" when "0011101000000", -- t[1856] = 0
      "000" when "0011101000001", -- t[1857] = 0
      "000" when "0011101000010", -- t[1858] = 0
      "000" when "0011101000011", -- t[1859] = 0
      "000" when "0011101000100", -- t[1860] = 0
      "000" when "0011101000101", -- t[1861] = 0
      "000" when "0011101000110", -- t[1862] = 0
      "000" when "0011101000111", -- t[1863] = 0
      "000" when "0011101001000", -- t[1864] = 0
      "000" when "0011101001001", -- t[1865] = 0
      "000" when "0011101001010", -- t[1866] = 0
      "000" when "0011101001011", -- t[1867] = 0
      "000" when "0011101001100", -- t[1868] = 0
      "000" when "0011101001101", -- t[1869] = 0
      "000" when "0011101001110", -- t[1870] = 0
      "000" when "0011101001111", -- t[1871] = 0
      "000" when "0011101010000", -- t[1872] = 0
      "000" when "0011101010001", -- t[1873] = 0
      "000" when "0011101010010", -- t[1874] = 0
      "000" when "0011101010011", -- t[1875] = 0
      "000" when "0011101010100", -- t[1876] = 0
      "000" when "0011101010101", -- t[1877] = 0
      "000" when "0011101010110", -- t[1878] = 0
      "000" when "0011101010111", -- t[1879] = 0
      "000" when "0011101011000", -- t[1880] = 0
      "000" when "0011101011001", -- t[1881] = 0
      "000" when "0011101011010", -- t[1882] = 0
      "000" when "0011101011011", -- t[1883] = 0
      "000" when "0011101011100", -- t[1884] = 0
      "000" when "0011101011101", -- t[1885] = 0
      "000" when "0011101011110", -- t[1886] = 0
      "000" when "0011101011111", -- t[1887] = 0
      "000" when "0011101100000", -- t[1888] = 0
      "000" when "0011101100001", -- t[1889] = 0
      "000" when "0011101100010", -- t[1890] = 0
      "000" when "0011101100011", -- t[1891] = 0
      "000" when "0011101100100", -- t[1892] = 0
      "000" when "0011101100101", -- t[1893] = 0
      "000" when "0011101100110", -- t[1894] = 0
      "000" when "0011101100111", -- t[1895] = 0
      "000" when "0011101101000", -- t[1896] = 0
      "000" when "0011101101001", -- t[1897] = 0
      "000" when "0011101101010", -- t[1898] = 0
      "000" when "0011101101011", -- t[1899] = 0
      "000" when "0011101101100", -- t[1900] = 0
      "000" when "0011101101101", -- t[1901] = 0
      "000" when "0011101101110", -- t[1902] = 0
      "000" when "0011101101111", -- t[1903] = 0
      "000" when "0011101110000", -- t[1904] = 0
      "000" when "0011101110001", -- t[1905] = 0
      "000" when "0011101110010", -- t[1906] = 0
      "000" when "0011101110011", -- t[1907] = 0
      "000" when "0011101110100", -- t[1908] = 0
      "000" when "0011101110101", -- t[1909] = 0
      "000" when "0011101110110", -- t[1910] = 0
      "000" when "0011101110111", -- t[1911] = 0
      "000" when "0011101111000", -- t[1912] = 0
      "000" when "0011101111001", -- t[1913] = 0
      "000" when "0011101111010", -- t[1914] = 0
      "000" when "0011101111011", -- t[1915] = 0
      "000" when "0011101111100", -- t[1916] = 0
      "000" when "0011101111101", -- t[1917] = 0
      "000" when "0011101111110", -- t[1918] = 0
      "000" when "0011101111111", -- t[1919] = 0
      "000" when "0011110000000", -- t[1920] = 0
      "000" when "0011110000001", -- t[1921] = 0
      "000" when "0011110000010", -- t[1922] = 0
      "000" when "0011110000011", -- t[1923] = 0
      "000" when "0011110000100", -- t[1924] = 0
      "000" when "0011110000101", -- t[1925] = 0
      "000" when "0011110000110", -- t[1926] = 0
      "000" when "0011110000111", -- t[1927] = 0
      "000" when "0011110001000", -- t[1928] = 0
      "000" when "0011110001001", -- t[1929] = 0
      "000" when "0011110001010", -- t[1930] = 0
      "000" when "0011110001011", -- t[1931] = 0
      "000" when "0011110001100", -- t[1932] = 0
      "000" when "0011110001101", -- t[1933] = 0
      "000" when "0011110001110", -- t[1934] = 0
      "000" when "0011110001111", -- t[1935] = 0
      "000" when "0011110010000", -- t[1936] = 0
      "000" when "0011110010001", -- t[1937] = 0
      "000" when "0011110010010", -- t[1938] = 0
      "000" when "0011110010011", -- t[1939] = 0
      "000" when "0011110010100", -- t[1940] = 0
      "000" when "0011110010101", -- t[1941] = 0
      "000" when "0011110010110", -- t[1942] = 0
      "000" when "0011110010111", -- t[1943] = 0
      "000" when "0011110011000", -- t[1944] = 0
      "000" when "0011110011001", -- t[1945] = 0
      "000" when "0011110011010", -- t[1946] = 0
      "000" when "0011110011011", -- t[1947] = 0
      "000" when "0011110011100", -- t[1948] = 0
      "000" when "0011110011101", -- t[1949] = 0
      "000" when "0011110011110", -- t[1950] = 0
      "000" when "0011110011111", -- t[1951] = 0
      "000" when "0011110100000", -- t[1952] = 0
      "000" when "0011110100001", -- t[1953] = 0
      "000" when "0011110100010", -- t[1954] = 0
      "000" when "0011110100011", -- t[1955] = 0
      "000" when "0011110100100", -- t[1956] = 0
      "000" when "0011110100101", -- t[1957] = 0
      "000" when "0011110100110", -- t[1958] = 0
      "000" when "0011110100111", -- t[1959] = 0
      "000" when "0011110101000", -- t[1960] = 0
      "000" when "0011110101001", -- t[1961] = 0
      "000" when "0011110101010", -- t[1962] = 0
      "000" when "0011110101011", -- t[1963] = 0
      "000" when "0011110101100", -- t[1964] = 0
      "000" when "0011110101101", -- t[1965] = 0
      "000" when "0011110101110", -- t[1966] = 0
      "000" when "0011110101111", -- t[1967] = 0
      "000" when "0011110110000", -- t[1968] = 0
      "000" when "0011110110001", -- t[1969] = 0
      "000" when "0011110110010", -- t[1970] = 0
      "000" when "0011110110011", -- t[1971] = 0
      "000" when "0011110110100", -- t[1972] = 0
      "000" when "0011110110101", -- t[1973] = 0
      "000" when "0011110110110", -- t[1974] = 0
      "000" when "0011110110111", -- t[1975] = 0
      "000" when "0011110111000", -- t[1976] = 0
      "000" when "0011110111001", -- t[1977] = 0
      "000" when "0011110111010", -- t[1978] = 0
      "000" when "0011110111011", -- t[1979] = 0
      "000" when "0011110111100", -- t[1980] = 0
      "000" when "0011110111101", -- t[1981] = 0
      "000" when "0011110111110", -- t[1982] = 0
      "000" when "0011110111111", -- t[1983] = 0
      "000" when "0011111000000", -- t[1984] = 0
      "000" when "0011111000001", -- t[1985] = 0
      "000" when "0011111000010", -- t[1986] = 0
      "000" when "0011111000011", -- t[1987] = 0
      "000" when "0011111000100", -- t[1988] = 0
      "000" when "0011111000101", -- t[1989] = 0
      "000" when "0011111000110", -- t[1990] = 0
      "000" when "0011111000111", -- t[1991] = 0
      "000" when "0011111001000", -- t[1992] = 0
      "000" when "0011111001001", -- t[1993] = 0
      "000" when "0011111001010", -- t[1994] = 0
      "000" when "0011111001011", -- t[1995] = 0
      "000" when "0011111001100", -- t[1996] = 0
      "000" when "0011111001101", -- t[1997] = 0
      "000" when "0011111001110", -- t[1998] = 0
      "000" when "0011111001111", -- t[1999] = 0
      "000" when "0011111010000", -- t[2000] = 0
      "000" when "0011111010001", -- t[2001] = 0
      "000" when "0011111010010", -- t[2002] = 0
      "000" when "0011111010011", -- t[2003] = 0
      "000" when "0011111010100", -- t[2004] = 0
      "000" when "0011111010101", -- t[2005] = 0
      "000" when "0011111010110", -- t[2006] = 0
      "000" when "0011111010111", -- t[2007] = 0
      "000" when "0011111011000", -- t[2008] = 0
      "000" when "0011111011001", -- t[2009] = 0
      "000" when "0011111011010", -- t[2010] = 0
      "000" when "0011111011011", -- t[2011] = 0
      "000" when "0011111011100", -- t[2012] = 0
      "000" when "0011111011101", -- t[2013] = 0
      "000" when "0011111011110", -- t[2014] = 0
      "000" when "0011111011111", -- t[2015] = 0
      "000" when "0011111100000", -- t[2016] = 0
      "000" when "0011111100001", -- t[2017] = 0
      "000" when "0011111100010", -- t[2018] = 0
      "000" when "0011111100011", -- t[2019] = 0
      "000" when "0011111100100", -- t[2020] = 0
      "000" when "0011111100101", -- t[2021] = 0
      "000" when "0011111100110", -- t[2022] = 0
      "000" when "0011111100111", -- t[2023] = 0
      "000" when "0011111101000", -- t[2024] = 0
      "000" when "0011111101001", -- t[2025] = 0
      "000" when "0011111101010", -- t[2026] = 0
      "000" when "0011111101011", -- t[2027] = 0
      "000" when "0011111101100", -- t[2028] = 0
      "000" when "0011111101101", -- t[2029] = 0
      "000" when "0011111101110", -- t[2030] = 0
      "000" when "0011111101111", -- t[2031] = 0
      "000" when "0011111110000", -- t[2032] = 0
      "000" when "0011111110001", -- t[2033] = 0
      "000" when "0011111110010", -- t[2034] = 0
      "000" when "0011111110011", -- t[2035] = 0
      "000" when "0011111110100", -- t[2036] = 0
      "000" when "0011111110101", -- t[2037] = 0
      "000" when "0011111110110", -- t[2038] = 0
      "000" when "0011111110111", -- t[2039] = 0
      "000" when "0011111111000", -- t[2040] = 0
      "000" when "0011111111001", -- t[2041] = 0
      "000" when "0011111111010", -- t[2042] = 0
      "000" when "0011111111011", -- t[2043] = 0
      "000" when "0011111111100", -- t[2044] = 0
      "000" when "0011111111101", -- t[2045] = 0
      "000" when "0011111111110", -- t[2046] = 0
      "000" when "0011111111111", -- t[2047] = 0
      "000" when "0100000000000", -- t[2048] = 0
      "000" when "0100000000001", -- t[2049] = 0
      "000" when "0100000000010", -- t[2050] = 0
      "000" when "0100000000011", -- t[2051] = 0
      "000" when "0100000000100", -- t[2052] = 0
      "000" when "0100000000101", -- t[2053] = 0
      "000" when "0100000000110", -- t[2054] = 0
      "000" when "0100000000111", -- t[2055] = 0
      "000" when "0100000001000", -- t[2056] = 0
      "000" when "0100000001001", -- t[2057] = 0
      "000" when "0100000001010", -- t[2058] = 0
      "000" when "0100000001011", -- t[2059] = 0
      "000" when "0100000001100", -- t[2060] = 0
      "000" when "0100000001101", -- t[2061] = 0
      "000" when "0100000001110", -- t[2062] = 0
      "000" when "0100000001111", -- t[2063] = 0
      "000" when "0100000010000", -- t[2064] = 0
      "000" when "0100000010001", -- t[2065] = 0
      "000" when "0100000010010", -- t[2066] = 0
      "000" when "0100000010011", -- t[2067] = 0
      "000" when "0100000010100", -- t[2068] = 0
      "000" when "0100000010101", -- t[2069] = 0
      "000" when "0100000010110", -- t[2070] = 0
      "000" when "0100000010111", -- t[2071] = 0
      "000" when "0100000011000", -- t[2072] = 0
      "000" when "0100000011001", -- t[2073] = 0
      "000" when "0100000011010", -- t[2074] = 0
      "000" when "0100000011011", -- t[2075] = 0
      "000" when "0100000011100", -- t[2076] = 0
      "000" when "0100000011101", -- t[2077] = 0
      "000" when "0100000011110", -- t[2078] = 0
      "000" when "0100000011111", -- t[2079] = 0
      "000" when "0100000100000", -- t[2080] = 0
      "000" when "0100000100001", -- t[2081] = 0
      "000" when "0100000100010", -- t[2082] = 0
      "000" when "0100000100011", -- t[2083] = 0
      "000" when "0100000100100", -- t[2084] = 0
      "000" when "0100000100101", -- t[2085] = 0
      "000" when "0100000100110", -- t[2086] = 0
      "000" when "0100000100111", -- t[2087] = 0
      "000" when "0100000101000", -- t[2088] = 0
      "000" when "0100000101001", -- t[2089] = 0
      "000" when "0100000101010", -- t[2090] = 0
      "000" when "0100000101011", -- t[2091] = 0
      "000" when "0100000101100", -- t[2092] = 0
      "000" when "0100000101101", -- t[2093] = 0
      "000" when "0100000101110", -- t[2094] = 0
      "000" when "0100000101111", -- t[2095] = 0
      "000" when "0100000110000", -- t[2096] = 0
      "000" when "0100000110001", -- t[2097] = 0
      "000" when "0100000110010", -- t[2098] = 0
      "000" when "0100000110011", -- t[2099] = 0
      "000" when "0100000110100", -- t[2100] = 0
      "000" when "0100000110101", -- t[2101] = 0
      "000" when "0100000110110", -- t[2102] = 0
      "000" when "0100000110111", -- t[2103] = 0
      "000" when "0100000111000", -- t[2104] = 0
      "000" when "0100000111001", -- t[2105] = 0
      "000" when "0100000111010", -- t[2106] = 0
      "000" when "0100000111011", -- t[2107] = 0
      "000" when "0100000111100", -- t[2108] = 0
      "000" when "0100000111101", -- t[2109] = 0
      "000" when "0100000111110", -- t[2110] = 0
      "000" when "0100000111111", -- t[2111] = 0
      "000" when "0100001000000", -- t[2112] = 0
      "000" when "0100001000001", -- t[2113] = 0
      "000" when "0100001000010", -- t[2114] = 0
      "000" when "0100001000011", -- t[2115] = 0
      "000" when "0100001000100", -- t[2116] = 0
      "000" when "0100001000101", -- t[2117] = 0
      "000" when "0100001000110", -- t[2118] = 0
      "000" when "0100001000111", -- t[2119] = 0
      "000" when "0100001001000", -- t[2120] = 0
      "000" when "0100001001001", -- t[2121] = 0
      "000" when "0100001001010", -- t[2122] = 0
      "000" when "0100001001011", -- t[2123] = 0
      "000" when "0100001001100", -- t[2124] = 0
      "000" when "0100001001101", -- t[2125] = 0
      "000" when "0100001001110", -- t[2126] = 0
      "000" when "0100001001111", -- t[2127] = 0
      "000" when "0100001010000", -- t[2128] = 0
      "000" when "0100001010001", -- t[2129] = 0
      "000" when "0100001010010", -- t[2130] = 0
      "000" when "0100001010011", -- t[2131] = 0
      "000" when "0100001010100", -- t[2132] = 0
      "000" when "0100001010101", -- t[2133] = 0
      "000" when "0100001010110", -- t[2134] = 0
      "000" when "0100001010111", -- t[2135] = 0
      "000" when "0100001011000", -- t[2136] = 0
      "000" when "0100001011001", -- t[2137] = 0
      "000" when "0100001011010", -- t[2138] = 0
      "000" when "0100001011011", -- t[2139] = 0
      "000" when "0100001011100", -- t[2140] = 0
      "000" when "0100001011101", -- t[2141] = 0
      "000" when "0100001011110", -- t[2142] = 0
      "000" when "0100001011111", -- t[2143] = 0
      "000" when "0100001100000", -- t[2144] = 0
      "000" when "0100001100001", -- t[2145] = 0
      "000" when "0100001100010", -- t[2146] = 0
      "000" when "0100001100011", -- t[2147] = 0
      "000" when "0100001100100", -- t[2148] = 0
      "000" when "0100001100101", -- t[2149] = 0
      "000" when "0100001100110", -- t[2150] = 0
      "000" when "0100001100111", -- t[2151] = 0
      "000" when "0100001101000", -- t[2152] = 0
      "000" when "0100001101001", -- t[2153] = 0
      "000" when "0100001101010", -- t[2154] = 0
      "000" when "0100001101011", -- t[2155] = 0
      "000" when "0100001101100", -- t[2156] = 0
      "000" when "0100001101101", -- t[2157] = 0
      "000" when "0100001101110", -- t[2158] = 0
      "000" when "0100001101111", -- t[2159] = 0
      "000" when "0100001110000", -- t[2160] = 0
      "000" when "0100001110001", -- t[2161] = 0
      "000" when "0100001110010", -- t[2162] = 0
      "000" when "0100001110011", -- t[2163] = 0
      "000" when "0100001110100", -- t[2164] = 0
      "000" when "0100001110101", -- t[2165] = 0
      "000" when "0100001110110", -- t[2166] = 0
      "000" when "0100001110111", -- t[2167] = 0
      "000" when "0100001111000", -- t[2168] = 0
      "000" when "0100001111001", -- t[2169] = 0
      "000" when "0100001111010", -- t[2170] = 0
      "000" when "0100001111011", -- t[2171] = 0
      "000" when "0100001111100", -- t[2172] = 0
      "000" when "0100001111101", -- t[2173] = 0
      "000" when "0100001111110", -- t[2174] = 0
      "000" when "0100001111111", -- t[2175] = 0
      "000" when "0100010000000", -- t[2176] = 0
      "000" when "0100010000001", -- t[2177] = 0
      "000" when "0100010000010", -- t[2178] = 0
      "000" when "0100010000011", -- t[2179] = 0
      "000" when "0100010000100", -- t[2180] = 0
      "000" when "0100010000101", -- t[2181] = 0
      "000" when "0100010000110", -- t[2182] = 0
      "000" when "0100010000111", -- t[2183] = 0
      "000" when "0100010001000", -- t[2184] = 0
      "000" when "0100010001001", -- t[2185] = 0
      "000" when "0100010001010", -- t[2186] = 0
      "000" when "0100010001011", -- t[2187] = 0
      "000" when "0100010001100", -- t[2188] = 0
      "000" when "0100010001101", -- t[2189] = 0
      "000" when "0100010001110", -- t[2190] = 0
      "000" when "0100010001111", -- t[2191] = 0
      "000" when "0100010010000", -- t[2192] = 0
      "000" when "0100010010001", -- t[2193] = 0
      "000" when "0100010010010", -- t[2194] = 0
      "000" when "0100010010011", -- t[2195] = 0
      "000" when "0100010010100", -- t[2196] = 0
      "000" when "0100010010101", -- t[2197] = 0
      "000" when "0100010010110", -- t[2198] = 0
      "000" when "0100010010111", -- t[2199] = 0
      "000" when "0100010011000", -- t[2200] = 0
      "000" when "0100010011001", -- t[2201] = 0
      "000" when "0100010011010", -- t[2202] = 0
      "000" when "0100010011011", -- t[2203] = 0
      "000" when "0100010011100", -- t[2204] = 0
      "000" when "0100010011101", -- t[2205] = 0
      "000" when "0100010011110", -- t[2206] = 0
      "000" when "0100010011111", -- t[2207] = 0
      "000" when "0100010100000", -- t[2208] = 0
      "000" when "0100010100001", -- t[2209] = 0
      "000" when "0100010100010", -- t[2210] = 0
      "000" when "0100010100011", -- t[2211] = 0
      "000" when "0100010100100", -- t[2212] = 0
      "000" when "0100010100101", -- t[2213] = 0
      "000" when "0100010100110", -- t[2214] = 0
      "000" when "0100010100111", -- t[2215] = 0
      "000" when "0100010101000", -- t[2216] = 0
      "000" when "0100010101001", -- t[2217] = 0
      "000" when "0100010101010", -- t[2218] = 0
      "000" when "0100010101011", -- t[2219] = 0
      "000" when "0100010101100", -- t[2220] = 0
      "000" when "0100010101101", -- t[2221] = 0
      "000" when "0100010101110", -- t[2222] = 0
      "000" when "0100010101111", -- t[2223] = 0
      "000" when "0100010110000", -- t[2224] = 0
      "000" when "0100010110001", -- t[2225] = 0
      "000" when "0100010110010", -- t[2226] = 0
      "000" when "0100010110011", -- t[2227] = 0
      "000" when "0100010110100", -- t[2228] = 0
      "000" when "0100010110101", -- t[2229] = 0
      "000" when "0100010110110", -- t[2230] = 0
      "000" when "0100010110111", -- t[2231] = 0
      "000" when "0100010111000", -- t[2232] = 0
      "000" when "0100010111001", -- t[2233] = 0
      "000" when "0100010111010", -- t[2234] = 0
      "000" when "0100010111011", -- t[2235] = 0
      "000" when "0100010111100", -- t[2236] = 0
      "000" when "0100010111101", -- t[2237] = 0
      "000" when "0100010111110", -- t[2238] = 0
      "000" when "0100010111111", -- t[2239] = 0
      "000" when "0100011000000", -- t[2240] = 0
      "000" when "0100011000001", -- t[2241] = 0
      "000" when "0100011000010", -- t[2242] = 0
      "000" when "0100011000011", -- t[2243] = 0
      "000" when "0100011000100", -- t[2244] = 0
      "000" when "0100011000101", -- t[2245] = 0
      "000" when "0100011000110", -- t[2246] = 0
      "000" when "0100011000111", -- t[2247] = 0
      "000" when "0100011001000", -- t[2248] = 0
      "000" when "0100011001001", -- t[2249] = 0
      "000" when "0100011001010", -- t[2250] = 0
      "000" when "0100011001011", -- t[2251] = 0
      "000" when "0100011001100", -- t[2252] = 0
      "000" when "0100011001101", -- t[2253] = 0
      "000" when "0100011001110", -- t[2254] = 0
      "000" when "0100011001111", -- t[2255] = 0
      "000" when "0100011010000", -- t[2256] = 0
      "000" when "0100011010001", -- t[2257] = 0
      "000" when "0100011010010", -- t[2258] = 0
      "000" when "0100011010011", -- t[2259] = 0
      "000" when "0100011010100", -- t[2260] = 0
      "000" when "0100011010101", -- t[2261] = 0
      "000" when "0100011010110", -- t[2262] = 0
      "000" when "0100011010111", -- t[2263] = 0
      "000" when "0100011011000", -- t[2264] = 0
      "000" when "0100011011001", -- t[2265] = 0
      "000" when "0100011011010", -- t[2266] = 0
      "000" when "0100011011011", -- t[2267] = 0
      "000" when "0100011011100", -- t[2268] = 0
      "000" when "0100011011101", -- t[2269] = 0
      "000" when "0100011011110", -- t[2270] = 0
      "000" when "0100011011111", -- t[2271] = 0
      "000" when "0100011100000", -- t[2272] = 0
      "000" when "0100011100001", -- t[2273] = 0
      "000" when "0100011100010", -- t[2274] = 0
      "000" when "0100011100011", -- t[2275] = 0
      "000" when "0100011100100", -- t[2276] = 0
      "000" when "0100011100101", -- t[2277] = 0
      "000" when "0100011100110", -- t[2278] = 0
      "000" when "0100011100111", -- t[2279] = 0
      "000" when "0100011101000", -- t[2280] = 0
      "000" when "0100011101001", -- t[2281] = 0
      "000" when "0100011101010", -- t[2282] = 0
      "000" when "0100011101011", -- t[2283] = 0
      "000" when "0100011101100", -- t[2284] = 0
      "000" when "0100011101101", -- t[2285] = 0
      "000" when "0100011101110", -- t[2286] = 0
      "000" when "0100011101111", -- t[2287] = 0
      "000" when "0100011110000", -- t[2288] = 0
      "000" when "0100011110001", -- t[2289] = 0
      "000" when "0100011110010", -- t[2290] = 0
      "000" when "0100011110011", -- t[2291] = 0
      "000" when "0100011110100", -- t[2292] = 0
      "000" when "0100011110101", -- t[2293] = 0
      "000" when "0100011110110", -- t[2294] = 0
      "000" when "0100011110111", -- t[2295] = 0
      "000" when "0100011111000", -- t[2296] = 0
      "000" when "0100011111001", -- t[2297] = 0
      "000" when "0100011111010", -- t[2298] = 0
      "000" when "0100011111011", -- t[2299] = 0
      "000" when "0100011111100", -- t[2300] = 0
      "000" when "0100011111101", -- t[2301] = 0
      "000" when "0100011111110", -- t[2302] = 0
      "000" when "0100011111111", -- t[2303] = 0
      "000" when "0100100000000", -- t[2304] = 0
      "000" when "0100100000001", -- t[2305] = 0
      "000" when "0100100000010", -- t[2306] = 0
      "000" when "0100100000011", -- t[2307] = 0
      "000" when "0100100000100", -- t[2308] = 0
      "000" when "0100100000101", -- t[2309] = 0
      "000" when "0100100000110", -- t[2310] = 0
      "000" when "0100100000111", -- t[2311] = 0
      "000" when "0100100001000", -- t[2312] = 0
      "000" when "0100100001001", -- t[2313] = 0
      "000" when "0100100001010", -- t[2314] = 0
      "000" when "0100100001011", -- t[2315] = 0
      "000" when "0100100001100", -- t[2316] = 0
      "000" when "0100100001101", -- t[2317] = 0
      "000" when "0100100001110", -- t[2318] = 0
      "000" when "0100100001111", -- t[2319] = 0
      "000" when "0100100010000", -- t[2320] = 0
      "000" when "0100100010001", -- t[2321] = 0
      "000" when "0100100010010", -- t[2322] = 0
      "000" when "0100100010011", -- t[2323] = 0
      "000" when "0100100010100", -- t[2324] = 0
      "000" when "0100100010101", -- t[2325] = 0
      "000" when "0100100010110", -- t[2326] = 0
      "000" when "0100100010111", -- t[2327] = 0
      "000" when "0100100011000", -- t[2328] = 0
      "000" when "0100100011001", -- t[2329] = 0
      "000" when "0100100011010", -- t[2330] = 0
      "000" when "0100100011011", -- t[2331] = 0
      "000" when "0100100011100", -- t[2332] = 0
      "000" when "0100100011101", -- t[2333] = 0
      "000" when "0100100011110", -- t[2334] = 0
      "000" when "0100100011111", -- t[2335] = 0
      "000" when "0100100100000", -- t[2336] = 0
      "000" when "0100100100001", -- t[2337] = 0
      "000" when "0100100100010", -- t[2338] = 0
      "000" when "0100100100011", -- t[2339] = 0
      "000" when "0100100100100", -- t[2340] = 0
      "000" when "0100100100101", -- t[2341] = 0
      "000" when "0100100100110", -- t[2342] = 0
      "000" when "0100100100111", -- t[2343] = 0
      "000" when "0100100101000", -- t[2344] = 0
      "000" when "0100100101001", -- t[2345] = 0
      "000" when "0100100101010", -- t[2346] = 0
      "000" when "0100100101011", -- t[2347] = 0
      "000" when "0100100101100", -- t[2348] = 0
      "000" when "0100100101101", -- t[2349] = 0
      "000" when "0100100101110", -- t[2350] = 0
      "000" when "0100100101111", -- t[2351] = 0
      "000" when "0100100110000", -- t[2352] = 0
      "000" when "0100100110001", -- t[2353] = 0
      "000" when "0100100110010", -- t[2354] = 0
      "000" when "0100100110011", -- t[2355] = 0
      "000" when "0100100110100", -- t[2356] = 0
      "000" when "0100100110101", -- t[2357] = 0
      "000" when "0100100110110", -- t[2358] = 0
      "000" when "0100100110111", -- t[2359] = 0
      "000" when "0100100111000", -- t[2360] = 0
      "000" when "0100100111001", -- t[2361] = 0
      "000" when "0100100111010", -- t[2362] = 0
      "000" when "0100100111011", -- t[2363] = 0
      "000" when "0100100111100", -- t[2364] = 0
      "000" when "0100100111101", -- t[2365] = 0
      "000" when "0100100111110", -- t[2366] = 0
      "000" when "0100100111111", -- t[2367] = 0
      "000" when "0100101000000", -- t[2368] = 0
      "000" when "0100101000001", -- t[2369] = 0
      "000" when "0100101000010", -- t[2370] = 0
      "000" when "0100101000011", -- t[2371] = 0
      "000" when "0100101000100", -- t[2372] = 0
      "000" when "0100101000101", -- t[2373] = 0
      "000" when "0100101000110", -- t[2374] = 0
      "000" when "0100101000111", -- t[2375] = 0
      "000" when "0100101001000", -- t[2376] = 0
      "000" when "0100101001001", -- t[2377] = 0
      "000" when "0100101001010", -- t[2378] = 0
      "000" when "0100101001011", -- t[2379] = 0
      "000" when "0100101001100", -- t[2380] = 0
      "000" when "0100101001101", -- t[2381] = 0
      "000" when "0100101001110", -- t[2382] = 0
      "000" when "0100101001111", -- t[2383] = 0
      "000" when "0100101010000", -- t[2384] = 0
      "000" when "0100101010001", -- t[2385] = 0
      "000" when "0100101010010", -- t[2386] = 0
      "000" when "0100101010011", -- t[2387] = 0
      "000" when "0100101010100", -- t[2388] = 0
      "000" when "0100101010101", -- t[2389] = 0
      "000" when "0100101010110", -- t[2390] = 0
      "000" when "0100101010111", -- t[2391] = 0
      "000" when "0100101011000", -- t[2392] = 0
      "000" when "0100101011001", -- t[2393] = 0
      "000" when "0100101011010", -- t[2394] = 0
      "000" when "0100101011011", -- t[2395] = 0
      "000" when "0100101011100", -- t[2396] = 0
      "000" when "0100101011101", -- t[2397] = 0
      "000" when "0100101011110", -- t[2398] = 0
      "000" when "0100101011111", -- t[2399] = 0
      "000" when "0100101100000", -- t[2400] = 0
      "000" when "0100101100001", -- t[2401] = 0
      "000" when "0100101100010", -- t[2402] = 0
      "000" when "0100101100011", -- t[2403] = 0
      "000" when "0100101100100", -- t[2404] = 0
      "000" when "0100101100101", -- t[2405] = 0
      "000" when "0100101100110", -- t[2406] = 0
      "000" when "0100101100111", -- t[2407] = 0
      "000" when "0100101101000", -- t[2408] = 0
      "000" when "0100101101001", -- t[2409] = 0
      "000" when "0100101101010", -- t[2410] = 0
      "000" when "0100101101011", -- t[2411] = 0
      "000" when "0100101101100", -- t[2412] = 0
      "000" when "0100101101101", -- t[2413] = 0
      "000" when "0100101101110", -- t[2414] = 0
      "000" when "0100101101111", -- t[2415] = 0
      "000" when "0100101110000", -- t[2416] = 0
      "000" when "0100101110001", -- t[2417] = 0
      "000" when "0100101110010", -- t[2418] = 0
      "000" when "0100101110011", -- t[2419] = 0
      "000" when "0100101110100", -- t[2420] = 0
      "000" when "0100101110101", -- t[2421] = 0
      "000" when "0100101110110", -- t[2422] = 0
      "000" when "0100101110111", -- t[2423] = 0
      "000" when "0100101111000", -- t[2424] = 0
      "000" when "0100101111001", -- t[2425] = 0
      "000" when "0100101111010", -- t[2426] = 0
      "000" when "0100101111011", -- t[2427] = 0
      "000" when "0100101111100", -- t[2428] = 0
      "000" when "0100101111101", -- t[2429] = 0
      "000" when "0100101111110", -- t[2430] = 0
      "000" when "0100101111111", -- t[2431] = 0
      "000" when "0100110000000", -- t[2432] = 0
      "000" when "0100110000001", -- t[2433] = 0
      "000" when "0100110000010", -- t[2434] = 0
      "000" when "0100110000011", -- t[2435] = 0
      "000" when "0100110000100", -- t[2436] = 0
      "000" when "0100110000101", -- t[2437] = 0
      "000" when "0100110000110", -- t[2438] = 0
      "000" when "0100110000111", -- t[2439] = 0
      "000" when "0100110001000", -- t[2440] = 0
      "000" when "0100110001001", -- t[2441] = 0
      "000" when "0100110001010", -- t[2442] = 0
      "000" when "0100110001011", -- t[2443] = 0
      "000" when "0100110001100", -- t[2444] = 0
      "000" when "0100110001101", -- t[2445] = 0
      "000" when "0100110001110", -- t[2446] = 0
      "000" when "0100110001111", -- t[2447] = 0
      "000" when "0100110010000", -- t[2448] = 0
      "000" when "0100110010001", -- t[2449] = 0
      "000" when "0100110010010", -- t[2450] = 0
      "000" when "0100110010011", -- t[2451] = 0
      "000" when "0100110010100", -- t[2452] = 0
      "000" when "0100110010101", -- t[2453] = 0
      "000" when "0100110010110", -- t[2454] = 0
      "000" when "0100110010111", -- t[2455] = 0
      "000" when "0100110011000", -- t[2456] = 0
      "000" when "0100110011001", -- t[2457] = 0
      "000" when "0100110011010", -- t[2458] = 0
      "000" when "0100110011011", -- t[2459] = 0
      "000" when "0100110011100", -- t[2460] = 0
      "000" when "0100110011101", -- t[2461] = 0
      "000" when "0100110011110", -- t[2462] = 0
      "000" when "0100110011111", -- t[2463] = 0
      "000" when "0100110100000", -- t[2464] = 0
      "000" when "0100110100001", -- t[2465] = 0
      "000" when "0100110100010", -- t[2466] = 0
      "000" when "0100110100011", -- t[2467] = 0
      "000" when "0100110100100", -- t[2468] = 0
      "000" when "0100110100101", -- t[2469] = 0
      "000" when "0100110100110", -- t[2470] = 0
      "000" when "0100110100111", -- t[2471] = 0
      "000" when "0100110101000", -- t[2472] = 0
      "000" when "0100110101001", -- t[2473] = 0
      "000" when "0100110101010", -- t[2474] = 0
      "000" when "0100110101011", -- t[2475] = 0
      "000" when "0100110101100", -- t[2476] = 0
      "000" when "0100110101101", -- t[2477] = 0
      "000" when "0100110101110", -- t[2478] = 0
      "000" when "0100110101111", -- t[2479] = 0
      "000" when "0100110110000", -- t[2480] = 0
      "000" when "0100110110001", -- t[2481] = 0
      "000" when "0100110110010", -- t[2482] = 0
      "000" when "0100110110011", -- t[2483] = 0
      "000" when "0100110110100", -- t[2484] = 0
      "000" when "0100110110101", -- t[2485] = 0
      "000" when "0100110110110", -- t[2486] = 0
      "000" when "0100110110111", -- t[2487] = 0
      "000" when "0100110111000", -- t[2488] = 0
      "000" when "0100110111001", -- t[2489] = 0
      "000" when "0100110111010", -- t[2490] = 0
      "000" when "0100110111011", -- t[2491] = 0
      "000" when "0100110111100", -- t[2492] = 0
      "000" when "0100110111101", -- t[2493] = 0
      "000" when "0100110111110", -- t[2494] = 0
      "000" when "0100110111111", -- t[2495] = 0
      "000" when "0100111000000", -- t[2496] = 0
      "000" when "0100111000001", -- t[2497] = 0
      "000" when "0100111000010", -- t[2498] = 0
      "000" when "0100111000011", -- t[2499] = 0
      "000" when "0100111000100", -- t[2500] = 0
      "000" when "0100111000101", -- t[2501] = 0
      "000" when "0100111000110", -- t[2502] = 0
      "000" when "0100111000111", -- t[2503] = 0
      "000" when "0100111001000", -- t[2504] = 0
      "000" when "0100111001001", -- t[2505] = 0
      "000" when "0100111001010", -- t[2506] = 0
      "000" when "0100111001011", -- t[2507] = 0
      "000" when "0100111001100", -- t[2508] = 0
      "000" when "0100111001101", -- t[2509] = 0
      "000" when "0100111001110", -- t[2510] = 0
      "000" when "0100111001111", -- t[2511] = 0
      "000" when "0100111010000", -- t[2512] = 0
      "000" when "0100111010001", -- t[2513] = 0
      "000" when "0100111010010", -- t[2514] = 0
      "000" when "0100111010011", -- t[2515] = 0
      "000" when "0100111010100", -- t[2516] = 0
      "000" when "0100111010101", -- t[2517] = 0
      "000" when "0100111010110", -- t[2518] = 0
      "000" when "0100111010111", -- t[2519] = 0
      "000" when "0100111011000", -- t[2520] = 0
      "000" when "0100111011001", -- t[2521] = 0
      "000" when "0100111011010", -- t[2522] = 0
      "000" when "0100111011011", -- t[2523] = 0
      "000" when "0100111011100", -- t[2524] = 0
      "000" when "0100111011101", -- t[2525] = 0
      "000" when "0100111011110", -- t[2526] = 0
      "000" when "0100111011111", -- t[2527] = 0
      "000" when "0100111100000", -- t[2528] = 0
      "000" when "0100111100001", -- t[2529] = 0
      "000" when "0100111100010", -- t[2530] = 0
      "000" when "0100111100011", -- t[2531] = 0
      "000" when "0100111100100", -- t[2532] = 0
      "000" when "0100111100101", -- t[2533] = 0
      "000" when "0100111100110", -- t[2534] = 0
      "000" when "0100111100111", -- t[2535] = 0
      "000" when "0100111101000", -- t[2536] = 0
      "000" when "0100111101001", -- t[2537] = 0
      "000" when "0100111101010", -- t[2538] = 0
      "000" when "0100111101011", -- t[2539] = 0
      "000" when "0100111101100", -- t[2540] = 0
      "000" when "0100111101101", -- t[2541] = 0
      "000" when "0100111101110", -- t[2542] = 0
      "000" when "0100111101111", -- t[2543] = 0
      "000" when "0100111110000", -- t[2544] = 0
      "000" when "0100111110001", -- t[2545] = 0
      "000" when "0100111110010", -- t[2546] = 0
      "000" when "0100111110011", -- t[2547] = 0
      "000" when "0100111110100", -- t[2548] = 0
      "000" when "0100111110101", -- t[2549] = 0
      "000" when "0100111110110", -- t[2550] = 0
      "000" when "0100111110111", -- t[2551] = 0
      "000" when "0100111111000", -- t[2552] = 0
      "000" when "0100111111001", -- t[2553] = 0
      "000" when "0100111111010", -- t[2554] = 0
      "000" when "0100111111011", -- t[2555] = 0
      "000" when "0100111111100", -- t[2556] = 0
      "000" when "0100111111101", -- t[2557] = 0
      "000" when "0100111111110", -- t[2558] = 0
      "000" when "0100111111111", -- t[2559] = 0
      "000" when "0101000000000", -- t[2560] = 0
      "000" when "0101000000001", -- t[2561] = 0
      "000" when "0101000000010", -- t[2562] = 0
      "000" when "0101000000011", -- t[2563] = 0
      "000" when "0101000000100", -- t[2564] = 0
      "000" when "0101000000101", -- t[2565] = 0
      "000" when "0101000000110", -- t[2566] = 0
      "000" when "0101000000111", -- t[2567] = 0
      "000" when "0101000001000", -- t[2568] = 0
      "000" when "0101000001001", -- t[2569] = 0
      "000" when "0101000001010", -- t[2570] = 0
      "000" when "0101000001011", -- t[2571] = 0
      "000" when "0101000001100", -- t[2572] = 0
      "000" when "0101000001101", -- t[2573] = 0
      "000" when "0101000001110", -- t[2574] = 0
      "000" when "0101000001111", -- t[2575] = 0
      "000" when "0101000010000", -- t[2576] = 0
      "000" when "0101000010001", -- t[2577] = 0
      "000" when "0101000010010", -- t[2578] = 0
      "000" when "0101000010011", -- t[2579] = 0
      "000" when "0101000010100", -- t[2580] = 0
      "000" when "0101000010101", -- t[2581] = 0
      "000" when "0101000010110", -- t[2582] = 0
      "000" when "0101000010111", -- t[2583] = 0
      "000" when "0101000011000", -- t[2584] = 0
      "000" when "0101000011001", -- t[2585] = 0
      "000" when "0101000011010", -- t[2586] = 0
      "000" when "0101000011011", -- t[2587] = 0
      "000" when "0101000011100", -- t[2588] = 0
      "000" when "0101000011101", -- t[2589] = 0
      "000" when "0101000011110", -- t[2590] = 0
      "000" when "0101000011111", -- t[2591] = 0
      "000" when "0101000100000", -- t[2592] = 0
      "000" when "0101000100001", -- t[2593] = 0
      "000" when "0101000100010", -- t[2594] = 0
      "000" when "0101000100011", -- t[2595] = 0
      "000" when "0101000100100", -- t[2596] = 0
      "000" when "0101000100101", -- t[2597] = 0
      "000" when "0101000100110", -- t[2598] = 0
      "000" when "0101000100111", -- t[2599] = 0
      "000" when "0101000101000", -- t[2600] = 0
      "000" when "0101000101001", -- t[2601] = 0
      "000" when "0101000101010", -- t[2602] = 0
      "000" when "0101000101011", -- t[2603] = 0
      "000" when "0101000101100", -- t[2604] = 0
      "000" when "0101000101101", -- t[2605] = 0
      "000" when "0101000101110", -- t[2606] = 0
      "000" when "0101000101111", -- t[2607] = 0
      "000" when "0101000110000", -- t[2608] = 0
      "000" when "0101000110001", -- t[2609] = 0
      "000" when "0101000110010", -- t[2610] = 0
      "000" when "0101000110011", -- t[2611] = 0
      "000" when "0101000110100", -- t[2612] = 0
      "000" when "0101000110101", -- t[2613] = 0
      "000" when "0101000110110", -- t[2614] = 0
      "000" when "0101000110111", -- t[2615] = 0
      "000" when "0101000111000", -- t[2616] = 0
      "000" when "0101000111001", -- t[2617] = 0
      "000" when "0101000111010", -- t[2618] = 0
      "000" when "0101000111011", -- t[2619] = 0
      "000" when "0101000111100", -- t[2620] = 0
      "000" when "0101000111101", -- t[2621] = 0
      "000" when "0101000111110", -- t[2622] = 0
      "000" when "0101000111111", -- t[2623] = 0
      "000" when "0101001000000", -- t[2624] = 0
      "000" when "0101001000001", -- t[2625] = 0
      "000" when "0101001000010", -- t[2626] = 0
      "000" when "0101001000011", -- t[2627] = 0
      "000" when "0101001000100", -- t[2628] = 0
      "000" when "0101001000101", -- t[2629] = 0
      "000" when "0101001000110", -- t[2630] = 0
      "000" when "0101001000111", -- t[2631] = 0
      "000" when "0101001001000", -- t[2632] = 0
      "000" when "0101001001001", -- t[2633] = 0
      "000" when "0101001001010", -- t[2634] = 0
      "000" when "0101001001011", -- t[2635] = 0
      "000" when "0101001001100", -- t[2636] = 0
      "000" when "0101001001101", -- t[2637] = 0
      "000" when "0101001001110", -- t[2638] = 0
      "000" when "0101001001111", -- t[2639] = 0
      "000" when "0101001010000", -- t[2640] = 0
      "000" when "0101001010001", -- t[2641] = 0
      "000" when "0101001010010", -- t[2642] = 0
      "000" when "0101001010011", -- t[2643] = 0
      "000" when "0101001010100", -- t[2644] = 0
      "000" when "0101001010101", -- t[2645] = 0
      "000" when "0101001010110", -- t[2646] = 0
      "000" when "0101001010111", -- t[2647] = 0
      "000" when "0101001011000", -- t[2648] = 0
      "000" when "0101001011001", -- t[2649] = 0
      "000" when "0101001011010", -- t[2650] = 0
      "000" when "0101001011011", -- t[2651] = 0
      "000" when "0101001011100", -- t[2652] = 0
      "000" when "0101001011101", -- t[2653] = 0
      "000" when "0101001011110", -- t[2654] = 0
      "000" when "0101001011111", -- t[2655] = 0
      "000" when "0101001100000", -- t[2656] = 0
      "000" when "0101001100001", -- t[2657] = 0
      "000" when "0101001100010", -- t[2658] = 0
      "000" when "0101001100011", -- t[2659] = 0
      "000" when "0101001100100", -- t[2660] = 0
      "000" when "0101001100101", -- t[2661] = 0
      "000" when "0101001100110", -- t[2662] = 0
      "000" when "0101001100111", -- t[2663] = 0
      "000" when "0101001101000", -- t[2664] = 0
      "000" when "0101001101001", -- t[2665] = 0
      "000" when "0101001101010", -- t[2666] = 0
      "000" when "0101001101011", -- t[2667] = 0
      "000" when "0101001101100", -- t[2668] = 0
      "000" when "0101001101101", -- t[2669] = 0
      "000" when "0101001101110", -- t[2670] = 0
      "000" when "0101001101111", -- t[2671] = 0
      "000" when "0101001110000", -- t[2672] = 0
      "000" when "0101001110001", -- t[2673] = 0
      "000" when "0101001110010", -- t[2674] = 0
      "000" when "0101001110011", -- t[2675] = 0
      "000" when "0101001110100", -- t[2676] = 0
      "000" when "0101001110101", -- t[2677] = 0
      "000" when "0101001110110", -- t[2678] = 0
      "000" when "0101001110111", -- t[2679] = 0
      "000" when "0101001111000", -- t[2680] = 0
      "000" when "0101001111001", -- t[2681] = 0
      "000" when "0101001111010", -- t[2682] = 0
      "000" when "0101001111011", -- t[2683] = 0
      "000" when "0101001111100", -- t[2684] = 0
      "000" when "0101001111101", -- t[2685] = 0
      "000" when "0101001111110", -- t[2686] = 0
      "000" when "0101001111111", -- t[2687] = 0
      "000" when "0101010000000", -- t[2688] = 0
      "000" when "0101010000001", -- t[2689] = 0
      "000" when "0101010000010", -- t[2690] = 0
      "000" when "0101010000011", -- t[2691] = 0
      "000" when "0101010000100", -- t[2692] = 0
      "000" when "0101010000101", -- t[2693] = 0
      "000" when "0101010000110", -- t[2694] = 0
      "000" when "0101010000111", -- t[2695] = 0
      "000" when "0101010001000", -- t[2696] = 0
      "000" when "0101010001001", -- t[2697] = 0
      "000" when "0101010001010", -- t[2698] = 0
      "000" when "0101010001011", -- t[2699] = 0
      "000" when "0101010001100", -- t[2700] = 0
      "000" when "0101010001101", -- t[2701] = 0
      "000" when "0101010001110", -- t[2702] = 0
      "000" when "0101010001111", -- t[2703] = 0
      "000" when "0101010010000", -- t[2704] = 0
      "000" when "0101010010001", -- t[2705] = 0
      "000" when "0101010010010", -- t[2706] = 0
      "000" when "0101010010011", -- t[2707] = 0
      "000" when "0101010010100", -- t[2708] = 0
      "000" when "0101010010101", -- t[2709] = 0
      "000" when "0101010010110", -- t[2710] = 0
      "000" when "0101010010111", -- t[2711] = 0
      "000" when "0101010011000", -- t[2712] = 0
      "000" when "0101010011001", -- t[2713] = 0
      "000" when "0101010011010", -- t[2714] = 0
      "000" when "0101010011011", -- t[2715] = 0
      "000" when "0101010011100", -- t[2716] = 0
      "000" when "0101010011101", -- t[2717] = 0
      "000" when "0101010011110", -- t[2718] = 0
      "000" when "0101010011111", -- t[2719] = 0
      "000" when "0101010100000", -- t[2720] = 0
      "000" when "0101010100001", -- t[2721] = 0
      "000" when "0101010100010", -- t[2722] = 0
      "000" when "0101010100011", -- t[2723] = 0
      "000" when "0101010100100", -- t[2724] = 0
      "000" when "0101010100101", -- t[2725] = 0
      "000" when "0101010100110", -- t[2726] = 0
      "000" when "0101010100111", -- t[2727] = 0
      "000" when "0101010101000", -- t[2728] = 0
      "000" when "0101010101001", -- t[2729] = 0
      "000" when "0101010101010", -- t[2730] = 0
      "000" when "0101010101011", -- t[2731] = 0
      "000" when "0101010101100", -- t[2732] = 0
      "000" when "0101010101101", -- t[2733] = 0
      "000" when "0101010101110", -- t[2734] = 0
      "000" when "0101010101111", -- t[2735] = 0
      "000" when "0101010110000", -- t[2736] = 0
      "000" when "0101010110001", -- t[2737] = 0
      "000" when "0101010110010", -- t[2738] = 0
      "000" when "0101010110011", -- t[2739] = 0
      "000" when "0101010110100", -- t[2740] = 0
      "000" when "0101010110101", -- t[2741] = 0
      "000" when "0101010110110", -- t[2742] = 0
      "000" when "0101010110111", -- t[2743] = 0
      "000" when "0101010111000", -- t[2744] = 0
      "000" when "0101010111001", -- t[2745] = 0
      "000" when "0101010111010", -- t[2746] = 0
      "000" when "0101010111011", -- t[2747] = 0
      "000" when "0101010111100", -- t[2748] = 0
      "000" when "0101010111101", -- t[2749] = 0
      "000" when "0101010111110", -- t[2750] = 0
      "000" when "0101010111111", -- t[2751] = 0
      "000" when "0101011000000", -- t[2752] = 0
      "000" when "0101011000001", -- t[2753] = 0
      "000" when "0101011000010", -- t[2754] = 0
      "000" when "0101011000011", -- t[2755] = 0
      "000" when "0101011000100", -- t[2756] = 0
      "000" when "0101011000101", -- t[2757] = 0
      "000" when "0101011000110", -- t[2758] = 0
      "000" when "0101011000111", -- t[2759] = 0
      "000" when "0101011001000", -- t[2760] = 0
      "000" when "0101011001001", -- t[2761] = 0
      "000" when "0101011001010", -- t[2762] = 0
      "000" when "0101011001011", -- t[2763] = 0
      "000" when "0101011001100", -- t[2764] = 0
      "000" when "0101011001101", -- t[2765] = 0
      "000" when "0101011001110", -- t[2766] = 0
      "000" when "0101011001111", -- t[2767] = 0
      "000" when "0101011010000", -- t[2768] = 0
      "000" when "0101011010001", -- t[2769] = 0
      "000" when "0101011010010", -- t[2770] = 0
      "000" when "0101011010011", -- t[2771] = 0
      "000" when "0101011010100", -- t[2772] = 0
      "000" when "0101011010101", -- t[2773] = 0
      "000" when "0101011010110", -- t[2774] = 0
      "000" when "0101011010111", -- t[2775] = 0
      "000" when "0101011011000", -- t[2776] = 0
      "000" when "0101011011001", -- t[2777] = 0
      "000" when "0101011011010", -- t[2778] = 0
      "000" when "0101011011011", -- t[2779] = 0
      "000" when "0101011011100", -- t[2780] = 0
      "000" when "0101011011101", -- t[2781] = 0
      "000" when "0101011011110", -- t[2782] = 0
      "000" when "0101011011111", -- t[2783] = 0
      "000" when "0101011100000", -- t[2784] = 0
      "000" when "0101011100001", -- t[2785] = 0
      "000" when "0101011100010", -- t[2786] = 0
      "000" when "0101011100011", -- t[2787] = 0
      "000" when "0101011100100", -- t[2788] = 0
      "000" when "0101011100101", -- t[2789] = 0
      "000" when "0101011100110", -- t[2790] = 0
      "000" when "0101011100111", -- t[2791] = 0
      "000" when "0101011101000", -- t[2792] = 0
      "000" when "0101011101001", -- t[2793] = 0
      "000" when "0101011101010", -- t[2794] = 0
      "000" when "0101011101011", -- t[2795] = 0
      "000" when "0101011101100", -- t[2796] = 0
      "000" when "0101011101101", -- t[2797] = 0
      "000" when "0101011101110", -- t[2798] = 0
      "000" when "0101011101111", -- t[2799] = 0
      "000" when "0101011110000", -- t[2800] = 0
      "000" when "0101011110001", -- t[2801] = 0
      "001" when "0101011110010", -- t[2802] = 1
      "001" when "0101011110011", -- t[2803] = 1
      "001" when "0101011110100", -- t[2804] = 1
      "001" when "0101011110101", -- t[2805] = 1
      "001" when "0101011110110", -- t[2806] = 1
      "001" when "0101011110111", -- t[2807] = 1
      "001" when "0101011111000", -- t[2808] = 1
      "001" when "0101011111001", -- t[2809] = 1
      "001" when "0101011111010", -- t[2810] = 1
      "001" when "0101011111011", -- t[2811] = 1
      "001" when "0101011111100", -- t[2812] = 1
      "001" when "0101011111101", -- t[2813] = 1
      "001" when "0101011111110", -- t[2814] = 1
      "001" when "0101011111111", -- t[2815] = 1
      "001" when "0101100000000", -- t[2816] = 1
      "001" when "0101100000001", -- t[2817] = 1
      "001" when "0101100000010", -- t[2818] = 1
      "001" when "0101100000011", -- t[2819] = 1
      "001" when "0101100000100", -- t[2820] = 1
      "001" when "0101100000101", -- t[2821] = 1
      "001" when "0101100000110", -- t[2822] = 1
      "001" when "0101100000111", -- t[2823] = 1
      "001" when "0101100001000", -- t[2824] = 1
      "001" when "0101100001001", -- t[2825] = 1
      "001" when "0101100001010", -- t[2826] = 1
      "001" when "0101100001011", -- t[2827] = 1
      "001" when "0101100001100", -- t[2828] = 1
      "001" when "0101100001101", -- t[2829] = 1
      "001" when "0101100001110", -- t[2830] = 1
      "001" when "0101100001111", -- t[2831] = 1
      "001" when "0101100010000", -- t[2832] = 1
      "001" when "0101100010001", -- t[2833] = 1
      "001" when "0101100010010", -- t[2834] = 1
      "001" when "0101100010011", -- t[2835] = 1
      "001" when "0101100010100", -- t[2836] = 1
      "001" when "0101100010101", -- t[2837] = 1
      "001" when "0101100010110", -- t[2838] = 1
      "001" when "0101100010111", -- t[2839] = 1
      "001" when "0101100011000", -- t[2840] = 1
      "001" when "0101100011001", -- t[2841] = 1
      "001" when "0101100011010", -- t[2842] = 1
      "001" when "0101100011011", -- t[2843] = 1
      "001" when "0101100011100", -- t[2844] = 1
      "001" when "0101100011101", -- t[2845] = 1
      "001" when "0101100011110", -- t[2846] = 1
      "001" when "0101100011111", -- t[2847] = 1
      "001" when "0101100100000", -- t[2848] = 1
      "001" when "0101100100001", -- t[2849] = 1
      "001" when "0101100100010", -- t[2850] = 1
      "001" when "0101100100011", -- t[2851] = 1
      "001" when "0101100100100", -- t[2852] = 1
      "001" when "0101100100101", -- t[2853] = 1
      "001" when "0101100100110", -- t[2854] = 1
      "001" when "0101100100111", -- t[2855] = 1
      "001" when "0101100101000", -- t[2856] = 1
      "001" when "0101100101001", -- t[2857] = 1
      "001" when "0101100101010", -- t[2858] = 1
      "001" when "0101100101011", -- t[2859] = 1
      "001" when "0101100101100", -- t[2860] = 1
      "001" when "0101100101101", -- t[2861] = 1
      "001" when "0101100101110", -- t[2862] = 1
      "001" when "0101100101111", -- t[2863] = 1
      "001" when "0101100110000", -- t[2864] = 1
      "001" when "0101100110001", -- t[2865] = 1
      "001" when "0101100110010", -- t[2866] = 1
      "001" when "0101100110011", -- t[2867] = 1
      "001" when "0101100110100", -- t[2868] = 1
      "001" when "0101100110101", -- t[2869] = 1
      "001" when "0101100110110", -- t[2870] = 1
      "001" when "0101100110111", -- t[2871] = 1
      "001" when "0101100111000", -- t[2872] = 1
      "001" when "0101100111001", -- t[2873] = 1
      "001" when "0101100111010", -- t[2874] = 1
      "001" when "0101100111011", -- t[2875] = 1
      "001" when "0101100111100", -- t[2876] = 1
      "001" when "0101100111101", -- t[2877] = 1
      "001" when "0101100111110", -- t[2878] = 1
      "001" when "0101100111111", -- t[2879] = 1
      "001" when "0101101000000", -- t[2880] = 1
      "001" when "0101101000001", -- t[2881] = 1
      "001" when "0101101000010", -- t[2882] = 1
      "001" when "0101101000011", -- t[2883] = 1
      "001" when "0101101000100", -- t[2884] = 1
      "001" when "0101101000101", -- t[2885] = 1
      "001" when "0101101000110", -- t[2886] = 1
      "001" when "0101101000111", -- t[2887] = 1
      "001" when "0101101001000", -- t[2888] = 1
      "001" when "0101101001001", -- t[2889] = 1
      "001" when "0101101001010", -- t[2890] = 1
      "001" when "0101101001011", -- t[2891] = 1
      "001" when "0101101001100", -- t[2892] = 1
      "001" when "0101101001101", -- t[2893] = 1
      "001" when "0101101001110", -- t[2894] = 1
      "001" when "0101101001111", -- t[2895] = 1
      "001" when "0101101010000", -- t[2896] = 1
      "001" when "0101101010001", -- t[2897] = 1
      "001" when "0101101010010", -- t[2898] = 1
      "001" when "0101101010011", -- t[2899] = 1
      "001" when "0101101010100", -- t[2900] = 1
      "001" when "0101101010101", -- t[2901] = 1
      "001" when "0101101010110", -- t[2902] = 1
      "001" when "0101101010111", -- t[2903] = 1
      "001" when "0101101011000", -- t[2904] = 1
      "001" when "0101101011001", -- t[2905] = 1
      "001" when "0101101011010", -- t[2906] = 1
      "001" when "0101101011011", -- t[2907] = 1
      "001" when "0101101011100", -- t[2908] = 1
      "001" when "0101101011101", -- t[2909] = 1
      "001" when "0101101011110", -- t[2910] = 1
      "001" when "0101101011111", -- t[2911] = 1
      "001" when "0101101100000", -- t[2912] = 1
      "001" when "0101101100001", -- t[2913] = 1
      "001" when "0101101100010", -- t[2914] = 1
      "001" when "0101101100011", -- t[2915] = 1
      "001" when "0101101100100", -- t[2916] = 1
      "001" when "0101101100101", -- t[2917] = 1
      "001" when "0101101100110", -- t[2918] = 1
      "001" when "0101101100111", -- t[2919] = 1
      "001" when "0101101101000", -- t[2920] = 1
      "001" when "0101101101001", -- t[2921] = 1
      "001" when "0101101101010", -- t[2922] = 1
      "001" when "0101101101011", -- t[2923] = 1
      "001" when "0101101101100", -- t[2924] = 1
      "001" when "0101101101101", -- t[2925] = 1
      "001" when "0101101101110", -- t[2926] = 1
      "001" when "0101101101111", -- t[2927] = 1
      "001" when "0101101110000", -- t[2928] = 1
      "001" when "0101101110001", -- t[2929] = 1
      "001" when "0101101110010", -- t[2930] = 1
      "001" when "0101101110011", -- t[2931] = 1
      "001" when "0101101110100", -- t[2932] = 1
      "001" when "0101101110101", -- t[2933] = 1
      "001" when "0101101110110", -- t[2934] = 1
      "001" when "0101101110111", -- t[2935] = 1
      "001" when "0101101111000", -- t[2936] = 1
      "001" when "0101101111001", -- t[2937] = 1
      "001" when "0101101111010", -- t[2938] = 1
      "001" when "0101101111011", -- t[2939] = 1
      "001" when "0101101111100", -- t[2940] = 1
      "001" when "0101101111101", -- t[2941] = 1
      "001" when "0101101111110", -- t[2942] = 1
      "001" when "0101101111111", -- t[2943] = 1
      "001" when "0101110000000", -- t[2944] = 1
      "001" when "0101110000001", -- t[2945] = 1
      "001" when "0101110000010", -- t[2946] = 1
      "001" when "0101110000011", -- t[2947] = 1
      "001" when "0101110000100", -- t[2948] = 1
      "001" when "0101110000101", -- t[2949] = 1
      "001" when "0101110000110", -- t[2950] = 1
      "001" when "0101110000111", -- t[2951] = 1
      "001" when "0101110001000", -- t[2952] = 1
      "001" when "0101110001001", -- t[2953] = 1
      "001" when "0101110001010", -- t[2954] = 1
      "001" when "0101110001011", -- t[2955] = 1
      "001" when "0101110001100", -- t[2956] = 1
      "001" when "0101110001101", -- t[2957] = 1
      "001" when "0101110001110", -- t[2958] = 1
      "001" when "0101110001111", -- t[2959] = 1
      "001" when "0101110010000", -- t[2960] = 1
      "001" when "0101110010001", -- t[2961] = 1
      "001" when "0101110010010", -- t[2962] = 1
      "001" when "0101110010011", -- t[2963] = 1
      "001" when "0101110010100", -- t[2964] = 1
      "001" when "0101110010101", -- t[2965] = 1
      "001" when "0101110010110", -- t[2966] = 1
      "001" when "0101110010111", -- t[2967] = 1
      "001" when "0101110011000", -- t[2968] = 1
      "001" when "0101110011001", -- t[2969] = 1
      "001" when "0101110011010", -- t[2970] = 1
      "001" when "0101110011011", -- t[2971] = 1
      "001" when "0101110011100", -- t[2972] = 1
      "001" when "0101110011101", -- t[2973] = 1
      "001" when "0101110011110", -- t[2974] = 1
      "001" when "0101110011111", -- t[2975] = 1
      "001" when "0101110100000", -- t[2976] = 1
      "001" when "0101110100001", -- t[2977] = 1
      "001" when "0101110100010", -- t[2978] = 1
      "001" when "0101110100011", -- t[2979] = 1
      "001" when "0101110100100", -- t[2980] = 1
      "001" when "0101110100101", -- t[2981] = 1
      "001" when "0101110100110", -- t[2982] = 1
      "001" when "0101110100111", -- t[2983] = 1
      "001" when "0101110101000", -- t[2984] = 1
      "001" when "0101110101001", -- t[2985] = 1
      "001" when "0101110101010", -- t[2986] = 1
      "001" when "0101110101011", -- t[2987] = 1
      "001" when "0101110101100", -- t[2988] = 1
      "001" when "0101110101101", -- t[2989] = 1
      "001" when "0101110101110", -- t[2990] = 1
      "001" when "0101110101111", -- t[2991] = 1
      "001" when "0101110110000", -- t[2992] = 1
      "001" when "0101110110001", -- t[2993] = 1
      "001" when "0101110110010", -- t[2994] = 1
      "001" when "0101110110011", -- t[2995] = 1
      "001" when "0101110110100", -- t[2996] = 1
      "001" when "0101110110101", -- t[2997] = 1
      "001" when "0101110110110", -- t[2998] = 1
      "001" when "0101110110111", -- t[2999] = 1
      "001" when "0101110111000", -- t[3000] = 1
      "001" when "0101110111001", -- t[3001] = 1
      "001" when "0101110111010", -- t[3002] = 1
      "001" when "0101110111011", -- t[3003] = 1
      "001" when "0101110111100", -- t[3004] = 1
      "001" when "0101110111101", -- t[3005] = 1
      "001" when "0101110111110", -- t[3006] = 1
      "001" when "0101110111111", -- t[3007] = 1
      "001" when "0101111000000", -- t[3008] = 1
      "001" when "0101111000001", -- t[3009] = 1
      "001" when "0101111000010", -- t[3010] = 1
      "001" when "0101111000011", -- t[3011] = 1
      "001" when "0101111000100", -- t[3012] = 1
      "001" when "0101111000101", -- t[3013] = 1
      "001" when "0101111000110", -- t[3014] = 1
      "001" when "0101111000111", -- t[3015] = 1
      "001" when "0101111001000", -- t[3016] = 1
      "001" when "0101111001001", -- t[3017] = 1
      "001" when "0101111001010", -- t[3018] = 1
      "001" when "0101111001011", -- t[3019] = 1
      "001" when "0101111001100", -- t[3020] = 1
      "001" when "0101111001101", -- t[3021] = 1
      "001" when "0101111001110", -- t[3022] = 1
      "001" when "0101111001111", -- t[3023] = 1
      "001" when "0101111010000", -- t[3024] = 1
      "001" when "0101111010001", -- t[3025] = 1
      "001" when "0101111010010", -- t[3026] = 1
      "001" when "0101111010011", -- t[3027] = 1
      "001" when "0101111010100", -- t[3028] = 1
      "001" when "0101111010101", -- t[3029] = 1
      "001" when "0101111010110", -- t[3030] = 1
      "001" when "0101111010111", -- t[3031] = 1
      "001" when "0101111011000", -- t[3032] = 1
      "001" when "0101111011001", -- t[3033] = 1
      "001" when "0101111011010", -- t[3034] = 1
      "001" when "0101111011011", -- t[3035] = 1
      "001" when "0101111011100", -- t[3036] = 1
      "001" when "0101111011101", -- t[3037] = 1
      "001" when "0101111011110", -- t[3038] = 1
      "001" when "0101111011111", -- t[3039] = 1
      "001" when "0101111100000", -- t[3040] = 1
      "001" when "0101111100001", -- t[3041] = 1
      "001" when "0101111100010", -- t[3042] = 1
      "001" when "0101111100011", -- t[3043] = 1
      "001" when "0101111100100", -- t[3044] = 1
      "001" when "0101111100101", -- t[3045] = 1
      "001" when "0101111100110", -- t[3046] = 1
      "001" when "0101111100111", -- t[3047] = 1
      "001" when "0101111101000", -- t[3048] = 1
      "001" when "0101111101001", -- t[3049] = 1
      "001" when "0101111101010", -- t[3050] = 1
      "001" when "0101111101011", -- t[3051] = 1
      "001" when "0101111101100", -- t[3052] = 1
      "001" when "0101111101101", -- t[3053] = 1
      "001" when "0101111101110", -- t[3054] = 1
      "001" when "0101111101111", -- t[3055] = 1
      "001" when "0101111110000", -- t[3056] = 1
      "001" when "0101111110001", -- t[3057] = 1
      "001" when "0101111110010", -- t[3058] = 1
      "001" when "0101111110011", -- t[3059] = 1
      "001" when "0101111110100", -- t[3060] = 1
      "001" when "0101111110101", -- t[3061] = 1
      "001" when "0101111110110", -- t[3062] = 1
      "001" when "0101111110111", -- t[3063] = 1
      "001" when "0101111111000", -- t[3064] = 1
      "001" when "0101111111001", -- t[3065] = 1
      "001" when "0101111111010", -- t[3066] = 1
      "001" when "0101111111011", -- t[3067] = 1
      "001" when "0101111111100", -- t[3068] = 1
      "001" when "0101111111101", -- t[3069] = 1
      "001" when "0101111111110", -- t[3070] = 1
      "001" when "0101111111111", -- t[3071] = 1
      "001" when "0110000000000", -- t[3072] = 1
      "001" when "0110000000001", -- t[3073] = 1
      "001" when "0110000000010", -- t[3074] = 1
      "001" when "0110000000011", -- t[3075] = 1
      "001" when "0110000000100", -- t[3076] = 1
      "001" when "0110000000101", -- t[3077] = 1
      "001" when "0110000000110", -- t[3078] = 1
      "001" when "0110000000111", -- t[3079] = 1
      "001" when "0110000001000", -- t[3080] = 1
      "001" when "0110000001001", -- t[3081] = 1
      "001" when "0110000001010", -- t[3082] = 1
      "001" when "0110000001011", -- t[3083] = 1
      "001" when "0110000001100", -- t[3084] = 1
      "001" when "0110000001101", -- t[3085] = 1
      "001" when "0110000001110", -- t[3086] = 1
      "001" when "0110000001111", -- t[3087] = 1
      "001" when "0110000010000", -- t[3088] = 1
      "001" when "0110000010001", -- t[3089] = 1
      "001" when "0110000010010", -- t[3090] = 1
      "001" when "0110000010011", -- t[3091] = 1
      "001" when "0110000010100", -- t[3092] = 1
      "001" when "0110000010101", -- t[3093] = 1
      "001" when "0110000010110", -- t[3094] = 1
      "001" when "0110000010111", -- t[3095] = 1
      "001" when "0110000011000", -- t[3096] = 1
      "001" when "0110000011001", -- t[3097] = 1
      "001" when "0110000011010", -- t[3098] = 1
      "001" when "0110000011011", -- t[3099] = 1
      "001" when "0110000011100", -- t[3100] = 1
      "001" when "0110000011101", -- t[3101] = 1
      "001" when "0110000011110", -- t[3102] = 1
      "001" when "0110000011111", -- t[3103] = 1
      "001" when "0110000100000", -- t[3104] = 1
      "001" when "0110000100001", -- t[3105] = 1
      "001" when "0110000100010", -- t[3106] = 1
      "001" when "0110000100011", -- t[3107] = 1
      "001" when "0110000100100", -- t[3108] = 1
      "001" when "0110000100101", -- t[3109] = 1
      "001" when "0110000100110", -- t[3110] = 1
      "001" when "0110000100111", -- t[3111] = 1
      "001" when "0110000101000", -- t[3112] = 1
      "001" when "0110000101001", -- t[3113] = 1
      "001" when "0110000101010", -- t[3114] = 1
      "001" when "0110000101011", -- t[3115] = 1
      "001" when "0110000101100", -- t[3116] = 1
      "001" when "0110000101101", -- t[3117] = 1
      "001" when "0110000101110", -- t[3118] = 1
      "001" when "0110000101111", -- t[3119] = 1
      "001" when "0110000110000", -- t[3120] = 1
      "001" when "0110000110001", -- t[3121] = 1
      "001" when "0110000110010", -- t[3122] = 1
      "001" when "0110000110011", -- t[3123] = 1
      "001" when "0110000110100", -- t[3124] = 1
      "001" when "0110000110101", -- t[3125] = 1
      "001" when "0110000110110", -- t[3126] = 1
      "001" when "0110000110111", -- t[3127] = 1
      "001" when "0110000111000", -- t[3128] = 1
      "001" when "0110000111001", -- t[3129] = 1
      "001" when "0110000111010", -- t[3130] = 1
      "001" when "0110000111011", -- t[3131] = 1
      "001" when "0110000111100", -- t[3132] = 1
      "001" when "0110000111101", -- t[3133] = 1
      "001" when "0110000111110", -- t[3134] = 1
      "001" when "0110000111111", -- t[3135] = 1
      "001" when "0110001000000", -- t[3136] = 1
      "001" when "0110001000001", -- t[3137] = 1
      "001" when "0110001000010", -- t[3138] = 1
      "001" when "0110001000011", -- t[3139] = 1
      "001" when "0110001000100", -- t[3140] = 1
      "001" when "0110001000101", -- t[3141] = 1
      "001" when "0110001000110", -- t[3142] = 1
      "001" when "0110001000111", -- t[3143] = 1
      "001" when "0110001001000", -- t[3144] = 1
      "001" when "0110001001001", -- t[3145] = 1
      "001" when "0110001001010", -- t[3146] = 1
      "001" when "0110001001011", -- t[3147] = 1
      "001" when "0110001001100", -- t[3148] = 1
      "001" when "0110001001101", -- t[3149] = 1
      "001" when "0110001001110", -- t[3150] = 1
      "001" when "0110001001111", -- t[3151] = 1
      "001" when "0110001010000", -- t[3152] = 1
      "001" when "0110001010001", -- t[3153] = 1
      "001" when "0110001010010", -- t[3154] = 1
      "001" when "0110001010011", -- t[3155] = 1
      "001" when "0110001010100", -- t[3156] = 1
      "001" when "0110001010101", -- t[3157] = 1
      "001" when "0110001010110", -- t[3158] = 1
      "001" when "0110001010111", -- t[3159] = 1
      "001" when "0110001011000", -- t[3160] = 1
      "001" when "0110001011001", -- t[3161] = 1
      "001" when "0110001011010", -- t[3162] = 1
      "001" when "0110001011011", -- t[3163] = 1
      "001" when "0110001011100", -- t[3164] = 1
      "001" when "0110001011101", -- t[3165] = 1
      "001" when "0110001011110", -- t[3166] = 1
      "001" when "0110001011111", -- t[3167] = 1
      "001" when "0110001100000", -- t[3168] = 1
      "001" when "0110001100001", -- t[3169] = 1
      "001" when "0110001100010", -- t[3170] = 1
      "001" when "0110001100011", -- t[3171] = 1
      "001" when "0110001100100", -- t[3172] = 1
      "001" when "0110001100101", -- t[3173] = 1
      "001" when "0110001100110", -- t[3174] = 1
      "001" when "0110001100111", -- t[3175] = 1
      "001" when "0110001101000", -- t[3176] = 1
      "001" when "0110001101001", -- t[3177] = 1
      "001" when "0110001101010", -- t[3178] = 1
      "001" when "0110001101011", -- t[3179] = 1
      "001" when "0110001101100", -- t[3180] = 1
      "001" when "0110001101101", -- t[3181] = 1
      "001" when "0110001101110", -- t[3182] = 1
      "001" when "0110001101111", -- t[3183] = 1
      "001" when "0110001110000", -- t[3184] = 1
      "001" when "0110001110001", -- t[3185] = 1
      "001" when "0110001110010", -- t[3186] = 1
      "001" when "0110001110011", -- t[3187] = 1
      "001" when "0110001110100", -- t[3188] = 1
      "001" when "0110001110101", -- t[3189] = 1
      "001" when "0110001110110", -- t[3190] = 1
      "001" when "0110001110111", -- t[3191] = 1
      "001" when "0110001111000", -- t[3192] = 1
      "001" when "0110001111001", -- t[3193] = 1
      "001" when "0110001111010", -- t[3194] = 1
      "001" when "0110001111011", -- t[3195] = 1
      "001" when "0110001111100", -- t[3196] = 1
      "001" when "0110001111101", -- t[3197] = 1
      "001" when "0110001111110", -- t[3198] = 1
      "001" when "0110001111111", -- t[3199] = 1
      "001" when "0110010000000", -- t[3200] = 1
      "001" when "0110010000001", -- t[3201] = 1
      "001" when "0110010000010", -- t[3202] = 1
      "001" when "0110010000011", -- t[3203] = 1
      "001" when "0110010000100", -- t[3204] = 1
      "001" when "0110010000101", -- t[3205] = 1
      "001" when "0110010000110", -- t[3206] = 1
      "001" when "0110010000111", -- t[3207] = 1
      "001" when "0110010001000", -- t[3208] = 1
      "001" when "0110010001001", -- t[3209] = 1
      "001" when "0110010001010", -- t[3210] = 1
      "001" when "0110010001011", -- t[3211] = 1
      "001" when "0110010001100", -- t[3212] = 1
      "001" when "0110010001101", -- t[3213] = 1
      "001" when "0110010001110", -- t[3214] = 1
      "001" when "0110010001111", -- t[3215] = 1
      "001" when "0110010010000", -- t[3216] = 1
      "001" when "0110010010001", -- t[3217] = 1
      "001" when "0110010010010", -- t[3218] = 1
      "001" when "0110010010011", -- t[3219] = 1
      "001" when "0110010010100", -- t[3220] = 1
      "001" when "0110010010101", -- t[3221] = 1
      "001" when "0110010010110", -- t[3222] = 1
      "001" when "0110010010111", -- t[3223] = 1
      "001" when "0110010011000", -- t[3224] = 1
      "001" when "0110010011001", -- t[3225] = 1
      "001" when "0110010011010", -- t[3226] = 1
      "001" when "0110010011011", -- t[3227] = 1
      "001" when "0110010011100", -- t[3228] = 1
      "001" when "0110010011101", -- t[3229] = 1
      "001" when "0110010011110", -- t[3230] = 1
      "001" when "0110010011111", -- t[3231] = 1
      "001" when "0110010100000", -- t[3232] = 1
      "001" when "0110010100001", -- t[3233] = 1
      "001" when "0110010100010", -- t[3234] = 1
      "001" when "0110010100011", -- t[3235] = 1
      "001" when "0110010100100", -- t[3236] = 1
      "001" when "0110010100101", -- t[3237] = 1
      "001" when "0110010100110", -- t[3238] = 1
      "001" when "0110010100111", -- t[3239] = 1
      "001" when "0110010101000", -- t[3240] = 1
      "001" when "0110010101001", -- t[3241] = 1
      "001" when "0110010101010", -- t[3242] = 1
      "001" when "0110010101011", -- t[3243] = 1
      "001" when "0110010101100", -- t[3244] = 1
      "001" when "0110010101101", -- t[3245] = 1
      "001" when "0110010101110", -- t[3246] = 1
      "001" when "0110010101111", -- t[3247] = 1
      "001" when "0110010110000", -- t[3248] = 1
      "001" when "0110010110001", -- t[3249] = 1
      "001" when "0110010110010", -- t[3250] = 1
      "001" when "0110010110011", -- t[3251] = 1
      "001" when "0110010110100", -- t[3252] = 1
      "001" when "0110010110101", -- t[3253] = 1
      "001" when "0110010110110", -- t[3254] = 1
      "001" when "0110010110111", -- t[3255] = 1
      "001" when "0110010111000", -- t[3256] = 1
      "001" when "0110010111001", -- t[3257] = 1
      "001" when "0110010111010", -- t[3258] = 1
      "001" when "0110010111011", -- t[3259] = 1
      "001" when "0110010111100", -- t[3260] = 1
      "001" when "0110010111101", -- t[3261] = 1
      "001" when "0110010111110", -- t[3262] = 1
      "001" when "0110010111111", -- t[3263] = 1
      "001" when "0110011000000", -- t[3264] = 1
      "001" when "0110011000001", -- t[3265] = 1
      "001" when "0110011000010", -- t[3266] = 1
      "001" when "0110011000011", -- t[3267] = 1
      "001" when "0110011000100", -- t[3268] = 1
      "001" when "0110011000101", -- t[3269] = 1
      "001" when "0110011000110", -- t[3270] = 1
      "001" when "0110011000111", -- t[3271] = 1
      "001" when "0110011001000", -- t[3272] = 1
      "001" when "0110011001001", -- t[3273] = 1
      "001" when "0110011001010", -- t[3274] = 1
      "001" when "0110011001011", -- t[3275] = 1
      "001" when "0110011001100", -- t[3276] = 1
      "001" when "0110011001101", -- t[3277] = 1
      "001" when "0110011001110", -- t[3278] = 1
      "001" when "0110011001111", -- t[3279] = 1
      "001" when "0110011010000", -- t[3280] = 1
      "001" when "0110011010001", -- t[3281] = 1
      "001" when "0110011010010", -- t[3282] = 1
      "001" when "0110011010011", -- t[3283] = 1
      "001" when "0110011010100", -- t[3284] = 1
      "001" when "0110011010101", -- t[3285] = 1
      "001" when "0110011010110", -- t[3286] = 1
      "001" when "0110011010111", -- t[3287] = 1
      "001" when "0110011011000", -- t[3288] = 1
      "001" when "0110011011001", -- t[3289] = 1
      "001" when "0110011011010", -- t[3290] = 1
      "001" when "0110011011011", -- t[3291] = 1
      "001" when "0110011011100", -- t[3292] = 1
      "001" when "0110011011101", -- t[3293] = 1
      "001" when "0110011011110", -- t[3294] = 1
      "001" when "0110011011111", -- t[3295] = 1
      "001" when "0110011100000", -- t[3296] = 1
      "001" when "0110011100001", -- t[3297] = 1
      "001" when "0110011100010", -- t[3298] = 1
      "001" when "0110011100011", -- t[3299] = 1
      "001" when "0110011100100", -- t[3300] = 1
      "001" when "0110011100101", -- t[3301] = 1
      "001" when "0110011100110", -- t[3302] = 1
      "001" when "0110011100111", -- t[3303] = 1
      "001" when "0110011101000", -- t[3304] = 1
      "001" when "0110011101001", -- t[3305] = 1
      "001" when "0110011101010", -- t[3306] = 1
      "001" when "0110011101011", -- t[3307] = 1
      "001" when "0110011101100", -- t[3308] = 1
      "001" when "0110011101101", -- t[3309] = 1
      "001" when "0110011101110", -- t[3310] = 1
      "001" when "0110011101111", -- t[3311] = 1
      "001" when "0110011110000", -- t[3312] = 1
      "001" when "0110011110001", -- t[3313] = 1
      "001" when "0110011110010", -- t[3314] = 1
      "001" when "0110011110011", -- t[3315] = 1
      "001" when "0110011110100", -- t[3316] = 1
      "001" when "0110011110101", -- t[3317] = 1
      "001" when "0110011110110", -- t[3318] = 1
      "001" when "0110011110111", -- t[3319] = 1
      "001" when "0110011111000", -- t[3320] = 1
      "001" when "0110011111001", -- t[3321] = 1
      "001" when "0110011111010", -- t[3322] = 1
      "001" when "0110011111011", -- t[3323] = 1
      "001" when "0110011111100", -- t[3324] = 1
      "001" when "0110011111101", -- t[3325] = 1
      "001" when "0110011111110", -- t[3326] = 1
      "001" when "0110011111111", -- t[3327] = 1
      "001" when "0110100000000", -- t[3328] = 1
      "001" when "0110100000001", -- t[3329] = 1
      "001" when "0110100000010", -- t[3330] = 1
      "001" when "0110100000011", -- t[3331] = 1
      "001" when "0110100000100", -- t[3332] = 1
      "001" when "0110100000101", -- t[3333] = 1
      "001" when "0110100000110", -- t[3334] = 1
      "001" when "0110100000111", -- t[3335] = 1
      "001" when "0110100001000", -- t[3336] = 1
      "001" when "0110100001001", -- t[3337] = 1
      "001" when "0110100001010", -- t[3338] = 1
      "001" when "0110100001011", -- t[3339] = 1
      "001" when "0110100001100", -- t[3340] = 1
      "001" when "0110100001101", -- t[3341] = 1
      "001" when "0110100001110", -- t[3342] = 1
      "001" when "0110100001111", -- t[3343] = 1
      "001" when "0110100010000", -- t[3344] = 1
      "001" when "0110100010001", -- t[3345] = 1
      "001" when "0110100010010", -- t[3346] = 1
      "001" when "0110100010011", -- t[3347] = 1
      "001" when "0110100010100", -- t[3348] = 1
      "001" when "0110100010101", -- t[3349] = 1
      "001" when "0110100010110", -- t[3350] = 1
      "001" when "0110100010111", -- t[3351] = 1
      "001" when "0110100011000", -- t[3352] = 1
      "001" when "0110100011001", -- t[3353] = 1
      "001" when "0110100011010", -- t[3354] = 1
      "001" when "0110100011011", -- t[3355] = 1
      "001" when "0110100011100", -- t[3356] = 1
      "001" when "0110100011101", -- t[3357] = 1
      "001" when "0110100011110", -- t[3358] = 1
      "001" when "0110100011111", -- t[3359] = 1
      "001" when "0110100100000", -- t[3360] = 1
      "001" when "0110100100001", -- t[3361] = 1
      "001" when "0110100100010", -- t[3362] = 1
      "001" when "0110100100011", -- t[3363] = 1
      "001" when "0110100100100", -- t[3364] = 1
      "001" when "0110100100101", -- t[3365] = 1
      "001" when "0110100100110", -- t[3366] = 1
      "001" when "0110100100111", -- t[3367] = 1
      "001" when "0110100101000", -- t[3368] = 1
      "001" when "0110100101001", -- t[3369] = 1
      "001" when "0110100101010", -- t[3370] = 1
      "001" when "0110100101011", -- t[3371] = 1
      "001" when "0110100101100", -- t[3372] = 1
      "001" when "0110100101101", -- t[3373] = 1
      "001" when "0110100101110", -- t[3374] = 1
      "001" when "0110100101111", -- t[3375] = 1
      "001" when "0110100110000", -- t[3376] = 1
      "001" when "0110100110001", -- t[3377] = 1
      "001" when "0110100110010", -- t[3378] = 1
      "001" when "0110100110011", -- t[3379] = 1
      "001" when "0110100110100", -- t[3380] = 1
      "001" when "0110100110101", -- t[3381] = 1
      "001" when "0110100110110", -- t[3382] = 1
      "001" when "0110100110111", -- t[3383] = 1
      "001" when "0110100111000", -- t[3384] = 1
      "001" when "0110100111001", -- t[3385] = 1
      "001" when "0110100111010", -- t[3386] = 1
      "001" when "0110100111011", -- t[3387] = 1
      "001" when "0110100111100", -- t[3388] = 1
      "001" when "0110100111101", -- t[3389] = 1
      "001" when "0110100111110", -- t[3390] = 1
      "001" when "0110100111111", -- t[3391] = 1
      "001" when "0110101000000", -- t[3392] = 1
      "001" when "0110101000001", -- t[3393] = 1
      "001" when "0110101000010", -- t[3394] = 1
      "001" when "0110101000011", -- t[3395] = 1
      "001" when "0110101000100", -- t[3396] = 1
      "001" when "0110101000101", -- t[3397] = 1
      "001" when "0110101000110", -- t[3398] = 1
      "001" when "0110101000111", -- t[3399] = 1
      "001" when "0110101001000", -- t[3400] = 1
      "001" when "0110101001001", -- t[3401] = 1
      "001" when "0110101001010", -- t[3402] = 1
      "001" when "0110101001011", -- t[3403] = 1
      "001" when "0110101001100", -- t[3404] = 1
      "001" when "0110101001101", -- t[3405] = 1
      "001" when "0110101001110", -- t[3406] = 1
      "001" when "0110101001111", -- t[3407] = 1
      "001" when "0110101010000", -- t[3408] = 1
      "001" when "0110101010001", -- t[3409] = 1
      "001" when "0110101010010", -- t[3410] = 1
      "001" when "0110101010011", -- t[3411] = 1
      "001" when "0110101010100", -- t[3412] = 1
      "001" when "0110101010101", -- t[3413] = 1
      "001" when "0110101010110", -- t[3414] = 1
      "001" when "0110101010111", -- t[3415] = 1
      "001" when "0110101011000", -- t[3416] = 1
      "001" when "0110101011001", -- t[3417] = 1
      "001" when "0110101011010", -- t[3418] = 1
      "001" when "0110101011011", -- t[3419] = 1
      "001" when "0110101011100", -- t[3420] = 1
      "001" when "0110101011101", -- t[3421] = 1
      "001" when "0110101011110", -- t[3422] = 1
      "001" when "0110101011111", -- t[3423] = 1
      "001" when "0110101100000", -- t[3424] = 1
      "001" when "0110101100001", -- t[3425] = 1
      "001" when "0110101100010", -- t[3426] = 1
      "001" when "0110101100011", -- t[3427] = 1
      "001" when "0110101100100", -- t[3428] = 1
      "001" when "0110101100101", -- t[3429] = 1
      "001" when "0110101100110", -- t[3430] = 1
      "001" when "0110101100111", -- t[3431] = 1
      "001" when "0110101101000", -- t[3432] = 1
      "001" when "0110101101001", -- t[3433] = 1
      "001" when "0110101101010", -- t[3434] = 1
      "001" when "0110101101011", -- t[3435] = 1
      "001" when "0110101101100", -- t[3436] = 1
      "001" when "0110101101101", -- t[3437] = 1
      "001" when "0110101101110", -- t[3438] = 1
      "001" when "0110101101111", -- t[3439] = 1
      "001" when "0110101110000", -- t[3440] = 1
      "001" when "0110101110001", -- t[3441] = 1
      "001" when "0110101110010", -- t[3442] = 1
      "001" when "0110101110011", -- t[3443] = 1
      "001" when "0110101110100", -- t[3444] = 1
      "001" when "0110101110101", -- t[3445] = 1
      "001" when "0110101110110", -- t[3446] = 1
      "001" when "0110101110111", -- t[3447] = 1
      "001" when "0110101111000", -- t[3448] = 1
      "001" when "0110101111001", -- t[3449] = 1
      "001" when "0110101111010", -- t[3450] = 1
      "001" when "0110101111011", -- t[3451] = 1
      "001" when "0110101111100", -- t[3452] = 1
      "001" when "0110101111101", -- t[3453] = 1
      "001" when "0110101111110", -- t[3454] = 1
      "001" when "0110101111111", -- t[3455] = 1
      "001" when "0110110000000", -- t[3456] = 1
      "001" when "0110110000001", -- t[3457] = 1
      "001" when "0110110000010", -- t[3458] = 1
      "001" when "0110110000011", -- t[3459] = 1
      "001" when "0110110000100", -- t[3460] = 1
      "001" when "0110110000101", -- t[3461] = 1
      "001" when "0110110000110", -- t[3462] = 1
      "001" when "0110110000111", -- t[3463] = 1
      "001" when "0110110001000", -- t[3464] = 1
      "001" when "0110110001001", -- t[3465] = 1
      "001" when "0110110001010", -- t[3466] = 1
      "001" when "0110110001011", -- t[3467] = 1
      "001" when "0110110001100", -- t[3468] = 1
      "001" when "0110110001101", -- t[3469] = 1
      "001" when "0110110001110", -- t[3470] = 1
      "001" when "0110110001111", -- t[3471] = 1
      "001" when "0110110010000", -- t[3472] = 1
      "001" when "0110110010001", -- t[3473] = 1
      "001" when "0110110010010", -- t[3474] = 1
      "001" when "0110110010011", -- t[3475] = 1
      "001" when "0110110010100", -- t[3476] = 1
      "001" when "0110110010101", -- t[3477] = 1
      "001" when "0110110010110", -- t[3478] = 1
      "001" when "0110110010111", -- t[3479] = 1
      "001" when "0110110011000", -- t[3480] = 1
      "001" when "0110110011001", -- t[3481] = 1
      "001" when "0110110011010", -- t[3482] = 1
      "001" when "0110110011011", -- t[3483] = 1
      "001" when "0110110011100", -- t[3484] = 1
      "001" when "0110110011101", -- t[3485] = 1
      "001" when "0110110011110", -- t[3486] = 1
      "001" when "0110110011111", -- t[3487] = 1
      "001" when "0110110100000", -- t[3488] = 1
      "001" when "0110110100001", -- t[3489] = 1
      "001" when "0110110100010", -- t[3490] = 1
      "001" when "0110110100011", -- t[3491] = 1
      "001" when "0110110100100", -- t[3492] = 1
      "001" when "0110110100101", -- t[3493] = 1
      "001" when "0110110100110", -- t[3494] = 1
      "001" when "0110110100111", -- t[3495] = 1
      "001" when "0110110101000", -- t[3496] = 1
      "001" when "0110110101001", -- t[3497] = 1
      "001" when "0110110101010", -- t[3498] = 1
      "001" when "0110110101011", -- t[3499] = 1
      "001" when "0110110101100", -- t[3500] = 1
      "001" when "0110110101101", -- t[3501] = 1
      "001" when "0110110101110", -- t[3502] = 1
      "001" when "0110110101111", -- t[3503] = 1
      "001" when "0110110110000", -- t[3504] = 1
      "001" when "0110110110001", -- t[3505] = 1
      "001" when "0110110110010", -- t[3506] = 1
      "001" when "0110110110011", -- t[3507] = 1
      "001" when "0110110110100", -- t[3508] = 1
      "001" when "0110110110101", -- t[3509] = 1
      "001" when "0110110110110", -- t[3510] = 1
      "001" when "0110110110111", -- t[3511] = 1
      "001" when "0110110111000", -- t[3512] = 1
      "001" when "0110110111001", -- t[3513] = 1
      "001" when "0110110111010", -- t[3514] = 1
      "001" when "0110110111011", -- t[3515] = 1
      "001" when "0110110111100", -- t[3516] = 1
      "001" when "0110110111101", -- t[3517] = 1
      "001" when "0110110111110", -- t[3518] = 1
      "001" when "0110110111111", -- t[3519] = 1
      "001" when "0110111000000", -- t[3520] = 1
      "001" when "0110111000001", -- t[3521] = 1
      "001" when "0110111000010", -- t[3522] = 1
      "001" when "0110111000011", -- t[3523] = 1
      "001" when "0110111000100", -- t[3524] = 1
      "001" when "0110111000101", -- t[3525] = 1
      "001" when "0110111000110", -- t[3526] = 1
      "001" when "0110111000111", -- t[3527] = 1
      "001" when "0110111001000", -- t[3528] = 1
      "001" when "0110111001001", -- t[3529] = 1
      "001" when "0110111001010", -- t[3530] = 1
      "001" when "0110111001011", -- t[3531] = 1
      "001" when "0110111001100", -- t[3532] = 1
      "001" when "0110111001101", -- t[3533] = 1
      "001" when "0110111001110", -- t[3534] = 1
      "001" when "0110111001111", -- t[3535] = 1
      "001" when "0110111010000", -- t[3536] = 1
      "001" when "0110111010001", -- t[3537] = 1
      "001" when "0110111010010", -- t[3538] = 1
      "001" when "0110111010011", -- t[3539] = 1
      "001" when "0110111010100", -- t[3540] = 1
      "001" when "0110111010101", -- t[3541] = 1
      "001" when "0110111010110", -- t[3542] = 1
      "001" when "0110111010111", -- t[3543] = 1
      "001" when "0110111011000", -- t[3544] = 1
      "001" when "0110111011001", -- t[3545] = 1
      "001" when "0110111011010", -- t[3546] = 1
      "001" when "0110111011011", -- t[3547] = 1
      "001" when "0110111011100", -- t[3548] = 1
      "001" when "0110111011101", -- t[3549] = 1
      "001" when "0110111011110", -- t[3550] = 1
      "001" when "0110111011111", -- t[3551] = 1
      "001" when "0110111100000", -- t[3552] = 1
      "001" when "0110111100001", -- t[3553] = 1
      "001" when "0110111100010", -- t[3554] = 1
      "001" when "0110111100011", -- t[3555] = 1
      "001" when "0110111100100", -- t[3556] = 1
      "001" when "0110111100101", -- t[3557] = 1
      "001" when "0110111100110", -- t[3558] = 1
      "001" when "0110111100111", -- t[3559] = 1
      "001" when "0110111101000", -- t[3560] = 1
      "001" when "0110111101001", -- t[3561] = 1
      "001" when "0110111101010", -- t[3562] = 1
      "001" when "0110111101011", -- t[3563] = 1
      "001" when "0110111101100", -- t[3564] = 1
      "001" when "0110111101101", -- t[3565] = 1
      "001" when "0110111101110", -- t[3566] = 1
      "001" when "0110111101111", -- t[3567] = 1
      "001" when "0110111110000", -- t[3568] = 1
      "001" when "0110111110001", -- t[3569] = 1
      "001" when "0110111110010", -- t[3570] = 1
      "001" when "0110111110011", -- t[3571] = 1
      "001" when "0110111110100", -- t[3572] = 1
      "001" when "0110111110101", -- t[3573] = 1
      "001" when "0110111110110", -- t[3574] = 1
      "001" when "0110111110111", -- t[3575] = 1
      "001" when "0110111111000", -- t[3576] = 1
      "001" when "0110111111001", -- t[3577] = 1
      "001" when "0110111111010", -- t[3578] = 1
      "001" when "0110111111011", -- t[3579] = 1
      "001" when "0110111111100", -- t[3580] = 1
      "001" when "0110111111101", -- t[3581] = 1
      "001" when "0110111111110", -- t[3582] = 1
      "001" when "0110111111111", -- t[3583] = 1
      "001" when "0111000000000", -- t[3584] = 1
      "001" when "0111000000001", -- t[3585] = 1
      "001" when "0111000000010", -- t[3586] = 1
      "001" when "0111000000011", -- t[3587] = 1
      "001" when "0111000000100", -- t[3588] = 1
      "001" when "0111000000101", -- t[3589] = 1
      "001" when "0111000000110", -- t[3590] = 1
      "001" when "0111000000111", -- t[3591] = 1
      "001" when "0111000001000", -- t[3592] = 1
      "001" when "0111000001001", -- t[3593] = 1
      "001" when "0111000001010", -- t[3594] = 1
      "001" when "0111000001011", -- t[3595] = 1
      "001" when "0111000001100", -- t[3596] = 1
      "001" when "0111000001101", -- t[3597] = 1
      "001" when "0111000001110", -- t[3598] = 1
      "001" when "0111000001111", -- t[3599] = 1
      "001" when "0111000010000", -- t[3600] = 1
      "001" when "0111000010001", -- t[3601] = 1
      "001" when "0111000010010", -- t[3602] = 1
      "001" when "0111000010011", -- t[3603] = 1
      "001" when "0111000010100", -- t[3604] = 1
      "001" when "0111000010101", -- t[3605] = 1
      "001" when "0111000010110", -- t[3606] = 1
      "001" when "0111000010111", -- t[3607] = 1
      "001" when "0111000011000", -- t[3608] = 1
      "001" when "0111000011001", -- t[3609] = 1
      "001" when "0111000011010", -- t[3610] = 1
      "001" when "0111000011011", -- t[3611] = 1
      "001" when "0111000011100", -- t[3612] = 1
      "001" when "0111000011101", -- t[3613] = 1
      "010" when "0111000011110", -- t[3614] = 2
      "010" when "0111000011111", -- t[3615] = 2
      "010" when "0111000100000", -- t[3616] = 2
      "010" when "0111000100001", -- t[3617] = 2
      "010" when "0111000100010", -- t[3618] = 2
      "010" when "0111000100011", -- t[3619] = 2
      "010" when "0111000100100", -- t[3620] = 2
      "010" when "0111000100101", -- t[3621] = 2
      "010" when "0111000100110", -- t[3622] = 2
      "010" when "0111000100111", -- t[3623] = 2
      "010" when "0111000101000", -- t[3624] = 2
      "010" when "0111000101001", -- t[3625] = 2
      "010" when "0111000101010", -- t[3626] = 2
      "010" when "0111000101011", -- t[3627] = 2
      "010" when "0111000101100", -- t[3628] = 2
      "010" when "0111000101101", -- t[3629] = 2
      "010" when "0111000101110", -- t[3630] = 2
      "010" when "0111000101111", -- t[3631] = 2
      "010" when "0111000110000", -- t[3632] = 2
      "010" when "0111000110001", -- t[3633] = 2
      "010" when "0111000110010", -- t[3634] = 2
      "010" when "0111000110011", -- t[3635] = 2
      "010" when "0111000110100", -- t[3636] = 2
      "010" when "0111000110101", -- t[3637] = 2
      "010" when "0111000110110", -- t[3638] = 2
      "010" when "0111000110111", -- t[3639] = 2
      "010" when "0111000111000", -- t[3640] = 2
      "010" when "0111000111001", -- t[3641] = 2
      "010" when "0111000111010", -- t[3642] = 2
      "010" when "0111000111011", -- t[3643] = 2
      "010" when "0111000111100", -- t[3644] = 2
      "010" when "0111000111101", -- t[3645] = 2
      "010" when "0111000111110", -- t[3646] = 2
      "010" when "0111000111111", -- t[3647] = 2
      "010" when "0111001000000", -- t[3648] = 2
      "010" when "0111001000001", -- t[3649] = 2
      "010" when "0111001000010", -- t[3650] = 2
      "010" when "0111001000011", -- t[3651] = 2
      "010" when "0111001000100", -- t[3652] = 2
      "010" when "0111001000101", -- t[3653] = 2
      "010" when "0111001000110", -- t[3654] = 2
      "010" when "0111001000111", -- t[3655] = 2
      "010" when "0111001001000", -- t[3656] = 2
      "010" when "0111001001001", -- t[3657] = 2
      "010" when "0111001001010", -- t[3658] = 2
      "010" when "0111001001011", -- t[3659] = 2
      "010" when "0111001001100", -- t[3660] = 2
      "010" when "0111001001101", -- t[3661] = 2
      "010" when "0111001001110", -- t[3662] = 2
      "010" when "0111001001111", -- t[3663] = 2
      "010" when "0111001010000", -- t[3664] = 2
      "010" when "0111001010001", -- t[3665] = 2
      "010" when "0111001010010", -- t[3666] = 2
      "010" when "0111001010011", -- t[3667] = 2
      "010" when "0111001010100", -- t[3668] = 2
      "010" when "0111001010101", -- t[3669] = 2
      "010" when "0111001010110", -- t[3670] = 2
      "010" when "0111001010111", -- t[3671] = 2
      "010" when "0111001011000", -- t[3672] = 2
      "010" when "0111001011001", -- t[3673] = 2
      "010" when "0111001011010", -- t[3674] = 2
      "010" when "0111001011011", -- t[3675] = 2
      "010" when "0111001011100", -- t[3676] = 2
      "010" when "0111001011101", -- t[3677] = 2
      "010" when "0111001011110", -- t[3678] = 2
      "010" when "0111001011111", -- t[3679] = 2
      "010" when "0111001100000", -- t[3680] = 2
      "010" when "0111001100001", -- t[3681] = 2
      "010" when "0111001100010", -- t[3682] = 2
      "010" when "0111001100011", -- t[3683] = 2
      "010" when "0111001100100", -- t[3684] = 2
      "010" when "0111001100101", -- t[3685] = 2
      "010" when "0111001100110", -- t[3686] = 2
      "010" when "0111001100111", -- t[3687] = 2
      "010" when "0111001101000", -- t[3688] = 2
      "010" when "0111001101001", -- t[3689] = 2
      "010" when "0111001101010", -- t[3690] = 2
      "010" when "0111001101011", -- t[3691] = 2
      "010" when "0111001101100", -- t[3692] = 2
      "010" when "0111001101101", -- t[3693] = 2
      "010" when "0111001101110", -- t[3694] = 2
      "010" when "0111001101111", -- t[3695] = 2
      "010" when "0111001110000", -- t[3696] = 2
      "010" when "0111001110001", -- t[3697] = 2
      "010" when "0111001110010", -- t[3698] = 2
      "010" when "0111001110011", -- t[3699] = 2
      "010" when "0111001110100", -- t[3700] = 2
      "010" when "0111001110101", -- t[3701] = 2
      "010" when "0111001110110", -- t[3702] = 2
      "010" when "0111001110111", -- t[3703] = 2
      "010" when "0111001111000", -- t[3704] = 2
      "010" when "0111001111001", -- t[3705] = 2
      "010" when "0111001111010", -- t[3706] = 2
      "010" when "0111001111011", -- t[3707] = 2
      "010" when "0111001111100", -- t[3708] = 2
      "010" when "0111001111101", -- t[3709] = 2
      "010" when "0111001111110", -- t[3710] = 2
      "010" when "0111001111111", -- t[3711] = 2
      "010" when "0111010000000", -- t[3712] = 2
      "010" when "0111010000001", -- t[3713] = 2
      "010" when "0111010000010", -- t[3714] = 2
      "010" when "0111010000011", -- t[3715] = 2
      "010" when "0111010000100", -- t[3716] = 2
      "010" when "0111010000101", -- t[3717] = 2
      "010" when "0111010000110", -- t[3718] = 2
      "010" when "0111010000111", -- t[3719] = 2
      "010" when "0111010001000", -- t[3720] = 2
      "010" when "0111010001001", -- t[3721] = 2
      "010" when "0111010001010", -- t[3722] = 2
      "010" when "0111010001011", -- t[3723] = 2
      "010" when "0111010001100", -- t[3724] = 2
      "010" when "0111010001101", -- t[3725] = 2
      "010" when "0111010001110", -- t[3726] = 2
      "010" when "0111010001111", -- t[3727] = 2
      "010" when "0111010010000", -- t[3728] = 2
      "010" when "0111010010001", -- t[3729] = 2
      "010" when "0111010010010", -- t[3730] = 2
      "010" when "0111010010011", -- t[3731] = 2
      "010" when "0111010010100", -- t[3732] = 2
      "010" when "0111010010101", -- t[3733] = 2
      "010" when "0111010010110", -- t[3734] = 2
      "010" when "0111010010111", -- t[3735] = 2
      "010" when "0111010011000", -- t[3736] = 2
      "010" when "0111010011001", -- t[3737] = 2
      "010" when "0111010011010", -- t[3738] = 2
      "010" when "0111010011011", -- t[3739] = 2
      "010" when "0111010011100", -- t[3740] = 2
      "010" when "0111010011101", -- t[3741] = 2
      "010" when "0111010011110", -- t[3742] = 2
      "010" when "0111010011111", -- t[3743] = 2
      "010" when "0111010100000", -- t[3744] = 2
      "010" when "0111010100001", -- t[3745] = 2
      "010" when "0111010100010", -- t[3746] = 2
      "010" when "0111010100011", -- t[3747] = 2
      "010" when "0111010100100", -- t[3748] = 2
      "010" when "0111010100101", -- t[3749] = 2
      "010" when "0111010100110", -- t[3750] = 2
      "010" when "0111010100111", -- t[3751] = 2
      "010" when "0111010101000", -- t[3752] = 2
      "010" when "0111010101001", -- t[3753] = 2
      "010" when "0111010101010", -- t[3754] = 2
      "010" when "0111010101011", -- t[3755] = 2
      "010" when "0111010101100", -- t[3756] = 2
      "010" when "0111010101101", -- t[3757] = 2
      "010" when "0111010101110", -- t[3758] = 2
      "010" when "0111010101111", -- t[3759] = 2
      "010" when "0111010110000", -- t[3760] = 2
      "010" when "0111010110001", -- t[3761] = 2
      "010" when "0111010110010", -- t[3762] = 2
      "010" when "0111010110011", -- t[3763] = 2
      "010" when "0111010110100", -- t[3764] = 2
      "010" when "0111010110101", -- t[3765] = 2
      "010" when "0111010110110", -- t[3766] = 2
      "010" when "0111010110111", -- t[3767] = 2
      "010" when "0111010111000", -- t[3768] = 2
      "010" when "0111010111001", -- t[3769] = 2
      "010" when "0111010111010", -- t[3770] = 2
      "010" when "0111010111011", -- t[3771] = 2
      "010" when "0111010111100", -- t[3772] = 2
      "010" when "0111010111101", -- t[3773] = 2
      "010" when "0111010111110", -- t[3774] = 2
      "010" when "0111010111111", -- t[3775] = 2
      "010" when "0111011000000", -- t[3776] = 2
      "010" when "0111011000001", -- t[3777] = 2
      "010" when "0111011000010", -- t[3778] = 2
      "010" when "0111011000011", -- t[3779] = 2
      "010" when "0111011000100", -- t[3780] = 2
      "010" when "0111011000101", -- t[3781] = 2
      "010" when "0111011000110", -- t[3782] = 2
      "010" when "0111011000111", -- t[3783] = 2
      "010" when "0111011001000", -- t[3784] = 2
      "010" when "0111011001001", -- t[3785] = 2
      "010" when "0111011001010", -- t[3786] = 2
      "010" when "0111011001011", -- t[3787] = 2
      "010" when "0111011001100", -- t[3788] = 2
      "010" when "0111011001101", -- t[3789] = 2
      "010" when "0111011001110", -- t[3790] = 2
      "010" when "0111011001111", -- t[3791] = 2
      "010" when "0111011010000", -- t[3792] = 2
      "010" when "0111011010001", -- t[3793] = 2
      "010" when "0111011010010", -- t[3794] = 2
      "010" when "0111011010011", -- t[3795] = 2
      "010" when "0111011010100", -- t[3796] = 2
      "010" when "0111011010101", -- t[3797] = 2
      "010" when "0111011010110", -- t[3798] = 2
      "010" when "0111011010111", -- t[3799] = 2
      "010" when "0111011011000", -- t[3800] = 2
      "010" when "0111011011001", -- t[3801] = 2
      "010" when "0111011011010", -- t[3802] = 2
      "010" when "0111011011011", -- t[3803] = 2
      "010" when "0111011011100", -- t[3804] = 2
      "010" when "0111011011101", -- t[3805] = 2
      "010" when "0111011011110", -- t[3806] = 2
      "010" when "0111011011111", -- t[3807] = 2
      "010" when "0111011100000", -- t[3808] = 2
      "010" when "0111011100001", -- t[3809] = 2
      "010" when "0111011100010", -- t[3810] = 2
      "010" when "0111011100011", -- t[3811] = 2
      "010" when "0111011100100", -- t[3812] = 2
      "010" when "0111011100101", -- t[3813] = 2
      "010" when "0111011100110", -- t[3814] = 2
      "010" when "0111011100111", -- t[3815] = 2
      "010" when "0111011101000", -- t[3816] = 2
      "010" when "0111011101001", -- t[3817] = 2
      "010" when "0111011101010", -- t[3818] = 2
      "010" when "0111011101011", -- t[3819] = 2
      "010" when "0111011101100", -- t[3820] = 2
      "010" when "0111011101101", -- t[3821] = 2
      "010" when "0111011101110", -- t[3822] = 2
      "010" when "0111011101111", -- t[3823] = 2
      "010" when "0111011110000", -- t[3824] = 2
      "010" when "0111011110001", -- t[3825] = 2
      "010" when "0111011110010", -- t[3826] = 2
      "010" when "0111011110011", -- t[3827] = 2
      "010" when "0111011110100", -- t[3828] = 2
      "010" when "0111011110101", -- t[3829] = 2
      "010" when "0111011110110", -- t[3830] = 2
      "010" when "0111011110111", -- t[3831] = 2
      "010" when "0111011111000", -- t[3832] = 2
      "010" when "0111011111001", -- t[3833] = 2
      "010" when "0111011111010", -- t[3834] = 2
      "010" when "0111011111011", -- t[3835] = 2
      "010" when "0111011111100", -- t[3836] = 2
      "010" when "0111011111101", -- t[3837] = 2
      "010" when "0111011111110", -- t[3838] = 2
      "010" when "0111011111111", -- t[3839] = 2
      "010" when "0111100000000", -- t[3840] = 2
      "010" when "0111100000001", -- t[3841] = 2
      "010" when "0111100000010", -- t[3842] = 2
      "010" when "0111100000011", -- t[3843] = 2
      "010" when "0111100000100", -- t[3844] = 2
      "010" when "0111100000101", -- t[3845] = 2
      "010" when "0111100000110", -- t[3846] = 2
      "010" when "0111100000111", -- t[3847] = 2
      "010" when "0111100001000", -- t[3848] = 2
      "010" when "0111100001001", -- t[3849] = 2
      "010" when "0111100001010", -- t[3850] = 2
      "010" when "0111100001011", -- t[3851] = 2
      "010" when "0111100001100", -- t[3852] = 2
      "010" when "0111100001101", -- t[3853] = 2
      "010" when "0111100001110", -- t[3854] = 2
      "010" when "0111100001111", -- t[3855] = 2
      "010" when "0111100010000", -- t[3856] = 2
      "010" when "0111100010001", -- t[3857] = 2
      "010" when "0111100010010", -- t[3858] = 2
      "010" when "0111100010011", -- t[3859] = 2
      "010" when "0111100010100", -- t[3860] = 2
      "010" when "0111100010101", -- t[3861] = 2
      "010" when "0111100010110", -- t[3862] = 2
      "010" when "0111100010111", -- t[3863] = 2
      "010" when "0111100011000", -- t[3864] = 2
      "010" when "0111100011001", -- t[3865] = 2
      "010" when "0111100011010", -- t[3866] = 2
      "010" when "0111100011011", -- t[3867] = 2
      "010" when "0111100011100", -- t[3868] = 2
      "010" when "0111100011101", -- t[3869] = 2
      "010" when "0111100011110", -- t[3870] = 2
      "010" when "0111100011111", -- t[3871] = 2
      "010" when "0111100100000", -- t[3872] = 2
      "010" when "0111100100001", -- t[3873] = 2
      "010" when "0111100100010", -- t[3874] = 2
      "010" when "0111100100011", -- t[3875] = 2
      "010" when "0111100100100", -- t[3876] = 2
      "010" when "0111100100101", -- t[3877] = 2
      "010" when "0111100100110", -- t[3878] = 2
      "010" when "0111100100111", -- t[3879] = 2
      "010" when "0111100101000", -- t[3880] = 2
      "010" when "0111100101001", -- t[3881] = 2
      "010" when "0111100101010", -- t[3882] = 2
      "010" when "0111100101011", -- t[3883] = 2
      "010" when "0111100101100", -- t[3884] = 2
      "010" when "0111100101101", -- t[3885] = 2
      "010" when "0111100101110", -- t[3886] = 2
      "010" when "0111100101111", -- t[3887] = 2
      "010" when "0111100110000", -- t[3888] = 2
      "010" when "0111100110001", -- t[3889] = 2
      "010" when "0111100110010", -- t[3890] = 2
      "010" when "0111100110011", -- t[3891] = 2
      "010" when "0111100110100", -- t[3892] = 2
      "010" when "0111100110101", -- t[3893] = 2
      "010" when "0111100110110", -- t[3894] = 2
      "010" when "0111100110111", -- t[3895] = 2
      "010" when "0111100111000", -- t[3896] = 2
      "010" when "0111100111001", -- t[3897] = 2
      "010" when "0111100111010", -- t[3898] = 2
      "010" when "0111100111011", -- t[3899] = 2
      "010" when "0111100111100", -- t[3900] = 2
      "010" when "0111100111101", -- t[3901] = 2
      "010" when "0111100111110", -- t[3902] = 2
      "010" when "0111100111111", -- t[3903] = 2
      "010" when "0111101000000", -- t[3904] = 2
      "010" when "0111101000001", -- t[3905] = 2
      "010" when "0111101000010", -- t[3906] = 2
      "010" when "0111101000011", -- t[3907] = 2
      "010" when "0111101000100", -- t[3908] = 2
      "010" when "0111101000101", -- t[3909] = 2
      "010" when "0111101000110", -- t[3910] = 2
      "010" when "0111101000111", -- t[3911] = 2
      "010" when "0111101001000", -- t[3912] = 2
      "010" when "0111101001001", -- t[3913] = 2
      "010" when "0111101001010", -- t[3914] = 2
      "010" when "0111101001011", -- t[3915] = 2
      "010" when "0111101001100", -- t[3916] = 2
      "010" when "0111101001101", -- t[3917] = 2
      "010" when "0111101001110", -- t[3918] = 2
      "010" when "0111101001111", -- t[3919] = 2
      "010" when "0111101010000", -- t[3920] = 2
      "010" when "0111101010001", -- t[3921] = 2
      "010" when "0111101010010", -- t[3922] = 2
      "010" when "0111101010011", -- t[3923] = 2
      "010" when "0111101010100", -- t[3924] = 2
      "010" when "0111101010101", -- t[3925] = 2
      "010" when "0111101010110", -- t[3926] = 2
      "010" when "0111101010111", -- t[3927] = 2
      "010" when "0111101011000", -- t[3928] = 2
      "010" when "0111101011001", -- t[3929] = 2
      "010" when "0111101011010", -- t[3930] = 2
      "010" when "0111101011011", -- t[3931] = 2
      "010" when "0111101011100", -- t[3932] = 2
      "010" when "0111101011101", -- t[3933] = 2
      "010" when "0111101011110", -- t[3934] = 2
      "010" when "0111101011111", -- t[3935] = 2
      "010" when "0111101100000", -- t[3936] = 2
      "010" when "0111101100001", -- t[3937] = 2
      "010" when "0111101100010", -- t[3938] = 2
      "010" when "0111101100011", -- t[3939] = 2
      "010" when "0111101100100", -- t[3940] = 2
      "010" when "0111101100101", -- t[3941] = 2
      "010" when "0111101100110", -- t[3942] = 2
      "010" when "0111101100111", -- t[3943] = 2
      "010" when "0111101101000", -- t[3944] = 2
      "010" when "0111101101001", -- t[3945] = 2
      "010" when "0111101101010", -- t[3946] = 2
      "010" when "0111101101011", -- t[3947] = 2
      "010" when "0111101101100", -- t[3948] = 2
      "010" when "0111101101101", -- t[3949] = 2
      "010" when "0111101101110", -- t[3950] = 2
      "010" when "0111101101111", -- t[3951] = 2
      "010" when "0111101110000", -- t[3952] = 2
      "010" when "0111101110001", -- t[3953] = 2
      "010" when "0111101110010", -- t[3954] = 2
      "010" when "0111101110011", -- t[3955] = 2
      "010" when "0111101110100", -- t[3956] = 2
      "010" when "0111101110101", -- t[3957] = 2
      "010" when "0111101110110", -- t[3958] = 2
      "010" when "0111101110111", -- t[3959] = 2
      "010" when "0111101111000", -- t[3960] = 2
      "010" when "0111101111001", -- t[3961] = 2
      "010" when "0111101111010", -- t[3962] = 2
      "010" when "0111101111011", -- t[3963] = 2
      "010" when "0111101111100", -- t[3964] = 2
      "010" when "0111101111101", -- t[3965] = 2
      "010" when "0111101111110", -- t[3966] = 2
      "010" when "0111101111111", -- t[3967] = 2
      "010" when "0111110000000", -- t[3968] = 2
      "010" when "0111110000001", -- t[3969] = 2
      "010" when "0111110000010", -- t[3970] = 2
      "010" when "0111110000011", -- t[3971] = 2
      "010" when "0111110000100", -- t[3972] = 2
      "010" when "0111110000101", -- t[3973] = 2
      "010" when "0111110000110", -- t[3974] = 2
      "010" when "0111110000111", -- t[3975] = 2
      "010" when "0111110001000", -- t[3976] = 2
      "010" when "0111110001001", -- t[3977] = 2
      "010" when "0111110001010", -- t[3978] = 2
      "010" when "0111110001011", -- t[3979] = 2
      "010" when "0111110001100", -- t[3980] = 2
      "010" when "0111110001101", -- t[3981] = 2
      "010" when "0111110001110", -- t[3982] = 2
      "010" when "0111110001111", -- t[3983] = 2
      "010" when "0111110010000", -- t[3984] = 2
      "010" when "0111110010001", -- t[3985] = 2
      "010" when "0111110010010", -- t[3986] = 2
      "010" when "0111110010011", -- t[3987] = 2
      "010" when "0111110010100", -- t[3988] = 2
      "010" when "0111110010101", -- t[3989] = 2
      "010" when "0111110010110", -- t[3990] = 2
      "010" when "0111110010111", -- t[3991] = 2
      "011" when "0111110011000", -- t[3992] = 3
      "011" when "0111110011001", -- t[3993] = 3
      "011" when "0111110011010", -- t[3994] = 3
      "011" when "0111110011011", -- t[3995] = 3
      "011" when "0111110011100", -- t[3996] = 3
      "011" when "0111110011101", -- t[3997] = 3
      "011" when "0111110011110", -- t[3998] = 3
      "011" when "0111110011111", -- t[3999] = 3
      "011" when "0111110100000", -- t[4000] = 3
      "011" when "0111110100001", -- t[4001] = 3
      "011" when "0111110100010", -- t[4002] = 3
      "011" when "0111110100011", -- t[4003] = 3
      "011" when "0111110100100", -- t[4004] = 3
      "011" when "0111110100101", -- t[4005] = 3
      "011" when "0111110100110", -- t[4006] = 3
      "011" when "0111110100111", -- t[4007] = 3
      "011" when "0111110101000", -- t[4008] = 3
      "011" when "0111110101001", -- t[4009] = 3
      "011" when "0111110101010", -- t[4010] = 3
      "011" when "0111110101011", -- t[4011] = 3
      "011" when "0111110101100", -- t[4012] = 3
      "011" when "0111110101101", -- t[4013] = 3
      "011" when "0111110101110", -- t[4014] = 3
      "011" when "0111110101111", -- t[4015] = 3
      "011" when "0111110110000", -- t[4016] = 3
      "011" when "0111110110001", -- t[4017] = 3
      "011" when "0111110110010", -- t[4018] = 3
      "011" when "0111110110011", -- t[4019] = 3
      "011" when "0111110110100", -- t[4020] = 3
      "011" when "0111110110101", -- t[4021] = 3
      "011" when "0111110110110", -- t[4022] = 3
      "011" when "0111110110111", -- t[4023] = 3
      "011" when "0111110111000", -- t[4024] = 3
      "011" when "0111110111001", -- t[4025] = 3
      "011" when "0111110111010", -- t[4026] = 3
      "011" when "0111110111011", -- t[4027] = 3
      "011" when "0111110111100", -- t[4028] = 3
      "011" when "0111110111101", -- t[4029] = 3
      "011" when "0111110111110", -- t[4030] = 3
      "011" when "0111110111111", -- t[4031] = 3
      "011" when "0111111000000", -- t[4032] = 3
      "011" when "0111111000001", -- t[4033] = 3
      "011" when "0111111000010", -- t[4034] = 3
      "011" when "0111111000011", -- t[4035] = 3
      "011" when "0111111000100", -- t[4036] = 3
      "011" when "0111111000101", -- t[4037] = 3
      "011" when "0111111000110", -- t[4038] = 3
      "011" when "0111111000111", -- t[4039] = 3
      "011" when "0111111001000", -- t[4040] = 3
      "011" when "0111111001001", -- t[4041] = 3
      "011" when "0111111001010", -- t[4042] = 3
      "011" when "0111111001011", -- t[4043] = 3
      "011" when "0111111001100", -- t[4044] = 3
      "011" when "0111111001101", -- t[4045] = 3
      "011" when "0111111001110", -- t[4046] = 3
      "011" when "0111111001111", -- t[4047] = 3
      "011" when "0111111010000", -- t[4048] = 3
      "011" when "0111111010001", -- t[4049] = 3
      "011" when "0111111010010", -- t[4050] = 3
      "011" when "0111111010011", -- t[4051] = 3
      "011" when "0111111010100", -- t[4052] = 3
      "011" when "0111111010101", -- t[4053] = 3
      "011" when "0111111010110", -- t[4054] = 3
      "011" when "0111111010111", -- t[4055] = 3
      "011" when "0111111011000", -- t[4056] = 3
      "011" when "0111111011001", -- t[4057] = 3
      "011" when "0111111011010", -- t[4058] = 3
      "011" when "0111111011011", -- t[4059] = 3
      "011" when "0111111011100", -- t[4060] = 3
      "011" when "0111111011101", -- t[4061] = 3
      "011" when "0111111011110", -- t[4062] = 3
      "011" when "0111111011111", -- t[4063] = 3
      "011" when "0111111100000", -- t[4064] = 3
      "011" when "0111111100001", -- t[4065] = 3
      "011" when "0111111100010", -- t[4066] = 3
      "011" when "0111111100011", -- t[4067] = 3
      "011" when "0111111100100", -- t[4068] = 3
      "011" when "0111111100101", -- t[4069] = 3
      "011" when "0111111100110", -- t[4070] = 3
      "011" when "0111111100111", -- t[4071] = 3
      "011" when "0111111101000", -- t[4072] = 3
      "011" when "0111111101001", -- t[4073] = 3
      "011" when "0111111101010", -- t[4074] = 3
      "011" when "0111111101011", -- t[4075] = 3
      "011" when "0111111101100", -- t[4076] = 3
      "011" when "0111111101101", -- t[4077] = 3
      "011" when "0111111101110", -- t[4078] = 3
      "011" when "0111111101111", -- t[4079] = 3
      "011" when "0111111110000", -- t[4080] = 3
      "011" when "0111111110001", -- t[4081] = 3
      "011" when "0111111110010", -- t[4082] = 3
      "011" when "0111111110011", -- t[4083] = 3
      "011" when "0111111110100", -- t[4084] = 3
      "011" when "0111111110101", -- t[4085] = 3
      "011" when "0111111110110", -- t[4086] = 3
      "011" when "0111111110111", -- t[4087] = 3
      "011" when "0111111111000", -- t[4088] = 3
      "011" when "0111111111001", -- t[4089] = 3
      "011" when "0111111111010", -- t[4090] = 3
      "011" when "0111111111011", -- t[4091] = 3
      "011" when "0111111111100", -- t[4092] = 3
      "011" when "0111111111101", -- t[4093] = 3
      "011" when "0111111111110", -- t[4094] = 3
      "011" when "0111111111111", -- t[4095] = 3
      "---" when others;
end architecture;


-- MultiPartite: LNS addition function: [-8.0 0.0[ -> [0.0 2.0[
-- wI = 12 bits
-- wO = 10 bits
-- Decomposition: 7, 5 / 6, 4 / 2, 3
-- Guard bits: 2
-- Size: 2368 = 12.2^7 + 5.2^7 + 3.2^6

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSAdd_MPT_T2_9 is
  component LNSAdd_MPT_T2_9_tiv is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9_to1 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9_to0 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9_to1_xor is
    port( a : in  std_logic_vector(5 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSAdd_MPT_T2_9_to0_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_9_tiv is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9_tiv is
begin
  with x select
    r <=
      "000000001110" when "0000000", -- t[0] = 14
      "000000001111" when "0000001", -- t[1] = 15
      "000000001111" when "0000010", -- t[2] = 15
      "000000010000" when "0000011", -- t[3] = 16
      "000000010000" when "0000100", -- t[4] = 16
      "000000010001" when "0000101", -- t[5] = 17
      "000000010010" when "0000110", -- t[6] = 18
      "000000010010" when "0000111", -- t[7] = 18
      "000000010011" when "0001000", -- t[8] = 19
      "000000010100" when "0001001", -- t[9] = 20
      "000000010101" when "0001010", -- t[10] = 21
      "000000010101" when "0001011", -- t[11] = 21
      "000000010110" when "0001100", -- t[12] = 22
      "000000010111" when "0001101", -- t[13] = 23
      "000000011000" when "0001110", -- t[14] = 24
      "000000011001" when "0001111", -- t[15] = 25
      "000000011010" when "0010000", -- t[16] = 26
      "000000011011" when "0010001", -- t[17] = 27
      "000000011100" when "0010010", -- t[18] = 28
      "000000011101" when "0010011", -- t[19] = 29
      "000000011110" when "0010100", -- t[20] = 30
      "000000100000" when "0010101", -- t[21] = 32
      "000000100001" when "0010110", -- t[22] = 33
      "000000100010" when "0010111", -- t[23] = 34
      "000000100100" when "0011000", -- t[24] = 36
      "000000100101" when "0011001", -- t[25] = 37
      "000000100111" when "0011010", -- t[26] = 39
      "000000101000" when "0011011", -- t[27] = 40
      "000000101010" when "0011100", -- t[28] = 42
      "000000101100" when "0011101", -- t[29] = 44
      "000000101101" when "0011110", -- t[30] = 45
      "000000101111" when "0011111", -- t[31] = 47
      "000000110001" when "0100000", -- t[32] = 49
      "000000110011" when "0100001", -- t[33] = 51
      "000000110101" when "0100010", -- t[34] = 53
      "000000111000" when "0100011", -- t[35] = 56
      "000000111010" when "0100100", -- t[36] = 58
      "000000111100" when "0100101", -- t[37] = 60
      "000000111111" when "0100110", -- t[38] = 63
      "000001000010" when "0100111", -- t[39] = 66
      "000001000100" when "0101000", -- t[40] = 68
      "000001000111" when "0101001", -- t[41] = 71
      "000001001010" when "0101010", -- t[42] = 74
      "000001001101" when "0101011", -- t[43] = 77
      "000001010001" when "0101100", -- t[44] = 81
      "000001010100" when "0101101", -- t[45] = 84
      "000001011000" when "0101110", -- t[46] = 88
      "000001011011" when "0101111", -- t[47] = 91
      "000001011111" when "0110000", -- t[48] = 95
      "000001100011" when "0110001", -- t[49] = 99
      "000001101000" when "0110010", -- t[50] = 104
      "000001101100" when "0110011", -- t[51] = 108
      "000001110001" when "0110100", -- t[52] = 113
      "000001110101" when "0110101", -- t[53] = 117
      "000001111010" when "0110110", -- t[54] = 122
      "000010000000" when "0110111", -- t[55] = 128
      "000010000101" when "0111000", -- t[56] = 133
      "000010001011" when "0111001", -- t[57] = 139
      "000010010000" when "0111010", -- t[58] = 144
      "000010010111" when "0111011", -- t[59] = 151
      "000010011101" when "0111100", -- t[60] = 157
      "000010100100" when "0111101", -- t[61] = 164
      "000010101011" when "0111110", -- t[62] = 171
      "000010110010" when "0111111", -- t[63] = 178
      "000010111001" when "1000000", -- t[64] = 185
      "000011000001" when "1000001", -- t[65] = 193
      "000011001001" when "1000010", -- t[66] = 201
      "000011010010" when "1000011", -- t[67] = 210
      "000011011011" when "1000100", -- t[68] = 219
      "000011100100" when "1000101", -- t[69] = 228
      "000011101110" when "1000110", -- t[70] = 238
      "000011110111" when "1000111", -- t[71] = 247
      "000100000010" when "1001000", -- t[72] = 258
      "000100001101" when "1001001", -- t[73] = 269
      "000100011000" when "1001010", -- t[74] = 280
      "000100100100" when "1001011", -- t[75] = 292
      "000100110000" when "1001100", -- t[76] = 304
      "000100111100" when "1001101", -- t[77] = 316
      "000101001010" when "1001110", -- t[78] = 330
      "000101010111" when "1001111", -- t[79] = 343
      "000101100110" when "1010000", -- t[80] = 358
      "000101110100" when "1010001", -- t[81] = 372
      "000110000100" when "1010010", -- t[82] = 388
      "000110010100" when "1010011", -- t[83] = 404
      "000110100100" when "1010100", -- t[84] = 420
      "000110110101" when "1010101", -- t[85] = 437
      "000111000111" when "1010110", -- t[86] = 455
      "000111011010" when "1010111", -- t[87] = 474
      "000111101101" when "1011000", -- t[88] = 493
      "001000000001" when "1011001", -- t[89] = 513
      "001000010110" when "1011010", -- t[90] = 534
      "001000101011" when "1011011", -- t[91] = 555
      "001001000001" when "1011100", -- t[92] = 577
      "001001011000" when "1011101", -- t[93] = 600
      "001001110000" when "1011110", -- t[94] = 624
      "001010001001" when "1011111", -- t[95] = 649
      "001010100010" when "1100000", -- t[96] = 674
      "001010111101" when "1100001", -- t[97] = 701
      "001011011000" when "1100010", -- t[98] = 728
      "001011110101" when "1100011", -- t[99] = 757
      "001100010010" when "1100100", -- t[100] = 786
      "001100110000" when "1100101", -- t[101] = 816
      "001101010000" when "1100110", -- t[102] = 848
      "001101110000" when "1100111", -- t[103] = 880
      "001110010001" when "1101000", -- t[104] = 913
      "001110110100" when "1101001", -- t[105] = 948
      "001111011000" when "1101010", -- t[106] = 984
      "001111111100" when "1101011", -- t[107] = 1020
      "010000100010" when "1101100", -- t[108] = 1058
      "010001001001" when "1101101", -- t[109] = 1097
      "010001110001" when "1101110", -- t[110] = 1137
      "010010011011" when "1101111", -- t[111] = 1179
      "010011000101" when "1110000", -- t[112] = 1221
      "010011110001" when "1110001", -- t[113] = 1265
      "010100011110" when "1110010", -- t[114] = 1310
      "010101001101" when "1110011", -- t[115] = 1357
      "010101111101" when "1110100", -- t[116] = 1405
      "010110101110" when "1110101", -- t[117] = 1454
      "010111100000" when "1110110", -- t[118] = 1504
      "011000010100" when "1110111", -- t[119] = 1556
      "011001001001" when "1111000", -- t[120] = 1609
      "011001111111" when "1111001", -- t[121] = 1663
      "011010110111" when "1111010", -- t[122] = 1719
      "011011110000" when "1111011", -- t[123] = 1776
      "011100101010" when "1111100", -- t[124] = 1834
      "011101100110" when "1111101", -- t[125] = 1894
      "011110100011" when "1111110", -- t[126] = 1955
      "011111100010" when "1111111", -- t[127] = 2018
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_9_to1 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9_to1 is
begin
  with x select
    r <=
      "00000" when "0000000", -- t[0] = 0
      "00000" when "0000001", -- t[1] = 0
      "00000" when "0000010", -- t[2] = 0
      "00000" when "0000011", -- t[3] = 0
      "00000" when "0000100", -- t[4] = 0
      "00000" when "0000101", -- t[5] = 0
      "00000" when "0000110", -- t[6] = 0
      "00000" when "0000111", -- t[7] = 0
      "00000" when "0001000", -- t[8] = 0
      "00000" when "0001001", -- t[9] = 0
      "00000" when "0001010", -- t[10] = 0
      "00000" when "0001011", -- t[11] = 0
      "00000" when "0001100", -- t[12] = 0
      "00000" when "0001101", -- t[13] = 0
      "00000" when "0001110", -- t[14] = 0
      "00000" when "0001111", -- t[15] = 0
      "00000" when "0010000", -- t[16] = 0
      "00000" when "0010001", -- t[17] = 0
      "00000" when "0010010", -- t[18] = 0
      "00000" when "0010011", -- t[19] = 0
      "00000" when "0010100", -- t[20] = 0
      "00000" when "0010101", -- t[21] = 0
      "00000" when "0010110", -- t[22] = 0
      "00000" when "0010111", -- t[23] = 0
      "00000" when "0011000", -- t[24] = 0
      "00000" when "0011001", -- t[25] = 0
      "00000" when "0011010", -- t[26] = 0
      "00000" when "0011011", -- t[27] = 0
      "00000" when "0011100", -- t[28] = 0
      "00000" when "0011101", -- t[29] = 0
      "00000" when "0011110", -- t[30] = 0
      "00000" when "0011111", -- t[31] = 0
      "00000" when "0100000", -- t[32] = 0
      "00000" when "0100001", -- t[33] = 0
      "00000" when "0100010", -- t[34] = 0
      "00000" when "0100011", -- t[35] = 0
      "00000" when "0100100", -- t[36] = 0
      "00000" when "0100101", -- t[37] = 0
      "00000" when "0100110", -- t[38] = 0
      "00000" when "0100111", -- t[39] = 0
      "00000" when "0101000", -- t[40] = 0
      "00001" when "0101001", -- t[41] = 1
      "00000" when "0101010", -- t[42] = 0
      "00001" when "0101011", -- t[43] = 1
      "00000" when "0101100", -- t[44] = 0
      "00001" when "0101101", -- t[45] = 1
      "00000" when "0101110", -- t[46] = 0
      "00001" when "0101111", -- t[47] = 1
      "00000" when "0110000", -- t[48] = 0
      "00001" when "0110001", -- t[49] = 1
      "00000" when "0110010", -- t[50] = 0
      "00001" when "0110011", -- t[51] = 1
      "00000" when "0110100", -- t[52] = 0
      "00001" when "0110101", -- t[53] = 1
      "00000" when "0110110", -- t[54] = 0
      "00001" when "0110111", -- t[55] = 1
      "00000" when "0111000", -- t[56] = 0
      "00010" when "0111001", -- t[57] = 2
      "00000" when "0111010", -- t[58] = 0
      "00010" when "0111011", -- t[59] = 2
      "00000" when "0111100", -- t[60] = 0
      "00010" when "0111101", -- t[61] = 2
      "00000" when "0111110", -- t[62] = 0
      "00010" when "0111111", -- t[63] = 2
      "00000" when "1000000", -- t[64] = 0
      "00010" when "1000001", -- t[65] = 2
      "00001" when "1000010", -- t[66] = 1
      "00011" when "1000011", -- t[67] = 3
      "00001" when "1000100", -- t[68] = 1
      "00011" when "1000101", -- t[69] = 3
      "00001" when "1000110", -- t[70] = 1
      "00011" when "1000111", -- t[71] = 3
      "00001" when "1001000", -- t[72] = 1
      "00100" when "1001001", -- t[73] = 4
      "00001" when "1001010", -- t[74] = 1
      "00100" when "1001011", -- t[75] = 4
      "00001" when "1001100", -- t[76] = 1
      "00100" when "1001101", -- t[77] = 4
      "00001" when "1001110", -- t[78] = 1
      "00101" when "1001111", -- t[79] = 5
      "00001" when "1010000", -- t[80] = 1
      "00101" when "1010001", -- t[81] = 5
      "00001" when "1010010", -- t[82] = 1
      "00101" when "1010011", -- t[83] = 5
      "00010" when "1010100", -- t[84] = 2
      "00110" when "1010101", -- t[85] = 6
      "00010" when "1010110", -- t[86] = 2
      "00110" when "1010111", -- t[87] = 6
      "00010" when "1011000", -- t[88] = 2
      "00111" when "1011001", -- t[89] = 7
      "00010" when "1011010", -- t[90] = 2
      "01000" when "1011011", -- t[91] = 8
      "00010" when "1011100", -- t[92] = 2
      "01000" when "1011101", -- t[93] = 8
      "00011" when "1011110", -- t[94] = 3
      "01001" when "1011111", -- t[95] = 9
      "00011" when "1100000", -- t[96] = 3
      "01001" when "1100001", -- t[97] = 9
      "00011" when "1100010", -- t[98] = 3
      "01010" when "1100011", -- t[99] = 10
      "00011" when "1100100", -- t[100] = 3
      "01011" when "1100101", -- t[101] = 11
      "00100" when "1100110", -- t[102] = 4
      "01100" when "1100111", -- t[103] = 12
      "00100" when "1101000", -- t[104] = 4
      "01100" when "1101001", -- t[105] = 12
      "00100" when "1101010", -- t[106] = 4
      "01101" when "1101011", -- t[107] = 13
      "00100" when "1101100", -- t[108] = 4
      "01110" when "1101101", -- t[109] = 14
      "00101" when "1101110", -- t[110] = 5
      "01111" when "1101111", -- t[111] = 15
      "00101" when "1110000", -- t[112] = 5
      "10000" when "1110001", -- t[113] = 16
      "00101" when "1110010", -- t[114] = 5
      "10001" when "1110011", -- t[115] = 17
      "00110" when "1110100", -- t[116] = 6
      "10010" when "1110101", -- t[117] = 18
      "00110" when "1110110", -- t[118] = 6
      "10011" when "1110111", -- t[119] = 19
      "00110" when "1111000", -- t[120] = 6
      "10100" when "1111001", -- t[121] = 20
      "00111" when "1111010", -- t[122] = 7
      "10101" when "1111011", -- t[123] = 21
      "00111" when "1111100", -- t[124] = 7
      "10110" when "1111101", -- t[125] = 22
      "00111" when "1111110", -- t[126] = 7
      "10111" when "1111111", -- t[127] = 23
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_9_to0 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9_to0 is
begin
  with x select
    r <=
      "000" when "000000", -- t[0] = 0
      "000" when "000001", -- t[1] = 0
      "000" when "000010", -- t[2] = 0
      "000" when "000011", -- t[3] = 0
      "000" when "000100", -- t[4] = 0
      "000" when "000101", -- t[5] = 0
      "000" when "000110", -- t[6] = 0
      "000" when "000111", -- t[7] = 0
      "000" when "001000", -- t[8] = 0
      "000" when "001001", -- t[9] = 0
      "000" when "001010", -- t[10] = 0
      "000" when "001011", -- t[11] = 0
      "000" when "001100", -- t[12] = 0
      "000" when "001101", -- t[13] = 0
      "000" when "001110", -- t[14] = 0
      "000" when "001111", -- t[15] = 0
      "000" when "010000", -- t[16] = 0
      "000" when "010001", -- t[17] = 0
      "000" when "010010", -- t[18] = 0
      "000" when "010011", -- t[19] = 0
      "000" when "010100", -- t[20] = 0
      "000" when "010101", -- t[21] = 0
      "000" when "010110", -- t[22] = 0
      "000" when "010111", -- t[23] = 0
      "000" when "011000", -- t[24] = 0
      "000" when "011001", -- t[25] = 0
      "000" when "011010", -- t[26] = 0
      "000" when "011011", -- t[27] = 0
      "000" when "011100", -- t[28] = 0
      "000" when "011101", -- t[29] = 0
      "000" when "011110", -- t[30] = 0
      "000" when "011111", -- t[31] = 0
      "000" when "100000", -- t[32] = 0
      "000" when "100001", -- t[33] = 0
      "000" when "100010", -- t[34] = 0
      "000" when "100011", -- t[35] = 0
      "000" when "100100", -- t[36] = 0
      "000" when "100101", -- t[37] = 0
      "000" when "100110", -- t[38] = 0
      "001" when "100111", -- t[39] = 1
      "000" when "101000", -- t[40] = 0
      "000" when "101001", -- t[41] = 0
      "001" when "101010", -- t[42] = 1
      "001" when "101011", -- t[43] = 1
      "000" when "101100", -- t[44] = 0
      "001" when "101101", -- t[45] = 1
      "001" when "101110", -- t[46] = 1
      "010" when "101111", -- t[47] = 2
      "000" when "110000", -- t[48] = 0
      "001" when "110001", -- t[49] = 1
      "010" when "110010", -- t[50] = 2
      "011" when "110011", -- t[51] = 3
      "000" when "110100", -- t[52] = 0
      "001" when "110101", -- t[53] = 1
      "010" when "110110", -- t[54] = 2
      "100" when "110111", -- t[55] = 4
      "000" when "111000", -- t[56] = 0
      "010" when "111001", -- t[57] = 2
      "011" when "111010", -- t[58] = 3
      "101" when "111011", -- t[59] = 5
      "000" when "111100", -- t[60] = 0
      "010" when "111101", -- t[61] = 2
      "100" when "111110", -- t[62] = 4
      "110" when "111111", -- t[63] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_9.all;

entity LNSAdd_MPT_T2_9_to1_xor is
  port( a : in  std_logic_vector(5 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(6 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(6 downto 1) <= a(5 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSAdd_MPT_T2_9_to1
    port map( x => in_t,
              r => out_t );

  r(11 downto 5) <= (11 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_9.all;

entity LNSAdd_MPT_T2_9_to0_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(2);
  in_t(5 downto 2) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSAdd_MPT_T2_9_to0
    port map( x => in_t,
              r => out_t );

  r(11 downto 3) <= (11 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_9.all;

entity LNSAdd_MPT_T2_9 is
  port( x : in  std_logic_vector(11 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_9 is
  signal in_tiv  : std_logic_vector(6 downto 0);
  signal out_tiv : std_logic_vector(11 downto 0);
  signal a1      : std_logic_vector(5 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(11 downto 0);
  signal a0      : std_logic_vector(3 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(11 downto 0);
  signal sum     : std_logic_vector(11 downto 0);
begin
  in_tiv <= x(11 downto 5);
  inst_tiv : LNSAdd_MPT_T2_9_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(11 downto 6);
  b1 <= x(4 downto 3);
  inst_to1_xor : LNSAdd_MPT_T2_9_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(11 downto 8);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSAdd_MPT_T2_9_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(11 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_9.all;
use fplib.pkg_misc.all;

entity LNSAdd_MPT_T2_9_Clk is
  port( x   : in  std_logic_vector(11 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSAdd_MPT_T2_9_Clk is
  signal in_tiv_1  : std_logic_vector(6 downto 0);
  signal out_tiv_1 : std_logic_vector(11 downto 0);
  signal out_tiv_2 : std_logic_vector(11 downto 0);
  signal a1_1      : std_logic_vector(5 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(11 downto 0);
  signal out1_2    : std_logic_vector(11 downto 0);
  signal a0_1      : std_logic_vector(3 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(11 downto 0);
  signal out0_2    : std_logic_vector(11 downto 0);
  signal psum1_2     : std_logic_vector(11 downto 0);
  signal psum1_3     : std_logic_vector(11 downto 0);
  signal psum2_2     : std_logic_vector(11 downto 0);
  signal psum2_3     : std_logic_vector(11 downto 0);
  signal sum_3     : std_logic_vector(11 downto 0);
begin
  in_tiv_1 <= x(11 downto 5);
  inst_tiv : LNSAdd_MPT_T2_9_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(11 downto 6);
  b1_1 <= x(4 downto 3);
  inst_to1_xor : LNSAdd_MPT_T2_9_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(11 downto 8);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSAdd_MPT_T2_9_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(11 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_9.all;

entity LNSAdd_MPT_9 is
  port( x : in  std_logic_vector(12 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_9 is
  signal out_t1 : std_logic_vector(2 downto 0);
  signal out_t2 : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSAdd_MPT_T1_9
    port map( x => x,
              r => out_t1 );

  inst_t2 : LNSAdd_MPT_T2_9
    port map( x => x(11 downto 0),
              r => out_t2 );

  r <= out_t2 when x(12 downto 12) = (12 downto 12 => '1') else
       (9 downto 3 => '0') & out_t1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_9.all;
use fplib.pkg_misc.all;

entity LNSAdd_MPT_9_Clk is
  port( x   : in  std_logic_vector(12 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSAdd_MPT_9_Clk is
  signal x_1  : std_logic_vector(12 downto 0);
  signal x_10 : std_logic_vector(12 downto 0);

  signal out_t1_1  : std_logic_vector(2 downto 0);
  signal out_t1_10 : std_logic_vector(2 downto 0);
  signal out_t2_10 : std_logic_vector(9 downto 0);
begin
  x_1 <= x;

  inst_t1 : LNSAdd_MPT_T1_9
    port map( x => x_1,
              r => out_t1_1 );

  out_t1_delay : Delay
    generic map ( w => 3,
                  n => 1 )
    port map ( input  => out_t1_1,
               output => out_t1_10,
               clk    => clk );

  inst_t2 : LNSAdd_MPT_T2_9_Clk
    port map( x   => x(11 downto 0),
              r   => out_t2_10,
              clk => clk );

  x_delay : Delay
    generic map ( w => 13,
                  n => 1 )
    port map ( input  => x_1,
               output => x_10,
               clk    => clk );

  r <= out_t2_10 when x_10(12 downto 12) = (12 downto 12 => '1') else
       (9 downto 3 => '0') & out_t1_10;
end architecture;
