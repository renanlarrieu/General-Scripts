library verilog;
use verilog.vl_types.all;
entity circuito_combinacional_vlg_vec_tst is
end circuito_combinacional_vlg_vec_tst;
