incantation

ABER
CAM
GAB
CAR
PUR