-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of MultiPartiteAdder object for LNS arithmetic in base 2.0 with 8-bit integer part and 8-bit fractional part
-- wI = 12 bits
-- wO = 9 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnsadd_mpt_8 is
  component LNSAdd_MPT_T1_8 is
    port( x : in  std_logic_vector(11 downto 0);
          r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8 is
    port( x : in  std_logic_vector(10 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8_Clk is
    port( x   : in  std_logic_vector(10 downto 0);
          r   : out std_logic_vector(8 downto 0);
          clk : in  std_logic );
  end component;
end package;


-- SimpleTable: LNS addition function: [-16.0 0.0[ -> [0.0 2.0[
-- (bounded to [-16.0; -8.0[)
-- wI = 12 bits
-- wO = 2 bits

library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T1_8 is
  port( x : in  std_logic_vector(11 downto 0);
        r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T1_8 is
begin
  with x select
    r <=
      "00" when "000000000000", -- t[0] = 0
      "00" when "000000000001", -- t[1] = 0
      "00" when "000000000010", -- t[2] = 0
      "00" when "000000000011", -- t[3] = 0
      "00" when "000000000100", -- t[4] = 0
      "00" when "000000000101", -- t[5] = 0
      "00" when "000000000110", -- t[6] = 0
      "00" when "000000000111", -- t[7] = 0
      "00" when "000000001000", -- t[8] = 0
      "00" when "000000001001", -- t[9] = 0
      "00" when "000000001010", -- t[10] = 0
      "00" when "000000001011", -- t[11] = 0
      "00" when "000000001100", -- t[12] = 0
      "00" when "000000001101", -- t[13] = 0
      "00" when "000000001110", -- t[14] = 0
      "00" when "000000001111", -- t[15] = 0
      "00" when "000000010000", -- t[16] = 0
      "00" when "000000010001", -- t[17] = 0
      "00" when "000000010010", -- t[18] = 0
      "00" when "000000010011", -- t[19] = 0
      "00" when "000000010100", -- t[20] = 0
      "00" when "000000010101", -- t[21] = 0
      "00" when "000000010110", -- t[22] = 0
      "00" when "000000010111", -- t[23] = 0
      "00" when "000000011000", -- t[24] = 0
      "00" when "000000011001", -- t[25] = 0
      "00" when "000000011010", -- t[26] = 0
      "00" when "000000011011", -- t[27] = 0
      "00" when "000000011100", -- t[28] = 0
      "00" when "000000011101", -- t[29] = 0
      "00" when "000000011110", -- t[30] = 0
      "00" when "000000011111", -- t[31] = 0
      "00" when "000000100000", -- t[32] = 0
      "00" when "000000100001", -- t[33] = 0
      "00" when "000000100010", -- t[34] = 0
      "00" when "000000100011", -- t[35] = 0
      "00" when "000000100100", -- t[36] = 0
      "00" when "000000100101", -- t[37] = 0
      "00" when "000000100110", -- t[38] = 0
      "00" when "000000100111", -- t[39] = 0
      "00" when "000000101000", -- t[40] = 0
      "00" when "000000101001", -- t[41] = 0
      "00" when "000000101010", -- t[42] = 0
      "00" when "000000101011", -- t[43] = 0
      "00" when "000000101100", -- t[44] = 0
      "00" when "000000101101", -- t[45] = 0
      "00" when "000000101110", -- t[46] = 0
      "00" when "000000101111", -- t[47] = 0
      "00" when "000000110000", -- t[48] = 0
      "00" when "000000110001", -- t[49] = 0
      "00" when "000000110010", -- t[50] = 0
      "00" when "000000110011", -- t[51] = 0
      "00" when "000000110100", -- t[52] = 0
      "00" when "000000110101", -- t[53] = 0
      "00" when "000000110110", -- t[54] = 0
      "00" when "000000110111", -- t[55] = 0
      "00" when "000000111000", -- t[56] = 0
      "00" when "000000111001", -- t[57] = 0
      "00" when "000000111010", -- t[58] = 0
      "00" when "000000111011", -- t[59] = 0
      "00" when "000000111100", -- t[60] = 0
      "00" when "000000111101", -- t[61] = 0
      "00" when "000000111110", -- t[62] = 0
      "00" when "000000111111", -- t[63] = 0
      "00" when "000001000000", -- t[64] = 0
      "00" when "000001000001", -- t[65] = 0
      "00" when "000001000010", -- t[66] = 0
      "00" when "000001000011", -- t[67] = 0
      "00" when "000001000100", -- t[68] = 0
      "00" when "000001000101", -- t[69] = 0
      "00" when "000001000110", -- t[70] = 0
      "00" when "000001000111", -- t[71] = 0
      "00" when "000001001000", -- t[72] = 0
      "00" when "000001001001", -- t[73] = 0
      "00" when "000001001010", -- t[74] = 0
      "00" when "000001001011", -- t[75] = 0
      "00" when "000001001100", -- t[76] = 0
      "00" when "000001001101", -- t[77] = 0
      "00" when "000001001110", -- t[78] = 0
      "00" when "000001001111", -- t[79] = 0
      "00" when "000001010000", -- t[80] = 0
      "00" when "000001010001", -- t[81] = 0
      "00" when "000001010010", -- t[82] = 0
      "00" when "000001010011", -- t[83] = 0
      "00" when "000001010100", -- t[84] = 0
      "00" when "000001010101", -- t[85] = 0
      "00" when "000001010110", -- t[86] = 0
      "00" when "000001010111", -- t[87] = 0
      "00" when "000001011000", -- t[88] = 0
      "00" when "000001011001", -- t[89] = 0
      "00" when "000001011010", -- t[90] = 0
      "00" when "000001011011", -- t[91] = 0
      "00" when "000001011100", -- t[92] = 0
      "00" when "000001011101", -- t[93] = 0
      "00" when "000001011110", -- t[94] = 0
      "00" when "000001011111", -- t[95] = 0
      "00" when "000001100000", -- t[96] = 0
      "00" when "000001100001", -- t[97] = 0
      "00" when "000001100010", -- t[98] = 0
      "00" when "000001100011", -- t[99] = 0
      "00" when "000001100100", -- t[100] = 0
      "00" when "000001100101", -- t[101] = 0
      "00" when "000001100110", -- t[102] = 0
      "00" when "000001100111", -- t[103] = 0
      "00" when "000001101000", -- t[104] = 0
      "00" when "000001101001", -- t[105] = 0
      "00" when "000001101010", -- t[106] = 0
      "00" when "000001101011", -- t[107] = 0
      "00" when "000001101100", -- t[108] = 0
      "00" when "000001101101", -- t[109] = 0
      "00" when "000001101110", -- t[110] = 0
      "00" when "000001101111", -- t[111] = 0
      "00" when "000001110000", -- t[112] = 0
      "00" when "000001110001", -- t[113] = 0
      "00" when "000001110010", -- t[114] = 0
      "00" when "000001110011", -- t[115] = 0
      "00" when "000001110100", -- t[116] = 0
      "00" when "000001110101", -- t[117] = 0
      "00" when "000001110110", -- t[118] = 0
      "00" when "000001110111", -- t[119] = 0
      "00" when "000001111000", -- t[120] = 0
      "00" when "000001111001", -- t[121] = 0
      "00" when "000001111010", -- t[122] = 0
      "00" when "000001111011", -- t[123] = 0
      "00" when "000001111100", -- t[124] = 0
      "00" when "000001111101", -- t[125] = 0
      "00" when "000001111110", -- t[126] = 0
      "00" when "000001111111", -- t[127] = 0
      "00" when "000010000000", -- t[128] = 0
      "00" when "000010000001", -- t[129] = 0
      "00" when "000010000010", -- t[130] = 0
      "00" when "000010000011", -- t[131] = 0
      "00" when "000010000100", -- t[132] = 0
      "00" when "000010000101", -- t[133] = 0
      "00" when "000010000110", -- t[134] = 0
      "00" when "000010000111", -- t[135] = 0
      "00" when "000010001000", -- t[136] = 0
      "00" when "000010001001", -- t[137] = 0
      "00" when "000010001010", -- t[138] = 0
      "00" when "000010001011", -- t[139] = 0
      "00" when "000010001100", -- t[140] = 0
      "00" when "000010001101", -- t[141] = 0
      "00" when "000010001110", -- t[142] = 0
      "00" when "000010001111", -- t[143] = 0
      "00" when "000010010000", -- t[144] = 0
      "00" when "000010010001", -- t[145] = 0
      "00" when "000010010010", -- t[146] = 0
      "00" when "000010010011", -- t[147] = 0
      "00" when "000010010100", -- t[148] = 0
      "00" when "000010010101", -- t[149] = 0
      "00" when "000010010110", -- t[150] = 0
      "00" when "000010010111", -- t[151] = 0
      "00" when "000010011000", -- t[152] = 0
      "00" when "000010011001", -- t[153] = 0
      "00" when "000010011010", -- t[154] = 0
      "00" when "000010011011", -- t[155] = 0
      "00" when "000010011100", -- t[156] = 0
      "00" when "000010011101", -- t[157] = 0
      "00" when "000010011110", -- t[158] = 0
      "00" when "000010011111", -- t[159] = 0
      "00" when "000010100000", -- t[160] = 0
      "00" when "000010100001", -- t[161] = 0
      "00" when "000010100010", -- t[162] = 0
      "00" when "000010100011", -- t[163] = 0
      "00" when "000010100100", -- t[164] = 0
      "00" when "000010100101", -- t[165] = 0
      "00" when "000010100110", -- t[166] = 0
      "00" when "000010100111", -- t[167] = 0
      "00" when "000010101000", -- t[168] = 0
      "00" when "000010101001", -- t[169] = 0
      "00" when "000010101010", -- t[170] = 0
      "00" when "000010101011", -- t[171] = 0
      "00" when "000010101100", -- t[172] = 0
      "00" when "000010101101", -- t[173] = 0
      "00" when "000010101110", -- t[174] = 0
      "00" when "000010101111", -- t[175] = 0
      "00" when "000010110000", -- t[176] = 0
      "00" when "000010110001", -- t[177] = 0
      "00" when "000010110010", -- t[178] = 0
      "00" when "000010110011", -- t[179] = 0
      "00" when "000010110100", -- t[180] = 0
      "00" when "000010110101", -- t[181] = 0
      "00" when "000010110110", -- t[182] = 0
      "00" when "000010110111", -- t[183] = 0
      "00" when "000010111000", -- t[184] = 0
      "00" when "000010111001", -- t[185] = 0
      "00" when "000010111010", -- t[186] = 0
      "00" when "000010111011", -- t[187] = 0
      "00" when "000010111100", -- t[188] = 0
      "00" when "000010111101", -- t[189] = 0
      "00" when "000010111110", -- t[190] = 0
      "00" when "000010111111", -- t[191] = 0
      "00" when "000011000000", -- t[192] = 0
      "00" when "000011000001", -- t[193] = 0
      "00" when "000011000010", -- t[194] = 0
      "00" when "000011000011", -- t[195] = 0
      "00" when "000011000100", -- t[196] = 0
      "00" when "000011000101", -- t[197] = 0
      "00" when "000011000110", -- t[198] = 0
      "00" when "000011000111", -- t[199] = 0
      "00" when "000011001000", -- t[200] = 0
      "00" when "000011001001", -- t[201] = 0
      "00" when "000011001010", -- t[202] = 0
      "00" when "000011001011", -- t[203] = 0
      "00" when "000011001100", -- t[204] = 0
      "00" when "000011001101", -- t[205] = 0
      "00" when "000011001110", -- t[206] = 0
      "00" when "000011001111", -- t[207] = 0
      "00" when "000011010000", -- t[208] = 0
      "00" when "000011010001", -- t[209] = 0
      "00" when "000011010010", -- t[210] = 0
      "00" when "000011010011", -- t[211] = 0
      "00" when "000011010100", -- t[212] = 0
      "00" when "000011010101", -- t[213] = 0
      "00" when "000011010110", -- t[214] = 0
      "00" when "000011010111", -- t[215] = 0
      "00" when "000011011000", -- t[216] = 0
      "00" when "000011011001", -- t[217] = 0
      "00" when "000011011010", -- t[218] = 0
      "00" when "000011011011", -- t[219] = 0
      "00" when "000011011100", -- t[220] = 0
      "00" when "000011011101", -- t[221] = 0
      "00" when "000011011110", -- t[222] = 0
      "00" when "000011011111", -- t[223] = 0
      "00" when "000011100000", -- t[224] = 0
      "00" when "000011100001", -- t[225] = 0
      "00" when "000011100010", -- t[226] = 0
      "00" when "000011100011", -- t[227] = 0
      "00" when "000011100100", -- t[228] = 0
      "00" when "000011100101", -- t[229] = 0
      "00" when "000011100110", -- t[230] = 0
      "00" when "000011100111", -- t[231] = 0
      "00" when "000011101000", -- t[232] = 0
      "00" when "000011101001", -- t[233] = 0
      "00" when "000011101010", -- t[234] = 0
      "00" when "000011101011", -- t[235] = 0
      "00" when "000011101100", -- t[236] = 0
      "00" when "000011101101", -- t[237] = 0
      "00" when "000011101110", -- t[238] = 0
      "00" when "000011101111", -- t[239] = 0
      "00" when "000011110000", -- t[240] = 0
      "00" when "000011110001", -- t[241] = 0
      "00" when "000011110010", -- t[242] = 0
      "00" when "000011110011", -- t[243] = 0
      "00" when "000011110100", -- t[244] = 0
      "00" when "000011110101", -- t[245] = 0
      "00" when "000011110110", -- t[246] = 0
      "00" when "000011110111", -- t[247] = 0
      "00" when "000011111000", -- t[248] = 0
      "00" when "000011111001", -- t[249] = 0
      "00" when "000011111010", -- t[250] = 0
      "00" when "000011111011", -- t[251] = 0
      "00" when "000011111100", -- t[252] = 0
      "00" when "000011111101", -- t[253] = 0
      "00" when "000011111110", -- t[254] = 0
      "00" when "000011111111", -- t[255] = 0
      "00" when "000100000000", -- t[256] = 0
      "00" when "000100000001", -- t[257] = 0
      "00" when "000100000010", -- t[258] = 0
      "00" when "000100000011", -- t[259] = 0
      "00" when "000100000100", -- t[260] = 0
      "00" when "000100000101", -- t[261] = 0
      "00" when "000100000110", -- t[262] = 0
      "00" when "000100000111", -- t[263] = 0
      "00" when "000100001000", -- t[264] = 0
      "00" when "000100001001", -- t[265] = 0
      "00" when "000100001010", -- t[266] = 0
      "00" when "000100001011", -- t[267] = 0
      "00" when "000100001100", -- t[268] = 0
      "00" when "000100001101", -- t[269] = 0
      "00" when "000100001110", -- t[270] = 0
      "00" when "000100001111", -- t[271] = 0
      "00" when "000100010000", -- t[272] = 0
      "00" when "000100010001", -- t[273] = 0
      "00" when "000100010010", -- t[274] = 0
      "00" when "000100010011", -- t[275] = 0
      "00" when "000100010100", -- t[276] = 0
      "00" when "000100010101", -- t[277] = 0
      "00" when "000100010110", -- t[278] = 0
      "00" when "000100010111", -- t[279] = 0
      "00" when "000100011000", -- t[280] = 0
      "00" when "000100011001", -- t[281] = 0
      "00" when "000100011010", -- t[282] = 0
      "00" when "000100011011", -- t[283] = 0
      "00" when "000100011100", -- t[284] = 0
      "00" when "000100011101", -- t[285] = 0
      "00" when "000100011110", -- t[286] = 0
      "00" when "000100011111", -- t[287] = 0
      "00" when "000100100000", -- t[288] = 0
      "00" when "000100100001", -- t[289] = 0
      "00" when "000100100010", -- t[290] = 0
      "00" when "000100100011", -- t[291] = 0
      "00" when "000100100100", -- t[292] = 0
      "00" when "000100100101", -- t[293] = 0
      "00" when "000100100110", -- t[294] = 0
      "00" when "000100100111", -- t[295] = 0
      "00" when "000100101000", -- t[296] = 0
      "00" when "000100101001", -- t[297] = 0
      "00" when "000100101010", -- t[298] = 0
      "00" when "000100101011", -- t[299] = 0
      "00" when "000100101100", -- t[300] = 0
      "00" when "000100101101", -- t[301] = 0
      "00" when "000100101110", -- t[302] = 0
      "00" when "000100101111", -- t[303] = 0
      "00" when "000100110000", -- t[304] = 0
      "00" when "000100110001", -- t[305] = 0
      "00" when "000100110010", -- t[306] = 0
      "00" when "000100110011", -- t[307] = 0
      "00" when "000100110100", -- t[308] = 0
      "00" when "000100110101", -- t[309] = 0
      "00" when "000100110110", -- t[310] = 0
      "00" when "000100110111", -- t[311] = 0
      "00" when "000100111000", -- t[312] = 0
      "00" when "000100111001", -- t[313] = 0
      "00" when "000100111010", -- t[314] = 0
      "00" when "000100111011", -- t[315] = 0
      "00" when "000100111100", -- t[316] = 0
      "00" when "000100111101", -- t[317] = 0
      "00" when "000100111110", -- t[318] = 0
      "00" when "000100111111", -- t[319] = 0
      "00" when "000101000000", -- t[320] = 0
      "00" when "000101000001", -- t[321] = 0
      "00" when "000101000010", -- t[322] = 0
      "00" when "000101000011", -- t[323] = 0
      "00" when "000101000100", -- t[324] = 0
      "00" when "000101000101", -- t[325] = 0
      "00" when "000101000110", -- t[326] = 0
      "00" when "000101000111", -- t[327] = 0
      "00" when "000101001000", -- t[328] = 0
      "00" when "000101001001", -- t[329] = 0
      "00" when "000101001010", -- t[330] = 0
      "00" when "000101001011", -- t[331] = 0
      "00" when "000101001100", -- t[332] = 0
      "00" when "000101001101", -- t[333] = 0
      "00" when "000101001110", -- t[334] = 0
      "00" when "000101001111", -- t[335] = 0
      "00" when "000101010000", -- t[336] = 0
      "00" when "000101010001", -- t[337] = 0
      "00" when "000101010010", -- t[338] = 0
      "00" when "000101010011", -- t[339] = 0
      "00" when "000101010100", -- t[340] = 0
      "00" when "000101010101", -- t[341] = 0
      "00" when "000101010110", -- t[342] = 0
      "00" when "000101010111", -- t[343] = 0
      "00" when "000101011000", -- t[344] = 0
      "00" when "000101011001", -- t[345] = 0
      "00" when "000101011010", -- t[346] = 0
      "00" when "000101011011", -- t[347] = 0
      "00" when "000101011100", -- t[348] = 0
      "00" when "000101011101", -- t[349] = 0
      "00" when "000101011110", -- t[350] = 0
      "00" when "000101011111", -- t[351] = 0
      "00" when "000101100000", -- t[352] = 0
      "00" when "000101100001", -- t[353] = 0
      "00" when "000101100010", -- t[354] = 0
      "00" when "000101100011", -- t[355] = 0
      "00" when "000101100100", -- t[356] = 0
      "00" when "000101100101", -- t[357] = 0
      "00" when "000101100110", -- t[358] = 0
      "00" when "000101100111", -- t[359] = 0
      "00" when "000101101000", -- t[360] = 0
      "00" when "000101101001", -- t[361] = 0
      "00" when "000101101010", -- t[362] = 0
      "00" when "000101101011", -- t[363] = 0
      "00" when "000101101100", -- t[364] = 0
      "00" when "000101101101", -- t[365] = 0
      "00" when "000101101110", -- t[366] = 0
      "00" when "000101101111", -- t[367] = 0
      "00" when "000101110000", -- t[368] = 0
      "00" when "000101110001", -- t[369] = 0
      "00" when "000101110010", -- t[370] = 0
      "00" when "000101110011", -- t[371] = 0
      "00" when "000101110100", -- t[372] = 0
      "00" when "000101110101", -- t[373] = 0
      "00" when "000101110110", -- t[374] = 0
      "00" when "000101110111", -- t[375] = 0
      "00" when "000101111000", -- t[376] = 0
      "00" when "000101111001", -- t[377] = 0
      "00" when "000101111010", -- t[378] = 0
      "00" when "000101111011", -- t[379] = 0
      "00" when "000101111100", -- t[380] = 0
      "00" when "000101111101", -- t[381] = 0
      "00" when "000101111110", -- t[382] = 0
      "00" when "000101111111", -- t[383] = 0
      "00" when "000110000000", -- t[384] = 0
      "00" when "000110000001", -- t[385] = 0
      "00" when "000110000010", -- t[386] = 0
      "00" when "000110000011", -- t[387] = 0
      "00" when "000110000100", -- t[388] = 0
      "00" when "000110000101", -- t[389] = 0
      "00" when "000110000110", -- t[390] = 0
      "00" when "000110000111", -- t[391] = 0
      "00" when "000110001000", -- t[392] = 0
      "00" when "000110001001", -- t[393] = 0
      "00" when "000110001010", -- t[394] = 0
      "00" when "000110001011", -- t[395] = 0
      "00" when "000110001100", -- t[396] = 0
      "00" when "000110001101", -- t[397] = 0
      "00" when "000110001110", -- t[398] = 0
      "00" when "000110001111", -- t[399] = 0
      "00" when "000110010000", -- t[400] = 0
      "00" when "000110010001", -- t[401] = 0
      "00" when "000110010010", -- t[402] = 0
      "00" when "000110010011", -- t[403] = 0
      "00" when "000110010100", -- t[404] = 0
      "00" when "000110010101", -- t[405] = 0
      "00" when "000110010110", -- t[406] = 0
      "00" when "000110010111", -- t[407] = 0
      "00" when "000110011000", -- t[408] = 0
      "00" when "000110011001", -- t[409] = 0
      "00" when "000110011010", -- t[410] = 0
      "00" when "000110011011", -- t[411] = 0
      "00" when "000110011100", -- t[412] = 0
      "00" when "000110011101", -- t[413] = 0
      "00" when "000110011110", -- t[414] = 0
      "00" when "000110011111", -- t[415] = 0
      "00" when "000110100000", -- t[416] = 0
      "00" when "000110100001", -- t[417] = 0
      "00" when "000110100010", -- t[418] = 0
      "00" when "000110100011", -- t[419] = 0
      "00" when "000110100100", -- t[420] = 0
      "00" when "000110100101", -- t[421] = 0
      "00" when "000110100110", -- t[422] = 0
      "00" when "000110100111", -- t[423] = 0
      "00" when "000110101000", -- t[424] = 0
      "00" when "000110101001", -- t[425] = 0
      "00" when "000110101010", -- t[426] = 0
      "00" when "000110101011", -- t[427] = 0
      "00" when "000110101100", -- t[428] = 0
      "00" when "000110101101", -- t[429] = 0
      "00" when "000110101110", -- t[430] = 0
      "00" when "000110101111", -- t[431] = 0
      "00" when "000110110000", -- t[432] = 0
      "00" when "000110110001", -- t[433] = 0
      "00" when "000110110010", -- t[434] = 0
      "00" when "000110110011", -- t[435] = 0
      "00" when "000110110100", -- t[436] = 0
      "00" when "000110110101", -- t[437] = 0
      "00" when "000110110110", -- t[438] = 0
      "00" when "000110110111", -- t[439] = 0
      "00" when "000110111000", -- t[440] = 0
      "00" when "000110111001", -- t[441] = 0
      "00" when "000110111010", -- t[442] = 0
      "00" when "000110111011", -- t[443] = 0
      "00" when "000110111100", -- t[444] = 0
      "00" when "000110111101", -- t[445] = 0
      "00" when "000110111110", -- t[446] = 0
      "00" when "000110111111", -- t[447] = 0
      "00" when "000111000000", -- t[448] = 0
      "00" when "000111000001", -- t[449] = 0
      "00" when "000111000010", -- t[450] = 0
      "00" when "000111000011", -- t[451] = 0
      "00" when "000111000100", -- t[452] = 0
      "00" when "000111000101", -- t[453] = 0
      "00" when "000111000110", -- t[454] = 0
      "00" when "000111000111", -- t[455] = 0
      "00" when "000111001000", -- t[456] = 0
      "00" when "000111001001", -- t[457] = 0
      "00" when "000111001010", -- t[458] = 0
      "00" when "000111001011", -- t[459] = 0
      "00" when "000111001100", -- t[460] = 0
      "00" when "000111001101", -- t[461] = 0
      "00" when "000111001110", -- t[462] = 0
      "00" when "000111001111", -- t[463] = 0
      "00" when "000111010000", -- t[464] = 0
      "00" when "000111010001", -- t[465] = 0
      "00" when "000111010010", -- t[466] = 0
      "00" when "000111010011", -- t[467] = 0
      "00" when "000111010100", -- t[468] = 0
      "00" when "000111010101", -- t[469] = 0
      "00" when "000111010110", -- t[470] = 0
      "00" when "000111010111", -- t[471] = 0
      "00" when "000111011000", -- t[472] = 0
      "00" when "000111011001", -- t[473] = 0
      "00" when "000111011010", -- t[474] = 0
      "00" when "000111011011", -- t[475] = 0
      "00" when "000111011100", -- t[476] = 0
      "00" when "000111011101", -- t[477] = 0
      "00" when "000111011110", -- t[478] = 0
      "00" when "000111011111", -- t[479] = 0
      "00" when "000111100000", -- t[480] = 0
      "00" when "000111100001", -- t[481] = 0
      "00" when "000111100010", -- t[482] = 0
      "00" when "000111100011", -- t[483] = 0
      "00" when "000111100100", -- t[484] = 0
      "00" when "000111100101", -- t[485] = 0
      "00" when "000111100110", -- t[486] = 0
      "00" when "000111100111", -- t[487] = 0
      "00" when "000111101000", -- t[488] = 0
      "00" when "000111101001", -- t[489] = 0
      "00" when "000111101010", -- t[490] = 0
      "00" when "000111101011", -- t[491] = 0
      "00" when "000111101100", -- t[492] = 0
      "00" when "000111101101", -- t[493] = 0
      "00" when "000111101110", -- t[494] = 0
      "00" when "000111101111", -- t[495] = 0
      "00" when "000111110000", -- t[496] = 0
      "00" when "000111110001", -- t[497] = 0
      "00" when "000111110010", -- t[498] = 0
      "00" when "000111110011", -- t[499] = 0
      "00" when "000111110100", -- t[500] = 0
      "00" when "000111110101", -- t[501] = 0
      "00" when "000111110110", -- t[502] = 0
      "00" when "000111110111", -- t[503] = 0
      "00" when "000111111000", -- t[504] = 0
      "00" when "000111111001", -- t[505] = 0
      "00" when "000111111010", -- t[506] = 0
      "00" when "000111111011", -- t[507] = 0
      "00" when "000111111100", -- t[508] = 0
      "00" when "000111111101", -- t[509] = 0
      "00" when "000111111110", -- t[510] = 0
      "00" when "000111111111", -- t[511] = 0
      "00" when "001000000000", -- t[512] = 0
      "00" when "001000000001", -- t[513] = 0
      "00" when "001000000010", -- t[514] = 0
      "00" when "001000000011", -- t[515] = 0
      "00" when "001000000100", -- t[516] = 0
      "00" when "001000000101", -- t[517] = 0
      "00" when "001000000110", -- t[518] = 0
      "00" when "001000000111", -- t[519] = 0
      "00" when "001000001000", -- t[520] = 0
      "00" when "001000001001", -- t[521] = 0
      "00" when "001000001010", -- t[522] = 0
      "00" when "001000001011", -- t[523] = 0
      "00" when "001000001100", -- t[524] = 0
      "00" when "001000001101", -- t[525] = 0
      "00" when "001000001110", -- t[526] = 0
      "00" when "001000001111", -- t[527] = 0
      "00" when "001000010000", -- t[528] = 0
      "00" when "001000010001", -- t[529] = 0
      "00" when "001000010010", -- t[530] = 0
      "00" when "001000010011", -- t[531] = 0
      "00" when "001000010100", -- t[532] = 0
      "00" when "001000010101", -- t[533] = 0
      "00" when "001000010110", -- t[534] = 0
      "00" when "001000010111", -- t[535] = 0
      "00" when "001000011000", -- t[536] = 0
      "00" when "001000011001", -- t[537] = 0
      "00" when "001000011010", -- t[538] = 0
      "00" when "001000011011", -- t[539] = 0
      "00" when "001000011100", -- t[540] = 0
      "00" when "001000011101", -- t[541] = 0
      "00" when "001000011110", -- t[542] = 0
      "00" when "001000011111", -- t[543] = 0
      "00" when "001000100000", -- t[544] = 0
      "00" when "001000100001", -- t[545] = 0
      "00" when "001000100010", -- t[546] = 0
      "00" when "001000100011", -- t[547] = 0
      "00" when "001000100100", -- t[548] = 0
      "00" when "001000100101", -- t[549] = 0
      "00" when "001000100110", -- t[550] = 0
      "00" when "001000100111", -- t[551] = 0
      "00" when "001000101000", -- t[552] = 0
      "00" when "001000101001", -- t[553] = 0
      "00" when "001000101010", -- t[554] = 0
      "00" when "001000101011", -- t[555] = 0
      "00" when "001000101100", -- t[556] = 0
      "00" when "001000101101", -- t[557] = 0
      "00" when "001000101110", -- t[558] = 0
      "00" when "001000101111", -- t[559] = 0
      "00" when "001000110000", -- t[560] = 0
      "00" when "001000110001", -- t[561] = 0
      "00" when "001000110010", -- t[562] = 0
      "00" when "001000110011", -- t[563] = 0
      "00" when "001000110100", -- t[564] = 0
      "00" when "001000110101", -- t[565] = 0
      "00" when "001000110110", -- t[566] = 0
      "00" when "001000110111", -- t[567] = 0
      "00" when "001000111000", -- t[568] = 0
      "00" when "001000111001", -- t[569] = 0
      "00" when "001000111010", -- t[570] = 0
      "00" when "001000111011", -- t[571] = 0
      "00" when "001000111100", -- t[572] = 0
      "00" when "001000111101", -- t[573] = 0
      "00" when "001000111110", -- t[574] = 0
      "00" when "001000111111", -- t[575] = 0
      "00" when "001001000000", -- t[576] = 0
      "00" when "001001000001", -- t[577] = 0
      "00" when "001001000010", -- t[578] = 0
      "00" when "001001000011", -- t[579] = 0
      "00" when "001001000100", -- t[580] = 0
      "00" when "001001000101", -- t[581] = 0
      "00" when "001001000110", -- t[582] = 0
      "00" when "001001000111", -- t[583] = 0
      "00" when "001001001000", -- t[584] = 0
      "00" when "001001001001", -- t[585] = 0
      "00" when "001001001010", -- t[586] = 0
      "00" when "001001001011", -- t[587] = 0
      "00" when "001001001100", -- t[588] = 0
      "00" when "001001001101", -- t[589] = 0
      "00" when "001001001110", -- t[590] = 0
      "00" when "001001001111", -- t[591] = 0
      "00" when "001001010000", -- t[592] = 0
      "00" when "001001010001", -- t[593] = 0
      "00" when "001001010010", -- t[594] = 0
      "00" when "001001010011", -- t[595] = 0
      "00" when "001001010100", -- t[596] = 0
      "00" when "001001010101", -- t[597] = 0
      "00" when "001001010110", -- t[598] = 0
      "00" when "001001010111", -- t[599] = 0
      "00" when "001001011000", -- t[600] = 0
      "00" when "001001011001", -- t[601] = 0
      "00" when "001001011010", -- t[602] = 0
      "00" when "001001011011", -- t[603] = 0
      "00" when "001001011100", -- t[604] = 0
      "00" when "001001011101", -- t[605] = 0
      "00" when "001001011110", -- t[606] = 0
      "00" when "001001011111", -- t[607] = 0
      "00" when "001001100000", -- t[608] = 0
      "00" when "001001100001", -- t[609] = 0
      "00" when "001001100010", -- t[610] = 0
      "00" when "001001100011", -- t[611] = 0
      "00" when "001001100100", -- t[612] = 0
      "00" when "001001100101", -- t[613] = 0
      "00" when "001001100110", -- t[614] = 0
      "00" when "001001100111", -- t[615] = 0
      "00" when "001001101000", -- t[616] = 0
      "00" when "001001101001", -- t[617] = 0
      "00" when "001001101010", -- t[618] = 0
      "00" when "001001101011", -- t[619] = 0
      "00" when "001001101100", -- t[620] = 0
      "00" when "001001101101", -- t[621] = 0
      "00" when "001001101110", -- t[622] = 0
      "00" when "001001101111", -- t[623] = 0
      "00" when "001001110000", -- t[624] = 0
      "00" when "001001110001", -- t[625] = 0
      "00" when "001001110010", -- t[626] = 0
      "00" when "001001110011", -- t[627] = 0
      "00" when "001001110100", -- t[628] = 0
      "00" when "001001110101", -- t[629] = 0
      "00" when "001001110110", -- t[630] = 0
      "00" when "001001110111", -- t[631] = 0
      "00" when "001001111000", -- t[632] = 0
      "00" when "001001111001", -- t[633] = 0
      "00" when "001001111010", -- t[634] = 0
      "00" when "001001111011", -- t[635] = 0
      "00" when "001001111100", -- t[636] = 0
      "00" when "001001111101", -- t[637] = 0
      "00" when "001001111110", -- t[638] = 0
      "00" when "001001111111", -- t[639] = 0
      "00" when "001010000000", -- t[640] = 0
      "00" when "001010000001", -- t[641] = 0
      "00" when "001010000010", -- t[642] = 0
      "00" when "001010000011", -- t[643] = 0
      "00" when "001010000100", -- t[644] = 0
      "00" when "001010000101", -- t[645] = 0
      "00" when "001010000110", -- t[646] = 0
      "00" when "001010000111", -- t[647] = 0
      "00" when "001010001000", -- t[648] = 0
      "00" when "001010001001", -- t[649] = 0
      "00" when "001010001010", -- t[650] = 0
      "00" when "001010001011", -- t[651] = 0
      "00" when "001010001100", -- t[652] = 0
      "00" when "001010001101", -- t[653] = 0
      "00" when "001010001110", -- t[654] = 0
      "00" when "001010001111", -- t[655] = 0
      "00" when "001010010000", -- t[656] = 0
      "00" when "001010010001", -- t[657] = 0
      "00" when "001010010010", -- t[658] = 0
      "00" when "001010010011", -- t[659] = 0
      "00" when "001010010100", -- t[660] = 0
      "00" when "001010010101", -- t[661] = 0
      "00" when "001010010110", -- t[662] = 0
      "00" when "001010010111", -- t[663] = 0
      "00" when "001010011000", -- t[664] = 0
      "00" when "001010011001", -- t[665] = 0
      "00" when "001010011010", -- t[666] = 0
      "00" when "001010011011", -- t[667] = 0
      "00" when "001010011100", -- t[668] = 0
      "00" when "001010011101", -- t[669] = 0
      "00" when "001010011110", -- t[670] = 0
      "00" when "001010011111", -- t[671] = 0
      "00" when "001010100000", -- t[672] = 0
      "00" when "001010100001", -- t[673] = 0
      "00" when "001010100010", -- t[674] = 0
      "00" when "001010100011", -- t[675] = 0
      "00" when "001010100100", -- t[676] = 0
      "00" when "001010100101", -- t[677] = 0
      "00" when "001010100110", -- t[678] = 0
      "00" when "001010100111", -- t[679] = 0
      "00" when "001010101000", -- t[680] = 0
      "00" when "001010101001", -- t[681] = 0
      "00" when "001010101010", -- t[682] = 0
      "00" when "001010101011", -- t[683] = 0
      "00" when "001010101100", -- t[684] = 0
      "00" when "001010101101", -- t[685] = 0
      "00" when "001010101110", -- t[686] = 0
      "00" when "001010101111", -- t[687] = 0
      "00" when "001010110000", -- t[688] = 0
      "00" when "001010110001", -- t[689] = 0
      "00" when "001010110010", -- t[690] = 0
      "00" when "001010110011", -- t[691] = 0
      "00" when "001010110100", -- t[692] = 0
      "00" when "001010110101", -- t[693] = 0
      "00" when "001010110110", -- t[694] = 0
      "00" when "001010110111", -- t[695] = 0
      "00" when "001010111000", -- t[696] = 0
      "00" when "001010111001", -- t[697] = 0
      "00" when "001010111010", -- t[698] = 0
      "00" when "001010111011", -- t[699] = 0
      "00" when "001010111100", -- t[700] = 0
      "00" when "001010111101", -- t[701] = 0
      "00" when "001010111110", -- t[702] = 0
      "00" when "001010111111", -- t[703] = 0
      "00" when "001011000000", -- t[704] = 0
      "00" when "001011000001", -- t[705] = 0
      "00" when "001011000010", -- t[706] = 0
      "00" when "001011000011", -- t[707] = 0
      "00" when "001011000100", -- t[708] = 0
      "00" when "001011000101", -- t[709] = 0
      "00" when "001011000110", -- t[710] = 0
      "00" when "001011000111", -- t[711] = 0
      "00" when "001011001000", -- t[712] = 0
      "00" when "001011001001", -- t[713] = 0
      "00" when "001011001010", -- t[714] = 0
      "00" when "001011001011", -- t[715] = 0
      "00" when "001011001100", -- t[716] = 0
      "00" when "001011001101", -- t[717] = 0
      "00" when "001011001110", -- t[718] = 0
      "00" when "001011001111", -- t[719] = 0
      "00" when "001011010000", -- t[720] = 0
      "00" when "001011010001", -- t[721] = 0
      "00" when "001011010010", -- t[722] = 0
      "00" when "001011010011", -- t[723] = 0
      "00" when "001011010100", -- t[724] = 0
      "00" when "001011010101", -- t[725] = 0
      "00" when "001011010110", -- t[726] = 0
      "00" when "001011010111", -- t[727] = 0
      "00" when "001011011000", -- t[728] = 0
      "00" when "001011011001", -- t[729] = 0
      "00" when "001011011010", -- t[730] = 0
      "00" when "001011011011", -- t[731] = 0
      "00" when "001011011100", -- t[732] = 0
      "00" when "001011011101", -- t[733] = 0
      "00" when "001011011110", -- t[734] = 0
      "00" when "001011011111", -- t[735] = 0
      "00" when "001011100000", -- t[736] = 0
      "00" when "001011100001", -- t[737] = 0
      "00" when "001011100010", -- t[738] = 0
      "00" when "001011100011", -- t[739] = 0
      "00" when "001011100100", -- t[740] = 0
      "00" when "001011100101", -- t[741] = 0
      "00" when "001011100110", -- t[742] = 0
      "00" when "001011100111", -- t[743] = 0
      "00" when "001011101000", -- t[744] = 0
      "00" when "001011101001", -- t[745] = 0
      "00" when "001011101010", -- t[746] = 0
      "00" when "001011101011", -- t[747] = 0
      "00" when "001011101100", -- t[748] = 0
      "00" when "001011101101", -- t[749] = 0
      "00" when "001011101110", -- t[750] = 0
      "00" when "001011101111", -- t[751] = 0
      "00" when "001011110000", -- t[752] = 0
      "00" when "001011110001", -- t[753] = 0
      "00" when "001011110010", -- t[754] = 0
      "00" when "001011110011", -- t[755] = 0
      "00" when "001011110100", -- t[756] = 0
      "00" when "001011110101", -- t[757] = 0
      "00" when "001011110110", -- t[758] = 0
      "00" when "001011110111", -- t[759] = 0
      "00" when "001011111000", -- t[760] = 0
      "00" when "001011111001", -- t[761] = 0
      "00" when "001011111010", -- t[762] = 0
      "00" when "001011111011", -- t[763] = 0
      "00" when "001011111100", -- t[764] = 0
      "00" when "001011111101", -- t[765] = 0
      "00" when "001011111110", -- t[766] = 0
      "00" when "001011111111", -- t[767] = 0
      "00" when "001100000000", -- t[768] = 0
      "00" when "001100000001", -- t[769] = 0
      "00" when "001100000010", -- t[770] = 0
      "00" when "001100000011", -- t[771] = 0
      "00" when "001100000100", -- t[772] = 0
      "00" when "001100000101", -- t[773] = 0
      "00" when "001100000110", -- t[774] = 0
      "00" when "001100000111", -- t[775] = 0
      "00" when "001100001000", -- t[776] = 0
      "00" when "001100001001", -- t[777] = 0
      "00" when "001100001010", -- t[778] = 0
      "00" when "001100001011", -- t[779] = 0
      "00" when "001100001100", -- t[780] = 0
      "00" when "001100001101", -- t[781] = 0
      "00" when "001100001110", -- t[782] = 0
      "00" when "001100001111", -- t[783] = 0
      "00" when "001100010000", -- t[784] = 0
      "00" when "001100010001", -- t[785] = 0
      "00" when "001100010010", -- t[786] = 0
      "00" when "001100010011", -- t[787] = 0
      "00" when "001100010100", -- t[788] = 0
      "00" when "001100010101", -- t[789] = 0
      "00" when "001100010110", -- t[790] = 0
      "00" when "001100010111", -- t[791] = 0
      "00" when "001100011000", -- t[792] = 0
      "00" when "001100011001", -- t[793] = 0
      "00" when "001100011010", -- t[794] = 0
      "00" when "001100011011", -- t[795] = 0
      "00" when "001100011100", -- t[796] = 0
      "00" when "001100011101", -- t[797] = 0
      "00" when "001100011110", -- t[798] = 0
      "00" when "001100011111", -- t[799] = 0
      "00" when "001100100000", -- t[800] = 0
      "00" when "001100100001", -- t[801] = 0
      "00" when "001100100010", -- t[802] = 0
      "00" when "001100100011", -- t[803] = 0
      "00" when "001100100100", -- t[804] = 0
      "00" when "001100100101", -- t[805] = 0
      "00" when "001100100110", -- t[806] = 0
      "00" when "001100100111", -- t[807] = 0
      "00" when "001100101000", -- t[808] = 0
      "00" when "001100101001", -- t[809] = 0
      "00" when "001100101010", -- t[810] = 0
      "00" when "001100101011", -- t[811] = 0
      "00" when "001100101100", -- t[812] = 0
      "00" when "001100101101", -- t[813] = 0
      "00" when "001100101110", -- t[814] = 0
      "00" when "001100101111", -- t[815] = 0
      "00" when "001100110000", -- t[816] = 0
      "00" when "001100110001", -- t[817] = 0
      "00" when "001100110010", -- t[818] = 0
      "00" when "001100110011", -- t[819] = 0
      "00" when "001100110100", -- t[820] = 0
      "00" when "001100110101", -- t[821] = 0
      "00" when "001100110110", -- t[822] = 0
      "00" when "001100110111", -- t[823] = 0
      "00" when "001100111000", -- t[824] = 0
      "00" when "001100111001", -- t[825] = 0
      "00" when "001100111010", -- t[826] = 0
      "00" when "001100111011", -- t[827] = 0
      "00" when "001100111100", -- t[828] = 0
      "00" when "001100111101", -- t[829] = 0
      "00" when "001100111110", -- t[830] = 0
      "00" when "001100111111", -- t[831] = 0
      "00" when "001101000000", -- t[832] = 0
      "00" when "001101000001", -- t[833] = 0
      "00" when "001101000010", -- t[834] = 0
      "00" when "001101000011", -- t[835] = 0
      "00" when "001101000100", -- t[836] = 0
      "00" when "001101000101", -- t[837] = 0
      "00" when "001101000110", -- t[838] = 0
      "00" when "001101000111", -- t[839] = 0
      "00" when "001101001000", -- t[840] = 0
      "00" when "001101001001", -- t[841] = 0
      "00" when "001101001010", -- t[842] = 0
      "00" when "001101001011", -- t[843] = 0
      "00" when "001101001100", -- t[844] = 0
      "00" when "001101001101", -- t[845] = 0
      "00" when "001101001110", -- t[846] = 0
      "00" when "001101001111", -- t[847] = 0
      "00" when "001101010000", -- t[848] = 0
      "00" when "001101010001", -- t[849] = 0
      "00" when "001101010010", -- t[850] = 0
      "00" when "001101010011", -- t[851] = 0
      "00" when "001101010100", -- t[852] = 0
      "00" when "001101010101", -- t[853] = 0
      "00" when "001101010110", -- t[854] = 0
      "00" when "001101010111", -- t[855] = 0
      "00" when "001101011000", -- t[856] = 0
      "00" when "001101011001", -- t[857] = 0
      "00" when "001101011010", -- t[858] = 0
      "00" when "001101011011", -- t[859] = 0
      "00" when "001101011100", -- t[860] = 0
      "00" when "001101011101", -- t[861] = 0
      "00" when "001101011110", -- t[862] = 0
      "00" when "001101011111", -- t[863] = 0
      "00" when "001101100000", -- t[864] = 0
      "00" when "001101100001", -- t[865] = 0
      "00" when "001101100010", -- t[866] = 0
      "00" when "001101100011", -- t[867] = 0
      "00" when "001101100100", -- t[868] = 0
      "00" when "001101100101", -- t[869] = 0
      "00" when "001101100110", -- t[870] = 0
      "00" when "001101100111", -- t[871] = 0
      "00" when "001101101000", -- t[872] = 0
      "00" when "001101101001", -- t[873] = 0
      "00" when "001101101010", -- t[874] = 0
      "00" when "001101101011", -- t[875] = 0
      "00" when "001101101100", -- t[876] = 0
      "00" when "001101101101", -- t[877] = 0
      "00" when "001101101110", -- t[878] = 0
      "00" when "001101101111", -- t[879] = 0
      "00" when "001101110000", -- t[880] = 0
      "00" when "001101110001", -- t[881] = 0
      "00" when "001101110010", -- t[882] = 0
      "00" when "001101110011", -- t[883] = 0
      "00" when "001101110100", -- t[884] = 0
      "00" when "001101110101", -- t[885] = 0
      "00" when "001101110110", -- t[886] = 0
      "00" when "001101110111", -- t[887] = 0
      "00" when "001101111000", -- t[888] = 0
      "00" when "001101111001", -- t[889] = 0
      "00" when "001101111010", -- t[890] = 0
      "00" when "001101111011", -- t[891] = 0
      "00" when "001101111100", -- t[892] = 0
      "00" when "001101111101", -- t[893] = 0
      "00" when "001101111110", -- t[894] = 0
      "00" when "001101111111", -- t[895] = 0
      "00" when "001110000000", -- t[896] = 0
      "00" when "001110000001", -- t[897] = 0
      "00" when "001110000010", -- t[898] = 0
      "00" when "001110000011", -- t[899] = 0
      "00" when "001110000100", -- t[900] = 0
      "00" when "001110000101", -- t[901] = 0
      "00" when "001110000110", -- t[902] = 0
      "00" when "001110000111", -- t[903] = 0
      "00" when "001110001000", -- t[904] = 0
      "00" when "001110001001", -- t[905] = 0
      "00" when "001110001010", -- t[906] = 0
      "00" when "001110001011", -- t[907] = 0
      "00" when "001110001100", -- t[908] = 0
      "00" when "001110001101", -- t[909] = 0
      "00" when "001110001110", -- t[910] = 0
      "00" when "001110001111", -- t[911] = 0
      "00" when "001110010000", -- t[912] = 0
      "00" when "001110010001", -- t[913] = 0
      "00" when "001110010010", -- t[914] = 0
      "00" when "001110010011", -- t[915] = 0
      "00" when "001110010100", -- t[916] = 0
      "00" when "001110010101", -- t[917] = 0
      "00" when "001110010110", -- t[918] = 0
      "00" when "001110010111", -- t[919] = 0
      "00" when "001110011000", -- t[920] = 0
      "00" when "001110011001", -- t[921] = 0
      "00" when "001110011010", -- t[922] = 0
      "00" when "001110011011", -- t[923] = 0
      "00" when "001110011100", -- t[924] = 0
      "00" when "001110011101", -- t[925] = 0
      "00" when "001110011110", -- t[926] = 0
      "00" when "001110011111", -- t[927] = 0
      "00" when "001110100000", -- t[928] = 0
      "00" when "001110100001", -- t[929] = 0
      "00" when "001110100010", -- t[930] = 0
      "00" when "001110100011", -- t[931] = 0
      "00" when "001110100100", -- t[932] = 0
      "00" when "001110100101", -- t[933] = 0
      "00" when "001110100110", -- t[934] = 0
      "00" when "001110100111", -- t[935] = 0
      "00" when "001110101000", -- t[936] = 0
      "00" when "001110101001", -- t[937] = 0
      "00" when "001110101010", -- t[938] = 0
      "00" when "001110101011", -- t[939] = 0
      "00" when "001110101100", -- t[940] = 0
      "00" when "001110101101", -- t[941] = 0
      "00" when "001110101110", -- t[942] = 0
      "00" when "001110101111", -- t[943] = 0
      "00" when "001110110000", -- t[944] = 0
      "00" when "001110110001", -- t[945] = 0
      "00" when "001110110010", -- t[946] = 0
      "00" when "001110110011", -- t[947] = 0
      "00" when "001110110100", -- t[948] = 0
      "00" when "001110110101", -- t[949] = 0
      "00" when "001110110110", -- t[950] = 0
      "00" when "001110110111", -- t[951] = 0
      "00" when "001110111000", -- t[952] = 0
      "00" when "001110111001", -- t[953] = 0
      "00" when "001110111010", -- t[954] = 0
      "00" when "001110111011", -- t[955] = 0
      "00" when "001110111100", -- t[956] = 0
      "00" when "001110111101", -- t[957] = 0
      "00" when "001110111110", -- t[958] = 0
      "00" when "001110111111", -- t[959] = 0
      "00" when "001111000000", -- t[960] = 0
      "00" when "001111000001", -- t[961] = 0
      "00" when "001111000010", -- t[962] = 0
      "00" when "001111000011", -- t[963] = 0
      "00" when "001111000100", -- t[964] = 0
      "00" when "001111000101", -- t[965] = 0
      "00" when "001111000110", -- t[966] = 0
      "00" when "001111000111", -- t[967] = 0
      "00" when "001111001000", -- t[968] = 0
      "00" when "001111001001", -- t[969] = 0
      "00" when "001111001010", -- t[970] = 0
      "00" when "001111001011", -- t[971] = 0
      "00" when "001111001100", -- t[972] = 0
      "00" when "001111001101", -- t[973] = 0
      "00" when "001111001110", -- t[974] = 0
      "00" when "001111001111", -- t[975] = 0
      "00" when "001111010000", -- t[976] = 0
      "00" when "001111010001", -- t[977] = 0
      "00" when "001111010010", -- t[978] = 0
      "00" when "001111010011", -- t[979] = 0
      "00" when "001111010100", -- t[980] = 0
      "00" when "001111010101", -- t[981] = 0
      "00" when "001111010110", -- t[982] = 0
      "00" when "001111010111", -- t[983] = 0
      "00" when "001111011000", -- t[984] = 0
      "00" when "001111011001", -- t[985] = 0
      "00" when "001111011010", -- t[986] = 0
      "00" when "001111011011", -- t[987] = 0
      "00" when "001111011100", -- t[988] = 0
      "00" when "001111011101", -- t[989] = 0
      "00" when "001111011110", -- t[990] = 0
      "00" when "001111011111", -- t[991] = 0
      "00" when "001111100000", -- t[992] = 0
      "00" when "001111100001", -- t[993] = 0
      "00" when "001111100010", -- t[994] = 0
      "00" when "001111100011", -- t[995] = 0
      "00" when "001111100100", -- t[996] = 0
      "00" when "001111100101", -- t[997] = 0
      "00" when "001111100110", -- t[998] = 0
      "00" when "001111100111", -- t[999] = 0
      "00" when "001111101000", -- t[1000] = 0
      "00" when "001111101001", -- t[1001] = 0
      "00" when "001111101010", -- t[1002] = 0
      "00" when "001111101011", -- t[1003] = 0
      "00" when "001111101100", -- t[1004] = 0
      "00" when "001111101101", -- t[1005] = 0
      "00" when "001111101110", -- t[1006] = 0
      "00" when "001111101111", -- t[1007] = 0
      "00" when "001111110000", -- t[1008] = 0
      "00" when "001111110001", -- t[1009] = 0
      "00" when "001111110010", -- t[1010] = 0
      "00" when "001111110011", -- t[1011] = 0
      "00" when "001111110100", -- t[1012] = 0
      "00" when "001111110101", -- t[1013] = 0
      "00" when "001111110110", -- t[1014] = 0
      "00" when "001111110111", -- t[1015] = 0
      "00" when "001111111000", -- t[1016] = 0
      "00" when "001111111001", -- t[1017] = 0
      "00" when "001111111010", -- t[1018] = 0
      "00" when "001111111011", -- t[1019] = 0
      "00" when "001111111100", -- t[1020] = 0
      "00" when "001111111101", -- t[1021] = 0
      "00" when "001111111110", -- t[1022] = 0
      "00" when "001111111111", -- t[1023] = 0
      "00" when "010000000000", -- t[1024] = 0
      "00" when "010000000001", -- t[1025] = 0
      "00" when "010000000010", -- t[1026] = 0
      "00" when "010000000011", -- t[1027] = 0
      "00" when "010000000100", -- t[1028] = 0
      "00" when "010000000101", -- t[1029] = 0
      "00" when "010000000110", -- t[1030] = 0
      "00" when "010000000111", -- t[1031] = 0
      "00" when "010000001000", -- t[1032] = 0
      "00" when "010000001001", -- t[1033] = 0
      "00" when "010000001010", -- t[1034] = 0
      "00" when "010000001011", -- t[1035] = 0
      "00" when "010000001100", -- t[1036] = 0
      "00" when "010000001101", -- t[1037] = 0
      "00" when "010000001110", -- t[1038] = 0
      "00" when "010000001111", -- t[1039] = 0
      "00" when "010000010000", -- t[1040] = 0
      "00" when "010000010001", -- t[1041] = 0
      "00" when "010000010010", -- t[1042] = 0
      "00" when "010000010011", -- t[1043] = 0
      "00" when "010000010100", -- t[1044] = 0
      "00" when "010000010101", -- t[1045] = 0
      "00" when "010000010110", -- t[1046] = 0
      "00" when "010000010111", -- t[1047] = 0
      "00" when "010000011000", -- t[1048] = 0
      "00" when "010000011001", -- t[1049] = 0
      "00" when "010000011010", -- t[1050] = 0
      "00" when "010000011011", -- t[1051] = 0
      "00" when "010000011100", -- t[1052] = 0
      "00" when "010000011101", -- t[1053] = 0
      "00" when "010000011110", -- t[1054] = 0
      "00" when "010000011111", -- t[1055] = 0
      "00" when "010000100000", -- t[1056] = 0
      "00" when "010000100001", -- t[1057] = 0
      "00" when "010000100010", -- t[1058] = 0
      "00" when "010000100011", -- t[1059] = 0
      "00" when "010000100100", -- t[1060] = 0
      "00" when "010000100101", -- t[1061] = 0
      "00" when "010000100110", -- t[1062] = 0
      "00" when "010000100111", -- t[1063] = 0
      "00" when "010000101000", -- t[1064] = 0
      "00" when "010000101001", -- t[1065] = 0
      "00" when "010000101010", -- t[1066] = 0
      "00" when "010000101011", -- t[1067] = 0
      "00" when "010000101100", -- t[1068] = 0
      "00" when "010000101101", -- t[1069] = 0
      "00" when "010000101110", -- t[1070] = 0
      "00" when "010000101111", -- t[1071] = 0
      "00" when "010000110000", -- t[1072] = 0
      "00" when "010000110001", -- t[1073] = 0
      "00" when "010000110010", -- t[1074] = 0
      "00" when "010000110011", -- t[1075] = 0
      "00" when "010000110100", -- t[1076] = 0
      "00" when "010000110101", -- t[1077] = 0
      "00" when "010000110110", -- t[1078] = 0
      "00" when "010000110111", -- t[1079] = 0
      "00" when "010000111000", -- t[1080] = 0
      "00" when "010000111001", -- t[1081] = 0
      "00" when "010000111010", -- t[1082] = 0
      "00" when "010000111011", -- t[1083] = 0
      "00" when "010000111100", -- t[1084] = 0
      "00" when "010000111101", -- t[1085] = 0
      "00" when "010000111110", -- t[1086] = 0
      "00" when "010000111111", -- t[1087] = 0
      "00" when "010001000000", -- t[1088] = 0
      "00" when "010001000001", -- t[1089] = 0
      "00" when "010001000010", -- t[1090] = 0
      "00" when "010001000011", -- t[1091] = 0
      "00" when "010001000100", -- t[1092] = 0
      "00" when "010001000101", -- t[1093] = 0
      "00" when "010001000110", -- t[1094] = 0
      "00" when "010001000111", -- t[1095] = 0
      "00" when "010001001000", -- t[1096] = 0
      "00" when "010001001001", -- t[1097] = 0
      "00" when "010001001010", -- t[1098] = 0
      "00" when "010001001011", -- t[1099] = 0
      "00" when "010001001100", -- t[1100] = 0
      "00" when "010001001101", -- t[1101] = 0
      "00" when "010001001110", -- t[1102] = 0
      "00" when "010001001111", -- t[1103] = 0
      "00" when "010001010000", -- t[1104] = 0
      "00" when "010001010001", -- t[1105] = 0
      "00" when "010001010010", -- t[1106] = 0
      "00" when "010001010011", -- t[1107] = 0
      "00" when "010001010100", -- t[1108] = 0
      "00" when "010001010101", -- t[1109] = 0
      "00" when "010001010110", -- t[1110] = 0
      "00" when "010001010111", -- t[1111] = 0
      "00" when "010001011000", -- t[1112] = 0
      "00" when "010001011001", -- t[1113] = 0
      "00" when "010001011010", -- t[1114] = 0
      "00" when "010001011011", -- t[1115] = 0
      "00" when "010001011100", -- t[1116] = 0
      "00" when "010001011101", -- t[1117] = 0
      "00" when "010001011110", -- t[1118] = 0
      "00" when "010001011111", -- t[1119] = 0
      "00" when "010001100000", -- t[1120] = 0
      "00" when "010001100001", -- t[1121] = 0
      "00" when "010001100010", -- t[1122] = 0
      "00" when "010001100011", -- t[1123] = 0
      "00" when "010001100100", -- t[1124] = 0
      "00" when "010001100101", -- t[1125] = 0
      "00" when "010001100110", -- t[1126] = 0
      "00" when "010001100111", -- t[1127] = 0
      "00" when "010001101000", -- t[1128] = 0
      "00" when "010001101001", -- t[1129] = 0
      "00" when "010001101010", -- t[1130] = 0
      "00" when "010001101011", -- t[1131] = 0
      "00" when "010001101100", -- t[1132] = 0
      "00" when "010001101101", -- t[1133] = 0
      "00" when "010001101110", -- t[1134] = 0
      "00" when "010001101111", -- t[1135] = 0
      "00" when "010001110000", -- t[1136] = 0
      "00" when "010001110001", -- t[1137] = 0
      "00" when "010001110010", -- t[1138] = 0
      "00" when "010001110011", -- t[1139] = 0
      "00" when "010001110100", -- t[1140] = 0
      "00" when "010001110101", -- t[1141] = 0
      "00" when "010001110110", -- t[1142] = 0
      "00" when "010001110111", -- t[1143] = 0
      "00" when "010001111000", -- t[1144] = 0
      "00" when "010001111001", -- t[1145] = 0
      "00" when "010001111010", -- t[1146] = 0
      "00" when "010001111011", -- t[1147] = 0
      "00" when "010001111100", -- t[1148] = 0
      "00" when "010001111101", -- t[1149] = 0
      "00" when "010001111110", -- t[1150] = 0
      "00" when "010001111111", -- t[1151] = 0
      "00" when "010010000000", -- t[1152] = 0
      "00" when "010010000001", -- t[1153] = 0
      "00" when "010010000010", -- t[1154] = 0
      "00" when "010010000011", -- t[1155] = 0
      "00" when "010010000100", -- t[1156] = 0
      "00" when "010010000101", -- t[1157] = 0
      "00" when "010010000110", -- t[1158] = 0
      "00" when "010010000111", -- t[1159] = 0
      "00" when "010010001000", -- t[1160] = 0
      "00" when "010010001001", -- t[1161] = 0
      "00" when "010010001010", -- t[1162] = 0
      "00" when "010010001011", -- t[1163] = 0
      "00" when "010010001100", -- t[1164] = 0
      "00" when "010010001101", -- t[1165] = 0
      "00" when "010010001110", -- t[1166] = 0
      "00" when "010010001111", -- t[1167] = 0
      "00" when "010010010000", -- t[1168] = 0
      "00" when "010010010001", -- t[1169] = 0
      "00" when "010010010010", -- t[1170] = 0
      "00" when "010010010011", -- t[1171] = 0
      "00" when "010010010100", -- t[1172] = 0
      "00" when "010010010101", -- t[1173] = 0
      "00" when "010010010110", -- t[1174] = 0
      "00" when "010010010111", -- t[1175] = 0
      "00" when "010010011000", -- t[1176] = 0
      "00" when "010010011001", -- t[1177] = 0
      "00" when "010010011010", -- t[1178] = 0
      "00" when "010010011011", -- t[1179] = 0
      "00" when "010010011100", -- t[1180] = 0
      "00" when "010010011101", -- t[1181] = 0
      "00" when "010010011110", -- t[1182] = 0
      "00" when "010010011111", -- t[1183] = 0
      "00" when "010010100000", -- t[1184] = 0
      "00" when "010010100001", -- t[1185] = 0
      "00" when "010010100010", -- t[1186] = 0
      "00" when "010010100011", -- t[1187] = 0
      "00" when "010010100100", -- t[1188] = 0
      "00" when "010010100101", -- t[1189] = 0
      "00" when "010010100110", -- t[1190] = 0
      "00" when "010010100111", -- t[1191] = 0
      "00" when "010010101000", -- t[1192] = 0
      "00" when "010010101001", -- t[1193] = 0
      "00" when "010010101010", -- t[1194] = 0
      "00" when "010010101011", -- t[1195] = 0
      "00" when "010010101100", -- t[1196] = 0
      "00" when "010010101101", -- t[1197] = 0
      "00" when "010010101110", -- t[1198] = 0
      "00" when "010010101111", -- t[1199] = 0
      "00" when "010010110000", -- t[1200] = 0
      "00" when "010010110001", -- t[1201] = 0
      "00" when "010010110010", -- t[1202] = 0
      "00" when "010010110011", -- t[1203] = 0
      "00" when "010010110100", -- t[1204] = 0
      "00" when "010010110101", -- t[1205] = 0
      "00" when "010010110110", -- t[1206] = 0
      "00" when "010010110111", -- t[1207] = 0
      "00" when "010010111000", -- t[1208] = 0
      "00" when "010010111001", -- t[1209] = 0
      "00" when "010010111010", -- t[1210] = 0
      "00" when "010010111011", -- t[1211] = 0
      "00" when "010010111100", -- t[1212] = 0
      "00" when "010010111101", -- t[1213] = 0
      "00" when "010010111110", -- t[1214] = 0
      "00" when "010010111111", -- t[1215] = 0
      "00" when "010011000000", -- t[1216] = 0
      "00" when "010011000001", -- t[1217] = 0
      "00" when "010011000010", -- t[1218] = 0
      "00" when "010011000011", -- t[1219] = 0
      "00" when "010011000100", -- t[1220] = 0
      "00" when "010011000101", -- t[1221] = 0
      "00" when "010011000110", -- t[1222] = 0
      "00" when "010011000111", -- t[1223] = 0
      "00" when "010011001000", -- t[1224] = 0
      "00" when "010011001001", -- t[1225] = 0
      "00" when "010011001010", -- t[1226] = 0
      "00" when "010011001011", -- t[1227] = 0
      "00" when "010011001100", -- t[1228] = 0
      "00" when "010011001101", -- t[1229] = 0
      "00" when "010011001110", -- t[1230] = 0
      "00" when "010011001111", -- t[1231] = 0
      "00" when "010011010000", -- t[1232] = 0
      "00" when "010011010001", -- t[1233] = 0
      "00" when "010011010010", -- t[1234] = 0
      "00" when "010011010011", -- t[1235] = 0
      "00" when "010011010100", -- t[1236] = 0
      "00" when "010011010101", -- t[1237] = 0
      "00" when "010011010110", -- t[1238] = 0
      "00" when "010011010111", -- t[1239] = 0
      "00" when "010011011000", -- t[1240] = 0
      "00" when "010011011001", -- t[1241] = 0
      "00" when "010011011010", -- t[1242] = 0
      "00" when "010011011011", -- t[1243] = 0
      "00" when "010011011100", -- t[1244] = 0
      "00" when "010011011101", -- t[1245] = 0
      "00" when "010011011110", -- t[1246] = 0
      "00" when "010011011111", -- t[1247] = 0
      "00" when "010011100000", -- t[1248] = 0
      "00" when "010011100001", -- t[1249] = 0
      "00" when "010011100010", -- t[1250] = 0
      "00" when "010011100011", -- t[1251] = 0
      "00" when "010011100100", -- t[1252] = 0
      "00" when "010011100101", -- t[1253] = 0
      "00" when "010011100110", -- t[1254] = 0
      "00" when "010011100111", -- t[1255] = 0
      "00" when "010011101000", -- t[1256] = 0
      "00" when "010011101001", -- t[1257] = 0
      "00" when "010011101010", -- t[1258] = 0
      "00" when "010011101011", -- t[1259] = 0
      "00" when "010011101100", -- t[1260] = 0
      "00" when "010011101101", -- t[1261] = 0
      "00" when "010011101110", -- t[1262] = 0
      "00" when "010011101111", -- t[1263] = 0
      "00" when "010011110000", -- t[1264] = 0
      "00" when "010011110001", -- t[1265] = 0
      "00" when "010011110010", -- t[1266] = 0
      "00" when "010011110011", -- t[1267] = 0
      "00" when "010011110100", -- t[1268] = 0
      "00" when "010011110101", -- t[1269] = 0
      "00" when "010011110110", -- t[1270] = 0
      "00" when "010011110111", -- t[1271] = 0
      "00" when "010011111000", -- t[1272] = 0
      "00" when "010011111001", -- t[1273] = 0
      "00" when "010011111010", -- t[1274] = 0
      "00" when "010011111011", -- t[1275] = 0
      "00" when "010011111100", -- t[1276] = 0
      "00" when "010011111101", -- t[1277] = 0
      "00" when "010011111110", -- t[1278] = 0
      "00" when "010011111111", -- t[1279] = 0
      "00" when "010100000000", -- t[1280] = 0
      "00" when "010100000001", -- t[1281] = 0
      "00" when "010100000010", -- t[1282] = 0
      "00" when "010100000011", -- t[1283] = 0
      "00" when "010100000100", -- t[1284] = 0
      "00" when "010100000101", -- t[1285] = 0
      "00" when "010100000110", -- t[1286] = 0
      "00" when "010100000111", -- t[1287] = 0
      "00" when "010100001000", -- t[1288] = 0
      "00" when "010100001001", -- t[1289] = 0
      "00" when "010100001010", -- t[1290] = 0
      "00" when "010100001011", -- t[1291] = 0
      "00" when "010100001100", -- t[1292] = 0
      "00" when "010100001101", -- t[1293] = 0
      "00" when "010100001110", -- t[1294] = 0
      "00" when "010100001111", -- t[1295] = 0
      "00" when "010100010000", -- t[1296] = 0
      "00" when "010100010001", -- t[1297] = 0
      "00" when "010100010010", -- t[1298] = 0
      "00" when "010100010011", -- t[1299] = 0
      "00" when "010100010100", -- t[1300] = 0
      "00" when "010100010101", -- t[1301] = 0
      "00" when "010100010110", -- t[1302] = 0
      "00" when "010100010111", -- t[1303] = 0
      "00" when "010100011000", -- t[1304] = 0
      "00" when "010100011001", -- t[1305] = 0
      "00" when "010100011010", -- t[1306] = 0
      "00" when "010100011011", -- t[1307] = 0
      "00" when "010100011100", -- t[1308] = 0
      "00" when "010100011101", -- t[1309] = 0
      "00" when "010100011110", -- t[1310] = 0
      "00" when "010100011111", -- t[1311] = 0
      "00" when "010100100000", -- t[1312] = 0
      "00" when "010100100001", -- t[1313] = 0
      "00" when "010100100010", -- t[1314] = 0
      "00" when "010100100011", -- t[1315] = 0
      "00" when "010100100100", -- t[1316] = 0
      "00" when "010100100101", -- t[1317] = 0
      "00" when "010100100110", -- t[1318] = 0
      "00" when "010100100111", -- t[1319] = 0
      "00" when "010100101000", -- t[1320] = 0
      "00" when "010100101001", -- t[1321] = 0
      "00" when "010100101010", -- t[1322] = 0
      "00" when "010100101011", -- t[1323] = 0
      "00" when "010100101100", -- t[1324] = 0
      "00" when "010100101101", -- t[1325] = 0
      "00" when "010100101110", -- t[1326] = 0
      "00" when "010100101111", -- t[1327] = 0
      "00" when "010100110000", -- t[1328] = 0
      "00" when "010100110001", -- t[1329] = 0
      "00" when "010100110010", -- t[1330] = 0
      "00" when "010100110011", -- t[1331] = 0
      "00" when "010100110100", -- t[1332] = 0
      "00" when "010100110101", -- t[1333] = 0
      "00" when "010100110110", -- t[1334] = 0
      "00" when "010100110111", -- t[1335] = 0
      "00" when "010100111000", -- t[1336] = 0
      "00" when "010100111001", -- t[1337] = 0
      "00" when "010100111010", -- t[1338] = 0
      "00" when "010100111011", -- t[1339] = 0
      "00" when "010100111100", -- t[1340] = 0
      "00" when "010100111101", -- t[1341] = 0
      "00" when "010100111110", -- t[1342] = 0
      "00" when "010100111111", -- t[1343] = 0
      "00" when "010101000000", -- t[1344] = 0
      "00" when "010101000001", -- t[1345] = 0
      "00" when "010101000010", -- t[1346] = 0
      "00" when "010101000011", -- t[1347] = 0
      "00" when "010101000100", -- t[1348] = 0
      "00" when "010101000101", -- t[1349] = 0
      "00" when "010101000110", -- t[1350] = 0
      "00" when "010101000111", -- t[1351] = 0
      "00" when "010101001000", -- t[1352] = 0
      "00" when "010101001001", -- t[1353] = 0
      "00" when "010101001010", -- t[1354] = 0
      "00" when "010101001011", -- t[1355] = 0
      "00" when "010101001100", -- t[1356] = 0
      "00" when "010101001101", -- t[1357] = 0
      "00" when "010101001110", -- t[1358] = 0
      "00" when "010101001111", -- t[1359] = 0
      "00" when "010101010000", -- t[1360] = 0
      "00" when "010101010001", -- t[1361] = 0
      "00" when "010101010010", -- t[1362] = 0
      "00" when "010101010011", -- t[1363] = 0
      "00" when "010101010100", -- t[1364] = 0
      "00" when "010101010101", -- t[1365] = 0
      "00" when "010101010110", -- t[1366] = 0
      "00" when "010101010111", -- t[1367] = 0
      "00" when "010101011000", -- t[1368] = 0
      "00" when "010101011001", -- t[1369] = 0
      "00" when "010101011010", -- t[1370] = 0
      "00" when "010101011011", -- t[1371] = 0
      "00" when "010101011100", -- t[1372] = 0
      "00" when "010101011101", -- t[1373] = 0
      "00" when "010101011110", -- t[1374] = 0
      "00" when "010101011111", -- t[1375] = 0
      "00" when "010101100000", -- t[1376] = 0
      "00" when "010101100001", -- t[1377] = 0
      "00" when "010101100010", -- t[1378] = 0
      "00" when "010101100011", -- t[1379] = 0
      "00" when "010101100100", -- t[1380] = 0
      "00" when "010101100101", -- t[1381] = 0
      "00" when "010101100110", -- t[1382] = 0
      "00" when "010101100111", -- t[1383] = 0
      "00" when "010101101000", -- t[1384] = 0
      "00" when "010101101001", -- t[1385] = 0
      "00" when "010101101010", -- t[1386] = 0
      "00" when "010101101011", -- t[1387] = 0
      "00" when "010101101100", -- t[1388] = 0
      "00" when "010101101101", -- t[1389] = 0
      "00" when "010101101110", -- t[1390] = 0
      "00" when "010101101111", -- t[1391] = 0
      "00" when "010101110000", -- t[1392] = 0
      "00" when "010101110001", -- t[1393] = 0
      "00" when "010101110010", -- t[1394] = 0
      "00" when "010101110011", -- t[1395] = 0
      "00" when "010101110100", -- t[1396] = 0
      "00" when "010101110101", -- t[1397] = 0
      "00" when "010101110110", -- t[1398] = 0
      "00" when "010101110111", -- t[1399] = 0
      "00" when "010101111000", -- t[1400] = 0
      "00" when "010101111001", -- t[1401] = 0
      "00" when "010101111010", -- t[1402] = 0
      "00" when "010101111011", -- t[1403] = 0
      "00" when "010101111100", -- t[1404] = 0
      "00" when "010101111101", -- t[1405] = 0
      "00" when "010101111110", -- t[1406] = 0
      "00" when "010101111111", -- t[1407] = 0
      "00" when "010110000000", -- t[1408] = 0
      "00" when "010110000001", -- t[1409] = 0
      "00" when "010110000010", -- t[1410] = 0
      "00" when "010110000011", -- t[1411] = 0
      "00" when "010110000100", -- t[1412] = 0
      "00" when "010110000101", -- t[1413] = 0
      "00" when "010110000110", -- t[1414] = 0
      "00" when "010110000111", -- t[1415] = 0
      "00" when "010110001000", -- t[1416] = 0
      "00" when "010110001001", -- t[1417] = 0
      "00" when "010110001010", -- t[1418] = 0
      "00" when "010110001011", -- t[1419] = 0
      "00" when "010110001100", -- t[1420] = 0
      "00" when "010110001101", -- t[1421] = 0
      "00" when "010110001110", -- t[1422] = 0
      "00" when "010110001111", -- t[1423] = 0
      "00" when "010110010000", -- t[1424] = 0
      "00" when "010110010001", -- t[1425] = 0
      "00" when "010110010010", -- t[1426] = 0
      "00" when "010110010011", -- t[1427] = 0
      "00" when "010110010100", -- t[1428] = 0
      "00" when "010110010101", -- t[1429] = 0
      "00" when "010110010110", -- t[1430] = 0
      "00" when "010110010111", -- t[1431] = 0
      "00" when "010110011000", -- t[1432] = 0
      "00" when "010110011001", -- t[1433] = 0
      "00" when "010110011010", -- t[1434] = 0
      "00" when "010110011011", -- t[1435] = 0
      "00" when "010110011100", -- t[1436] = 0
      "00" when "010110011101", -- t[1437] = 0
      "00" when "010110011110", -- t[1438] = 0
      "00" when "010110011111", -- t[1439] = 0
      "00" when "010110100000", -- t[1440] = 0
      "00" when "010110100001", -- t[1441] = 0
      "00" when "010110100010", -- t[1442] = 0
      "00" when "010110100011", -- t[1443] = 0
      "00" when "010110100100", -- t[1444] = 0
      "00" when "010110100101", -- t[1445] = 0
      "00" when "010110100110", -- t[1446] = 0
      "00" when "010110100111", -- t[1447] = 0
      "00" when "010110101000", -- t[1448] = 0
      "00" when "010110101001", -- t[1449] = 0
      "00" when "010110101010", -- t[1450] = 0
      "00" when "010110101011", -- t[1451] = 0
      "00" when "010110101100", -- t[1452] = 0
      "00" when "010110101101", -- t[1453] = 0
      "00" when "010110101110", -- t[1454] = 0
      "00" when "010110101111", -- t[1455] = 0
      "00" when "010110110000", -- t[1456] = 0
      "00" when "010110110001", -- t[1457] = 0
      "00" when "010110110010", -- t[1458] = 0
      "00" when "010110110011", -- t[1459] = 0
      "00" when "010110110100", -- t[1460] = 0
      "00" when "010110110101", -- t[1461] = 0
      "00" when "010110110110", -- t[1462] = 0
      "00" when "010110110111", -- t[1463] = 0
      "00" when "010110111000", -- t[1464] = 0
      "00" when "010110111001", -- t[1465] = 0
      "00" when "010110111010", -- t[1466] = 0
      "00" when "010110111011", -- t[1467] = 0
      "00" when "010110111100", -- t[1468] = 0
      "00" when "010110111101", -- t[1469] = 0
      "00" when "010110111110", -- t[1470] = 0
      "00" when "010110111111", -- t[1471] = 0
      "00" when "010111000000", -- t[1472] = 0
      "00" when "010111000001", -- t[1473] = 0
      "00" when "010111000010", -- t[1474] = 0
      "00" when "010111000011", -- t[1475] = 0
      "00" when "010111000100", -- t[1476] = 0
      "00" when "010111000101", -- t[1477] = 0
      "00" when "010111000110", -- t[1478] = 0
      "00" when "010111000111", -- t[1479] = 0
      "00" when "010111001000", -- t[1480] = 0
      "00" when "010111001001", -- t[1481] = 0
      "00" when "010111001010", -- t[1482] = 0
      "00" when "010111001011", -- t[1483] = 0
      "00" when "010111001100", -- t[1484] = 0
      "00" when "010111001101", -- t[1485] = 0
      "00" when "010111001110", -- t[1486] = 0
      "00" when "010111001111", -- t[1487] = 0
      "00" when "010111010000", -- t[1488] = 0
      "00" when "010111010001", -- t[1489] = 0
      "00" when "010111010010", -- t[1490] = 0
      "00" when "010111010011", -- t[1491] = 0
      "00" when "010111010100", -- t[1492] = 0
      "00" when "010111010101", -- t[1493] = 0
      "00" when "010111010110", -- t[1494] = 0
      "00" when "010111010111", -- t[1495] = 0
      "00" when "010111011000", -- t[1496] = 0
      "00" when "010111011001", -- t[1497] = 0
      "00" when "010111011010", -- t[1498] = 0
      "00" when "010111011011", -- t[1499] = 0
      "00" when "010111011100", -- t[1500] = 0
      "00" when "010111011101", -- t[1501] = 0
      "00" when "010111011110", -- t[1502] = 0
      "00" when "010111011111", -- t[1503] = 0
      "00" when "010111100000", -- t[1504] = 0
      "00" when "010111100001", -- t[1505] = 0
      "00" when "010111100010", -- t[1506] = 0
      "00" when "010111100011", -- t[1507] = 0
      "00" when "010111100100", -- t[1508] = 0
      "00" when "010111100101", -- t[1509] = 0
      "00" when "010111100110", -- t[1510] = 0
      "00" when "010111100111", -- t[1511] = 0
      "00" when "010111101000", -- t[1512] = 0
      "00" when "010111101001", -- t[1513] = 0
      "00" when "010111101010", -- t[1514] = 0
      "00" when "010111101011", -- t[1515] = 0
      "00" when "010111101100", -- t[1516] = 0
      "00" when "010111101101", -- t[1517] = 0
      "00" when "010111101110", -- t[1518] = 0
      "00" when "010111101111", -- t[1519] = 0
      "00" when "010111110000", -- t[1520] = 0
      "00" when "010111110001", -- t[1521] = 0
      "00" when "010111110010", -- t[1522] = 0
      "00" when "010111110011", -- t[1523] = 0
      "00" when "010111110100", -- t[1524] = 0
      "00" when "010111110101", -- t[1525] = 0
      "00" when "010111110110", -- t[1526] = 0
      "00" when "010111110111", -- t[1527] = 0
      "00" when "010111111000", -- t[1528] = 0
      "00" when "010111111001", -- t[1529] = 0
      "00" when "010111111010", -- t[1530] = 0
      "00" when "010111111011", -- t[1531] = 0
      "00" when "010111111100", -- t[1532] = 0
      "00" when "010111111101", -- t[1533] = 0
      "00" when "010111111110", -- t[1534] = 0
      "00" when "010111111111", -- t[1535] = 0
      "00" when "011000000000", -- t[1536] = 0
      "00" when "011000000001", -- t[1537] = 0
      "00" when "011000000010", -- t[1538] = 0
      "00" when "011000000011", -- t[1539] = 0
      "00" when "011000000100", -- t[1540] = 0
      "00" when "011000000101", -- t[1541] = 0
      "00" when "011000000110", -- t[1542] = 0
      "00" when "011000000111", -- t[1543] = 0
      "00" when "011000001000", -- t[1544] = 0
      "00" when "011000001001", -- t[1545] = 0
      "00" when "011000001010", -- t[1546] = 0
      "00" when "011000001011", -- t[1547] = 0
      "00" when "011000001100", -- t[1548] = 0
      "00" when "011000001101", -- t[1549] = 0
      "00" when "011000001110", -- t[1550] = 0
      "00" when "011000001111", -- t[1551] = 0
      "00" when "011000010000", -- t[1552] = 0
      "00" when "011000010001", -- t[1553] = 0
      "00" when "011000010010", -- t[1554] = 0
      "00" when "011000010011", -- t[1555] = 0
      "00" when "011000010100", -- t[1556] = 0
      "00" when "011000010101", -- t[1557] = 0
      "00" when "011000010110", -- t[1558] = 0
      "00" when "011000010111", -- t[1559] = 0
      "00" when "011000011000", -- t[1560] = 0
      "00" when "011000011001", -- t[1561] = 0
      "00" when "011000011010", -- t[1562] = 0
      "00" when "011000011011", -- t[1563] = 0
      "00" when "011000011100", -- t[1564] = 0
      "00" when "011000011101", -- t[1565] = 0
      "00" when "011000011110", -- t[1566] = 0
      "00" when "011000011111", -- t[1567] = 0
      "00" when "011000100000", -- t[1568] = 0
      "00" when "011000100001", -- t[1569] = 0
      "00" when "011000100010", -- t[1570] = 0
      "00" when "011000100011", -- t[1571] = 0
      "00" when "011000100100", -- t[1572] = 0
      "00" when "011000100101", -- t[1573] = 0
      "00" when "011000100110", -- t[1574] = 0
      "00" when "011000100111", -- t[1575] = 0
      "00" when "011000101000", -- t[1576] = 0
      "00" when "011000101001", -- t[1577] = 0
      "00" when "011000101010", -- t[1578] = 0
      "00" when "011000101011", -- t[1579] = 0
      "00" when "011000101100", -- t[1580] = 0
      "00" when "011000101101", -- t[1581] = 0
      "00" when "011000101110", -- t[1582] = 0
      "00" when "011000101111", -- t[1583] = 0
      "00" when "011000110000", -- t[1584] = 0
      "00" when "011000110001", -- t[1585] = 0
      "00" when "011000110010", -- t[1586] = 0
      "00" when "011000110011", -- t[1587] = 0
      "00" when "011000110100", -- t[1588] = 0
      "00" when "011000110101", -- t[1589] = 0
      "00" when "011000110110", -- t[1590] = 0
      "00" when "011000110111", -- t[1591] = 0
      "00" when "011000111000", -- t[1592] = 0
      "00" when "011000111001", -- t[1593] = 0
      "00" when "011000111010", -- t[1594] = 0
      "00" when "011000111011", -- t[1595] = 0
      "00" when "011000111100", -- t[1596] = 0
      "00" when "011000111101", -- t[1597] = 0
      "00" when "011000111110", -- t[1598] = 0
      "00" when "011000111111", -- t[1599] = 0
      "00" when "011001000000", -- t[1600] = 0
      "00" when "011001000001", -- t[1601] = 0
      "00" when "011001000010", -- t[1602] = 0
      "00" when "011001000011", -- t[1603] = 0
      "00" when "011001000100", -- t[1604] = 0
      "00" when "011001000101", -- t[1605] = 0
      "00" when "011001000110", -- t[1606] = 0
      "00" when "011001000111", -- t[1607] = 0
      "00" when "011001001000", -- t[1608] = 0
      "00" when "011001001001", -- t[1609] = 0
      "00" when "011001001010", -- t[1610] = 0
      "00" when "011001001011", -- t[1611] = 0
      "00" when "011001001100", -- t[1612] = 0
      "00" when "011001001101", -- t[1613] = 0
      "00" when "011001001110", -- t[1614] = 0
      "00" when "011001001111", -- t[1615] = 0
      "00" when "011001010000", -- t[1616] = 0
      "00" when "011001010001", -- t[1617] = 0
      "00" when "011001010010", -- t[1618] = 0
      "00" when "011001010011", -- t[1619] = 0
      "00" when "011001010100", -- t[1620] = 0
      "00" when "011001010101", -- t[1621] = 0
      "00" when "011001010110", -- t[1622] = 0
      "00" when "011001010111", -- t[1623] = 0
      "00" when "011001011000", -- t[1624] = 0
      "00" when "011001011001", -- t[1625] = 0
      "00" when "011001011010", -- t[1626] = 0
      "00" when "011001011011", -- t[1627] = 0
      "00" when "011001011100", -- t[1628] = 0
      "00" when "011001011101", -- t[1629] = 0
      "00" when "011001011110", -- t[1630] = 0
      "00" when "011001011111", -- t[1631] = 0
      "00" when "011001100000", -- t[1632] = 0
      "00" when "011001100001", -- t[1633] = 0
      "00" when "011001100010", -- t[1634] = 0
      "00" when "011001100011", -- t[1635] = 0
      "00" when "011001100100", -- t[1636] = 0
      "00" when "011001100101", -- t[1637] = 0
      "00" when "011001100110", -- t[1638] = 0
      "00" when "011001100111", -- t[1639] = 0
      "00" when "011001101000", -- t[1640] = 0
      "00" when "011001101001", -- t[1641] = 0
      "00" when "011001101010", -- t[1642] = 0
      "00" when "011001101011", -- t[1643] = 0
      "00" when "011001101100", -- t[1644] = 0
      "00" when "011001101101", -- t[1645] = 0
      "00" when "011001101110", -- t[1646] = 0
      "00" when "011001101111", -- t[1647] = 0
      "00" when "011001110000", -- t[1648] = 0
      "00" when "011001110001", -- t[1649] = 0
      "00" when "011001110010", -- t[1650] = 0
      "00" when "011001110011", -- t[1651] = 0
      "00" when "011001110100", -- t[1652] = 0
      "00" when "011001110101", -- t[1653] = 0
      "00" when "011001110110", -- t[1654] = 0
      "00" when "011001110111", -- t[1655] = 0
      "00" when "011001111000", -- t[1656] = 0
      "01" when "011001111001", -- t[1657] = 1
      "01" when "011001111010", -- t[1658] = 1
      "01" when "011001111011", -- t[1659] = 1
      "01" when "011001111100", -- t[1660] = 1
      "01" when "011001111101", -- t[1661] = 1
      "01" when "011001111110", -- t[1662] = 1
      "01" when "011001111111", -- t[1663] = 1
      "01" when "011010000000", -- t[1664] = 1
      "01" when "011010000001", -- t[1665] = 1
      "01" when "011010000010", -- t[1666] = 1
      "01" when "011010000011", -- t[1667] = 1
      "01" when "011010000100", -- t[1668] = 1
      "01" when "011010000101", -- t[1669] = 1
      "01" when "011010000110", -- t[1670] = 1
      "01" when "011010000111", -- t[1671] = 1
      "01" when "011010001000", -- t[1672] = 1
      "01" when "011010001001", -- t[1673] = 1
      "01" when "011010001010", -- t[1674] = 1
      "01" when "011010001011", -- t[1675] = 1
      "01" when "011010001100", -- t[1676] = 1
      "01" when "011010001101", -- t[1677] = 1
      "01" when "011010001110", -- t[1678] = 1
      "01" when "011010001111", -- t[1679] = 1
      "01" when "011010010000", -- t[1680] = 1
      "01" when "011010010001", -- t[1681] = 1
      "01" when "011010010010", -- t[1682] = 1
      "01" when "011010010011", -- t[1683] = 1
      "01" when "011010010100", -- t[1684] = 1
      "01" when "011010010101", -- t[1685] = 1
      "01" when "011010010110", -- t[1686] = 1
      "01" when "011010010111", -- t[1687] = 1
      "01" when "011010011000", -- t[1688] = 1
      "01" when "011010011001", -- t[1689] = 1
      "01" when "011010011010", -- t[1690] = 1
      "01" when "011010011011", -- t[1691] = 1
      "01" when "011010011100", -- t[1692] = 1
      "01" when "011010011101", -- t[1693] = 1
      "01" when "011010011110", -- t[1694] = 1
      "01" when "011010011111", -- t[1695] = 1
      "01" when "011010100000", -- t[1696] = 1
      "01" when "011010100001", -- t[1697] = 1
      "01" when "011010100010", -- t[1698] = 1
      "01" when "011010100011", -- t[1699] = 1
      "01" when "011010100100", -- t[1700] = 1
      "01" when "011010100101", -- t[1701] = 1
      "01" when "011010100110", -- t[1702] = 1
      "01" when "011010100111", -- t[1703] = 1
      "01" when "011010101000", -- t[1704] = 1
      "01" when "011010101001", -- t[1705] = 1
      "01" when "011010101010", -- t[1706] = 1
      "01" when "011010101011", -- t[1707] = 1
      "01" when "011010101100", -- t[1708] = 1
      "01" when "011010101101", -- t[1709] = 1
      "01" when "011010101110", -- t[1710] = 1
      "01" when "011010101111", -- t[1711] = 1
      "01" when "011010110000", -- t[1712] = 1
      "01" when "011010110001", -- t[1713] = 1
      "01" when "011010110010", -- t[1714] = 1
      "01" when "011010110011", -- t[1715] = 1
      "01" when "011010110100", -- t[1716] = 1
      "01" when "011010110101", -- t[1717] = 1
      "01" when "011010110110", -- t[1718] = 1
      "01" when "011010110111", -- t[1719] = 1
      "01" when "011010111000", -- t[1720] = 1
      "01" when "011010111001", -- t[1721] = 1
      "01" when "011010111010", -- t[1722] = 1
      "01" when "011010111011", -- t[1723] = 1
      "01" when "011010111100", -- t[1724] = 1
      "01" when "011010111101", -- t[1725] = 1
      "01" when "011010111110", -- t[1726] = 1
      "01" when "011010111111", -- t[1727] = 1
      "01" when "011011000000", -- t[1728] = 1
      "01" when "011011000001", -- t[1729] = 1
      "01" when "011011000010", -- t[1730] = 1
      "01" when "011011000011", -- t[1731] = 1
      "01" when "011011000100", -- t[1732] = 1
      "01" when "011011000101", -- t[1733] = 1
      "01" when "011011000110", -- t[1734] = 1
      "01" when "011011000111", -- t[1735] = 1
      "01" when "011011001000", -- t[1736] = 1
      "01" when "011011001001", -- t[1737] = 1
      "01" when "011011001010", -- t[1738] = 1
      "01" when "011011001011", -- t[1739] = 1
      "01" when "011011001100", -- t[1740] = 1
      "01" when "011011001101", -- t[1741] = 1
      "01" when "011011001110", -- t[1742] = 1
      "01" when "011011001111", -- t[1743] = 1
      "01" when "011011010000", -- t[1744] = 1
      "01" when "011011010001", -- t[1745] = 1
      "01" when "011011010010", -- t[1746] = 1
      "01" when "011011010011", -- t[1747] = 1
      "01" when "011011010100", -- t[1748] = 1
      "01" when "011011010101", -- t[1749] = 1
      "01" when "011011010110", -- t[1750] = 1
      "01" when "011011010111", -- t[1751] = 1
      "01" when "011011011000", -- t[1752] = 1
      "01" when "011011011001", -- t[1753] = 1
      "01" when "011011011010", -- t[1754] = 1
      "01" when "011011011011", -- t[1755] = 1
      "01" when "011011011100", -- t[1756] = 1
      "01" when "011011011101", -- t[1757] = 1
      "01" when "011011011110", -- t[1758] = 1
      "01" when "011011011111", -- t[1759] = 1
      "01" when "011011100000", -- t[1760] = 1
      "01" when "011011100001", -- t[1761] = 1
      "01" when "011011100010", -- t[1762] = 1
      "01" when "011011100011", -- t[1763] = 1
      "01" when "011011100100", -- t[1764] = 1
      "01" when "011011100101", -- t[1765] = 1
      "01" when "011011100110", -- t[1766] = 1
      "01" when "011011100111", -- t[1767] = 1
      "01" when "011011101000", -- t[1768] = 1
      "01" when "011011101001", -- t[1769] = 1
      "01" when "011011101010", -- t[1770] = 1
      "01" when "011011101011", -- t[1771] = 1
      "01" when "011011101100", -- t[1772] = 1
      "01" when "011011101101", -- t[1773] = 1
      "01" when "011011101110", -- t[1774] = 1
      "01" when "011011101111", -- t[1775] = 1
      "01" when "011011110000", -- t[1776] = 1
      "01" when "011011110001", -- t[1777] = 1
      "01" when "011011110010", -- t[1778] = 1
      "01" when "011011110011", -- t[1779] = 1
      "01" when "011011110100", -- t[1780] = 1
      "01" when "011011110101", -- t[1781] = 1
      "01" when "011011110110", -- t[1782] = 1
      "01" when "011011110111", -- t[1783] = 1
      "01" when "011011111000", -- t[1784] = 1
      "01" when "011011111001", -- t[1785] = 1
      "01" when "011011111010", -- t[1786] = 1
      "01" when "011011111011", -- t[1787] = 1
      "01" when "011011111100", -- t[1788] = 1
      "01" when "011011111101", -- t[1789] = 1
      "01" when "011011111110", -- t[1790] = 1
      "01" when "011011111111", -- t[1791] = 1
      "01" when "011100000000", -- t[1792] = 1
      "01" when "011100000001", -- t[1793] = 1
      "01" when "011100000010", -- t[1794] = 1
      "01" when "011100000011", -- t[1795] = 1
      "01" when "011100000100", -- t[1796] = 1
      "01" when "011100000101", -- t[1797] = 1
      "01" when "011100000110", -- t[1798] = 1
      "01" when "011100000111", -- t[1799] = 1
      "01" when "011100001000", -- t[1800] = 1
      "01" when "011100001001", -- t[1801] = 1
      "01" when "011100001010", -- t[1802] = 1
      "01" when "011100001011", -- t[1803] = 1
      "01" when "011100001100", -- t[1804] = 1
      "01" when "011100001101", -- t[1805] = 1
      "01" when "011100001110", -- t[1806] = 1
      "01" when "011100001111", -- t[1807] = 1
      "01" when "011100010000", -- t[1808] = 1
      "01" when "011100010001", -- t[1809] = 1
      "01" when "011100010010", -- t[1810] = 1
      "01" when "011100010011", -- t[1811] = 1
      "01" when "011100010100", -- t[1812] = 1
      "01" when "011100010101", -- t[1813] = 1
      "01" when "011100010110", -- t[1814] = 1
      "01" when "011100010111", -- t[1815] = 1
      "01" when "011100011000", -- t[1816] = 1
      "01" when "011100011001", -- t[1817] = 1
      "01" when "011100011010", -- t[1818] = 1
      "01" when "011100011011", -- t[1819] = 1
      "01" when "011100011100", -- t[1820] = 1
      "01" when "011100011101", -- t[1821] = 1
      "01" when "011100011110", -- t[1822] = 1
      "01" when "011100011111", -- t[1823] = 1
      "01" when "011100100000", -- t[1824] = 1
      "01" when "011100100001", -- t[1825] = 1
      "01" when "011100100010", -- t[1826] = 1
      "01" when "011100100011", -- t[1827] = 1
      "01" when "011100100100", -- t[1828] = 1
      "01" when "011100100101", -- t[1829] = 1
      "01" when "011100100110", -- t[1830] = 1
      "01" when "011100100111", -- t[1831] = 1
      "01" when "011100101000", -- t[1832] = 1
      "01" when "011100101001", -- t[1833] = 1
      "01" when "011100101010", -- t[1834] = 1
      "01" when "011100101011", -- t[1835] = 1
      "01" when "011100101100", -- t[1836] = 1
      "01" when "011100101101", -- t[1837] = 1
      "01" when "011100101110", -- t[1838] = 1
      "01" when "011100101111", -- t[1839] = 1
      "01" when "011100110000", -- t[1840] = 1
      "01" when "011100110001", -- t[1841] = 1
      "01" when "011100110010", -- t[1842] = 1
      "01" when "011100110011", -- t[1843] = 1
      "01" when "011100110100", -- t[1844] = 1
      "01" when "011100110101", -- t[1845] = 1
      "01" when "011100110110", -- t[1846] = 1
      "01" when "011100110111", -- t[1847] = 1
      "01" when "011100111000", -- t[1848] = 1
      "01" when "011100111001", -- t[1849] = 1
      "01" when "011100111010", -- t[1850] = 1
      "01" when "011100111011", -- t[1851] = 1
      "01" when "011100111100", -- t[1852] = 1
      "01" when "011100111101", -- t[1853] = 1
      "01" when "011100111110", -- t[1854] = 1
      "01" when "011100111111", -- t[1855] = 1
      "01" when "011101000000", -- t[1856] = 1
      "01" when "011101000001", -- t[1857] = 1
      "01" when "011101000010", -- t[1858] = 1
      "01" when "011101000011", -- t[1859] = 1
      "01" when "011101000100", -- t[1860] = 1
      "01" when "011101000101", -- t[1861] = 1
      "01" when "011101000110", -- t[1862] = 1
      "01" when "011101000111", -- t[1863] = 1
      "01" when "011101001000", -- t[1864] = 1
      "01" when "011101001001", -- t[1865] = 1
      "01" when "011101001010", -- t[1866] = 1
      "01" when "011101001011", -- t[1867] = 1
      "01" when "011101001100", -- t[1868] = 1
      "01" when "011101001101", -- t[1869] = 1
      "01" when "011101001110", -- t[1870] = 1
      "01" when "011101001111", -- t[1871] = 1
      "01" when "011101010000", -- t[1872] = 1
      "01" when "011101010001", -- t[1873] = 1
      "01" when "011101010010", -- t[1874] = 1
      "01" when "011101010011", -- t[1875] = 1
      "01" when "011101010100", -- t[1876] = 1
      "01" when "011101010101", -- t[1877] = 1
      "01" when "011101010110", -- t[1878] = 1
      "01" when "011101010111", -- t[1879] = 1
      "01" when "011101011000", -- t[1880] = 1
      "01" when "011101011001", -- t[1881] = 1
      "01" when "011101011010", -- t[1882] = 1
      "01" when "011101011011", -- t[1883] = 1
      "01" when "011101011100", -- t[1884] = 1
      "01" when "011101011101", -- t[1885] = 1
      "01" when "011101011110", -- t[1886] = 1
      "01" when "011101011111", -- t[1887] = 1
      "01" when "011101100000", -- t[1888] = 1
      "01" when "011101100001", -- t[1889] = 1
      "01" when "011101100010", -- t[1890] = 1
      "01" when "011101100011", -- t[1891] = 1
      "01" when "011101100100", -- t[1892] = 1
      "01" when "011101100101", -- t[1893] = 1
      "01" when "011101100110", -- t[1894] = 1
      "01" when "011101100111", -- t[1895] = 1
      "01" when "011101101000", -- t[1896] = 1
      "01" when "011101101001", -- t[1897] = 1
      "01" when "011101101010", -- t[1898] = 1
      "01" when "011101101011", -- t[1899] = 1
      "01" when "011101101100", -- t[1900] = 1
      "01" when "011101101101", -- t[1901] = 1
      "01" when "011101101110", -- t[1902] = 1
      "01" when "011101101111", -- t[1903] = 1
      "01" when "011101110000", -- t[1904] = 1
      "01" when "011101110001", -- t[1905] = 1
      "01" when "011101110010", -- t[1906] = 1
      "01" when "011101110011", -- t[1907] = 1
      "01" when "011101110100", -- t[1908] = 1
      "01" when "011101110101", -- t[1909] = 1
      "01" when "011101110110", -- t[1910] = 1
      "01" when "011101110111", -- t[1911] = 1
      "01" when "011101111000", -- t[1912] = 1
      "01" when "011101111001", -- t[1913] = 1
      "01" when "011101111010", -- t[1914] = 1
      "01" when "011101111011", -- t[1915] = 1
      "01" when "011101111100", -- t[1916] = 1
      "01" when "011101111101", -- t[1917] = 1
      "01" when "011101111110", -- t[1918] = 1
      "01" when "011101111111", -- t[1919] = 1
      "01" when "011110000000", -- t[1920] = 1
      "01" when "011110000001", -- t[1921] = 1
      "01" when "011110000010", -- t[1922] = 1
      "01" when "011110000011", -- t[1923] = 1
      "01" when "011110000100", -- t[1924] = 1
      "01" when "011110000101", -- t[1925] = 1
      "01" when "011110000110", -- t[1926] = 1
      "01" when "011110000111", -- t[1927] = 1
      "01" when "011110001000", -- t[1928] = 1
      "01" when "011110001001", -- t[1929] = 1
      "01" when "011110001010", -- t[1930] = 1
      "01" when "011110001011", -- t[1931] = 1
      "01" when "011110001100", -- t[1932] = 1
      "01" when "011110001101", -- t[1933] = 1
      "01" when "011110001110", -- t[1934] = 1
      "01" when "011110001111", -- t[1935] = 1
      "01" when "011110010000", -- t[1936] = 1
      "01" when "011110010001", -- t[1937] = 1
      "01" when "011110010010", -- t[1938] = 1
      "01" when "011110010011", -- t[1939] = 1
      "01" when "011110010100", -- t[1940] = 1
      "01" when "011110010101", -- t[1941] = 1
      "01" when "011110010110", -- t[1942] = 1
      "01" when "011110010111", -- t[1943] = 1
      "01" when "011110011000", -- t[1944] = 1
      "01" when "011110011001", -- t[1945] = 1
      "01" when "011110011010", -- t[1946] = 1
      "01" when "011110011011", -- t[1947] = 1
      "01" when "011110011100", -- t[1948] = 1
      "01" when "011110011101", -- t[1949] = 1
      "01" when "011110011110", -- t[1950] = 1
      "01" when "011110011111", -- t[1951] = 1
      "01" when "011110100000", -- t[1952] = 1
      "01" when "011110100001", -- t[1953] = 1
      "01" when "011110100010", -- t[1954] = 1
      "01" when "011110100011", -- t[1955] = 1
      "01" when "011110100100", -- t[1956] = 1
      "01" when "011110100101", -- t[1957] = 1
      "01" when "011110100110", -- t[1958] = 1
      "01" when "011110100111", -- t[1959] = 1
      "01" when "011110101000", -- t[1960] = 1
      "01" when "011110101001", -- t[1961] = 1
      "01" when "011110101010", -- t[1962] = 1
      "01" when "011110101011", -- t[1963] = 1
      "01" when "011110101100", -- t[1964] = 1
      "01" when "011110101101", -- t[1965] = 1
      "01" when "011110101110", -- t[1966] = 1
      "01" when "011110101111", -- t[1967] = 1
      "01" when "011110110000", -- t[1968] = 1
      "01" when "011110110001", -- t[1969] = 1
      "01" when "011110110010", -- t[1970] = 1
      "01" when "011110110011", -- t[1971] = 1
      "01" when "011110110100", -- t[1972] = 1
      "01" when "011110110101", -- t[1973] = 1
      "01" when "011110110110", -- t[1974] = 1
      "01" when "011110110111", -- t[1975] = 1
      "01" when "011110111000", -- t[1976] = 1
      "01" when "011110111001", -- t[1977] = 1
      "01" when "011110111010", -- t[1978] = 1
      "01" when "011110111011", -- t[1979] = 1
      "01" when "011110111100", -- t[1980] = 1
      "01" when "011110111101", -- t[1981] = 1
      "01" when "011110111110", -- t[1982] = 1
      "01" when "011110111111", -- t[1983] = 1
      "01" when "011111000000", -- t[1984] = 1
      "01" when "011111000001", -- t[1985] = 1
      "01" when "011111000010", -- t[1986] = 1
      "01" when "011111000011", -- t[1987] = 1
      "01" when "011111000100", -- t[1988] = 1
      "01" when "011111000101", -- t[1989] = 1
      "01" when "011111000110", -- t[1990] = 1
      "01" when "011111000111", -- t[1991] = 1
      "01" when "011111001000", -- t[1992] = 1
      "01" when "011111001001", -- t[1993] = 1
      "01" when "011111001010", -- t[1994] = 1
      "01" when "011111001011", -- t[1995] = 1
      "01" when "011111001100", -- t[1996] = 1
      "01" when "011111001101", -- t[1997] = 1
      "01" when "011111001110", -- t[1998] = 1
      "01" when "011111001111", -- t[1999] = 1
      "01" when "011111010000", -- t[2000] = 1
      "01" when "011111010001", -- t[2001] = 1
      "01" when "011111010010", -- t[2002] = 1
      "01" when "011111010011", -- t[2003] = 1
      "01" when "011111010100", -- t[2004] = 1
      "01" when "011111010101", -- t[2005] = 1
      "01" when "011111010110", -- t[2006] = 1
      "01" when "011111010111", -- t[2007] = 1
      "01" when "011111011000", -- t[2008] = 1
      "01" when "011111011001", -- t[2009] = 1
      "01" when "011111011010", -- t[2010] = 1
      "01" when "011111011011", -- t[2011] = 1
      "01" when "011111011100", -- t[2012] = 1
      "01" when "011111011101", -- t[2013] = 1
      "01" when "011111011110", -- t[2014] = 1
      "01" when "011111011111", -- t[2015] = 1
      "01" when "011111100000", -- t[2016] = 1
      "01" when "011111100001", -- t[2017] = 1
      "01" when "011111100010", -- t[2018] = 1
      "01" when "011111100011", -- t[2019] = 1
      "01" when "011111100100", -- t[2020] = 1
      "01" when "011111100101", -- t[2021] = 1
      "01" when "011111100110", -- t[2022] = 1
      "01" when "011111100111", -- t[2023] = 1
      "01" when "011111101000", -- t[2024] = 1
      "01" when "011111101001", -- t[2025] = 1
      "01" when "011111101010", -- t[2026] = 1
      "01" when "011111101011", -- t[2027] = 1
      "01" when "011111101100", -- t[2028] = 1
      "01" when "011111101101", -- t[2029] = 1
      "01" when "011111101110", -- t[2030] = 1
      "01" when "011111101111", -- t[2031] = 1
      "01" when "011111110000", -- t[2032] = 1
      "01" when "011111110001", -- t[2033] = 1
      "01" when "011111110010", -- t[2034] = 1
      "01" when "011111110011", -- t[2035] = 1
      "01" when "011111110100", -- t[2036] = 1
      "01" when "011111110101", -- t[2037] = 1
      "01" when "011111110110", -- t[2038] = 1
      "01" when "011111110111", -- t[2039] = 1
      "01" when "011111111000", -- t[2040] = 1
      "01" when "011111111001", -- t[2041] = 1
      "01" when "011111111010", -- t[2042] = 1
      "01" when "011111111011", -- t[2043] = 1
      "01" when "011111111100", -- t[2044] = 1
      "01" when "011111111101", -- t[2045] = 1
      "01" when "011111111110", -- t[2046] = 1
      "01" when "011111111111", -- t[2047] = 1
      "--" when others;
end architecture;


-- MultiPartite: LNS addition function: [-8.0 0.0[ -> [0.0 2.0[
-- wI = 11 bits
-- wO = 9 bits
-- Decomposition: 7, 4 / 5, 3 / 2, 2
-- Guard bits: 3
-- Size: 1904 = 12.2^7 + 5.2^6 + 3.2^4

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSAdd_MPT_T2_8 is
  component LNSAdd_MPT_T2_8_tiv is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8_to1 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8_to0 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8_to1_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSAdd_MPT_T2_8_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_8_tiv is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8_tiv is
begin
  with x select
    r <=
      "000000010000" when "0000000", -- t[0] = 16
      "000000010001" when "0000001", -- t[1] = 17
      "000000010001" when "0000010", -- t[2] = 17
      "000000010010" when "0000011", -- t[3] = 18
      "000000010010" when "0000100", -- t[4] = 18
      "000000010011" when "0000101", -- t[5] = 19
      "000000010100" when "0000110", -- t[6] = 20
      "000000010100" when "0000111", -- t[7] = 20
      "000000010101" when "0001000", -- t[8] = 21
      "000000010110" when "0001001", -- t[9] = 22
      "000000010111" when "0001010", -- t[10] = 23
      "000000010111" when "0001011", -- t[11] = 23
      "000000011000" when "0001100", -- t[12] = 24
      "000000011001" when "0001101", -- t[13] = 25
      "000000011010" when "0001110", -- t[14] = 26
      "000000011011" when "0001111", -- t[15] = 27
      "000000011100" when "0010000", -- t[16] = 28
      "000000011101" when "0010001", -- t[17] = 29
      "000000011110" when "0010010", -- t[18] = 30
      "000000011111" when "0010011", -- t[19] = 31
      "000000100000" when "0010100", -- t[20] = 32
      "000000100010" when "0010101", -- t[21] = 34
      "000000100011" when "0010110", -- t[22] = 35
      "000000100100" when "0010111", -- t[23] = 36
      "000000100110" when "0011000", -- t[24] = 38
      "000000100111" when "0011001", -- t[25] = 39
      "000000101001" when "0011010", -- t[26] = 41
      "000000101010" when "0011011", -- t[27] = 42
      "000000101100" when "0011100", -- t[28] = 44
      "000000101110" when "0011101", -- t[29] = 46
      "000000101111" when "0011110", -- t[30] = 47
      "000000110001" when "0011111", -- t[31] = 49
      "000000110011" when "0100000", -- t[32] = 51
      "000000110101" when "0100001", -- t[33] = 53
      "000000110111" when "0100010", -- t[34] = 55
      "000000111010" when "0100011", -- t[35] = 58
      "000000111100" when "0100100", -- t[36] = 60
      "000000111110" when "0100101", -- t[37] = 62
      "000001000001" when "0100110", -- t[38] = 65
      "000001000100" when "0100111", -- t[39] = 68
      "000001000110" when "0101000", -- t[40] = 70
      "000001001001" when "0101001", -- t[41] = 73
      "000001001100" when "0101010", -- t[42] = 76
      "000001001111" when "0101011", -- t[43] = 79
      "000001010011" when "0101100", -- t[44] = 83
      "000001010110" when "0101101", -- t[45] = 86
      "000001011010" when "0101110", -- t[46] = 90
      "000001011101" when "0101111", -- t[47] = 93
      "000001100001" when "0110000", -- t[48] = 97
      "000001100101" when "0110001", -- t[49] = 101
      "000001101010" when "0110010", -- t[50] = 106
      "000001101110" when "0110011", -- t[51] = 110
      "000001110011" when "0110100", -- t[52] = 115
      "000001110111" when "0110101", -- t[53] = 119
      "000001111100" when "0110110", -- t[54] = 124
      "000010000001" when "0110111", -- t[55] = 129
      "000010000111" when "0111000", -- t[56] = 135
      "000010001101" when "0111001", -- t[57] = 141
      "000010010010" when "0111010", -- t[58] = 146
      "000010011001" when "0111011", -- t[59] = 153
      "000010011111" when "0111100", -- t[60] = 159
      "000010100110" when "0111101", -- t[61] = 166
      "000010101100" when "0111110", -- t[62] = 172
      "000010110100" when "0111111", -- t[63] = 180
      "000010111011" when "1000000", -- t[64] = 187
      "000011000011" when "1000001", -- t[65] = 195
      "000011001011" when "1000010", -- t[66] = 203
      "000011010100" when "1000011", -- t[67] = 212
      "000011011101" when "1000100", -- t[68] = 221
      "000011100110" when "1000101", -- t[69] = 230
      "000011101111" when "1000110", -- t[70] = 239
      "000011111001" when "1000111", -- t[71] = 249
      "000100000100" when "1001000", -- t[72] = 260
      "000100001111" when "1001001", -- t[73] = 271
      "000100011010" when "1001010", -- t[74] = 282
      "000100100101" when "1001011", -- t[75] = 293
      "000100110010" when "1001100", -- t[76] = 306
      "000100111110" when "1001101", -- t[77] = 318
      "000101001011" when "1001110", -- t[78] = 331
      "000101011001" when "1001111", -- t[79] = 345
      "000101100111" when "1010000", -- t[80] = 359
      "000101110110" when "1010001", -- t[81] = 374
      "000110000101" when "1010010", -- t[82] = 389
      "000110010101" when "1010011", -- t[83] = 405
      "000110100110" when "1010100", -- t[84] = 422
      "000110110111" when "1010101", -- t[85] = 439
      "000111001001" when "1010110", -- t[86] = 457
      "000111011011" when "1010111", -- t[87] = 475
      "000111101111" when "1011000", -- t[88] = 495
      "001000000011" when "1011001", -- t[89] = 515
      "001000010111" when "1011010", -- t[90] = 535
      "001000101101" when "1011011", -- t[91] = 557
      "001001000011" when "1011100", -- t[92] = 579
      "001001011010" when "1011101", -- t[93] = 602
      "001001110010" when "1011110", -- t[94] = 626
      "001010001010" when "1011111", -- t[95] = 650
      "001010100100" when "1100000", -- t[96] = 676
      "001010111110" when "1100001", -- t[97] = 702
      "001011011010" when "1100010", -- t[98] = 730
      "001011110110" when "1100011", -- t[99] = 758
      "001100010100" when "1100100", -- t[100] = 788
      "001100110010" when "1100101", -- t[101] = 818
      "001101010001" when "1100110", -- t[102] = 849
      "001101110001" when "1100111", -- t[103] = 881
      "001110010011" when "1101000", -- t[104] = 915
      "001110110101" when "1101001", -- t[105] = 949
      "001111011001" when "1101010", -- t[106] = 985
      "001111111110" when "1101011", -- t[107] = 1022
      "010000100100" when "1101100", -- t[108] = 1060
      "010001001011" when "1101101", -- t[109] = 1099
      "010001110011" when "1101110", -- t[110] = 1139
      "010010011100" when "1101111", -- t[111] = 1180
      "010011000111" when "1110000", -- t[112] = 1223
      "010011110011" when "1110001", -- t[113] = 1267
      "010100100000" when "1110010", -- t[114] = 1312
      "010101001110" when "1110011", -- t[115] = 1358
      "010101111110" when "1110100", -- t[116] = 1406
      "010110101111" when "1110101", -- t[117] = 1455
      "010111100001" when "1110110", -- t[118] = 1505
      "011000010101" when "1110111", -- t[119] = 1557
      "011001001010" when "1111000", -- t[120] = 1610
      "011010000000" when "1111001", -- t[121] = 1664
      "011010111000" when "1111010", -- t[122] = 1720
      "011011110001" when "1111011", -- t[123] = 1777
      "011100101011" when "1111100", -- t[124] = 1835
      "011101100111" when "1111101", -- t[125] = 1895
      "011110100100" when "1111110", -- t[126] = 1956
      "011111100011" when "1111111", -- t[127] = 2019
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_8_to1 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8_to1 is
begin
  with x select
    r <=
      "00000" when "000000", -- t[0] = 0
      "00000" when "000001", -- t[1] = 0
      "00000" when "000010", -- t[2] = 0
      "00000" when "000011", -- t[3] = 0
      "00000" when "000100", -- t[4] = 0
      "00000" when "000101", -- t[5] = 0
      "00000" when "000110", -- t[6] = 0
      "00000" when "000111", -- t[7] = 0
      "00000" when "001000", -- t[8] = 0
      "00000" when "001001", -- t[9] = 0
      "00000" when "001010", -- t[10] = 0
      "00000" when "001011", -- t[11] = 0
      "00000" when "001100", -- t[12] = 0
      "00000" when "001101", -- t[13] = 0
      "00000" when "001110", -- t[14] = 0
      "00000" when "001111", -- t[15] = 0
      "00000" when "010000", -- t[16] = 0
      "00000" when "010001", -- t[17] = 0
      "00000" when "010010", -- t[18] = 0
      "00000" when "010011", -- t[19] = 0
      "00000" when "010100", -- t[20] = 0
      "00001" when "010101", -- t[21] = 1
      "00000" when "010110", -- t[22] = 0
      "00001" when "010111", -- t[23] = 1
      "00000" when "011000", -- t[24] = 0
      "00001" when "011001", -- t[25] = 1
      "00000" when "011010", -- t[26] = 0
      "00001" when "011011", -- t[27] = 1
      "00000" when "011100", -- t[28] = 0
      "00010" when "011101", -- t[29] = 2
      "00000" when "011110", -- t[30] = 0
      "00010" when "011111", -- t[31] = 2
      "00001" when "100000", -- t[32] = 1
      "00011" when "100001", -- t[33] = 3
      "00001" when "100010", -- t[34] = 1
      "00011" when "100011", -- t[35] = 3
      "00001" when "100100", -- t[36] = 1
      "00100" when "100101", -- t[37] = 4
      "00001" when "100110", -- t[38] = 1
      "00100" when "100111", -- t[39] = 4
      "00001" when "101000", -- t[40] = 1
      "00101" when "101001", -- t[41] = 5
      "00010" when "101010", -- t[42] = 2
      "00110" when "101011", -- t[43] = 6
      "00010" when "101100", -- t[44] = 2
      "00111" when "101101", -- t[45] = 7
      "00010" when "101110", -- t[46] = 2
      "01000" when "101111", -- t[47] = 8
      "00011" when "110000", -- t[48] = 3
      "01010" when "110001", -- t[49] = 10
      "00011" when "110010", -- t[50] = 3
      "01011" when "110011", -- t[51] = 11
      "00100" when "110100", -- t[52] = 4
      "01101" when "110101", -- t[53] = 13
      "00101" when "110110", -- t[54] = 5
      "01111" when "110111", -- t[55] = 15
      "00101" when "111000", -- t[56] = 5
      "10000" when "111001", -- t[57] = 16
      "00110" when "111010", -- t[58] = 6
      "10010" when "111011", -- t[59] = 18
      "00110" when "111100", -- t[60] = 6
      "10100" when "111101", -- t[61] = 20
      "00111" when "111110", -- t[62] = 7
      "10110" when "111111", -- t[63] = 22
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_8_to0 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8_to0 is
begin
  with x select
    r <=
      "000" when "0000", -- t[0] = 0
      "000" when "0001", -- t[1] = 0
      "000" when "0010", -- t[2] = 0
      "000" when "0011", -- t[3] = 0
      "000" when "0100", -- t[4] = 0
      "000" when "0101", -- t[5] = 0
      "000" when "0110", -- t[6] = 0
      "000" when "0111", -- t[7] = 0
      "000" when "1000", -- t[8] = 0
      "001" when "1001", -- t[9] = 1
      "000" when "1010", -- t[10] = 0
      "001" when "1011", -- t[11] = 1
      "001" when "1100", -- t[12] = 1
      "011" when "1101", -- t[13] = 3
      "001" when "1110", -- t[14] = 1
      "100" when "1111", -- t[15] = 4
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_8.all;

entity LNSAdd_MPT_T2_8_to1_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSAdd_MPT_T2_8_to1
    port map( x => in_t,
              r => out_t );

  r(11 downto 5) <= (11 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_8.all;

entity LNSAdd_MPT_T2_8_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSAdd_MPT_T2_8_to0
    port map( x => in_t,
              r => out_t );

  r(11 downto 3) <= (11 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_8.all;

entity LNSAdd_MPT_T2_8 is
  port( x : in  std_logic_vector(10 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_8 is
  signal in_tiv  : std_logic_vector(6 downto 0);
  signal out_tiv : std_logic_vector(11 downto 0);
  signal a1      : std_logic_vector(4 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(11 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(11 downto 0);
  signal sum     : std_logic_vector(11 downto 0);
begin
  in_tiv <= x(10 downto 4);
  inst_tiv : LNSAdd_MPT_T2_8_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(10 downto 6);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSAdd_MPT_T2_8_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(10 downto 8);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSAdd_MPT_T2_8_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(11 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_8.all;
use fplib.pkg_misc.all;

entity LNSAdd_MPT_T2_8_Clk is
  port( x   : in  std_logic_vector(10 downto 0);
        r   : out std_logic_vector(8 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSAdd_MPT_T2_8_Clk is
  signal in_tiv_1  : std_logic_vector(6 downto 0);
  signal out_tiv_1 : std_logic_vector(11 downto 0);
  signal out_tiv_2 : std_logic_vector(11 downto 0);
  signal a1_1      : std_logic_vector(4 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(11 downto 0);
  signal out1_2    : std_logic_vector(11 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(11 downto 0);
  signal out0_2    : std_logic_vector(11 downto 0);
  signal psum1_2     : std_logic_vector(11 downto 0);
  signal psum1_3     : std_logic_vector(11 downto 0);
  signal psum2_2     : std_logic_vector(11 downto 0);
  signal psum2_3     : std_logic_vector(11 downto 0);
  signal sum_3     : std_logic_vector(11 downto 0);
begin
  in_tiv_1 <= x(10 downto 4);
  inst_tiv : LNSAdd_MPT_T2_8_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(10 downto 6);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSAdd_MPT_T2_8_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(10 downto 8);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSAdd_MPT_T2_8_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(11 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_8.all;

entity LNSAdd_MPT_8 is
  port( x : in  std_logic_vector(11 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_8 is
  signal out_t1 : std_logic_vector(1 downto 0);
  signal out_t2 : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSAdd_MPT_T1_8
    port map( x => x,
              r => out_t1 );

  inst_t2 : LNSAdd_MPT_T2_8
    port map( x => x(10 downto 0),
              r => out_t2 );

  r <= out_t2 when x(11 downto 11) = (11 downto 11 => '1') else
       (8 downto 2 => '0') & out_t1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_8.all;
use fplib.pkg_misc.all;

entity LNSAdd_MPT_8_Clk is
  port( x   : in  std_logic_vector(11 downto 0);
        r   : out std_logic_vector(8 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSAdd_MPT_8_Clk is
  signal x_1  : std_logic_vector(11 downto 0);
  signal x_10 : std_logic_vector(11 downto 0);

  signal out_t1_1  : std_logic_vector(1 downto 0);
  signal out_t1_10 : std_logic_vector(1 downto 0);
  signal out_t2_10 : std_logic_vector(8 downto 0);
begin
  x_1 <= x;

  inst_t1 : LNSAdd_MPT_T1_8
    port map( x => x_1,
              r => out_t1_1 );

  out_t1_delay : Delay
    generic map ( w => 2,
                  n => 1 )
    port map ( input  => out_t1_1,
               output => out_t1_10,
               clk    => clk );

  inst_t2 : LNSAdd_MPT_T2_8_Clk
    port map( x   => x(10 downto 0),
              r   => out_t2_10,
              clk => clk );

  x_delay : Delay
    generic map ( w => 12,
                  n => 1 )
    port map ( input  => x_1,
               output => x_10,
               clk    => clk );

  r <= out_t2_10 when x_10(11 downto 11) = (11 downto 11 => '1') else
       (8 downto 2 => '0') & out_t1_10;
end architecture;
