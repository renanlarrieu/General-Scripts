-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of MultiPartiteAdder object for LNS arithmetic in base 2.0 with 8-bit integer part and 7-bit fractional part
-- wI = 11 bits
-- wO = 8 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnsadd_mpt_7 is
  component LNSAdd_MPT_T1_7 is
    port( x : in  std_logic_vector(10 downto 0);
          r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSAdd_MPT_T2_7 is
    port( x : in  std_logic_vector(9 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;
end package;


-- SimpleTable: LNS addition function: [-16.0 0.0[ -> [0.0 2.0[
-- (bounded to [-16.0; -8.0[)
-- wI = 11 bits
-- wO = 1 bits

library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T1_7 is
  port( x : in  std_logic_vector(10 downto 0);
        r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T1_7 is
begin
  with x select
    r <=
      "0" when "00000000000", -- t[0] = 0
      "0" when "00000000001", -- t[1] = 0
      "0" when "00000000010", -- t[2] = 0
      "0" when "00000000011", -- t[3] = 0
      "0" when "00000000100", -- t[4] = 0
      "0" when "00000000101", -- t[5] = 0
      "0" when "00000000110", -- t[6] = 0
      "0" when "00000000111", -- t[7] = 0
      "0" when "00000001000", -- t[8] = 0
      "0" when "00000001001", -- t[9] = 0
      "0" when "00000001010", -- t[10] = 0
      "0" when "00000001011", -- t[11] = 0
      "0" when "00000001100", -- t[12] = 0
      "0" when "00000001101", -- t[13] = 0
      "0" when "00000001110", -- t[14] = 0
      "0" when "00000001111", -- t[15] = 0
      "0" when "00000010000", -- t[16] = 0
      "0" when "00000010001", -- t[17] = 0
      "0" when "00000010010", -- t[18] = 0
      "0" when "00000010011", -- t[19] = 0
      "0" when "00000010100", -- t[20] = 0
      "0" when "00000010101", -- t[21] = 0
      "0" when "00000010110", -- t[22] = 0
      "0" when "00000010111", -- t[23] = 0
      "0" when "00000011000", -- t[24] = 0
      "0" when "00000011001", -- t[25] = 0
      "0" when "00000011010", -- t[26] = 0
      "0" when "00000011011", -- t[27] = 0
      "0" when "00000011100", -- t[28] = 0
      "0" when "00000011101", -- t[29] = 0
      "0" when "00000011110", -- t[30] = 0
      "0" when "00000011111", -- t[31] = 0
      "0" when "00000100000", -- t[32] = 0
      "0" when "00000100001", -- t[33] = 0
      "0" when "00000100010", -- t[34] = 0
      "0" when "00000100011", -- t[35] = 0
      "0" when "00000100100", -- t[36] = 0
      "0" when "00000100101", -- t[37] = 0
      "0" when "00000100110", -- t[38] = 0
      "0" when "00000100111", -- t[39] = 0
      "0" when "00000101000", -- t[40] = 0
      "0" when "00000101001", -- t[41] = 0
      "0" when "00000101010", -- t[42] = 0
      "0" when "00000101011", -- t[43] = 0
      "0" when "00000101100", -- t[44] = 0
      "0" when "00000101101", -- t[45] = 0
      "0" when "00000101110", -- t[46] = 0
      "0" when "00000101111", -- t[47] = 0
      "0" when "00000110000", -- t[48] = 0
      "0" when "00000110001", -- t[49] = 0
      "0" when "00000110010", -- t[50] = 0
      "0" when "00000110011", -- t[51] = 0
      "0" when "00000110100", -- t[52] = 0
      "0" when "00000110101", -- t[53] = 0
      "0" when "00000110110", -- t[54] = 0
      "0" when "00000110111", -- t[55] = 0
      "0" when "00000111000", -- t[56] = 0
      "0" when "00000111001", -- t[57] = 0
      "0" when "00000111010", -- t[58] = 0
      "0" when "00000111011", -- t[59] = 0
      "0" when "00000111100", -- t[60] = 0
      "0" when "00000111101", -- t[61] = 0
      "0" when "00000111110", -- t[62] = 0
      "0" when "00000111111", -- t[63] = 0
      "0" when "00001000000", -- t[64] = 0
      "0" when "00001000001", -- t[65] = 0
      "0" when "00001000010", -- t[66] = 0
      "0" when "00001000011", -- t[67] = 0
      "0" when "00001000100", -- t[68] = 0
      "0" when "00001000101", -- t[69] = 0
      "0" when "00001000110", -- t[70] = 0
      "0" when "00001000111", -- t[71] = 0
      "0" when "00001001000", -- t[72] = 0
      "0" when "00001001001", -- t[73] = 0
      "0" when "00001001010", -- t[74] = 0
      "0" when "00001001011", -- t[75] = 0
      "0" when "00001001100", -- t[76] = 0
      "0" when "00001001101", -- t[77] = 0
      "0" when "00001001110", -- t[78] = 0
      "0" when "00001001111", -- t[79] = 0
      "0" when "00001010000", -- t[80] = 0
      "0" when "00001010001", -- t[81] = 0
      "0" when "00001010010", -- t[82] = 0
      "0" when "00001010011", -- t[83] = 0
      "0" when "00001010100", -- t[84] = 0
      "0" when "00001010101", -- t[85] = 0
      "0" when "00001010110", -- t[86] = 0
      "0" when "00001010111", -- t[87] = 0
      "0" when "00001011000", -- t[88] = 0
      "0" when "00001011001", -- t[89] = 0
      "0" when "00001011010", -- t[90] = 0
      "0" when "00001011011", -- t[91] = 0
      "0" when "00001011100", -- t[92] = 0
      "0" when "00001011101", -- t[93] = 0
      "0" when "00001011110", -- t[94] = 0
      "0" when "00001011111", -- t[95] = 0
      "0" when "00001100000", -- t[96] = 0
      "0" when "00001100001", -- t[97] = 0
      "0" when "00001100010", -- t[98] = 0
      "0" when "00001100011", -- t[99] = 0
      "0" when "00001100100", -- t[100] = 0
      "0" when "00001100101", -- t[101] = 0
      "0" when "00001100110", -- t[102] = 0
      "0" when "00001100111", -- t[103] = 0
      "0" when "00001101000", -- t[104] = 0
      "0" when "00001101001", -- t[105] = 0
      "0" when "00001101010", -- t[106] = 0
      "0" when "00001101011", -- t[107] = 0
      "0" when "00001101100", -- t[108] = 0
      "0" when "00001101101", -- t[109] = 0
      "0" when "00001101110", -- t[110] = 0
      "0" when "00001101111", -- t[111] = 0
      "0" when "00001110000", -- t[112] = 0
      "0" when "00001110001", -- t[113] = 0
      "0" when "00001110010", -- t[114] = 0
      "0" when "00001110011", -- t[115] = 0
      "0" when "00001110100", -- t[116] = 0
      "0" when "00001110101", -- t[117] = 0
      "0" when "00001110110", -- t[118] = 0
      "0" when "00001110111", -- t[119] = 0
      "0" when "00001111000", -- t[120] = 0
      "0" when "00001111001", -- t[121] = 0
      "0" when "00001111010", -- t[122] = 0
      "0" when "00001111011", -- t[123] = 0
      "0" when "00001111100", -- t[124] = 0
      "0" when "00001111101", -- t[125] = 0
      "0" when "00001111110", -- t[126] = 0
      "0" when "00001111111", -- t[127] = 0
      "0" when "00010000000", -- t[128] = 0
      "0" when "00010000001", -- t[129] = 0
      "0" when "00010000010", -- t[130] = 0
      "0" when "00010000011", -- t[131] = 0
      "0" when "00010000100", -- t[132] = 0
      "0" when "00010000101", -- t[133] = 0
      "0" when "00010000110", -- t[134] = 0
      "0" when "00010000111", -- t[135] = 0
      "0" when "00010001000", -- t[136] = 0
      "0" when "00010001001", -- t[137] = 0
      "0" when "00010001010", -- t[138] = 0
      "0" when "00010001011", -- t[139] = 0
      "0" when "00010001100", -- t[140] = 0
      "0" when "00010001101", -- t[141] = 0
      "0" when "00010001110", -- t[142] = 0
      "0" when "00010001111", -- t[143] = 0
      "0" when "00010010000", -- t[144] = 0
      "0" when "00010010001", -- t[145] = 0
      "0" when "00010010010", -- t[146] = 0
      "0" when "00010010011", -- t[147] = 0
      "0" when "00010010100", -- t[148] = 0
      "0" when "00010010101", -- t[149] = 0
      "0" when "00010010110", -- t[150] = 0
      "0" when "00010010111", -- t[151] = 0
      "0" when "00010011000", -- t[152] = 0
      "0" when "00010011001", -- t[153] = 0
      "0" when "00010011010", -- t[154] = 0
      "0" when "00010011011", -- t[155] = 0
      "0" when "00010011100", -- t[156] = 0
      "0" when "00010011101", -- t[157] = 0
      "0" when "00010011110", -- t[158] = 0
      "0" when "00010011111", -- t[159] = 0
      "0" when "00010100000", -- t[160] = 0
      "0" when "00010100001", -- t[161] = 0
      "0" when "00010100010", -- t[162] = 0
      "0" when "00010100011", -- t[163] = 0
      "0" when "00010100100", -- t[164] = 0
      "0" when "00010100101", -- t[165] = 0
      "0" when "00010100110", -- t[166] = 0
      "0" when "00010100111", -- t[167] = 0
      "0" when "00010101000", -- t[168] = 0
      "0" when "00010101001", -- t[169] = 0
      "0" when "00010101010", -- t[170] = 0
      "0" when "00010101011", -- t[171] = 0
      "0" when "00010101100", -- t[172] = 0
      "0" when "00010101101", -- t[173] = 0
      "0" when "00010101110", -- t[174] = 0
      "0" when "00010101111", -- t[175] = 0
      "0" when "00010110000", -- t[176] = 0
      "0" when "00010110001", -- t[177] = 0
      "0" when "00010110010", -- t[178] = 0
      "0" when "00010110011", -- t[179] = 0
      "0" when "00010110100", -- t[180] = 0
      "0" when "00010110101", -- t[181] = 0
      "0" when "00010110110", -- t[182] = 0
      "0" when "00010110111", -- t[183] = 0
      "0" when "00010111000", -- t[184] = 0
      "0" when "00010111001", -- t[185] = 0
      "0" when "00010111010", -- t[186] = 0
      "0" when "00010111011", -- t[187] = 0
      "0" when "00010111100", -- t[188] = 0
      "0" when "00010111101", -- t[189] = 0
      "0" when "00010111110", -- t[190] = 0
      "0" when "00010111111", -- t[191] = 0
      "0" when "00011000000", -- t[192] = 0
      "0" when "00011000001", -- t[193] = 0
      "0" when "00011000010", -- t[194] = 0
      "0" when "00011000011", -- t[195] = 0
      "0" when "00011000100", -- t[196] = 0
      "0" when "00011000101", -- t[197] = 0
      "0" when "00011000110", -- t[198] = 0
      "0" when "00011000111", -- t[199] = 0
      "0" when "00011001000", -- t[200] = 0
      "0" when "00011001001", -- t[201] = 0
      "0" when "00011001010", -- t[202] = 0
      "0" when "00011001011", -- t[203] = 0
      "0" when "00011001100", -- t[204] = 0
      "0" when "00011001101", -- t[205] = 0
      "0" when "00011001110", -- t[206] = 0
      "0" when "00011001111", -- t[207] = 0
      "0" when "00011010000", -- t[208] = 0
      "0" when "00011010001", -- t[209] = 0
      "0" when "00011010010", -- t[210] = 0
      "0" when "00011010011", -- t[211] = 0
      "0" when "00011010100", -- t[212] = 0
      "0" when "00011010101", -- t[213] = 0
      "0" when "00011010110", -- t[214] = 0
      "0" when "00011010111", -- t[215] = 0
      "0" when "00011011000", -- t[216] = 0
      "0" when "00011011001", -- t[217] = 0
      "0" when "00011011010", -- t[218] = 0
      "0" when "00011011011", -- t[219] = 0
      "0" when "00011011100", -- t[220] = 0
      "0" when "00011011101", -- t[221] = 0
      "0" when "00011011110", -- t[222] = 0
      "0" when "00011011111", -- t[223] = 0
      "0" when "00011100000", -- t[224] = 0
      "0" when "00011100001", -- t[225] = 0
      "0" when "00011100010", -- t[226] = 0
      "0" when "00011100011", -- t[227] = 0
      "0" when "00011100100", -- t[228] = 0
      "0" when "00011100101", -- t[229] = 0
      "0" when "00011100110", -- t[230] = 0
      "0" when "00011100111", -- t[231] = 0
      "0" when "00011101000", -- t[232] = 0
      "0" when "00011101001", -- t[233] = 0
      "0" when "00011101010", -- t[234] = 0
      "0" when "00011101011", -- t[235] = 0
      "0" when "00011101100", -- t[236] = 0
      "0" when "00011101101", -- t[237] = 0
      "0" when "00011101110", -- t[238] = 0
      "0" when "00011101111", -- t[239] = 0
      "0" when "00011110000", -- t[240] = 0
      "0" when "00011110001", -- t[241] = 0
      "0" when "00011110010", -- t[242] = 0
      "0" when "00011110011", -- t[243] = 0
      "0" when "00011110100", -- t[244] = 0
      "0" when "00011110101", -- t[245] = 0
      "0" when "00011110110", -- t[246] = 0
      "0" when "00011110111", -- t[247] = 0
      "0" when "00011111000", -- t[248] = 0
      "0" when "00011111001", -- t[249] = 0
      "0" when "00011111010", -- t[250] = 0
      "0" when "00011111011", -- t[251] = 0
      "0" when "00011111100", -- t[252] = 0
      "0" when "00011111101", -- t[253] = 0
      "0" when "00011111110", -- t[254] = 0
      "0" when "00011111111", -- t[255] = 0
      "0" when "00100000000", -- t[256] = 0
      "0" when "00100000001", -- t[257] = 0
      "0" when "00100000010", -- t[258] = 0
      "0" when "00100000011", -- t[259] = 0
      "0" when "00100000100", -- t[260] = 0
      "0" when "00100000101", -- t[261] = 0
      "0" when "00100000110", -- t[262] = 0
      "0" when "00100000111", -- t[263] = 0
      "0" when "00100001000", -- t[264] = 0
      "0" when "00100001001", -- t[265] = 0
      "0" when "00100001010", -- t[266] = 0
      "0" when "00100001011", -- t[267] = 0
      "0" when "00100001100", -- t[268] = 0
      "0" when "00100001101", -- t[269] = 0
      "0" when "00100001110", -- t[270] = 0
      "0" when "00100001111", -- t[271] = 0
      "0" when "00100010000", -- t[272] = 0
      "0" when "00100010001", -- t[273] = 0
      "0" when "00100010010", -- t[274] = 0
      "0" when "00100010011", -- t[275] = 0
      "0" when "00100010100", -- t[276] = 0
      "0" when "00100010101", -- t[277] = 0
      "0" when "00100010110", -- t[278] = 0
      "0" when "00100010111", -- t[279] = 0
      "0" when "00100011000", -- t[280] = 0
      "0" when "00100011001", -- t[281] = 0
      "0" when "00100011010", -- t[282] = 0
      "0" when "00100011011", -- t[283] = 0
      "0" when "00100011100", -- t[284] = 0
      "0" when "00100011101", -- t[285] = 0
      "0" when "00100011110", -- t[286] = 0
      "0" when "00100011111", -- t[287] = 0
      "0" when "00100100000", -- t[288] = 0
      "0" when "00100100001", -- t[289] = 0
      "0" when "00100100010", -- t[290] = 0
      "0" when "00100100011", -- t[291] = 0
      "0" when "00100100100", -- t[292] = 0
      "0" when "00100100101", -- t[293] = 0
      "0" when "00100100110", -- t[294] = 0
      "0" when "00100100111", -- t[295] = 0
      "0" when "00100101000", -- t[296] = 0
      "0" when "00100101001", -- t[297] = 0
      "0" when "00100101010", -- t[298] = 0
      "0" when "00100101011", -- t[299] = 0
      "0" when "00100101100", -- t[300] = 0
      "0" when "00100101101", -- t[301] = 0
      "0" when "00100101110", -- t[302] = 0
      "0" when "00100101111", -- t[303] = 0
      "0" when "00100110000", -- t[304] = 0
      "0" when "00100110001", -- t[305] = 0
      "0" when "00100110010", -- t[306] = 0
      "0" when "00100110011", -- t[307] = 0
      "0" when "00100110100", -- t[308] = 0
      "0" when "00100110101", -- t[309] = 0
      "0" when "00100110110", -- t[310] = 0
      "0" when "00100110111", -- t[311] = 0
      "0" when "00100111000", -- t[312] = 0
      "0" when "00100111001", -- t[313] = 0
      "0" when "00100111010", -- t[314] = 0
      "0" when "00100111011", -- t[315] = 0
      "0" when "00100111100", -- t[316] = 0
      "0" when "00100111101", -- t[317] = 0
      "0" when "00100111110", -- t[318] = 0
      "0" when "00100111111", -- t[319] = 0
      "0" when "00101000000", -- t[320] = 0
      "0" when "00101000001", -- t[321] = 0
      "0" when "00101000010", -- t[322] = 0
      "0" when "00101000011", -- t[323] = 0
      "0" when "00101000100", -- t[324] = 0
      "0" when "00101000101", -- t[325] = 0
      "0" when "00101000110", -- t[326] = 0
      "0" when "00101000111", -- t[327] = 0
      "0" when "00101001000", -- t[328] = 0
      "0" when "00101001001", -- t[329] = 0
      "0" when "00101001010", -- t[330] = 0
      "0" when "00101001011", -- t[331] = 0
      "0" when "00101001100", -- t[332] = 0
      "0" when "00101001101", -- t[333] = 0
      "0" when "00101001110", -- t[334] = 0
      "0" when "00101001111", -- t[335] = 0
      "0" when "00101010000", -- t[336] = 0
      "0" when "00101010001", -- t[337] = 0
      "0" when "00101010010", -- t[338] = 0
      "0" when "00101010011", -- t[339] = 0
      "0" when "00101010100", -- t[340] = 0
      "0" when "00101010101", -- t[341] = 0
      "0" when "00101010110", -- t[342] = 0
      "0" when "00101010111", -- t[343] = 0
      "0" when "00101011000", -- t[344] = 0
      "0" when "00101011001", -- t[345] = 0
      "0" when "00101011010", -- t[346] = 0
      "0" when "00101011011", -- t[347] = 0
      "0" when "00101011100", -- t[348] = 0
      "0" when "00101011101", -- t[349] = 0
      "0" when "00101011110", -- t[350] = 0
      "0" when "00101011111", -- t[351] = 0
      "0" when "00101100000", -- t[352] = 0
      "0" when "00101100001", -- t[353] = 0
      "0" when "00101100010", -- t[354] = 0
      "0" when "00101100011", -- t[355] = 0
      "0" when "00101100100", -- t[356] = 0
      "0" when "00101100101", -- t[357] = 0
      "0" when "00101100110", -- t[358] = 0
      "0" when "00101100111", -- t[359] = 0
      "0" when "00101101000", -- t[360] = 0
      "0" when "00101101001", -- t[361] = 0
      "0" when "00101101010", -- t[362] = 0
      "0" when "00101101011", -- t[363] = 0
      "0" when "00101101100", -- t[364] = 0
      "0" when "00101101101", -- t[365] = 0
      "0" when "00101101110", -- t[366] = 0
      "0" when "00101101111", -- t[367] = 0
      "0" when "00101110000", -- t[368] = 0
      "0" when "00101110001", -- t[369] = 0
      "0" when "00101110010", -- t[370] = 0
      "0" when "00101110011", -- t[371] = 0
      "0" when "00101110100", -- t[372] = 0
      "0" when "00101110101", -- t[373] = 0
      "0" when "00101110110", -- t[374] = 0
      "0" when "00101110111", -- t[375] = 0
      "0" when "00101111000", -- t[376] = 0
      "0" when "00101111001", -- t[377] = 0
      "0" when "00101111010", -- t[378] = 0
      "0" when "00101111011", -- t[379] = 0
      "0" when "00101111100", -- t[380] = 0
      "0" when "00101111101", -- t[381] = 0
      "0" when "00101111110", -- t[382] = 0
      "0" when "00101111111", -- t[383] = 0
      "0" when "00110000000", -- t[384] = 0
      "0" when "00110000001", -- t[385] = 0
      "0" when "00110000010", -- t[386] = 0
      "0" when "00110000011", -- t[387] = 0
      "0" when "00110000100", -- t[388] = 0
      "0" when "00110000101", -- t[389] = 0
      "0" when "00110000110", -- t[390] = 0
      "0" when "00110000111", -- t[391] = 0
      "0" when "00110001000", -- t[392] = 0
      "0" when "00110001001", -- t[393] = 0
      "0" when "00110001010", -- t[394] = 0
      "0" when "00110001011", -- t[395] = 0
      "0" when "00110001100", -- t[396] = 0
      "0" when "00110001101", -- t[397] = 0
      "0" when "00110001110", -- t[398] = 0
      "0" when "00110001111", -- t[399] = 0
      "0" when "00110010000", -- t[400] = 0
      "0" when "00110010001", -- t[401] = 0
      "0" when "00110010010", -- t[402] = 0
      "0" when "00110010011", -- t[403] = 0
      "0" when "00110010100", -- t[404] = 0
      "0" when "00110010101", -- t[405] = 0
      "0" when "00110010110", -- t[406] = 0
      "0" when "00110010111", -- t[407] = 0
      "0" when "00110011000", -- t[408] = 0
      "0" when "00110011001", -- t[409] = 0
      "0" when "00110011010", -- t[410] = 0
      "0" when "00110011011", -- t[411] = 0
      "0" when "00110011100", -- t[412] = 0
      "0" when "00110011101", -- t[413] = 0
      "0" when "00110011110", -- t[414] = 0
      "0" when "00110011111", -- t[415] = 0
      "0" when "00110100000", -- t[416] = 0
      "0" when "00110100001", -- t[417] = 0
      "0" when "00110100010", -- t[418] = 0
      "0" when "00110100011", -- t[419] = 0
      "0" when "00110100100", -- t[420] = 0
      "0" when "00110100101", -- t[421] = 0
      "0" when "00110100110", -- t[422] = 0
      "0" when "00110100111", -- t[423] = 0
      "0" when "00110101000", -- t[424] = 0
      "0" when "00110101001", -- t[425] = 0
      "0" when "00110101010", -- t[426] = 0
      "0" when "00110101011", -- t[427] = 0
      "0" when "00110101100", -- t[428] = 0
      "0" when "00110101101", -- t[429] = 0
      "0" when "00110101110", -- t[430] = 0
      "0" when "00110101111", -- t[431] = 0
      "0" when "00110110000", -- t[432] = 0
      "0" when "00110110001", -- t[433] = 0
      "0" when "00110110010", -- t[434] = 0
      "0" when "00110110011", -- t[435] = 0
      "0" when "00110110100", -- t[436] = 0
      "0" when "00110110101", -- t[437] = 0
      "0" when "00110110110", -- t[438] = 0
      "0" when "00110110111", -- t[439] = 0
      "0" when "00110111000", -- t[440] = 0
      "0" when "00110111001", -- t[441] = 0
      "0" when "00110111010", -- t[442] = 0
      "0" when "00110111011", -- t[443] = 0
      "0" when "00110111100", -- t[444] = 0
      "0" when "00110111101", -- t[445] = 0
      "0" when "00110111110", -- t[446] = 0
      "0" when "00110111111", -- t[447] = 0
      "0" when "00111000000", -- t[448] = 0
      "0" when "00111000001", -- t[449] = 0
      "0" when "00111000010", -- t[450] = 0
      "0" when "00111000011", -- t[451] = 0
      "0" when "00111000100", -- t[452] = 0
      "0" when "00111000101", -- t[453] = 0
      "0" when "00111000110", -- t[454] = 0
      "0" when "00111000111", -- t[455] = 0
      "0" when "00111001000", -- t[456] = 0
      "0" when "00111001001", -- t[457] = 0
      "0" when "00111001010", -- t[458] = 0
      "0" when "00111001011", -- t[459] = 0
      "0" when "00111001100", -- t[460] = 0
      "0" when "00111001101", -- t[461] = 0
      "0" when "00111001110", -- t[462] = 0
      "0" when "00111001111", -- t[463] = 0
      "0" when "00111010000", -- t[464] = 0
      "0" when "00111010001", -- t[465] = 0
      "0" when "00111010010", -- t[466] = 0
      "0" when "00111010011", -- t[467] = 0
      "0" when "00111010100", -- t[468] = 0
      "0" when "00111010101", -- t[469] = 0
      "0" when "00111010110", -- t[470] = 0
      "0" when "00111010111", -- t[471] = 0
      "0" when "00111011000", -- t[472] = 0
      "0" when "00111011001", -- t[473] = 0
      "0" when "00111011010", -- t[474] = 0
      "0" when "00111011011", -- t[475] = 0
      "0" when "00111011100", -- t[476] = 0
      "0" when "00111011101", -- t[477] = 0
      "0" when "00111011110", -- t[478] = 0
      "0" when "00111011111", -- t[479] = 0
      "0" when "00111100000", -- t[480] = 0
      "0" when "00111100001", -- t[481] = 0
      "0" when "00111100010", -- t[482] = 0
      "0" when "00111100011", -- t[483] = 0
      "0" when "00111100100", -- t[484] = 0
      "0" when "00111100101", -- t[485] = 0
      "0" when "00111100110", -- t[486] = 0
      "0" when "00111100111", -- t[487] = 0
      "0" when "00111101000", -- t[488] = 0
      "0" when "00111101001", -- t[489] = 0
      "0" when "00111101010", -- t[490] = 0
      "0" when "00111101011", -- t[491] = 0
      "0" when "00111101100", -- t[492] = 0
      "0" when "00111101101", -- t[493] = 0
      "0" when "00111101110", -- t[494] = 0
      "0" when "00111101111", -- t[495] = 0
      "0" when "00111110000", -- t[496] = 0
      "0" when "00111110001", -- t[497] = 0
      "0" when "00111110010", -- t[498] = 0
      "0" when "00111110011", -- t[499] = 0
      "0" when "00111110100", -- t[500] = 0
      "0" when "00111110101", -- t[501] = 0
      "0" when "00111110110", -- t[502] = 0
      "0" when "00111110111", -- t[503] = 0
      "0" when "00111111000", -- t[504] = 0
      "0" when "00111111001", -- t[505] = 0
      "0" when "00111111010", -- t[506] = 0
      "0" when "00111111011", -- t[507] = 0
      "0" when "00111111100", -- t[508] = 0
      "0" when "00111111101", -- t[509] = 0
      "0" when "00111111110", -- t[510] = 0
      "0" when "00111111111", -- t[511] = 0
      "0" when "01000000000", -- t[512] = 0
      "0" when "01000000001", -- t[513] = 0
      "0" when "01000000010", -- t[514] = 0
      "0" when "01000000011", -- t[515] = 0
      "0" when "01000000100", -- t[516] = 0
      "0" when "01000000101", -- t[517] = 0
      "0" when "01000000110", -- t[518] = 0
      "0" when "01000000111", -- t[519] = 0
      "0" when "01000001000", -- t[520] = 0
      "0" when "01000001001", -- t[521] = 0
      "0" when "01000001010", -- t[522] = 0
      "0" when "01000001011", -- t[523] = 0
      "0" when "01000001100", -- t[524] = 0
      "0" when "01000001101", -- t[525] = 0
      "0" when "01000001110", -- t[526] = 0
      "0" when "01000001111", -- t[527] = 0
      "0" when "01000010000", -- t[528] = 0
      "0" when "01000010001", -- t[529] = 0
      "0" when "01000010010", -- t[530] = 0
      "0" when "01000010011", -- t[531] = 0
      "0" when "01000010100", -- t[532] = 0
      "0" when "01000010101", -- t[533] = 0
      "0" when "01000010110", -- t[534] = 0
      "0" when "01000010111", -- t[535] = 0
      "0" when "01000011000", -- t[536] = 0
      "0" when "01000011001", -- t[537] = 0
      "0" when "01000011010", -- t[538] = 0
      "0" when "01000011011", -- t[539] = 0
      "0" when "01000011100", -- t[540] = 0
      "0" when "01000011101", -- t[541] = 0
      "0" when "01000011110", -- t[542] = 0
      "0" when "01000011111", -- t[543] = 0
      "0" when "01000100000", -- t[544] = 0
      "0" when "01000100001", -- t[545] = 0
      "0" when "01000100010", -- t[546] = 0
      "0" when "01000100011", -- t[547] = 0
      "0" when "01000100100", -- t[548] = 0
      "0" when "01000100101", -- t[549] = 0
      "0" when "01000100110", -- t[550] = 0
      "0" when "01000100111", -- t[551] = 0
      "0" when "01000101000", -- t[552] = 0
      "0" when "01000101001", -- t[553] = 0
      "0" when "01000101010", -- t[554] = 0
      "0" when "01000101011", -- t[555] = 0
      "0" when "01000101100", -- t[556] = 0
      "0" when "01000101101", -- t[557] = 0
      "0" when "01000101110", -- t[558] = 0
      "0" when "01000101111", -- t[559] = 0
      "0" when "01000110000", -- t[560] = 0
      "0" when "01000110001", -- t[561] = 0
      "0" when "01000110010", -- t[562] = 0
      "0" when "01000110011", -- t[563] = 0
      "0" when "01000110100", -- t[564] = 0
      "0" when "01000110101", -- t[565] = 0
      "0" when "01000110110", -- t[566] = 0
      "0" when "01000110111", -- t[567] = 0
      "0" when "01000111000", -- t[568] = 0
      "0" when "01000111001", -- t[569] = 0
      "0" when "01000111010", -- t[570] = 0
      "0" when "01000111011", -- t[571] = 0
      "0" when "01000111100", -- t[572] = 0
      "0" when "01000111101", -- t[573] = 0
      "0" when "01000111110", -- t[574] = 0
      "0" when "01000111111", -- t[575] = 0
      "0" when "01001000000", -- t[576] = 0
      "0" when "01001000001", -- t[577] = 0
      "0" when "01001000010", -- t[578] = 0
      "0" when "01001000011", -- t[579] = 0
      "0" when "01001000100", -- t[580] = 0
      "0" when "01001000101", -- t[581] = 0
      "0" when "01001000110", -- t[582] = 0
      "0" when "01001000111", -- t[583] = 0
      "0" when "01001001000", -- t[584] = 0
      "0" when "01001001001", -- t[585] = 0
      "0" when "01001001010", -- t[586] = 0
      "0" when "01001001011", -- t[587] = 0
      "0" when "01001001100", -- t[588] = 0
      "0" when "01001001101", -- t[589] = 0
      "0" when "01001001110", -- t[590] = 0
      "0" when "01001001111", -- t[591] = 0
      "0" when "01001010000", -- t[592] = 0
      "0" when "01001010001", -- t[593] = 0
      "0" when "01001010010", -- t[594] = 0
      "0" when "01001010011", -- t[595] = 0
      "0" when "01001010100", -- t[596] = 0
      "0" when "01001010101", -- t[597] = 0
      "0" when "01001010110", -- t[598] = 0
      "0" when "01001010111", -- t[599] = 0
      "0" when "01001011000", -- t[600] = 0
      "0" when "01001011001", -- t[601] = 0
      "0" when "01001011010", -- t[602] = 0
      "0" when "01001011011", -- t[603] = 0
      "0" when "01001011100", -- t[604] = 0
      "0" when "01001011101", -- t[605] = 0
      "0" when "01001011110", -- t[606] = 0
      "0" when "01001011111", -- t[607] = 0
      "0" when "01001100000", -- t[608] = 0
      "0" when "01001100001", -- t[609] = 0
      "0" when "01001100010", -- t[610] = 0
      "0" when "01001100011", -- t[611] = 0
      "0" when "01001100100", -- t[612] = 0
      "0" when "01001100101", -- t[613] = 0
      "0" when "01001100110", -- t[614] = 0
      "0" when "01001100111", -- t[615] = 0
      "0" when "01001101000", -- t[616] = 0
      "0" when "01001101001", -- t[617] = 0
      "0" when "01001101010", -- t[618] = 0
      "0" when "01001101011", -- t[619] = 0
      "0" when "01001101100", -- t[620] = 0
      "0" when "01001101101", -- t[621] = 0
      "0" when "01001101110", -- t[622] = 0
      "0" when "01001101111", -- t[623] = 0
      "0" when "01001110000", -- t[624] = 0
      "0" when "01001110001", -- t[625] = 0
      "0" when "01001110010", -- t[626] = 0
      "0" when "01001110011", -- t[627] = 0
      "0" when "01001110100", -- t[628] = 0
      "0" when "01001110101", -- t[629] = 0
      "0" when "01001110110", -- t[630] = 0
      "0" when "01001110111", -- t[631] = 0
      "0" when "01001111000", -- t[632] = 0
      "0" when "01001111001", -- t[633] = 0
      "0" when "01001111010", -- t[634] = 0
      "0" when "01001111011", -- t[635] = 0
      "0" when "01001111100", -- t[636] = 0
      "0" when "01001111101", -- t[637] = 0
      "0" when "01001111110", -- t[638] = 0
      "0" when "01001111111", -- t[639] = 0
      "0" when "01010000000", -- t[640] = 0
      "0" when "01010000001", -- t[641] = 0
      "0" when "01010000010", -- t[642] = 0
      "0" when "01010000011", -- t[643] = 0
      "0" when "01010000100", -- t[644] = 0
      "0" when "01010000101", -- t[645] = 0
      "0" when "01010000110", -- t[646] = 0
      "0" when "01010000111", -- t[647] = 0
      "0" when "01010001000", -- t[648] = 0
      "0" when "01010001001", -- t[649] = 0
      "0" when "01010001010", -- t[650] = 0
      "0" when "01010001011", -- t[651] = 0
      "0" when "01010001100", -- t[652] = 0
      "0" when "01010001101", -- t[653] = 0
      "0" when "01010001110", -- t[654] = 0
      "0" when "01010001111", -- t[655] = 0
      "0" when "01010010000", -- t[656] = 0
      "0" when "01010010001", -- t[657] = 0
      "0" when "01010010010", -- t[658] = 0
      "0" when "01010010011", -- t[659] = 0
      "0" when "01010010100", -- t[660] = 0
      "0" when "01010010101", -- t[661] = 0
      "0" when "01010010110", -- t[662] = 0
      "0" when "01010010111", -- t[663] = 0
      "0" when "01010011000", -- t[664] = 0
      "0" when "01010011001", -- t[665] = 0
      "0" when "01010011010", -- t[666] = 0
      "0" when "01010011011", -- t[667] = 0
      "0" when "01010011100", -- t[668] = 0
      "0" when "01010011101", -- t[669] = 0
      "0" when "01010011110", -- t[670] = 0
      "0" when "01010011111", -- t[671] = 0
      "0" when "01010100000", -- t[672] = 0
      "0" when "01010100001", -- t[673] = 0
      "0" when "01010100010", -- t[674] = 0
      "0" when "01010100011", -- t[675] = 0
      "0" when "01010100100", -- t[676] = 0
      "0" when "01010100101", -- t[677] = 0
      "0" when "01010100110", -- t[678] = 0
      "0" when "01010100111", -- t[679] = 0
      "0" when "01010101000", -- t[680] = 0
      "0" when "01010101001", -- t[681] = 0
      "0" when "01010101010", -- t[682] = 0
      "0" when "01010101011", -- t[683] = 0
      "0" when "01010101100", -- t[684] = 0
      "0" when "01010101101", -- t[685] = 0
      "0" when "01010101110", -- t[686] = 0
      "0" when "01010101111", -- t[687] = 0
      "0" when "01010110000", -- t[688] = 0
      "0" when "01010110001", -- t[689] = 0
      "0" when "01010110010", -- t[690] = 0
      "0" when "01010110011", -- t[691] = 0
      "0" when "01010110100", -- t[692] = 0
      "0" when "01010110101", -- t[693] = 0
      "0" when "01010110110", -- t[694] = 0
      "0" when "01010110111", -- t[695] = 0
      "0" when "01010111000", -- t[696] = 0
      "0" when "01010111001", -- t[697] = 0
      "0" when "01010111010", -- t[698] = 0
      "0" when "01010111011", -- t[699] = 0
      "0" when "01010111100", -- t[700] = 0
      "0" when "01010111101", -- t[701] = 0
      "0" when "01010111110", -- t[702] = 0
      "0" when "01010111111", -- t[703] = 0
      "0" when "01011000000", -- t[704] = 0
      "0" when "01011000001", -- t[705] = 0
      "0" when "01011000010", -- t[706] = 0
      "0" when "01011000011", -- t[707] = 0
      "0" when "01011000100", -- t[708] = 0
      "0" when "01011000101", -- t[709] = 0
      "0" when "01011000110", -- t[710] = 0
      "0" when "01011000111", -- t[711] = 0
      "0" when "01011001000", -- t[712] = 0
      "0" when "01011001001", -- t[713] = 0
      "0" when "01011001010", -- t[714] = 0
      "0" when "01011001011", -- t[715] = 0
      "0" when "01011001100", -- t[716] = 0
      "0" when "01011001101", -- t[717] = 0
      "0" when "01011001110", -- t[718] = 0
      "0" when "01011001111", -- t[719] = 0
      "0" when "01011010000", -- t[720] = 0
      "0" when "01011010001", -- t[721] = 0
      "0" when "01011010010", -- t[722] = 0
      "0" when "01011010011", -- t[723] = 0
      "0" when "01011010100", -- t[724] = 0
      "0" when "01011010101", -- t[725] = 0
      "0" when "01011010110", -- t[726] = 0
      "0" when "01011010111", -- t[727] = 0
      "0" when "01011011000", -- t[728] = 0
      "0" when "01011011001", -- t[729] = 0
      "0" when "01011011010", -- t[730] = 0
      "0" when "01011011011", -- t[731] = 0
      "0" when "01011011100", -- t[732] = 0
      "0" when "01011011101", -- t[733] = 0
      "0" when "01011011110", -- t[734] = 0
      "0" when "01011011111", -- t[735] = 0
      "0" when "01011100000", -- t[736] = 0
      "0" when "01011100001", -- t[737] = 0
      "0" when "01011100010", -- t[738] = 0
      "0" when "01011100011", -- t[739] = 0
      "0" when "01011100100", -- t[740] = 0
      "0" when "01011100101", -- t[741] = 0
      "0" when "01011100110", -- t[742] = 0
      "0" when "01011100111", -- t[743] = 0
      "0" when "01011101000", -- t[744] = 0
      "0" when "01011101001", -- t[745] = 0
      "0" when "01011101010", -- t[746] = 0
      "0" when "01011101011", -- t[747] = 0
      "0" when "01011101100", -- t[748] = 0
      "0" when "01011101101", -- t[749] = 0
      "0" when "01011101110", -- t[750] = 0
      "0" when "01011101111", -- t[751] = 0
      "0" when "01011110000", -- t[752] = 0
      "0" when "01011110001", -- t[753] = 0
      "0" when "01011110010", -- t[754] = 0
      "0" when "01011110011", -- t[755] = 0
      "0" when "01011110100", -- t[756] = 0
      "0" when "01011110101", -- t[757] = 0
      "0" when "01011110110", -- t[758] = 0
      "0" when "01011110111", -- t[759] = 0
      "0" when "01011111000", -- t[760] = 0
      "0" when "01011111001", -- t[761] = 0
      "0" when "01011111010", -- t[762] = 0
      "0" when "01011111011", -- t[763] = 0
      "0" when "01011111100", -- t[764] = 0
      "0" when "01011111101", -- t[765] = 0
      "0" when "01011111110", -- t[766] = 0
      "0" when "01011111111", -- t[767] = 0
      "0" when "01100000000", -- t[768] = 0
      "0" when "01100000001", -- t[769] = 0
      "0" when "01100000010", -- t[770] = 0
      "0" when "01100000011", -- t[771] = 0
      "0" when "01100000100", -- t[772] = 0
      "0" when "01100000101", -- t[773] = 0
      "0" when "01100000110", -- t[774] = 0
      "0" when "01100000111", -- t[775] = 0
      "0" when "01100001000", -- t[776] = 0
      "0" when "01100001001", -- t[777] = 0
      "0" when "01100001010", -- t[778] = 0
      "0" when "01100001011", -- t[779] = 0
      "0" when "01100001100", -- t[780] = 0
      "0" when "01100001101", -- t[781] = 0
      "0" when "01100001110", -- t[782] = 0
      "0" when "01100001111", -- t[783] = 0
      "0" when "01100010000", -- t[784] = 0
      "0" when "01100010001", -- t[785] = 0
      "0" when "01100010010", -- t[786] = 0
      "0" when "01100010011", -- t[787] = 0
      "0" when "01100010100", -- t[788] = 0
      "0" when "01100010101", -- t[789] = 0
      "0" when "01100010110", -- t[790] = 0
      "0" when "01100010111", -- t[791] = 0
      "0" when "01100011000", -- t[792] = 0
      "0" when "01100011001", -- t[793] = 0
      "0" when "01100011010", -- t[794] = 0
      "0" when "01100011011", -- t[795] = 0
      "0" when "01100011100", -- t[796] = 0
      "0" when "01100011101", -- t[797] = 0
      "0" when "01100011110", -- t[798] = 0
      "0" when "01100011111", -- t[799] = 0
      "0" when "01100100000", -- t[800] = 0
      "0" when "01100100001", -- t[801] = 0
      "0" when "01100100010", -- t[802] = 0
      "0" when "01100100011", -- t[803] = 0
      "0" when "01100100100", -- t[804] = 0
      "0" when "01100100101", -- t[805] = 0
      "0" when "01100100110", -- t[806] = 0
      "0" when "01100100111", -- t[807] = 0
      "0" when "01100101000", -- t[808] = 0
      "0" when "01100101001", -- t[809] = 0
      "0" when "01100101010", -- t[810] = 0
      "0" when "01100101011", -- t[811] = 0
      "0" when "01100101100", -- t[812] = 0
      "0" when "01100101101", -- t[813] = 0
      "0" when "01100101110", -- t[814] = 0
      "0" when "01100101111", -- t[815] = 0
      "0" when "01100110000", -- t[816] = 0
      "0" when "01100110001", -- t[817] = 0
      "0" when "01100110010", -- t[818] = 0
      "0" when "01100110011", -- t[819] = 0
      "0" when "01100110100", -- t[820] = 0
      "0" when "01100110101", -- t[821] = 0
      "0" when "01100110110", -- t[822] = 0
      "0" when "01100110111", -- t[823] = 0
      "0" when "01100111000", -- t[824] = 0
      "0" when "01100111001", -- t[825] = 0
      "0" when "01100111010", -- t[826] = 0
      "0" when "01100111011", -- t[827] = 0
      "0" when "01100111100", -- t[828] = 0
      "0" when "01100111101", -- t[829] = 0
      "0" when "01100111110", -- t[830] = 0
      "0" when "01100111111", -- t[831] = 0
      "0" when "01101000000", -- t[832] = 0
      "0" when "01101000001", -- t[833] = 0
      "0" when "01101000010", -- t[834] = 0
      "0" when "01101000011", -- t[835] = 0
      "0" when "01101000100", -- t[836] = 0
      "0" when "01101000101", -- t[837] = 0
      "0" when "01101000110", -- t[838] = 0
      "0" when "01101000111", -- t[839] = 0
      "0" when "01101001000", -- t[840] = 0
      "0" when "01101001001", -- t[841] = 0
      "0" when "01101001010", -- t[842] = 0
      "0" when "01101001011", -- t[843] = 0
      "0" when "01101001100", -- t[844] = 0
      "0" when "01101001101", -- t[845] = 0
      "0" when "01101001110", -- t[846] = 0
      "0" when "01101001111", -- t[847] = 0
      "0" when "01101010000", -- t[848] = 0
      "0" when "01101010001", -- t[849] = 0
      "0" when "01101010010", -- t[850] = 0
      "0" when "01101010011", -- t[851] = 0
      "0" when "01101010100", -- t[852] = 0
      "0" when "01101010101", -- t[853] = 0
      "0" when "01101010110", -- t[854] = 0
      "0" when "01101010111", -- t[855] = 0
      "0" when "01101011000", -- t[856] = 0
      "0" when "01101011001", -- t[857] = 0
      "0" when "01101011010", -- t[858] = 0
      "0" when "01101011011", -- t[859] = 0
      "0" when "01101011100", -- t[860] = 0
      "0" when "01101011101", -- t[861] = 0
      "0" when "01101011110", -- t[862] = 0
      "0" when "01101011111", -- t[863] = 0
      "0" when "01101100000", -- t[864] = 0
      "0" when "01101100001", -- t[865] = 0
      "0" when "01101100010", -- t[866] = 0
      "0" when "01101100011", -- t[867] = 0
      "0" when "01101100100", -- t[868] = 0
      "0" when "01101100101", -- t[869] = 0
      "0" when "01101100110", -- t[870] = 0
      "0" when "01101100111", -- t[871] = 0
      "0" when "01101101000", -- t[872] = 0
      "0" when "01101101001", -- t[873] = 0
      "0" when "01101101010", -- t[874] = 0
      "0" when "01101101011", -- t[875] = 0
      "0" when "01101101100", -- t[876] = 0
      "0" when "01101101101", -- t[877] = 0
      "0" when "01101101110", -- t[878] = 0
      "0" when "01101101111", -- t[879] = 0
      "0" when "01101110000", -- t[880] = 0
      "0" when "01101110001", -- t[881] = 0
      "0" when "01101110010", -- t[882] = 0
      "0" when "01101110011", -- t[883] = 0
      "0" when "01101110100", -- t[884] = 0
      "0" when "01101110101", -- t[885] = 0
      "0" when "01101110110", -- t[886] = 0
      "0" when "01101110111", -- t[887] = 0
      "0" when "01101111000", -- t[888] = 0
      "0" when "01101111001", -- t[889] = 0
      "0" when "01101111010", -- t[890] = 0
      "0" when "01101111011", -- t[891] = 0
      "0" when "01101111100", -- t[892] = 0
      "0" when "01101111101", -- t[893] = 0
      "0" when "01101111110", -- t[894] = 0
      "0" when "01101111111", -- t[895] = 0
      "0" when "01110000000", -- t[896] = 0
      "0" when "01110000001", -- t[897] = 0
      "0" when "01110000010", -- t[898] = 0
      "0" when "01110000011", -- t[899] = 0
      "0" when "01110000100", -- t[900] = 0
      "0" when "01110000101", -- t[901] = 0
      "0" when "01110000110", -- t[902] = 0
      "0" when "01110000111", -- t[903] = 0
      "0" when "01110001000", -- t[904] = 0
      "0" when "01110001001", -- t[905] = 0
      "0" when "01110001010", -- t[906] = 0
      "0" when "01110001011", -- t[907] = 0
      "0" when "01110001100", -- t[908] = 0
      "0" when "01110001101", -- t[909] = 0
      "0" when "01110001110", -- t[910] = 0
      "0" when "01110001111", -- t[911] = 0
      "0" when "01110010000", -- t[912] = 0
      "0" when "01110010001", -- t[913] = 0
      "0" when "01110010010", -- t[914] = 0
      "0" when "01110010011", -- t[915] = 0
      "0" when "01110010100", -- t[916] = 0
      "0" when "01110010101", -- t[917] = 0
      "0" when "01110010110", -- t[918] = 0
      "0" when "01110010111", -- t[919] = 0
      "0" when "01110011000", -- t[920] = 0
      "0" when "01110011001", -- t[921] = 0
      "0" when "01110011010", -- t[922] = 0
      "0" when "01110011011", -- t[923] = 0
      "0" when "01110011100", -- t[924] = 0
      "0" when "01110011101", -- t[925] = 0
      "0" when "01110011110", -- t[926] = 0
      "0" when "01110011111", -- t[927] = 0
      "0" when "01110100000", -- t[928] = 0
      "0" when "01110100001", -- t[929] = 0
      "0" when "01110100010", -- t[930] = 0
      "0" when "01110100011", -- t[931] = 0
      "0" when "01110100100", -- t[932] = 0
      "0" when "01110100101", -- t[933] = 0
      "0" when "01110100110", -- t[934] = 0
      "0" when "01110100111", -- t[935] = 0
      "0" when "01110101000", -- t[936] = 0
      "0" when "01110101001", -- t[937] = 0
      "0" when "01110101010", -- t[938] = 0
      "0" when "01110101011", -- t[939] = 0
      "0" when "01110101100", -- t[940] = 0
      "0" when "01110101101", -- t[941] = 0
      "0" when "01110101110", -- t[942] = 0
      "0" when "01110101111", -- t[943] = 0
      "0" when "01110110000", -- t[944] = 0
      "0" when "01110110001", -- t[945] = 0
      "0" when "01110110010", -- t[946] = 0
      "0" when "01110110011", -- t[947] = 0
      "0" when "01110110100", -- t[948] = 0
      "0" when "01110110101", -- t[949] = 0
      "0" when "01110110110", -- t[950] = 0
      "0" when "01110110111", -- t[951] = 0
      "0" when "01110111000", -- t[952] = 0
      "0" when "01110111001", -- t[953] = 0
      "0" when "01110111010", -- t[954] = 0
      "0" when "01110111011", -- t[955] = 0
      "0" when "01110111100", -- t[956] = 0
      "1" when "01110111101", -- t[957] = 1
      "1" when "01110111110", -- t[958] = 1
      "1" when "01110111111", -- t[959] = 1
      "1" when "01111000000", -- t[960] = 1
      "1" when "01111000001", -- t[961] = 1
      "1" when "01111000010", -- t[962] = 1
      "1" when "01111000011", -- t[963] = 1
      "1" when "01111000100", -- t[964] = 1
      "1" when "01111000101", -- t[965] = 1
      "1" when "01111000110", -- t[966] = 1
      "1" when "01111000111", -- t[967] = 1
      "1" when "01111001000", -- t[968] = 1
      "1" when "01111001001", -- t[969] = 1
      "1" when "01111001010", -- t[970] = 1
      "1" when "01111001011", -- t[971] = 1
      "1" when "01111001100", -- t[972] = 1
      "1" when "01111001101", -- t[973] = 1
      "1" when "01111001110", -- t[974] = 1
      "1" when "01111001111", -- t[975] = 1
      "1" when "01111010000", -- t[976] = 1
      "1" when "01111010001", -- t[977] = 1
      "1" when "01111010010", -- t[978] = 1
      "1" when "01111010011", -- t[979] = 1
      "1" when "01111010100", -- t[980] = 1
      "1" when "01111010101", -- t[981] = 1
      "1" when "01111010110", -- t[982] = 1
      "1" when "01111010111", -- t[983] = 1
      "1" when "01111011000", -- t[984] = 1
      "1" when "01111011001", -- t[985] = 1
      "1" when "01111011010", -- t[986] = 1
      "1" when "01111011011", -- t[987] = 1
      "1" when "01111011100", -- t[988] = 1
      "1" when "01111011101", -- t[989] = 1
      "1" when "01111011110", -- t[990] = 1
      "1" when "01111011111", -- t[991] = 1
      "1" when "01111100000", -- t[992] = 1
      "1" when "01111100001", -- t[993] = 1
      "1" when "01111100010", -- t[994] = 1
      "1" when "01111100011", -- t[995] = 1
      "1" when "01111100100", -- t[996] = 1
      "1" when "01111100101", -- t[997] = 1
      "1" when "01111100110", -- t[998] = 1
      "1" when "01111100111", -- t[999] = 1
      "1" when "01111101000", -- t[1000] = 1
      "1" when "01111101001", -- t[1001] = 1
      "1" when "01111101010", -- t[1002] = 1
      "1" when "01111101011", -- t[1003] = 1
      "1" when "01111101100", -- t[1004] = 1
      "1" when "01111101101", -- t[1005] = 1
      "1" when "01111101110", -- t[1006] = 1
      "1" when "01111101111", -- t[1007] = 1
      "1" when "01111110000", -- t[1008] = 1
      "1" when "01111110001", -- t[1009] = 1
      "1" when "01111110010", -- t[1010] = 1
      "1" when "01111110011", -- t[1011] = 1
      "1" when "01111110100", -- t[1012] = 1
      "1" when "01111110101", -- t[1013] = 1
      "1" when "01111110110", -- t[1014] = 1
      "1" when "01111110111", -- t[1015] = 1
      "1" when "01111111000", -- t[1016] = 1
      "1" when "01111111001", -- t[1017] = 1
      "1" when "01111111010", -- t[1018] = 1
      "1" when "01111111011", -- t[1019] = 1
      "1" when "01111111100", -- t[1020] = 1
      "1" when "01111111101", -- t[1021] = 1
      "1" when "01111111110", -- t[1022] = 1
      "1" when "01111111111", -- t[1023] = 1
      "-" when others;
end architecture;


-- MultiPartite: LNS addition function: [-8.0 0.0[ -> [0.0 2.0[
-- wI = 10 bits
-- wO = 8 bits
-- Decomposition: 6, 4 / 5, 3 / 2, 2
-- Guard bits: 3
-- Size: 1072 = 11.2^6 + 5.2^6 + 3.2^4

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSAdd_MPT_T2_7 is
  component LNSAdd_MPT_T2_7_tiv is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSAdd_MPT_T2_7_to1 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSAdd_MPT_T2_7_to0 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSAdd_MPT_T2_7_to1_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSAdd_MPT_T2_7_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_7_tiv is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7_tiv is
begin
  with x select
    r <=
      "00000001011" when "000000", -- t[0] = 11
      "00000001011" when "000001", -- t[1] = 11
      "00000001100" when "000010", -- t[2] = 12
      "00000001100" when "000011", -- t[3] = 12
      "00000001101" when "000100", -- t[4] = 13
      "00000001110" when "000101", -- t[5] = 14
      "00000001111" when "000110", -- t[6] = 15
      "00000001111" when "000111", -- t[7] = 15
      "00000010000" when "001000", -- t[8] = 16
      "00000010010" when "001001", -- t[9] = 18
      "00000010011" when "001010", -- t[10] = 19
      "00000010100" when "001011", -- t[11] = 20
      "00000010101" when "001100", -- t[12] = 21
      "00000010111" when "001101", -- t[13] = 23
      "00000011001" when "001110", -- t[14] = 25
      "00000011010" when "001111", -- t[15] = 26
      "00000011100" when "010000", -- t[16] = 28
      "00000011111" when "010001", -- t[17] = 31
      "00000100001" when "010010", -- t[18] = 33
      "00000100011" when "010011", -- t[19] = 35
      "00000100110" when "010100", -- t[20] = 38
      "00000101001" when "010101", -- t[21] = 41
      "00000101100" when "010110", -- t[22] = 44
      "00000110000" when "010111", -- t[23] = 48
      "00000110100" when "011000", -- t[24] = 52
      "00000111000" when "011001", -- t[25] = 56
      "00000111101" when "011010", -- t[26] = 61
      "00001000010" when "011011", -- t[27] = 66
      "00001000111" when "011100", -- t[28] = 71
      "00001001101" when "011101", -- t[29] = 77
      "00001010011" when "011110", -- t[30] = 83
      "00001011010" when "011111", -- t[31] = 90
      "00001100010" when "100000", -- t[32] = 98
      "00001101010" when "100001", -- t[33] = 106
      "00001110011" when "100010", -- t[34] = 115
      "00001111100" when "100011", -- t[35] = 124
      "00010000111" when "100100", -- t[36] = 135
      "00010010010" when "100101", -- t[37] = 146
      "00010011110" when "100110", -- t[38] = 158
      "00010101011" when "100111", -- t[39] = 171
      "00010111001" when "101000", -- t[40] = 185
      "00011001001" when "101001", -- t[41] = 201
      "00011011001" when "101010", -- t[42] = 217
      "00011101011" when "101011", -- t[43] = 235
      "00011111110" when "101100", -- t[44] = 254
      "00100010011" when "101101", -- t[45] = 275
      "00100101001" when "101110", -- t[46] = 297
      "00101000001" when "101111", -- t[47] = 321
      "00101011011" when "110000", -- t[48] = 347
      "00101110110" when "110001", -- t[49] = 374
      "00110010011" when "110010", -- t[50] = 403
      "00110110011" when "110011", -- t[51] = 435
      "00111010100" when "110100", -- t[52] = 468
      "00111110111" when "110101", -- t[53] = 503
      "01000011101" when "110110", -- t[54] = 541
      "01001000101" when "110111", -- t[55] = 581
      "01001110000" when "111000", -- t[56] = 624
      "01010011101" when "111001", -- t[57] = 669
      "01011001101" when "111010", -- t[58] = 717
      "01011111111" when "111011", -- t[59] = 767
      "01100110100" when "111100", -- t[60] = 820
      "01101101100" when "111101", -- t[61] = 876
      "01110100110" when "111110", -- t[62] = 934
      "01111100011" when "111111", -- t[63] = 995
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_7_to1 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7_to1 is
begin
  with x select
    r <=
      "00000" when "000000", -- t[0] = 0
      "00000" when "000001", -- t[1] = 0
      "00000" when "000010", -- t[2] = 0
      "00000" when "000011", -- t[3] = 0
      "00000" when "000100", -- t[4] = 0
      "00000" when "000101", -- t[5] = 0
      "00000" when "000110", -- t[6] = 0
      "00000" when "000111", -- t[7] = 0
      "00000" when "001000", -- t[8] = 0
      "00000" when "001001", -- t[9] = 0
      "00000" when "001010", -- t[10] = 0
      "00000" when "001011", -- t[11] = 0
      "00000" when "001100", -- t[12] = 0
      "00000" when "001101", -- t[13] = 0
      "00000" when "001110", -- t[14] = 0
      "00000" when "001111", -- t[15] = 0
      "00000" when "010000", -- t[16] = 0
      "00000" when "010001", -- t[17] = 0
      "00000" when "010010", -- t[18] = 0
      "00000" when "010011", -- t[19] = 0
      "00000" when "010100", -- t[20] = 0
      "00001" when "010101", -- t[21] = 1
      "00000" when "010110", -- t[22] = 0
      "00001" when "010111", -- t[23] = 1
      "00000" when "011000", -- t[24] = 0
      "00001" when "011001", -- t[25] = 1
      "00000" when "011010", -- t[26] = 0
      "00001" when "011011", -- t[27] = 1
      "00000" when "011100", -- t[28] = 0
      "00010" when "011101", -- t[29] = 2
      "00000" when "011110", -- t[30] = 0
      "00010" when "011111", -- t[31] = 2
      "00001" when "100000", -- t[32] = 1
      "00011" when "100001", -- t[33] = 3
      "00001" when "100010", -- t[34] = 1
      "00011" when "100011", -- t[35] = 3
      "00001" when "100100", -- t[36] = 1
      "00100" when "100101", -- t[37] = 4
      "00001" when "100110", -- t[38] = 1
      "00100" when "100111", -- t[39] = 4
      "00001" when "101000", -- t[40] = 1
      "00101" when "101001", -- t[41] = 5
      "00010" when "101010", -- t[42] = 2
      "00110" when "101011", -- t[43] = 6
      "00010" when "101100", -- t[44] = 2
      "00111" when "101101", -- t[45] = 7
      "00010" when "101110", -- t[46] = 2
      "01000" when "101111", -- t[47] = 8
      "00011" when "110000", -- t[48] = 3
      "01010" when "110001", -- t[49] = 10
      "00011" when "110010", -- t[50] = 3
      "01011" when "110011", -- t[51] = 11
      "00100" when "110100", -- t[52] = 4
      "01101" when "110101", -- t[53] = 13
      "00100" when "110110", -- t[54] = 4
      "01110" when "110111", -- t[55] = 14
      "00101" when "111000", -- t[56] = 5
      "10000" when "111001", -- t[57] = 16
      "00110" when "111010", -- t[58] = 6
      "10010" when "111011", -- t[59] = 18
      "00110" when "111100", -- t[60] = 6
      "10100" when "111101", -- t[61] = 20
      "00111" when "111110", -- t[62] = 7
      "10110" when "111111", -- t[63] = 22
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSAdd_MPT_T2_7_to0 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7_to0 is
begin
  with x select
    r <=
      "000" when "0000", -- t[0] = 0
      "000" when "0001", -- t[1] = 0
      "000" when "0010", -- t[2] = 0
      "000" when "0011", -- t[3] = 0
      "000" when "0100", -- t[4] = 0
      "000" when "0101", -- t[5] = 0
      "000" when "0110", -- t[6] = 0
      "000" when "0111", -- t[7] = 0
      "000" when "1000", -- t[8] = 0
      "001" when "1001", -- t[9] = 1
      "000" when "1010", -- t[10] = 0
      "001" when "1011", -- t[11] = 1
      "001" when "1100", -- t[12] = 1
      "011" when "1101", -- t[13] = 3
      "001" when "1110", -- t[14] = 1
      "100" when "1111", -- t[15] = 4
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_7.all;

entity LNSAdd_MPT_T2_7_to1_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSAdd_MPT_T2_7_to1
    port map( x => in_t,
              r => out_t );

  r(10 downto 5) <= (10 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_7.all;

entity LNSAdd_MPT_T2_7_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSAdd_MPT_T2_7_to0
    port map( x => in_t,
              r => out_t );

  r(10 downto 3) <= (10 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSAdd_MPT_T2_7.all;

entity LNSAdd_MPT_T2_7 is
  port( x : in  std_logic_vector(9 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_T2_7 is
  signal in_tiv  : std_logic_vector(5 downto 0);
  signal out_tiv : std_logic_vector(10 downto 0);
  signal a1      : std_logic_vector(4 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(10 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(10 downto 0);
  signal sum     : std_logic_vector(10 downto 0);
begin
  in_tiv <= x(9 downto 4);
  inst_tiv : LNSAdd_MPT_T2_7_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(9 downto 5);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSAdd_MPT_T2_7_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(9 downto 7);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSAdd_MPT_T2_7_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(10 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_7.all;

entity LNSAdd_MPT_7 is
  port( x : in  std_logic_vector(10 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSAdd_MPT_7 is
  signal out_t1 : std_logic_vector(0 downto 0);
  signal out_t2 : std_logic_vector(7 downto 0);
begin
  inst_t1 : LNSAdd_MPT_T1_7
    port map( x => x,
              r => out_t1 );

  inst_t2 : LNSAdd_MPT_T2_7
    port map( x => x(9 downto 0),
              r => out_t2 );

  r <= out_t2 when x(10 downto 10) = (10 downto 10 => '1') else
       (7 downto 1 => '0') & out_t1;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnsadd_mpt_7.all;
use fplib.pkg_misc.all;

entity LNSAdd_MPT_7_Clk is
  port( x   : in  std_logic_vector(10 downto 0);
        r   : out std_logic_vector(7 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSAdd_MPT_7_Clk is
  signal x_1  : std_logic_vector(10 downto 0);
  signal x_10 : std_logic_vector(10 downto 0);

  signal out_t1_1  : std_logic_vector(0 downto 0);
  signal out_t1_10 : std_logic_vector(0 downto 0);
  signal out_t2_10 : std_logic_vector(7 downto 0);
begin
  x_1 <= x;

  inst_t1 : LNSAdd_MPT_T1_7
    port map( x => x_1,
              r => out_t1_1 );

  out_t1_delay : Delay
    generic map ( w => 1,
                  n => 0 )
    port map ( input  => out_t1_1,
               output => out_t1_10,
               clk    => clk );

  inst_t2 : LNSAdd_MPT_T2_7
    port map( x => x(9 downto 0),
              r => out_t2_10 );

  x_delay : Delay
    generic map ( w => 11,
                  n => 0 )
    port map ( input  => x_1,
               output => x_10,
               clk    => clk );

  r <= out_t2_10 when x_10(10 downto 10) = (10 downto 10 => '1') else
       (7 downto 1 => '0') & out_t1_10;
end architecture;
