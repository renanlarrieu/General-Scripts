-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of MultiPartiteSubtracter object for LNS arithmetic in base 2.0 with 8-bit integer part and 13-bit fractional part
-- wI = 17 bits
-- wO = 17 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnssub_mpt_13 is
  component LNSSub_MPT_T0_13 is
    port( x : in  std_logic_vector(16 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T1_13 is
    port( x : in  std_logic_vector(14 downto 0);
          r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_Clk is
    port( x   : in  std_logic_vector(14 downto 0);
          r   : out std_logic_vector(9 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T2_13 is
    port( x : in  std_logic_vector(13 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_Clk is
    port( x   : in  std_logic_vector(13 downto 0);
          r   : out std_logic_vector(11 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T3_13 is
    port( x : in  std_logic_vector(12 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_Clk is
    port( x   : in  std_logic_vector(12 downto 0);
          r   : out std_logic_vector(11 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T4_13 is
    port( x : in  std_logic_vector(11 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_Clk is
    port( x   : in  std_logic_vector(11 downto 0);
          r   : out std_logic_vector(11 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T5_13 is
    port( x : in  std_logic_vector(10 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T5_13_Clk is
    port( x   : in  std_logic_vector(10 downto 0);
          r   : out std_logic_vector(11 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T6_13 is
    port( x : in  std_logic_vector(9 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T6_13_Clk is
    port( x   : in  std_logic_vector(9 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T7_13 is
    port( x : in  std_logic_vector(8 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T7_13_Clk is
    port( x   : in  std_logic_vector(8 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T8_13 is
    port( x : in  std_logic_vector(7 downto 0);
          r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MPT_T8_13_Clk is
    port( x   : in  std_logic_vector(7 downto 0);
          r   : out std_logic_vector(9 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T9_13 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T9_13_Clk is
    port( x   : in  std_logic_vector(6 downto 0);
          r   : out std_logic_vector(8 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T10_13 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T10_13_Clk is
    port( x   : in  std_logic_vector(5 downto 0);
          r   : out std_logic_vector(7 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T11_13 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T11_13_Clk is
    port( x   : in  std_logic_vector(4 downto 0);
          r   : out std_logic_vector(7 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T12_13 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T12_13_Clk is
    port( x   : in  std_logic_vector(3 downto 0);
          r   : out std_logic_vector(6 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T13_13 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T13_13_Clk is
    port( x   : in  std_logic_vector(3 downto 0);
          r   : out std_logic_vector(6 downto 0);
          clk : in  std_logic );
  end component;
end package;


-- SimpleTable: LNS subtraction function: [-16.0 0.0[ -> [0.0 1.0[
-- (bounded to [-16.0; -8.0[)
-- wI = 17 bits
-- wO = 7 bits

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T0_13 is
  port( x : in  std_logic_vector(16 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T0_13 is
begin
  with x select
    r <=
      "0000000" when "00000000000000000", -- t[0] = 0
      "0000000" when "00000000000000001", -- t[1] = 0
      "0000000" when "00000000000000010", -- t[2] = 0
      "0000000" when "00000000000000011", -- t[3] = 0
      "0000000" when "00000000000000100", -- t[4] = 0
      "0000000" when "00000000000000101", -- t[5] = 0
      "0000000" when "00000000000000110", -- t[6] = 0
      "0000000" when "00000000000000111", -- t[7] = 0
      "0000000" when "00000000000001000", -- t[8] = 0
      "0000000" when "00000000000001001", -- t[9] = 0
      "0000000" when "00000000000001010", -- t[10] = 0
      "0000000" when "00000000000001011", -- t[11] = 0
      "0000000" when "00000000000001100", -- t[12] = 0
      "0000000" when "00000000000001101", -- t[13] = 0
      "0000000" when "00000000000001110", -- t[14] = 0
      "0000000" when "00000000000001111", -- t[15] = 0
      "0000000" when "00000000000010000", -- t[16] = 0
      "0000000" when "00000000000010001", -- t[17] = 0
      "0000000" when "00000000000010010", -- t[18] = 0
      "0000000" when "00000000000010011", -- t[19] = 0
      "0000000" when "00000000000010100", -- t[20] = 0
      "0000000" when "00000000000010101", -- t[21] = 0
      "0000000" when "00000000000010110", -- t[22] = 0
      "0000000" when "00000000000010111", -- t[23] = 0
      "0000000" when "00000000000011000", -- t[24] = 0
      "0000000" when "00000000000011001", -- t[25] = 0
      "0000000" when "00000000000011010", -- t[26] = 0
      "0000000" when "00000000000011011", -- t[27] = 0
      "0000000" when "00000000000011100", -- t[28] = 0
      "0000000" when "00000000000011101", -- t[29] = 0
      "0000000" when "00000000000011110", -- t[30] = 0
      "0000000" when "00000000000011111", -- t[31] = 0
      "0000000" when "00000000000100000", -- t[32] = 0
      "0000000" when "00000000000100001", -- t[33] = 0
      "0000000" when "00000000000100010", -- t[34] = 0
      "0000000" when "00000000000100011", -- t[35] = 0
      "0000000" when "00000000000100100", -- t[36] = 0
      "0000000" when "00000000000100101", -- t[37] = 0
      "0000000" when "00000000000100110", -- t[38] = 0
      "0000000" when "00000000000100111", -- t[39] = 0
      "0000000" when "00000000000101000", -- t[40] = 0
      "0000000" when "00000000000101001", -- t[41] = 0
      "0000000" when "00000000000101010", -- t[42] = 0
      "0000000" when "00000000000101011", -- t[43] = 0
      "0000000" when "00000000000101100", -- t[44] = 0
      "0000000" when "00000000000101101", -- t[45] = 0
      "0000000" when "00000000000101110", -- t[46] = 0
      "0000000" when "00000000000101111", -- t[47] = 0
      "0000000" when "00000000000110000", -- t[48] = 0
      "0000000" when "00000000000110001", -- t[49] = 0
      "0000000" when "00000000000110010", -- t[50] = 0
      "0000000" when "00000000000110011", -- t[51] = 0
      "0000000" when "00000000000110100", -- t[52] = 0
      "0000000" when "00000000000110101", -- t[53] = 0
      "0000000" when "00000000000110110", -- t[54] = 0
      "0000000" when "00000000000110111", -- t[55] = 0
      "0000000" when "00000000000111000", -- t[56] = 0
      "0000000" when "00000000000111001", -- t[57] = 0
      "0000000" when "00000000000111010", -- t[58] = 0
      "0000000" when "00000000000111011", -- t[59] = 0
      "0000000" when "00000000000111100", -- t[60] = 0
      "0000000" when "00000000000111101", -- t[61] = 0
      "0000000" when "00000000000111110", -- t[62] = 0
      "0000000" when "00000000000111111", -- t[63] = 0
      "0000000" when "00000000001000000", -- t[64] = 0
      "0000000" when "00000000001000001", -- t[65] = 0
      "0000000" when "00000000001000010", -- t[66] = 0
      "0000000" when "00000000001000011", -- t[67] = 0
      "0000000" when "00000000001000100", -- t[68] = 0
      "0000000" when "00000000001000101", -- t[69] = 0
      "0000000" when "00000000001000110", -- t[70] = 0
      "0000000" when "00000000001000111", -- t[71] = 0
      "0000000" when "00000000001001000", -- t[72] = 0
      "0000000" when "00000000001001001", -- t[73] = 0
      "0000000" when "00000000001001010", -- t[74] = 0
      "0000000" when "00000000001001011", -- t[75] = 0
      "0000000" when "00000000001001100", -- t[76] = 0
      "0000000" when "00000000001001101", -- t[77] = 0
      "0000000" when "00000000001001110", -- t[78] = 0
      "0000000" when "00000000001001111", -- t[79] = 0
      "0000000" when "00000000001010000", -- t[80] = 0
      "0000000" when "00000000001010001", -- t[81] = 0
      "0000000" when "00000000001010010", -- t[82] = 0
      "0000000" when "00000000001010011", -- t[83] = 0
      "0000000" when "00000000001010100", -- t[84] = 0
      "0000000" when "00000000001010101", -- t[85] = 0
      "0000000" when "00000000001010110", -- t[86] = 0
      "0000000" when "00000000001010111", -- t[87] = 0
      "0000000" when "00000000001011000", -- t[88] = 0
      "0000000" when "00000000001011001", -- t[89] = 0
      "0000000" when "00000000001011010", -- t[90] = 0
      "0000000" when "00000000001011011", -- t[91] = 0
      "0000000" when "00000000001011100", -- t[92] = 0
      "0000000" when "00000000001011101", -- t[93] = 0
      "0000000" when "00000000001011110", -- t[94] = 0
      "0000000" when "00000000001011111", -- t[95] = 0
      "0000000" when "00000000001100000", -- t[96] = 0
      "0000000" when "00000000001100001", -- t[97] = 0
      "0000000" when "00000000001100010", -- t[98] = 0
      "0000000" when "00000000001100011", -- t[99] = 0
      "0000000" when "00000000001100100", -- t[100] = 0
      "0000000" when "00000000001100101", -- t[101] = 0
      "0000000" when "00000000001100110", -- t[102] = 0
      "0000000" when "00000000001100111", -- t[103] = 0
      "0000000" when "00000000001101000", -- t[104] = 0
      "0000000" when "00000000001101001", -- t[105] = 0
      "0000000" when "00000000001101010", -- t[106] = 0
      "0000000" when "00000000001101011", -- t[107] = 0
      "0000000" when "00000000001101100", -- t[108] = 0
      "0000000" when "00000000001101101", -- t[109] = 0
      "0000000" when "00000000001101110", -- t[110] = 0
      "0000000" when "00000000001101111", -- t[111] = 0
      "0000000" when "00000000001110000", -- t[112] = 0
      "0000000" when "00000000001110001", -- t[113] = 0
      "0000000" when "00000000001110010", -- t[114] = 0
      "0000000" when "00000000001110011", -- t[115] = 0
      "0000000" when "00000000001110100", -- t[116] = 0
      "0000000" when "00000000001110101", -- t[117] = 0
      "0000000" when "00000000001110110", -- t[118] = 0
      "0000000" when "00000000001110111", -- t[119] = 0
      "0000000" when "00000000001111000", -- t[120] = 0
      "0000000" when "00000000001111001", -- t[121] = 0
      "0000000" when "00000000001111010", -- t[122] = 0
      "0000000" when "00000000001111011", -- t[123] = 0
      "0000000" when "00000000001111100", -- t[124] = 0
      "0000000" when "00000000001111101", -- t[125] = 0
      "0000000" when "00000000001111110", -- t[126] = 0
      "0000000" when "00000000001111111", -- t[127] = 0
      "0000000" when "00000000010000000", -- t[128] = 0
      "0000000" when "00000000010000001", -- t[129] = 0
      "0000000" when "00000000010000010", -- t[130] = 0
      "0000000" when "00000000010000011", -- t[131] = 0
      "0000000" when "00000000010000100", -- t[132] = 0
      "0000000" when "00000000010000101", -- t[133] = 0
      "0000000" when "00000000010000110", -- t[134] = 0
      "0000000" when "00000000010000111", -- t[135] = 0
      "0000000" when "00000000010001000", -- t[136] = 0
      "0000000" when "00000000010001001", -- t[137] = 0
      "0000000" when "00000000010001010", -- t[138] = 0
      "0000000" when "00000000010001011", -- t[139] = 0
      "0000000" when "00000000010001100", -- t[140] = 0
      "0000000" when "00000000010001101", -- t[141] = 0
      "0000000" when "00000000010001110", -- t[142] = 0
      "0000000" when "00000000010001111", -- t[143] = 0
      "0000000" when "00000000010010000", -- t[144] = 0
      "0000000" when "00000000010010001", -- t[145] = 0
      "0000000" when "00000000010010010", -- t[146] = 0
      "0000000" when "00000000010010011", -- t[147] = 0
      "0000000" when "00000000010010100", -- t[148] = 0
      "0000000" when "00000000010010101", -- t[149] = 0
      "0000000" when "00000000010010110", -- t[150] = 0
      "0000000" when "00000000010010111", -- t[151] = 0
      "0000000" when "00000000010011000", -- t[152] = 0
      "0000000" when "00000000010011001", -- t[153] = 0
      "0000000" when "00000000010011010", -- t[154] = 0
      "0000000" when "00000000010011011", -- t[155] = 0
      "0000000" when "00000000010011100", -- t[156] = 0
      "0000000" when "00000000010011101", -- t[157] = 0
      "0000000" when "00000000010011110", -- t[158] = 0
      "0000000" when "00000000010011111", -- t[159] = 0
      "0000000" when "00000000010100000", -- t[160] = 0
      "0000000" when "00000000010100001", -- t[161] = 0
      "0000000" when "00000000010100010", -- t[162] = 0
      "0000000" when "00000000010100011", -- t[163] = 0
      "0000000" when "00000000010100100", -- t[164] = 0
      "0000000" when "00000000010100101", -- t[165] = 0
      "0000000" when "00000000010100110", -- t[166] = 0
      "0000000" when "00000000010100111", -- t[167] = 0
      "0000000" when "00000000010101000", -- t[168] = 0
      "0000000" when "00000000010101001", -- t[169] = 0
      "0000000" when "00000000010101010", -- t[170] = 0
      "0000000" when "00000000010101011", -- t[171] = 0
      "0000000" when "00000000010101100", -- t[172] = 0
      "0000000" when "00000000010101101", -- t[173] = 0
      "0000000" when "00000000010101110", -- t[174] = 0
      "0000000" when "00000000010101111", -- t[175] = 0
      "0000000" when "00000000010110000", -- t[176] = 0
      "0000000" when "00000000010110001", -- t[177] = 0
      "0000000" when "00000000010110010", -- t[178] = 0
      "0000000" when "00000000010110011", -- t[179] = 0
      "0000000" when "00000000010110100", -- t[180] = 0
      "0000000" when "00000000010110101", -- t[181] = 0
      "0000000" when "00000000010110110", -- t[182] = 0
      "0000000" when "00000000010110111", -- t[183] = 0
      "0000000" when "00000000010111000", -- t[184] = 0
      "0000000" when "00000000010111001", -- t[185] = 0
      "0000000" when "00000000010111010", -- t[186] = 0
      "0000000" when "00000000010111011", -- t[187] = 0
      "0000000" when "00000000010111100", -- t[188] = 0
      "0000000" when "00000000010111101", -- t[189] = 0
      "0000000" when "00000000010111110", -- t[190] = 0
      "0000000" when "00000000010111111", -- t[191] = 0
      "0000000" when "00000000011000000", -- t[192] = 0
      "0000000" when "00000000011000001", -- t[193] = 0
      "0000000" when "00000000011000010", -- t[194] = 0
      "0000000" when "00000000011000011", -- t[195] = 0
      "0000000" when "00000000011000100", -- t[196] = 0
      "0000000" when "00000000011000101", -- t[197] = 0
      "0000000" when "00000000011000110", -- t[198] = 0
      "0000000" when "00000000011000111", -- t[199] = 0
      "0000000" when "00000000011001000", -- t[200] = 0
      "0000000" when "00000000011001001", -- t[201] = 0
      "0000000" when "00000000011001010", -- t[202] = 0
      "0000000" when "00000000011001011", -- t[203] = 0
      "0000000" when "00000000011001100", -- t[204] = 0
      "0000000" when "00000000011001101", -- t[205] = 0
      "0000000" when "00000000011001110", -- t[206] = 0
      "0000000" when "00000000011001111", -- t[207] = 0
      "0000000" when "00000000011010000", -- t[208] = 0
      "0000000" when "00000000011010001", -- t[209] = 0
      "0000000" when "00000000011010010", -- t[210] = 0
      "0000000" when "00000000011010011", -- t[211] = 0
      "0000000" when "00000000011010100", -- t[212] = 0
      "0000000" when "00000000011010101", -- t[213] = 0
      "0000000" when "00000000011010110", -- t[214] = 0
      "0000000" when "00000000011010111", -- t[215] = 0
      "0000000" when "00000000011011000", -- t[216] = 0
      "0000000" when "00000000011011001", -- t[217] = 0
      "0000000" when "00000000011011010", -- t[218] = 0
      "0000000" when "00000000011011011", -- t[219] = 0
      "0000000" when "00000000011011100", -- t[220] = 0
      "0000000" when "00000000011011101", -- t[221] = 0
      "0000000" when "00000000011011110", -- t[222] = 0
      "0000000" when "00000000011011111", -- t[223] = 0
      "0000000" when "00000000011100000", -- t[224] = 0
      "0000000" when "00000000011100001", -- t[225] = 0
      "0000000" when "00000000011100010", -- t[226] = 0
      "0000000" when "00000000011100011", -- t[227] = 0
      "0000000" when "00000000011100100", -- t[228] = 0
      "0000000" when "00000000011100101", -- t[229] = 0
      "0000000" when "00000000011100110", -- t[230] = 0
      "0000000" when "00000000011100111", -- t[231] = 0
      "0000000" when "00000000011101000", -- t[232] = 0
      "0000000" when "00000000011101001", -- t[233] = 0
      "0000000" when "00000000011101010", -- t[234] = 0
      "0000000" when "00000000011101011", -- t[235] = 0
      "0000000" when "00000000011101100", -- t[236] = 0
      "0000000" when "00000000011101101", -- t[237] = 0
      "0000000" when "00000000011101110", -- t[238] = 0
      "0000000" when "00000000011101111", -- t[239] = 0
      "0000000" when "00000000011110000", -- t[240] = 0
      "0000000" when "00000000011110001", -- t[241] = 0
      "0000000" when "00000000011110010", -- t[242] = 0
      "0000000" when "00000000011110011", -- t[243] = 0
      "0000000" when "00000000011110100", -- t[244] = 0
      "0000000" when "00000000011110101", -- t[245] = 0
      "0000000" when "00000000011110110", -- t[246] = 0
      "0000000" when "00000000011110111", -- t[247] = 0
      "0000000" when "00000000011111000", -- t[248] = 0
      "0000000" when "00000000011111001", -- t[249] = 0
      "0000000" when "00000000011111010", -- t[250] = 0
      "0000000" when "00000000011111011", -- t[251] = 0
      "0000000" when "00000000011111100", -- t[252] = 0
      "0000000" when "00000000011111101", -- t[253] = 0
      "0000000" when "00000000011111110", -- t[254] = 0
      "0000000" when "00000000011111111", -- t[255] = 0
      "0000000" when "00000000100000000", -- t[256] = 0
      "0000000" when "00000000100000001", -- t[257] = 0
      "0000000" when "00000000100000010", -- t[258] = 0
      "0000000" when "00000000100000011", -- t[259] = 0
      "0000000" when "00000000100000100", -- t[260] = 0
      "0000000" when "00000000100000101", -- t[261] = 0
      "0000000" when "00000000100000110", -- t[262] = 0
      "0000000" when "00000000100000111", -- t[263] = 0
      "0000000" when "00000000100001000", -- t[264] = 0
      "0000000" when "00000000100001001", -- t[265] = 0
      "0000000" when "00000000100001010", -- t[266] = 0
      "0000000" when "00000000100001011", -- t[267] = 0
      "0000000" when "00000000100001100", -- t[268] = 0
      "0000000" when "00000000100001101", -- t[269] = 0
      "0000000" when "00000000100001110", -- t[270] = 0
      "0000000" when "00000000100001111", -- t[271] = 0
      "0000000" when "00000000100010000", -- t[272] = 0
      "0000000" when "00000000100010001", -- t[273] = 0
      "0000000" when "00000000100010010", -- t[274] = 0
      "0000000" when "00000000100010011", -- t[275] = 0
      "0000000" when "00000000100010100", -- t[276] = 0
      "0000000" when "00000000100010101", -- t[277] = 0
      "0000000" when "00000000100010110", -- t[278] = 0
      "0000000" when "00000000100010111", -- t[279] = 0
      "0000000" when "00000000100011000", -- t[280] = 0
      "0000000" when "00000000100011001", -- t[281] = 0
      "0000000" when "00000000100011010", -- t[282] = 0
      "0000000" when "00000000100011011", -- t[283] = 0
      "0000000" when "00000000100011100", -- t[284] = 0
      "0000000" when "00000000100011101", -- t[285] = 0
      "0000000" when "00000000100011110", -- t[286] = 0
      "0000000" when "00000000100011111", -- t[287] = 0
      "0000000" when "00000000100100000", -- t[288] = 0
      "0000000" when "00000000100100001", -- t[289] = 0
      "0000000" when "00000000100100010", -- t[290] = 0
      "0000000" when "00000000100100011", -- t[291] = 0
      "0000000" when "00000000100100100", -- t[292] = 0
      "0000000" when "00000000100100101", -- t[293] = 0
      "0000000" when "00000000100100110", -- t[294] = 0
      "0000000" when "00000000100100111", -- t[295] = 0
      "0000000" when "00000000100101000", -- t[296] = 0
      "0000000" when "00000000100101001", -- t[297] = 0
      "0000000" when "00000000100101010", -- t[298] = 0
      "0000000" when "00000000100101011", -- t[299] = 0
      "0000000" when "00000000100101100", -- t[300] = 0
      "0000000" when "00000000100101101", -- t[301] = 0
      "0000000" when "00000000100101110", -- t[302] = 0
      "0000000" when "00000000100101111", -- t[303] = 0
      "0000000" when "00000000100110000", -- t[304] = 0
      "0000000" when "00000000100110001", -- t[305] = 0
      "0000000" when "00000000100110010", -- t[306] = 0
      "0000000" when "00000000100110011", -- t[307] = 0
      "0000000" when "00000000100110100", -- t[308] = 0
      "0000000" when "00000000100110101", -- t[309] = 0
      "0000000" when "00000000100110110", -- t[310] = 0
      "0000000" when "00000000100110111", -- t[311] = 0
      "0000000" when "00000000100111000", -- t[312] = 0
      "0000000" when "00000000100111001", -- t[313] = 0
      "0000000" when "00000000100111010", -- t[314] = 0
      "0000000" when "00000000100111011", -- t[315] = 0
      "0000000" when "00000000100111100", -- t[316] = 0
      "0000000" when "00000000100111101", -- t[317] = 0
      "0000000" when "00000000100111110", -- t[318] = 0
      "0000000" when "00000000100111111", -- t[319] = 0
      "0000000" when "00000000101000000", -- t[320] = 0
      "0000000" when "00000000101000001", -- t[321] = 0
      "0000000" when "00000000101000010", -- t[322] = 0
      "0000000" when "00000000101000011", -- t[323] = 0
      "0000000" when "00000000101000100", -- t[324] = 0
      "0000000" when "00000000101000101", -- t[325] = 0
      "0000000" when "00000000101000110", -- t[326] = 0
      "0000000" when "00000000101000111", -- t[327] = 0
      "0000000" when "00000000101001000", -- t[328] = 0
      "0000000" when "00000000101001001", -- t[329] = 0
      "0000000" when "00000000101001010", -- t[330] = 0
      "0000000" when "00000000101001011", -- t[331] = 0
      "0000000" when "00000000101001100", -- t[332] = 0
      "0000000" when "00000000101001101", -- t[333] = 0
      "0000000" when "00000000101001110", -- t[334] = 0
      "0000000" when "00000000101001111", -- t[335] = 0
      "0000000" when "00000000101010000", -- t[336] = 0
      "0000000" when "00000000101010001", -- t[337] = 0
      "0000000" when "00000000101010010", -- t[338] = 0
      "0000000" when "00000000101010011", -- t[339] = 0
      "0000000" when "00000000101010100", -- t[340] = 0
      "0000000" when "00000000101010101", -- t[341] = 0
      "0000000" when "00000000101010110", -- t[342] = 0
      "0000000" when "00000000101010111", -- t[343] = 0
      "0000000" when "00000000101011000", -- t[344] = 0
      "0000000" when "00000000101011001", -- t[345] = 0
      "0000000" when "00000000101011010", -- t[346] = 0
      "0000000" when "00000000101011011", -- t[347] = 0
      "0000000" when "00000000101011100", -- t[348] = 0
      "0000000" when "00000000101011101", -- t[349] = 0
      "0000000" when "00000000101011110", -- t[350] = 0
      "0000000" when "00000000101011111", -- t[351] = 0
      "0000000" when "00000000101100000", -- t[352] = 0
      "0000000" when "00000000101100001", -- t[353] = 0
      "0000000" when "00000000101100010", -- t[354] = 0
      "0000000" when "00000000101100011", -- t[355] = 0
      "0000000" when "00000000101100100", -- t[356] = 0
      "0000000" when "00000000101100101", -- t[357] = 0
      "0000000" when "00000000101100110", -- t[358] = 0
      "0000000" when "00000000101100111", -- t[359] = 0
      "0000000" when "00000000101101000", -- t[360] = 0
      "0000000" when "00000000101101001", -- t[361] = 0
      "0000000" when "00000000101101010", -- t[362] = 0
      "0000000" when "00000000101101011", -- t[363] = 0
      "0000000" when "00000000101101100", -- t[364] = 0
      "0000000" when "00000000101101101", -- t[365] = 0
      "0000000" when "00000000101101110", -- t[366] = 0
      "0000000" when "00000000101101111", -- t[367] = 0
      "0000000" when "00000000101110000", -- t[368] = 0
      "0000000" when "00000000101110001", -- t[369] = 0
      "0000000" when "00000000101110010", -- t[370] = 0
      "0000000" when "00000000101110011", -- t[371] = 0
      "0000000" when "00000000101110100", -- t[372] = 0
      "0000000" when "00000000101110101", -- t[373] = 0
      "0000000" when "00000000101110110", -- t[374] = 0
      "0000000" when "00000000101110111", -- t[375] = 0
      "0000000" when "00000000101111000", -- t[376] = 0
      "0000000" when "00000000101111001", -- t[377] = 0
      "0000000" when "00000000101111010", -- t[378] = 0
      "0000000" when "00000000101111011", -- t[379] = 0
      "0000000" when "00000000101111100", -- t[380] = 0
      "0000000" when "00000000101111101", -- t[381] = 0
      "0000000" when "00000000101111110", -- t[382] = 0
      "0000000" when "00000000101111111", -- t[383] = 0
      "0000000" when "00000000110000000", -- t[384] = 0
      "0000000" when "00000000110000001", -- t[385] = 0
      "0000000" when "00000000110000010", -- t[386] = 0
      "0000000" when "00000000110000011", -- t[387] = 0
      "0000000" when "00000000110000100", -- t[388] = 0
      "0000000" when "00000000110000101", -- t[389] = 0
      "0000000" when "00000000110000110", -- t[390] = 0
      "0000000" when "00000000110000111", -- t[391] = 0
      "0000000" when "00000000110001000", -- t[392] = 0
      "0000000" when "00000000110001001", -- t[393] = 0
      "0000000" when "00000000110001010", -- t[394] = 0
      "0000000" when "00000000110001011", -- t[395] = 0
      "0000000" when "00000000110001100", -- t[396] = 0
      "0000000" when "00000000110001101", -- t[397] = 0
      "0000000" when "00000000110001110", -- t[398] = 0
      "0000000" when "00000000110001111", -- t[399] = 0
      "0000000" when "00000000110010000", -- t[400] = 0
      "0000000" when "00000000110010001", -- t[401] = 0
      "0000000" when "00000000110010010", -- t[402] = 0
      "0000000" when "00000000110010011", -- t[403] = 0
      "0000000" when "00000000110010100", -- t[404] = 0
      "0000000" when "00000000110010101", -- t[405] = 0
      "0000000" when "00000000110010110", -- t[406] = 0
      "0000000" when "00000000110010111", -- t[407] = 0
      "0000000" when "00000000110011000", -- t[408] = 0
      "0000000" when "00000000110011001", -- t[409] = 0
      "0000000" when "00000000110011010", -- t[410] = 0
      "0000000" when "00000000110011011", -- t[411] = 0
      "0000000" when "00000000110011100", -- t[412] = 0
      "0000000" when "00000000110011101", -- t[413] = 0
      "0000000" when "00000000110011110", -- t[414] = 0
      "0000000" when "00000000110011111", -- t[415] = 0
      "0000000" when "00000000110100000", -- t[416] = 0
      "0000000" when "00000000110100001", -- t[417] = 0
      "0000000" when "00000000110100010", -- t[418] = 0
      "0000000" when "00000000110100011", -- t[419] = 0
      "0000000" when "00000000110100100", -- t[420] = 0
      "0000000" when "00000000110100101", -- t[421] = 0
      "0000000" when "00000000110100110", -- t[422] = 0
      "0000000" when "00000000110100111", -- t[423] = 0
      "0000000" when "00000000110101000", -- t[424] = 0
      "0000000" when "00000000110101001", -- t[425] = 0
      "0000000" when "00000000110101010", -- t[426] = 0
      "0000000" when "00000000110101011", -- t[427] = 0
      "0000000" when "00000000110101100", -- t[428] = 0
      "0000000" when "00000000110101101", -- t[429] = 0
      "0000000" when "00000000110101110", -- t[430] = 0
      "0000000" when "00000000110101111", -- t[431] = 0
      "0000000" when "00000000110110000", -- t[432] = 0
      "0000000" when "00000000110110001", -- t[433] = 0
      "0000000" when "00000000110110010", -- t[434] = 0
      "0000000" when "00000000110110011", -- t[435] = 0
      "0000000" when "00000000110110100", -- t[436] = 0
      "0000000" when "00000000110110101", -- t[437] = 0
      "0000000" when "00000000110110110", -- t[438] = 0
      "0000000" when "00000000110110111", -- t[439] = 0
      "0000000" when "00000000110111000", -- t[440] = 0
      "0000000" when "00000000110111001", -- t[441] = 0
      "0000000" when "00000000110111010", -- t[442] = 0
      "0000000" when "00000000110111011", -- t[443] = 0
      "0000000" when "00000000110111100", -- t[444] = 0
      "0000000" when "00000000110111101", -- t[445] = 0
      "0000000" when "00000000110111110", -- t[446] = 0
      "0000000" when "00000000110111111", -- t[447] = 0
      "0000000" when "00000000111000000", -- t[448] = 0
      "0000000" when "00000000111000001", -- t[449] = 0
      "0000000" when "00000000111000010", -- t[450] = 0
      "0000000" when "00000000111000011", -- t[451] = 0
      "0000000" when "00000000111000100", -- t[452] = 0
      "0000000" when "00000000111000101", -- t[453] = 0
      "0000000" when "00000000111000110", -- t[454] = 0
      "0000000" when "00000000111000111", -- t[455] = 0
      "0000000" when "00000000111001000", -- t[456] = 0
      "0000000" when "00000000111001001", -- t[457] = 0
      "0000000" when "00000000111001010", -- t[458] = 0
      "0000000" when "00000000111001011", -- t[459] = 0
      "0000000" when "00000000111001100", -- t[460] = 0
      "0000000" when "00000000111001101", -- t[461] = 0
      "0000000" when "00000000111001110", -- t[462] = 0
      "0000000" when "00000000111001111", -- t[463] = 0
      "0000000" when "00000000111010000", -- t[464] = 0
      "0000000" when "00000000111010001", -- t[465] = 0
      "0000000" when "00000000111010010", -- t[466] = 0
      "0000000" when "00000000111010011", -- t[467] = 0
      "0000000" when "00000000111010100", -- t[468] = 0
      "0000000" when "00000000111010101", -- t[469] = 0
      "0000000" when "00000000111010110", -- t[470] = 0
      "0000000" when "00000000111010111", -- t[471] = 0
      "0000000" when "00000000111011000", -- t[472] = 0
      "0000000" when "00000000111011001", -- t[473] = 0
      "0000000" when "00000000111011010", -- t[474] = 0
      "0000000" when "00000000111011011", -- t[475] = 0
      "0000000" when "00000000111011100", -- t[476] = 0
      "0000000" when "00000000111011101", -- t[477] = 0
      "0000000" when "00000000111011110", -- t[478] = 0
      "0000000" when "00000000111011111", -- t[479] = 0
      "0000000" when "00000000111100000", -- t[480] = 0
      "0000000" when "00000000111100001", -- t[481] = 0
      "0000000" when "00000000111100010", -- t[482] = 0
      "0000000" when "00000000111100011", -- t[483] = 0
      "0000000" when "00000000111100100", -- t[484] = 0
      "0000000" when "00000000111100101", -- t[485] = 0
      "0000000" when "00000000111100110", -- t[486] = 0
      "0000000" when "00000000111100111", -- t[487] = 0
      "0000000" when "00000000111101000", -- t[488] = 0
      "0000000" when "00000000111101001", -- t[489] = 0
      "0000000" when "00000000111101010", -- t[490] = 0
      "0000000" when "00000000111101011", -- t[491] = 0
      "0000000" when "00000000111101100", -- t[492] = 0
      "0000000" when "00000000111101101", -- t[493] = 0
      "0000000" when "00000000111101110", -- t[494] = 0
      "0000000" when "00000000111101111", -- t[495] = 0
      "0000000" when "00000000111110000", -- t[496] = 0
      "0000000" when "00000000111110001", -- t[497] = 0
      "0000000" when "00000000111110010", -- t[498] = 0
      "0000000" when "00000000111110011", -- t[499] = 0
      "0000000" when "00000000111110100", -- t[500] = 0
      "0000000" when "00000000111110101", -- t[501] = 0
      "0000000" when "00000000111110110", -- t[502] = 0
      "0000000" when "00000000111110111", -- t[503] = 0
      "0000000" when "00000000111111000", -- t[504] = 0
      "0000000" when "00000000111111001", -- t[505] = 0
      "0000000" when "00000000111111010", -- t[506] = 0
      "0000000" when "00000000111111011", -- t[507] = 0
      "0000000" when "00000000111111100", -- t[508] = 0
      "0000000" when "00000000111111101", -- t[509] = 0
      "0000000" when "00000000111111110", -- t[510] = 0
      "0000000" when "00000000111111111", -- t[511] = 0
      "0000000" when "00000001000000000", -- t[512] = 0
      "0000000" when "00000001000000001", -- t[513] = 0
      "0000000" when "00000001000000010", -- t[514] = 0
      "0000000" when "00000001000000011", -- t[515] = 0
      "0000000" when "00000001000000100", -- t[516] = 0
      "0000000" when "00000001000000101", -- t[517] = 0
      "0000000" when "00000001000000110", -- t[518] = 0
      "0000000" when "00000001000000111", -- t[519] = 0
      "0000000" when "00000001000001000", -- t[520] = 0
      "0000000" when "00000001000001001", -- t[521] = 0
      "0000000" when "00000001000001010", -- t[522] = 0
      "0000000" when "00000001000001011", -- t[523] = 0
      "0000000" when "00000001000001100", -- t[524] = 0
      "0000000" when "00000001000001101", -- t[525] = 0
      "0000000" when "00000001000001110", -- t[526] = 0
      "0000000" when "00000001000001111", -- t[527] = 0
      "0000000" when "00000001000010000", -- t[528] = 0
      "0000000" when "00000001000010001", -- t[529] = 0
      "0000000" when "00000001000010010", -- t[530] = 0
      "0000000" when "00000001000010011", -- t[531] = 0
      "0000000" when "00000001000010100", -- t[532] = 0
      "0000000" when "00000001000010101", -- t[533] = 0
      "0000000" when "00000001000010110", -- t[534] = 0
      "0000000" when "00000001000010111", -- t[535] = 0
      "0000000" when "00000001000011000", -- t[536] = 0
      "0000000" when "00000001000011001", -- t[537] = 0
      "0000000" when "00000001000011010", -- t[538] = 0
      "0000000" when "00000001000011011", -- t[539] = 0
      "0000000" when "00000001000011100", -- t[540] = 0
      "0000000" when "00000001000011101", -- t[541] = 0
      "0000000" when "00000001000011110", -- t[542] = 0
      "0000000" when "00000001000011111", -- t[543] = 0
      "0000000" when "00000001000100000", -- t[544] = 0
      "0000000" when "00000001000100001", -- t[545] = 0
      "0000000" when "00000001000100010", -- t[546] = 0
      "0000000" when "00000001000100011", -- t[547] = 0
      "0000000" when "00000001000100100", -- t[548] = 0
      "0000000" when "00000001000100101", -- t[549] = 0
      "0000000" when "00000001000100110", -- t[550] = 0
      "0000000" when "00000001000100111", -- t[551] = 0
      "0000000" when "00000001000101000", -- t[552] = 0
      "0000000" when "00000001000101001", -- t[553] = 0
      "0000000" when "00000001000101010", -- t[554] = 0
      "0000000" when "00000001000101011", -- t[555] = 0
      "0000000" when "00000001000101100", -- t[556] = 0
      "0000000" when "00000001000101101", -- t[557] = 0
      "0000000" when "00000001000101110", -- t[558] = 0
      "0000000" when "00000001000101111", -- t[559] = 0
      "0000000" when "00000001000110000", -- t[560] = 0
      "0000000" when "00000001000110001", -- t[561] = 0
      "0000000" when "00000001000110010", -- t[562] = 0
      "0000000" when "00000001000110011", -- t[563] = 0
      "0000000" when "00000001000110100", -- t[564] = 0
      "0000000" when "00000001000110101", -- t[565] = 0
      "0000000" when "00000001000110110", -- t[566] = 0
      "0000000" when "00000001000110111", -- t[567] = 0
      "0000000" when "00000001000111000", -- t[568] = 0
      "0000000" when "00000001000111001", -- t[569] = 0
      "0000000" when "00000001000111010", -- t[570] = 0
      "0000000" when "00000001000111011", -- t[571] = 0
      "0000000" when "00000001000111100", -- t[572] = 0
      "0000000" when "00000001000111101", -- t[573] = 0
      "0000000" when "00000001000111110", -- t[574] = 0
      "0000000" when "00000001000111111", -- t[575] = 0
      "0000000" when "00000001001000000", -- t[576] = 0
      "0000000" when "00000001001000001", -- t[577] = 0
      "0000000" when "00000001001000010", -- t[578] = 0
      "0000000" when "00000001001000011", -- t[579] = 0
      "0000000" when "00000001001000100", -- t[580] = 0
      "0000000" when "00000001001000101", -- t[581] = 0
      "0000000" when "00000001001000110", -- t[582] = 0
      "0000000" when "00000001001000111", -- t[583] = 0
      "0000000" when "00000001001001000", -- t[584] = 0
      "0000000" when "00000001001001001", -- t[585] = 0
      "0000000" when "00000001001001010", -- t[586] = 0
      "0000000" when "00000001001001011", -- t[587] = 0
      "0000000" when "00000001001001100", -- t[588] = 0
      "0000000" when "00000001001001101", -- t[589] = 0
      "0000000" when "00000001001001110", -- t[590] = 0
      "0000000" when "00000001001001111", -- t[591] = 0
      "0000000" when "00000001001010000", -- t[592] = 0
      "0000000" when "00000001001010001", -- t[593] = 0
      "0000000" when "00000001001010010", -- t[594] = 0
      "0000000" when "00000001001010011", -- t[595] = 0
      "0000000" when "00000001001010100", -- t[596] = 0
      "0000000" when "00000001001010101", -- t[597] = 0
      "0000000" when "00000001001010110", -- t[598] = 0
      "0000000" when "00000001001010111", -- t[599] = 0
      "0000000" when "00000001001011000", -- t[600] = 0
      "0000000" when "00000001001011001", -- t[601] = 0
      "0000000" when "00000001001011010", -- t[602] = 0
      "0000000" when "00000001001011011", -- t[603] = 0
      "0000000" when "00000001001011100", -- t[604] = 0
      "0000000" when "00000001001011101", -- t[605] = 0
      "0000000" when "00000001001011110", -- t[606] = 0
      "0000000" when "00000001001011111", -- t[607] = 0
      "0000000" when "00000001001100000", -- t[608] = 0
      "0000000" when "00000001001100001", -- t[609] = 0
      "0000000" when "00000001001100010", -- t[610] = 0
      "0000000" when "00000001001100011", -- t[611] = 0
      "0000000" when "00000001001100100", -- t[612] = 0
      "0000000" when "00000001001100101", -- t[613] = 0
      "0000000" when "00000001001100110", -- t[614] = 0
      "0000000" when "00000001001100111", -- t[615] = 0
      "0000000" when "00000001001101000", -- t[616] = 0
      "0000000" when "00000001001101001", -- t[617] = 0
      "0000000" when "00000001001101010", -- t[618] = 0
      "0000000" when "00000001001101011", -- t[619] = 0
      "0000000" when "00000001001101100", -- t[620] = 0
      "0000000" when "00000001001101101", -- t[621] = 0
      "0000000" when "00000001001101110", -- t[622] = 0
      "0000000" when "00000001001101111", -- t[623] = 0
      "0000000" when "00000001001110000", -- t[624] = 0
      "0000000" when "00000001001110001", -- t[625] = 0
      "0000000" when "00000001001110010", -- t[626] = 0
      "0000000" when "00000001001110011", -- t[627] = 0
      "0000000" when "00000001001110100", -- t[628] = 0
      "0000000" when "00000001001110101", -- t[629] = 0
      "0000000" when "00000001001110110", -- t[630] = 0
      "0000000" when "00000001001110111", -- t[631] = 0
      "0000000" when "00000001001111000", -- t[632] = 0
      "0000000" when "00000001001111001", -- t[633] = 0
      "0000000" when "00000001001111010", -- t[634] = 0
      "0000000" when "00000001001111011", -- t[635] = 0
      "0000000" when "00000001001111100", -- t[636] = 0
      "0000000" when "00000001001111101", -- t[637] = 0
      "0000000" when "00000001001111110", -- t[638] = 0
      "0000000" when "00000001001111111", -- t[639] = 0
      "0000000" when "00000001010000000", -- t[640] = 0
      "0000000" when "00000001010000001", -- t[641] = 0
      "0000000" when "00000001010000010", -- t[642] = 0
      "0000000" when "00000001010000011", -- t[643] = 0
      "0000000" when "00000001010000100", -- t[644] = 0
      "0000000" when "00000001010000101", -- t[645] = 0
      "0000000" when "00000001010000110", -- t[646] = 0
      "0000000" when "00000001010000111", -- t[647] = 0
      "0000000" when "00000001010001000", -- t[648] = 0
      "0000000" when "00000001010001001", -- t[649] = 0
      "0000000" when "00000001010001010", -- t[650] = 0
      "0000000" when "00000001010001011", -- t[651] = 0
      "0000000" when "00000001010001100", -- t[652] = 0
      "0000000" when "00000001010001101", -- t[653] = 0
      "0000000" when "00000001010001110", -- t[654] = 0
      "0000000" when "00000001010001111", -- t[655] = 0
      "0000000" when "00000001010010000", -- t[656] = 0
      "0000000" when "00000001010010001", -- t[657] = 0
      "0000000" when "00000001010010010", -- t[658] = 0
      "0000000" when "00000001010010011", -- t[659] = 0
      "0000000" when "00000001010010100", -- t[660] = 0
      "0000000" when "00000001010010101", -- t[661] = 0
      "0000000" when "00000001010010110", -- t[662] = 0
      "0000000" when "00000001010010111", -- t[663] = 0
      "0000000" when "00000001010011000", -- t[664] = 0
      "0000000" when "00000001010011001", -- t[665] = 0
      "0000000" when "00000001010011010", -- t[666] = 0
      "0000000" when "00000001010011011", -- t[667] = 0
      "0000000" when "00000001010011100", -- t[668] = 0
      "0000000" when "00000001010011101", -- t[669] = 0
      "0000000" when "00000001010011110", -- t[670] = 0
      "0000000" when "00000001010011111", -- t[671] = 0
      "0000000" when "00000001010100000", -- t[672] = 0
      "0000000" when "00000001010100001", -- t[673] = 0
      "0000000" when "00000001010100010", -- t[674] = 0
      "0000000" when "00000001010100011", -- t[675] = 0
      "0000000" when "00000001010100100", -- t[676] = 0
      "0000000" when "00000001010100101", -- t[677] = 0
      "0000000" when "00000001010100110", -- t[678] = 0
      "0000000" when "00000001010100111", -- t[679] = 0
      "0000000" when "00000001010101000", -- t[680] = 0
      "0000000" when "00000001010101001", -- t[681] = 0
      "0000000" when "00000001010101010", -- t[682] = 0
      "0000000" when "00000001010101011", -- t[683] = 0
      "0000000" when "00000001010101100", -- t[684] = 0
      "0000000" when "00000001010101101", -- t[685] = 0
      "0000000" when "00000001010101110", -- t[686] = 0
      "0000000" when "00000001010101111", -- t[687] = 0
      "0000000" when "00000001010110000", -- t[688] = 0
      "0000000" when "00000001010110001", -- t[689] = 0
      "0000000" when "00000001010110010", -- t[690] = 0
      "0000000" when "00000001010110011", -- t[691] = 0
      "0000000" when "00000001010110100", -- t[692] = 0
      "0000000" when "00000001010110101", -- t[693] = 0
      "0000000" when "00000001010110110", -- t[694] = 0
      "0000000" when "00000001010110111", -- t[695] = 0
      "0000000" when "00000001010111000", -- t[696] = 0
      "0000000" when "00000001010111001", -- t[697] = 0
      "0000000" when "00000001010111010", -- t[698] = 0
      "0000000" when "00000001010111011", -- t[699] = 0
      "0000000" when "00000001010111100", -- t[700] = 0
      "0000000" when "00000001010111101", -- t[701] = 0
      "0000000" when "00000001010111110", -- t[702] = 0
      "0000000" when "00000001010111111", -- t[703] = 0
      "0000000" when "00000001011000000", -- t[704] = 0
      "0000000" when "00000001011000001", -- t[705] = 0
      "0000000" when "00000001011000010", -- t[706] = 0
      "0000000" when "00000001011000011", -- t[707] = 0
      "0000000" when "00000001011000100", -- t[708] = 0
      "0000000" when "00000001011000101", -- t[709] = 0
      "0000000" when "00000001011000110", -- t[710] = 0
      "0000000" when "00000001011000111", -- t[711] = 0
      "0000000" when "00000001011001000", -- t[712] = 0
      "0000000" when "00000001011001001", -- t[713] = 0
      "0000000" when "00000001011001010", -- t[714] = 0
      "0000000" when "00000001011001011", -- t[715] = 0
      "0000000" when "00000001011001100", -- t[716] = 0
      "0000000" when "00000001011001101", -- t[717] = 0
      "0000000" when "00000001011001110", -- t[718] = 0
      "0000000" when "00000001011001111", -- t[719] = 0
      "0000000" when "00000001011010000", -- t[720] = 0
      "0000000" when "00000001011010001", -- t[721] = 0
      "0000000" when "00000001011010010", -- t[722] = 0
      "0000000" when "00000001011010011", -- t[723] = 0
      "0000000" when "00000001011010100", -- t[724] = 0
      "0000000" when "00000001011010101", -- t[725] = 0
      "0000000" when "00000001011010110", -- t[726] = 0
      "0000000" when "00000001011010111", -- t[727] = 0
      "0000000" when "00000001011011000", -- t[728] = 0
      "0000000" when "00000001011011001", -- t[729] = 0
      "0000000" when "00000001011011010", -- t[730] = 0
      "0000000" when "00000001011011011", -- t[731] = 0
      "0000000" when "00000001011011100", -- t[732] = 0
      "0000000" when "00000001011011101", -- t[733] = 0
      "0000000" when "00000001011011110", -- t[734] = 0
      "0000000" when "00000001011011111", -- t[735] = 0
      "0000000" when "00000001011100000", -- t[736] = 0
      "0000000" when "00000001011100001", -- t[737] = 0
      "0000000" when "00000001011100010", -- t[738] = 0
      "0000000" when "00000001011100011", -- t[739] = 0
      "0000000" when "00000001011100100", -- t[740] = 0
      "0000000" when "00000001011100101", -- t[741] = 0
      "0000000" when "00000001011100110", -- t[742] = 0
      "0000000" when "00000001011100111", -- t[743] = 0
      "0000000" when "00000001011101000", -- t[744] = 0
      "0000000" when "00000001011101001", -- t[745] = 0
      "0000000" when "00000001011101010", -- t[746] = 0
      "0000000" when "00000001011101011", -- t[747] = 0
      "0000000" when "00000001011101100", -- t[748] = 0
      "0000000" when "00000001011101101", -- t[749] = 0
      "0000000" when "00000001011101110", -- t[750] = 0
      "0000000" when "00000001011101111", -- t[751] = 0
      "0000000" when "00000001011110000", -- t[752] = 0
      "0000000" when "00000001011110001", -- t[753] = 0
      "0000000" when "00000001011110010", -- t[754] = 0
      "0000000" when "00000001011110011", -- t[755] = 0
      "0000000" when "00000001011110100", -- t[756] = 0
      "0000000" when "00000001011110101", -- t[757] = 0
      "0000000" when "00000001011110110", -- t[758] = 0
      "0000000" when "00000001011110111", -- t[759] = 0
      "0000000" when "00000001011111000", -- t[760] = 0
      "0000000" when "00000001011111001", -- t[761] = 0
      "0000000" when "00000001011111010", -- t[762] = 0
      "0000000" when "00000001011111011", -- t[763] = 0
      "0000000" when "00000001011111100", -- t[764] = 0
      "0000000" when "00000001011111101", -- t[765] = 0
      "0000000" when "00000001011111110", -- t[766] = 0
      "0000000" when "00000001011111111", -- t[767] = 0
      "0000000" when "00000001100000000", -- t[768] = 0
      "0000000" when "00000001100000001", -- t[769] = 0
      "0000000" when "00000001100000010", -- t[770] = 0
      "0000000" when "00000001100000011", -- t[771] = 0
      "0000000" when "00000001100000100", -- t[772] = 0
      "0000000" when "00000001100000101", -- t[773] = 0
      "0000000" when "00000001100000110", -- t[774] = 0
      "0000000" when "00000001100000111", -- t[775] = 0
      "0000000" when "00000001100001000", -- t[776] = 0
      "0000000" when "00000001100001001", -- t[777] = 0
      "0000000" when "00000001100001010", -- t[778] = 0
      "0000000" when "00000001100001011", -- t[779] = 0
      "0000000" when "00000001100001100", -- t[780] = 0
      "0000000" when "00000001100001101", -- t[781] = 0
      "0000000" when "00000001100001110", -- t[782] = 0
      "0000000" when "00000001100001111", -- t[783] = 0
      "0000000" when "00000001100010000", -- t[784] = 0
      "0000000" when "00000001100010001", -- t[785] = 0
      "0000000" when "00000001100010010", -- t[786] = 0
      "0000000" when "00000001100010011", -- t[787] = 0
      "0000000" when "00000001100010100", -- t[788] = 0
      "0000000" when "00000001100010101", -- t[789] = 0
      "0000000" when "00000001100010110", -- t[790] = 0
      "0000000" when "00000001100010111", -- t[791] = 0
      "0000000" when "00000001100011000", -- t[792] = 0
      "0000000" when "00000001100011001", -- t[793] = 0
      "0000000" when "00000001100011010", -- t[794] = 0
      "0000000" when "00000001100011011", -- t[795] = 0
      "0000000" when "00000001100011100", -- t[796] = 0
      "0000000" when "00000001100011101", -- t[797] = 0
      "0000000" when "00000001100011110", -- t[798] = 0
      "0000000" when "00000001100011111", -- t[799] = 0
      "0000000" when "00000001100100000", -- t[800] = 0
      "0000000" when "00000001100100001", -- t[801] = 0
      "0000000" when "00000001100100010", -- t[802] = 0
      "0000000" when "00000001100100011", -- t[803] = 0
      "0000000" when "00000001100100100", -- t[804] = 0
      "0000000" when "00000001100100101", -- t[805] = 0
      "0000000" when "00000001100100110", -- t[806] = 0
      "0000000" when "00000001100100111", -- t[807] = 0
      "0000000" when "00000001100101000", -- t[808] = 0
      "0000000" when "00000001100101001", -- t[809] = 0
      "0000000" when "00000001100101010", -- t[810] = 0
      "0000000" when "00000001100101011", -- t[811] = 0
      "0000000" when "00000001100101100", -- t[812] = 0
      "0000000" when "00000001100101101", -- t[813] = 0
      "0000000" when "00000001100101110", -- t[814] = 0
      "0000000" when "00000001100101111", -- t[815] = 0
      "0000000" when "00000001100110000", -- t[816] = 0
      "0000000" when "00000001100110001", -- t[817] = 0
      "0000000" when "00000001100110010", -- t[818] = 0
      "0000000" when "00000001100110011", -- t[819] = 0
      "0000000" when "00000001100110100", -- t[820] = 0
      "0000000" when "00000001100110101", -- t[821] = 0
      "0000000" when "00000001100110110", -- t[822] = 0
      "0000000" when "00000001100110111", -- t[823] = 0
      "0000000" when "00000001100111000", -- t[824] = 0
      "0000000" when "00000001100111001", -- t[825] = 0
      "0000000" when "00000001100111010", -- t[826] = 0
      "0000000" when "00000001100111011", -- t[827] = 0
      "0000000" when "00000001100111100", -- t[828] = 0
      "0000000" when "00000001100111101", -- t[829] = 0
      "0000000" when "00000001100111110", -- t[830] = 0
      "0000000" when "00000001100111111", -- t[831] = 0
      "0000000" when "00000001101000000", -- t[832] = 0
      "0000000" when "00000001101000001", -- t[833] = 0
      "0000000" when "00000001101000010", -- t[834] = 0
      "0000000" when "00000001101000011", -- t[835] = 0
      "0000000" when "00000001101000100", -- t[836] = 0
      "0000000" when "00000001101000101", -- t[837] = 0
      "0000000" when "00000001101000110", -- t[838] = 0
      "0000000" when "00000001101000111", -- t[839] = 0
      "0000000" when "00000001101001000", -- t[840] = 0
      "0000000" when "00000001101001001", -- t[841] = 0
      "0000000" when "00000001101001010", -- t[842] = 0
      "0000000" when "00000001101001011", -- t[843] = 0
      "0000000" when "00000001101001100", -- t[844] = 0
      "0000000" when "00000001101001101", -- t[845] = 0
      "0000000" when "00000001101001110", -- t[846] = 0
      "0000000" when "00000001101001111", -- t[847] = 0
      "0000000" when "00000001101010000", -- t[848] = 0
      "0000000" when "00000001101010001", -- t[849] = 0
      "0000000" when "00000001101010010", -- t[850] = 0
      "0000000" when "00000001101010011", -- t[851] = 0
      "0000000" when "00000001101010100", -- t[852] = 0
      "0000000" when "00000001101010101", -- t[853] = 0
      "0000000" when "00000001101010110", -- t[854] = 0
      "0000000" when "00000001101010111", -- t[855] = 0
      "0000000" when "00000001101011000", -- t[856] = 0
      "0000000" when "00000001101011001", -- t[857] = 0
      "0000000" when "00000001101011010", -- t[858] = 0
      "0000000" when "00000001101011011", -- t[859] = 0
      "0000000" when "00000001101011100", -- t[860] = 0
      "0000000" when "00000001101011101", -- t[861] = 0
      "0000000" when "00000001101011110", -- t[862] = 0
      "0000000" when "00000001101011111", -- t[863] = 0
      "0000000" when "00000001101100000", -- t[864] = 0
      "0000000" when "00000001101100001", -- t[865] = 0
      "0000000" when "00000001101100010", -- t[866] = 0
      "0000000" when "00000001101100011", -- t[867] = 0
      "0000000" when "00000001101100100", -- t[868] = 0
      "0000000" when "00000001101100101", -- t[869] = 0
      "0000000" when "00000001101100110", -- t[870] = 0
      "0000000" when "00000001101100111", -- t[871] = 0
      "0000000" when "00000001101101000", -- t[872] = 0
      "0000000" when "00000001101101001", -- t[873] = 0
      "0000000" when "00000001101101010", -- t[874] = 0
      "0000000" when "00000001101101011", -- t[875] = 0
      "0000000" when "00000001101101100", -- t[876] = 0
      "0000000" when "00000001101101101", -- t[877] = 0
      "0000000" when "00000001101101110", -- t[878] = 0
      "0000000" when "00000001101101111", -- t[879] = 0
      "0000000" when "00000001101110000", -- t[880] = 0
      "0000000" when "00000001101110001", -- t[881] = 0
      "0000000" when "00000001101110010", -- t[882] = 0
      "0000000" when "00000001101110011", -- t[883] = 0
      "0000000" when "00000001101110100", -- t[884] = 0
      "0000000" when "00000001101110101", -- t[885] = 0
      "0000000" when "00000001101110110", -- t[886] = 0
      "0000000" when "00000001101110111", -- t[887] = 0
      "0000000" when "00000001101111000", -- t[888] = 0
      "0000000" when "00000001101111001", -- t[889] = 0
      "0000000" when "00000001101111010", -- t[890] = 0
      "0000000" when "00000001101111011", -- t[891] = 0
      "0000000" when "00000001101111100", -- t[892] = 0
      "0000000" when "00000001101111101", -- t[893] = 0
      "0000000" when "00000001101111110", -- t[894] = 0
      "0000000" when "00000001101111111", -- t[895] = 0
      "0000000" when "00000001110000000", -- t[896] = 0
      "0000000" when "00000001110000001", -- t[897] = 0
      "0000000" when "00000001110000010", -- t[898] = 0
      "0000000" when "00000001110000011", -- t[899] = 0
      "0000000" when "00000001110000100", -- t[900] = 0
      "0000000" when "00000001110000101", -- t[901] = 0
      "0000000" when "00000001110000110", -- t[902] = 0
      "0000000" when "00000001110000111", -- t[903] = 0
      "0000000" when "00000001110001000", -- t[904] = 0
      "0000000" when "00000001110001001", -- t[905] = 0
      "0000000" when "00000001110001010", -- t[906] = 0
      "0000000" when "00000001110001011", -- t[907] = 0
      "0000000" when "00000001110001100", -- t[908] = 0
      "0000000" when "00000001110001101", -- t[909] = 0
      "0000000" when "00000001110001110", -- t[910] = 0
      "0000000" when "00000001110001111", -- t[911] = 0
      "0000000" when "00000001110010000", -- t[912] = 0
      "0000000" when "00000001110010001", -- t[913] = 0
      "0000000" when "00000001110010010", -- t[914] = 0
      "0000000" when "00000001110010011", -- t[915] = 0
      "0000000" when "00000001110010100", -- t[916] = 0
      "0000000" when "00000001110010101", -- t[917] = 0
      "0000000" when "00000001110010110", -- t[918] = 0
      "0000000" when "00000001110010111", -- t[919] = 0
      "0000000" when "00000001110011000", -- t[920] = 0
      "0000000" when "00000001110011001", -- t[921] = 0
      "0000000" when "00000001110011010", -- t[922] = 0
      "0000000" when "00000001110011011", -- t[923] = 0
      "0000000" when "00000001110011100", -- t[924] = 0
      "0000000" when "00000001110011101", -- t[925] = 0
      "0000000" when "00000001110011110", -- t[926] = 0
      "0000000" when "00000001110011111", -- t[927] = 0
      "0000000" when "00000001110100000", -- t[928] = 0
      "0000000" when "00000001110100001", -- t[929] = 0
      "0000000" when "00000001110100010", -- t[930] = 0
      "0000000" when "00000001110100011", -- t[931] = 0
      "0000000" when "00000001110100100", -- t[932] = 0
      "0000000" when "00000001110100101", -- t[933] = 0
      "0000000" when "00000001110100110", -- t[934] = 0
      "0000000" when "00000001110100111", -- t[935] = 0
      "0000000" when "00000001110101000", -- t[936] = 0
      "0000000" when "00000001110101001", -- t[937] = 0
      "0000000" when "00000001110101010", -- t[938] = 0
      "0000000" when "00000001110101011", -- t[939] = 0
      "0000000" when "00000001110101100", -- t[940] = 0
      "0000000" when "00000001110101101", -- t[941] = 0
      "0000000" when "00000001110101110", -- t[942] = 0
      "0000000" when "00000001110101111", -- t[943] = 0
      "0000000" when "00000001110110000", -- t[944] = 0
      "0000000" when "00000001110110001", -- t[945] = 0
      "0000000" when "00000001110110010", -- t[946] = 0
      "0000000" when "00000001110110011", -- t[947] = 0
      "0000000" when "00000001110110100", -- t[948] = 0
      "0000000" when "00000001110110101", -- t[949] = 0
      "0000000" when "00000001110110110", -- t[950] = 0
      "0000000" when "00000001110110111", -- t[951] = 0
      "0000000" when "00000001110111000", -- t[952] = 0
      "0000000" when "00000001110111001", -- t[953] = 0
      "0000000" when "00000001110111010", -- t[954] = 0
      "0000000" when "00000001110111011", -- t[955] = 0
      "0000000" when "00000001110111100", -- t[956] = 0
      "0000000" when "00000001110111101", -- t[957] = 0
      "0000000" when "00000001110111110", -- t[958] = 0
      "0000000" when "00000001110111111", -- t[959] = 0
      "0000000" when "00000001111000000", -- t[960] = 0
      "0000000" when "00000001111000001", -- t[961] = 0
      "0000000" when "00000001111000010", -- t[962] = 0
      "0000000" when "00000001111000011", -- t[963] = 0
      "0000000" when "00000001111000100", -- t[964] = 0
      "0000000" when "00000001111000101", -- t[965] = 0
      "0000000" when "00000001111000110", -- t[966] = 0
      "0000000" when "00000001111000111", -- t[967] = 0
      "0000000" when "00000001111001000", -- t[968] = 0
      "0000000" when "00000001111001001", -- t[969] = 0
      "0000000" when "00000001111001010", -- t[970] = 0
      "0000000" when "00000001111001011", -- t[971] = 0
      "0000000" when "00000001111001100", -- t[972] = 0
      "0000000" when "00000001111001101", -- t[973] = 0
      "0000000" when "00000001111001110", -- t[974] = 0
      "0000000" when "00000001111001111", -- t[975] = 0
      "0000000" when "00000001111010000", -- t[976] = 0
      "0000000" when "00000001111010001", -- t[977] = 0
      "0000000" when "00000001111010010", -- t[978] = 0
      "0000000" when "00000001111010011", -- t[979] = 0
      "0000000" when "00000001111010100", -- t[980] = 0
      "0000000" when "00000001111010101", -- t[981] = 0
      "0000000" when "00000001111010110", -- t[982] = 0
      "0000000" when "00000001111010111", -- t[983] = 0
      "0000000" when "00000001111011000", -- t[984] = 0
      "0000000" when "00000001111011001", -- t[985] = 0
      "0000000" when "00000001111011010", -- t[986] = 0
      "0000000" when "00000001111011011", -- t[987] = 0
      "0000000" when "00000001111011100", -- t[988] = 0
      "0000000" when "00000001111011101", -- t[989] = 0
      "0000000" when "00000001111011110", -- t[990] = 0
      "0000000" when "00000001111011111", -- t[991] = 0
      "0000000" when "00000001111100000", -- t[992] = 0
      "0000000" when "00000001111100001", -- t[993] = 0
      "0000000" when "00000001111100010", -- t[994] = 0
      "0000000" when "00000001111100011", -- t[995] = 0
      "0000000" when "00000001111100100", -- t[996] = 0
      "0000000" when "00000001111100101", -- t[997] = 0
      "0000000" when "00000001111100110", -- t[998] = 0
      "0000000" when "00000001111100111", -- t[999] = 0
      "0000000" when "00000001111101000", -- t[1000] = 0
      "0000000" when "00000001111101001", -- t[1001] = 0
      "0000000" when "00000001111101010", -- t[1002] = 0
      "0000000" when "00000001111101011", -- t[1003] = 0
      "0000000" when "00000001111101100", -- t[1004] = 0
      "0000000" when "00000001111101101", -- t[1005] = 0
      "0000000" when "00000001111101110", -- t[1006] = 0
      "0000000" when "00000001111101111", -- t[1007] = 0
      "0000000" when "00000001111110000", -- t[1008] = 0
      "0000000" when "00000001111110001", -- t[1009] = 0
      "0000000" when "00000001111110010", -- t[1010] = 0
      "0000000" when "00000001111110011", -- t[1011] = 0
      "0000000" when "00000001111110100", -- t[1012] = 0
      "0000000" when "00000001111110101", -- t[1013] = 0
      "0000000" when "00000001111110110", -- t[1014] = 0
      "0000000" when "00000001111110111", -- t[1015] = 0
      "0000000" when "00000001111111000", -- t[1016] = 0
      "0000000" when "00000001111111001", -- t[1017] = 0
      "0000000" when "00000001111111010", -- t[1018] = 0
      "0000000" when "00000001111111011", -- t[1019] = 0
      "0000000" when "00000001111111100", -- t[1020] = 0
      "0000000" when "00000001111111101", -- t[1021] = 0
      "0000000" when "00000001111111110", -- t[1022] = 0
      "0000000" when "00000001111111111", -- t[1023] = 0
      "0000000" when "00000010000000000", -- t[1024] = 0
      "0000000" when "00000010000000001", -- t[1025] = 0
      "0000000" when "00000010000000010", -- t[1026] = 0
      "0000000" when "00000010000000011", -- t[1027] = 0
      "0000000" when "00000010000000100", -- t[1028] = 0
      "0000000" when "00000010000000101", -- t[1029] = 0
      "0000000" when "00000010000000110", -- t[1030] = 0
      "0000000" when "00000010000000111", -- t[1031] = 0
      "0000000" when "00000010000001000", -- t[1032] = 0
      "0000000" when "00000010000001001", -- t[1033] = 0
      "0000000" when "00000010000001010", -- t[1034] = 0
      "0000000" when "00000010000001011", -- t[1035] = 0
      "0000000" when "00000010000001100", -- t[1036] = 0
      "0000000" when "00000010000001101", -- t[1037] = 0
      "0000000" when "00000010000001110", -- t[1038] = 0
      "0000000" when "00000010000001111", -- t[1039] = 0
      "0000000" when "00000010000010000", -- t[1040] = 0
      "0000000" when "00000010000010001", -- t[1041] = 0
      "0000000" when "00000010000010010", -- t[1042] = 0
      "0000000" when "00000010000010011", -- t[1043] = 0
      "0000000" when "00000010000010100", -- t[1044] = 0
      "0000000" when "00000010000010101", -- t[1045] = 0
      "0000000" when "00000010000010110", -- t[1046] = 0
      "0000000" when "00000010000010111", -- t[1047] = 0
      "0000000" when "00000010000011000", -- t[1048] = 0
      "0000000" when "00000010000011001", -- t[1049] = 0
      "0000000" when "00000010000011010", -- t[1050] = 0
      "0000000" when "00000010000011011", -- t[1051] = 0
      "0000000" when "00000010000011100", -- t[1052] = 0
      "0000000" when "00000010000011101", -- t[1053] = 0
      "0000000" when "00000010000011110", -- t[1054] = 0
      "0000000" when "00000010000011111", -- t[1055] = 0
      "0000000" when "00000010000100000", -- t[1056] = 0
      "0000000" when "00000010000100001", -- t[1057] = 0
      "0000000" when "00000010000100010", -- t[1058] = 0
      "0000000" when "00000010000100011", -- t[1059] = 0
      "0000000" when "00000010000100100", -- t[1060] = 0
      "0000000" when "00000010000100101", -- t[1061] = 0
      "0000000" when "00000010000100110", -- t[1062] = 0
      "0000000" when "00000010000100111", -- t[1063] = 0
      "0000000" when "00000010000101000", -- t[1064] = 0
      "0000000" when "00000010000101001", -- t[1065] = 0
      "0000000" when "00000010000101010", -- t[1066] = 0
      "0000000" when "00000010000101011", -- t[1067] = 0
      "0000000" when "00000010000101100", -- t[1068] = 0
      "0000000" when "00000010000101101", -- t[1069] = 0
      "0000000" when "00000010000101110", -- t[1070] = 0
      "0000000" when "00000010000101111", -- t[1071] = 0
      "0000000" when "00000010000110000", -- t[1072] = 0
      "0000000" when "00000010000110001", -- t[1073] = 0
      "0000000" when "00000010000110010", -- t[1074] = 0
      "0000000" when "00000010000110011", -- t[1075] = 0
      "0000000" when "00000010000110100", -- t[1076] = 0
      "0000000" when "00000010000110101", -- t[1077] = 0
      "0000000" when "00000010000110110", -- t[1078] = 0
      "0000000" when "00000010000110111", -- t[1079] = 0
      "0000000" when "00000010000111000", -- t[1080] = 0
      "0000000" when "00000010000111001", -- t[1081] = 0
      "0000000" when "00000010000111010", -- t[1082] = 0
      "0000000" when "00000010000111011", -- t[1083] = 0
      "0000000" when "00000010000111100", -- t[1084] = 0
      "0000000" when "00000010000111101", -- t[1085] = 0
      "0000000" when "00000010000111110", -- t[1086] = 0
      "0000000" when "00000010000111111", -- t[1087] = 0
      "0000000" when "00000010001000000", -- t[1088] = 0
      "0000000" when "00000010001000001", -- t[1089] = 0
      "0000000" when "00000010001000010", -- t[1090] = 0
      "0000000" when "00000010001000011", -- t[1091] = 0
      "0000000" when "00000010001000100", -- t[1092] = 0
      "0000000" when "00000010001000101", -- t[1093] = 0
      "0000000" when "00000010001000110", -- t[1094] = 0
      "0000000" when "00000010001000111", -- t[1095] = 0
      "0000000" when "00000010001001000", -- t[1096] = 0
      "0000000" when "00000010001001001", -- t[1097] = 0
      "0000000" when "00000010001001010", -- t[1098] = 0
      "0000000" when "00000010001001011", -- t[1099] = 0
      "0000000" when "00000010001001100", -- t[1100] = 0
      "0000000" when "00000010001001101", -- t[1101] = 0
      "0000000" when "00000010001001110", -- t[1102] = 0
      "0000000" when "00000010001001111", -- t[1103] = 0
      "0000000" when "00000010001010000", -- t[1104] = 0
      "0000000" when "00000010001010001", -- t[1105] = 0
      "0000000" when "00000010001010010", -- t[1106] = 0
      "0000000" when "00000010001010011", -- t[1107] = 0
      "0000000" when "00000010001010100", -- t[1108] = 0
      "0000000" when "00000010001010101", -- t[1109] = 0
      "0000000" when "00000010001010110", -- t[1110] = 0
      "0000000" when "00000010001010111", -- t[1111] = 0
      "0000000" when "00000010001011000", -- t[1112] = 0
      "0000000" when "00000010001011001", -- t[1113] = 0
      "0000000" when "00000010001011010", -- t[1114] = 0
      "0000000" when "00000010001011011", -- t[1115] = 0
      "0000000" when "00000010001011100", -- t[1116] = 0
      "0000000" when "00000010001011101", -- t[1117] = 0
      "0000000" when "00000010001011110", -- t[1118] = 0
      "0000000" when "00000010001011111", -- t[1119] = 0
      "0000000" when "00000010001100000", -- t[1120] = 0
      "0000000" when "00000010001100001", -- t[1121] = 0
      "0000000" when "00000010001100010", -- t[1122] = 0
      "0000000" when "00000010001100011", -- t[1123] = 0
      "0000000" when "00000010001100100", -- t[1124] = 0
      "0000000" when "00000010001100101", -- t[1125] = 0
      "0000000" when "00000010001100110", -- t[1126] = 0
      "0000000" when "00000010001100111", -- t[1127] = 0
      "0000000" when "00000010001101000", -- t[1128] = 0
      "0000000" when "00000010001101001", -- t[1129] = 0
      "0000000" when "00000010001101010", -- t[1130] = 0
      "0000000" when "00000010001101011", -- t[1131] = 0
      "0000000" when "00000010001101100", -- t[1132] = 0
      "0000000" when "00000010001101101", -- t[1133] = 0
      "0000000" when "00000010001101110", -- t[1134] = 0
      "0000000" when "00000010001101111", -- t[1135] = 0
      "0000000" when "00000010001110000", -- t[1136] = 0
      "0000000" when "00000010001110001", -- t[1137] = 0
      "0000000" when "00000010001110010", -- t[1138] = 0
      "0000000" when "00000010001110011", -- t[1139] = 0
      "0000000" when "00000010001110100", -- t[1140] = 0
      "0000000" when "00000010001110101", -- t[1141] = 0
      "0000000" when "00000010001110110", -- t[1142] = 0
      "0000000" when "00000010001110111", -- t[1143] = 0
      "0000000" when "00000010001111000", -- t[1144] = 0
      "0000000" when "00000010001111001", -- t[1145] = 0
      "0000000" when "00000010001111010", -- t[1146] = 0
      "0000000" when "00000010001111011", -- t[1147] = 0
      "0000000" when "00000010001111100", -- t[1148] = 0
      "0000000" when "00000010001111101", -- t[1149] = 0
      "0000000" when "00000010001111110", -- t[1150] = 0
      "0000000" when "00000010001111111", -- t[1151] = 0
      "0000000" when "00000010010000000", -- t[1152] = 0
      "0000000" when "00000010010000001", -- t[1153] = 0
      "0000000" when "00000010010000010", -- t[1154] = 0
      "0000000" when "00000010010000011", -- t[1155] = 0
      "0000000" when "00000010010000100", -- t[1156] = 0
      "0000000" when "00000010010000101", -- t[1157] = 0
      "0000000" when "00000010010000110", -- t[1158] = 0
      "0000000" when "00000010010000111", -- t[1159] = 0
      "0000000" when "00000010010001000", -- t[1160] = 0
      "0000000" when "00000010010001001", -- t[1161] = 0
      "0000000" when "00000010010001010", -- t[1162] = 0
      "0000000" when "00000010010001011", -- t[1163] = 0
      "0000000" when "00000010010001100", -- t[1164] = 0
      "0000000" when "00000010010001101", -- t[1165] = 0
      "0000000" when "00000010010001110", -- t[1166] = 0
      "0000000" when "00000010010001111", -- t[1167] = 0
      "0000000" when "00000010010010000", -- t[1168] = 0
      "0000000" when "00000010010010001", -- t[1169] = 0
      "0000000" when "00000010010010010", -- t[1170] = 0
      "0000000" when "00000010010010011", -- t[1171] = 0
      "0000000" when "00000010010010100", -- t[1172] = 0
      "0000000" when "00000010010010101", -- t[1173] = 0
      "0000000" when "00000010010010110", -- t[1174] = 0
      "0000000" when "00000010010010111", -- t[1175] = 0
      "0000000" when "00000010010011000", -- t[1176] = 0
      "0000000" when "00000010010011001", -- t[1177] = 0
      "0000000" when "00000010010011010", -- t[1178] = 0
      "0000000" when "00000010010011011", -- t[1179] = 0
      "0000000" when "00000010010011100", -- t[1180] = 0
      "0000000" when "00000010010011101", -- t[1181] = 0
      "0000000" when "00000010010011110", -- t[1182] = 0
      "0000000" when "00000010010011111", -- t[1183] = 0
      "0000000" when "00000010010100000", -- t[1184] = 0
      "0000000" when "00000010010100001", -- t[1185] = 0
      "0000000" when "00000010010100010", -- t[1186] = 0
      "0000000" when "00000010010100011", -- t[1187] = 0
      "0000000" when "00000010010100100", -- t[1188] = 0
      "0000000" when "00000010010100101", -- t[1189] = 0
      "0000000" when "00000010010100110", -- t[1190] = 0
      "0000000" when "00000010010100111", -- t[1191] = 0
      "0000000" when "00000010010101000", -- t[1192] = 0
      "0000000" when "00000010010101001", -- t[1193] = 0
      "0000000" when "00000010010101010", -- t[1194] = 0
      "0000000" when "00000010010101011", -- t[1195] = 0
      "0000000" when "00000010010101100", -- t[1196] = 0
      "0000000" when "00000010010101101", -- t[1197] = 0
      "0000000" when "00000010010101110", -- t[1198] = 0
      "0000000" when "00000010010101111", -- t[1199] = 0
      "0000000" when "00000010010110000", -- t[1200] = 0
      "0000000" when "00000010010110001", -- t[1201] = 0
      "0000000" when "00000010010110010", -- t[1202] = 0
      "0000000" when "00000010010110011", -- t[1203] = 0
      "0000000" when "00000010010110100", -- t[1204] = 0
      "0000000" when "00000010010110101", -- t[1205] = 0
      "0000000" when "00000010010110110", -- t[1206] = 0
      "0000000" when "00000010010110111", -- t[1207] = 0
      "0000000" when "00000010010111000", -- t[1208] = 0
      "0000000" when "00000010010111001", -- t[1209] = 0
      "0000000" when "00000010010111010", -- t[1210] = 0
      "0000000" when "00000010010111011", -- t[1211] = 0
      "0000000" when "00000010010111100", -- t[1212] = 0
      "0000000" when "00000010010111101", -- t[1213] = 0
      "0000000" when "00000010010111110", -- t[1214] = 0
      "0000000" when "00000010010111111", -- t[1215] = 0
      "0000000" when "00000010011000000", -- t[1216] = 0
      "0000000" when "00000010011000001", -- t[1217] = 0
      "0000000" when "00000010011000010", -- t[1218] = 0
      "0000000" when "00000010011000011", -- t[1219] = 0
      "0000000" when "00000010011000100", -- t[1220] = 0
      "0000000" when "00000010011000101", -- t[1221] = 0
      "0000000" when "00000010011000110", -- t[1222] = 0
      "0000000" when "00000010011000111", -- t[1223] = 0
      "0000000" when "00000010011001000", -- t[1224] = 0
      "0000000" when "00000010011001001", -- t[1225] = 0
      "0000000" when "00000010011001010", -- t[1226] = 0
      "0000000" when "00000010011001011", -- t[1227] = 0
      "0000000" when "00000010011001100", -- t[1228] = 0
      "0000000" when "00000010011001101", -- t[1229] = 0
      "0000000" when "00000010011001110", -- t[1230] = 0
      "0000000" when "00000010011001111", -- t[1231] = 0
      "0000000" when "00000010011010000", -- t[1232] = 0
      "0000000" when "00000010011010001", -- t[1233] = 0
      "0000000" when "00000010011010010", -- t[1234] = 0
      "0000000" when "00000010011010011", -- t[1235] = 0
      "0000000" when "00000010011010100", -- t[1236] = 0
      "0000000" when "00000010011010101", -- t[1237] = 0
      "0000000" when "00000010011010110", -- t[1238] = 0
      "0000000" when "00000010011010111", -- t[1239] = 0
      "0000000" when "00000010011011000", -- t[1240] = 0
      "0000000" when "00000010011011001", -- t[1241] = 0
      "0000000" when "00000010011011010", -- t[1242] = 0
      "0000000" when "00000010011011011", -- t[1243] = 0
      "0000000" when "00000010011011100", -- t[1244] = 0
      "0000000" when "00000010011011101", -- t[1245] = 0
      "0000000" when "00000010011011110", -- t[1246] = 0
      "0000000" when "00000010011011111", -- t[1247] = 0
      "0000000" when "00000010011100000", -- t[1248] = 0
      "0000000" when "00000010011100001", -- t[1249] = 0
      "0000000" when "00000010011100010", -- t[1250] = 0
      "0000000" when "00000010011100011", -- t[1251] = 0
      "0000000" when "00000010011100100", -- t[1252] = 0
      "0000000" when "00000010011100101", -- t[1253] = 0
      "0000000" when "00000010011100110", -- t[1254] = 0
      "0000000" when "00000010011100111", -- t[1255] = 0
      "0000000" when "00000010011101000", -- t[1256] = 0
      "0000000" when "00000010011101001", -- t[1257] = 0
      "0000000" when "00000010011101010", -- t[1258] = 0
      "0000000" when "00000010011101011", -- t[1259] = 0
      "0000000" when "00000010011101100", -- t[1260] = 0
      "0000000" when "00000010011101101", -- t[1261] = 0
      "0000000" when "00000010011101110", -- t[1262] = 0
      "0000000" when "00000010011101111", -- t[1263] = 0
      "0000000" when "00000010011110000", -- t[1264] = 0
      "0000000" when "00000010011110001", -- t[1265] = 0
      "0000000" when "00000010011110010", -- t[1266] = 0
      "0000000" when "00000010011110011", -- t[1267] = 0
      "0000000" when "00000010011110100", -- t[1268] = 0
      "0000000" when "00000010011110101", -- t[1269] = 0
      "0000000" when "00000010011110110", -- t[1270] = 0
      "0000000" when "00000010011110111", -- t[1271] = 0
      "0000000" when "00000010011111000", -- t[1272] = 0
      "0000000" when "00000010011111001", -- t[1273] = 0
      "0000000" when "00000010011111010", -- t[1274] = 0
      "0000000" when "00000010011111011", -- t[1275] = 0
      "0000000" when "00000010011111100", -- t[1276] = 0
      "0000000" when "00000010011111101", -- t[1277] = 0
      "0000000" when "00000010011111110", -- t[1278] = 0
      "0000000" when "00000010011111111", -- t[1279] = 0
      "0000000" when "00000010100000000", -- t[1280] = 0
      "0000000" when "00000010100000001", -- t[1281] = 0
      "0000000" when "00000010100000010", -- t[1282] = 0
      "0000000" when "00000010100000011", -- t[1283] = 0
      "0000000" when "00000010100000100", -- t[1284] = 0
      "0000000" when "00000010100000101", -- t[1285] = 0
      "0000000" when "00000010100000110", -- t[1286] = 0
      "0000000" when "00000010100000111", -- t[1287] = 0
      "0000000" when "00000010100001000", -- t[1288] = 0
      "0000000" when "00000010100001001", -- t[1289] = 0
      "0000000" when "00000010100001010", -- t[1290] = 0
      "0000000" when "00000010100001011", -- t[1291] = 0
      "0000000" when "00000010100001100", -- t[1292] = 0
      "0000000" when "00000010100001101", -- t[1293] = 0
      "0000000" when "00000010100001110", -- t[1294] = 0
      "0000000" when "00000010100001111", -- t[1295] = 0
      "0000000" when "00000010100010000", -- t[1296] = 0
      "0000000" when "00000010100010001", -- t[1297] = 0
      "0000000" when "00000010100010010", -- t[1298] = 0
      "0000000" when "00000010100010011", -- t[1299] = 0
      "0000000" when "00000010100010100", -- t[1300] = 0
      "0000000" when "00000010100010101", -- t[1301] = 0
      "0000000" when "00000010100010110", -- t[1302] = 0
      "0000000" when "00000010100010111", -- t[1303] = 0
      "0000000" when "00000010100011000", -- t[1304] = 0
      "0000000" when "00000010100011001", -- t[1305] = 0
      "0000000" when "00000010100011010", -- t[1306] = 0
      "0000000" when "00000010100011011", -- t[1307] = 0
      "0000000" when "00000010100011100", -- t[1308] = 0
      "0000000" when "00000010100011101", -- t[1309] = 0
      "0000000" when "00000010100011110", -- t[1310] = 0
      "0000000" when "00000010100011111", -- t[1311] = 0
      "0000000" when "00000010100100000", -- t[1312] = 0
      "0000000" when "00000010100100001", -- t[1313] = 0
      "0000000" when "00000010100100010", -- t[1314] = 0
      "0000000" when "00000010100100011", -- t[1315] = 0
      "0000000" when "00000010100100100", -- t[1316] = 0
      "0000000" when "00000010100100101", -- t[1317] = 0
      "0000000" when "00000010100100110", -- t[1318] = 0
      "0000000" when "00000010100100111", -- t[1319] = 0
      "0000000" when "00000010100101000", -- t[1320] = 0
      "0000000" when "00000010100101001", -- t[1321] = 0
      "0000000" when "00000010100101010", -- t[1322] = 0
      "0000000" when "00000010100101011", -- t[1323] = 0
      "0000000" when "00000010100101100", -- t[1324] = 0
      "0000000" when "00000010100101101", -- t[1325] = 0
      "0000000" when "00000010100101110", -- t[1326] = 0
      "0000000" when "00000010100101111", -- t[1327] = 0
      "0000000" when "00000010100110000", -- t[1328] = 0
      "0000000" when "00000010100110001", -- t[1329] = 0
      "0000000" when "00000010100110010", -- t[1330] = 0
      "0000000" when "00000010100110011", -- t[1331] = 0
      "0000000" when "00000010100110100", -- t[1332] = 0
      "0000000" when "00000010100110101", -- t[1333] = 0
      "0000000" when "00000010100110110", -- t[1334] = 0
      "0000000" when "00000010100110111", -- t[1335] = 0
      "0000000" when "00000010100111000", -- t[1336] = 0
      "0000000" when "00000010100111001", -- t[1337] = 0
      "0000000" when "00000010100111010", -- t[1338] = 0
      "0000000" when "00000010100111011", -- t[1339] = 0
      "0000000" when "00000010100111100", -- t[1340] = 0
      "0000000" when "00000010100111101", -- t[1341] = 0
      "0000000" when "00000010100111110", -- t[1342] = 0
      "0000000" when "00000010100111111", -- t[1343] = 0
      "0000000" when "00000010101000000", -- t[1344] = 0
      "0000000" when "00000010101000001", -- t[1345] = 0
      "0000000" when "00000010101000010", -- t[1346] = 0
      "0000000" when "00000010101000011", -- t[1347] = 0
      "0000000" when "00000010101000100", -- t[1348] = 0
      "0000000" when "00000010101000101", -- t[1349] = 0
      "0000000" when "00000010101000110", -- t[1350] = 0
      "0000000" when "00000010101000111", -- t[1351] = 0
      "0000000" when "00000010101001000", -- t[1352] = 0
      "0000000" when "00000010101001001", -- t[1353] = 0
      "0000000" when "00000010101001010", -- t[1354] = 0
      "0000000" when "00000010101001011", -- t[1355] = 0
      "0000000" when "00000010101001100", -- t[1356] = 0
      "0000000" when "00000010101001101", -- t[1357] = 0
      "0000000" when "00000010101001110", -- t[1358] = 0
      "0000000" when "00000010101001111", -- t[1359] = 0
      "0000000" when "00000010101010000", -- t[1360] = 0
      "0000000" when "00000010101010001", -- t[1361] = 0
      "0000000" when "00000010101010010", -- t[1362] = 0
      "0000000" when "00000010101010011", -- t[1363] = 0
      "0000000" when "00000010101010100", -- t[1364] = 0
      "0000000" when "00000010101010101", -- t[1365] = 0
      "0000000" when "00000010101010110", -- t[1366] = 0
      "0000000" when "00000010101010111", -- t[1367] = 0
      "0000000" when "00000010101011000", -- t[1368] = 0
      "0000000" when "00000010101011001", -- t[1369] = 0
      "0000000" when "00000010101011010", -- t[1370] = 0
      "0000000" when "00000010101011011", -- t[1371] = 0
      "0000000" when "00000010101011100", -- t[1372] = 0
      "0000000" when "00000010101011101", -- t[1373] = 0
      "0000000" when "00000010101011110", -- t[1374] = 0
      "0000000" when "00000010101011111", -- t[1375] = 0
      "0000000" when "00000010101100000", -- t[1376] = 0
      "0000000" when "00000010101100001", -- t[1377] = 0
      "0000000" when "00000010101100010", -- t[1378] = 0
      "0000000" when "00000010101100011", -- t[1379] = 0
      "0000000" when "00000010101100100", -- t[1380] = 0
      "0000000" when "00000010101100101", -- t[1381] = 0
      "0000000" when "00000010101100110", -- t[1382] = 0
      "0000000" when "00000010101100111", -- t[1383] = 0
      "0000000" when "00000010101101000", -- t[1384] = 0
      "0000000" when "00000010101101001", -- t[1385] = 0
      "0000000" when "00000010101101010", -- t[1386] = 0
      "0000000" when "00000010101101011", -- t[1387] = 0
      "0000000" when "00000010101101100", -- t[1388] = 0
      "0000000" when "00000010101101101", -- t[1389] = 0
      "0000000" when "00000010101101110", -- t[1390] = 0
      "0000000" when "00000010101101111", -- t[1391] = 0
      "0000000" when "00000010101110000", -- t[1392] = 0
      "0000000" when "00000010101110001", -- t[1393] = 0
      "0000000" when "00000010101110010", -- t[1394] = 0
      "0000000" when "00000010101110011", -- t[1395] = 0
      "0000000" when "00000010101110100", -- t[1396] = 0
      "0000000" when "00000010101110101", -- t[1397] = 0
      "0000000" when "00000010101110110", -- t[1398] = 0
      "0000000" when "00000010101110111", -- t[1399] = 0
      "0000000" when "00000010101111000", -- t[1400] = 0
      "0000000" when "00000010101111001", -- t[1401] = 0
      "0000000" when "00000010101111010", -- t[1402] = 0
      "0000000" when "00000010101111011", -- t[1403] = 0
      "0000000" when "00000010101111100", -- t[1404] = 0
      "0000000" when "00000010101111101", -- t[1405] = 0
      "0000000" when "00000010101111110", -- t[1406] = 0
      "0000000" when "00000010101111111", -- t[1407] = 0
      "0000000" when "00000010110000000", -- t[1408] = 0
      "0000000" when "00000010110000001", -- t[1409] = 0
      "0000000" when "00000010110000010", -- t[1410] = 0
      "0000000" when "00000010110000011", -- t[1411] = 0
      "0000000" when "00000010110000100", -- t[1412] = 0
      "0000000" when "00000010110000101", -- t[1413] = 0
      "0000000" when "00000010110000110", -- t[1414] = 0
      "0000000" when "00000010110000111", -- t[1415] = 0
      "0000000" when "00000010110001000", -- t[1416] = 0
      "0000000" when "00000010110001001", -- t[1417] = 0
      "0000000" when "00000010110001010", -- t[1418] = 0
      "0000000" when "00000010110001011", -- t[1419] = 0
      "0000000" when "00000010110001100", -- t[1420] = 0
      "0000000" when "00000010110001101", -- t[1421] = 0
      "0000000" when "00000010110001110", -- t[1422] = 0
      "0000000" when "00000010110001111", -- t[1423] = 0
      "0000000" when "00000010110010000", -- t[1424] = 0
      "0000000" when "00000010110010001", -- t[1425] = 0
      "0000000" when "00000010110010010", -- t[1426] = 0
      "0000000" when "00000010110010011", -- t[1427] = 0
      "0000000" when "00000010110010100", -- t[1428] = 0
      "0000000" when "00000010110010101", -- t[1429] = 0
      "0000000" when "00000010110010110", -- t[1430] = 0
      "0000000" when "00000010110010111", -- t[1431] = 0
      "0000000" when "00000010110011000", -- t[1432] = 0
      "0000000" when "00000010110011001", -- t[1433] = 0
      "0000000" when "00000010110011010", -- t[1434] = 0
      "0000000" when "00000010110011011", -- t[1435] = 0
      "0000000" when "00000010110011100", -- t[1436] = 0
      "0000000" when "00000010110011101", -- t[1437] = 0
      "0000000" when "00000010110011110", -- t[1438] = 0
      "0000000" when "00000010110011111", -- t[1439] = 0
      "0000000" when "00000010110100000", -- t[1440] = 0
      "0000000" when "00000010110100001", -- t[1441] = 0
      "0000000" when "00000010110100010", -- t[1442] = 0
      "0000000" when "00000010110100011", -- t[1443] = 0
      "0000000" when "00000010110100100", -- t[1444] = 0
      "0000000" when "00000010110100101", -- t[1445] = 0
      "0000000" when "00000010110100110", -- t[1446] = 0
      "0000000" when "00000010110100111", -- t[1447] = 0
      "0000000" when "00000010110101000", -- t[1448] = 0
      "0000000" when "00000010110101001", -- t[1449] = 0
      "0000000" when "00000010110101010", -- t[1450] = 0
      "0000000" when "00000010110101011", -- t[1451] = 0
      "0000000" when "00000010110101100", -- t[1452] = 0
      "0000000" when "00000010110101101", -- t[1453] = 0
      "0000000" when "00000010110101110", -- t[1454] = 0
      "0000000" when "00000010110101111", -- t[1455] = 0
      "0000000" when "00000010110110000", -- t[1456] = 0
      "0000000" when "00000010110110001", -- t[1457] = 0
      "0000000" when "00000010110110010", -- t[1458] = 0
      "0000000" when "00000010110110011", -- t[1459] = 0
      "0000000" when "00000010110110100", -- t[1460] = 0
      "0000000" when "00000010110110101", -- t[1461] = 0
      "0000000" when "00000010110110110", -- t[1462] = 0
      "0000000" when "00000010110110111", -- t[1463] = 0
      "0000000" when "00000010110111000", -- t[1464] = 0
      "0000000" when "00000010110111001", -- t[1465] = 0
      "0000000" when "00000010110111010", -- t[1466] = 0
      "0000000" when "00000010110111011", -- t[1467] = 0
      "0000000" when "00000010110111100", -- t[1468] = 0
      "0000000" when "00000010110111101", -- t[1469] = 0
      "0000000" when "00000010110111110", -- t[1470] = 0
      "0000000" when "00000010110111111", -- t[1471] = 0
      "0000000" when "00000010111000000", -- t[1472] = 0
      "0000000" when "00000010111000001", -- t[1473] = 0
      "0000000" when "00000010111000010", -- t[1474] = 0
      "0000000" when "00000010111000011", -- t[1475] = 0
      "0000000" when "00000010111000100", -- t[1476] = 0
      "0000000" when "00000010111000101", -- t[1477] = 0
      "0000000" when "00000010111000110", -- t[1478] = 0
      "0000000" when "00000010111000111", -- t[1479] = 0
      "0000000" when "00000010111001000", -- t[1480] = 0
      "0000000" when "00000010111001001", -- t[1481] = 0
      "0000000" when "00000010111001010", -- t[1482] = 0
      "0000000" when "00000010111001011", -- t[1483] = 0
      "0000000" when "00000010111001100", -- t[1484] = 0
      "0000000" when "00000010111001101", -- t[1485] = 0
      "0000000" when "00000010111001110", -- t[1486] = 0
      "0000000" when "00000010111001111", -- t[1487] = 0
      "0000000" when "00000010111010000", -- t[1488] = 0
      "0000000" when "00000010111010001", -- t[1489] = 0
      "0000000" when "00000010111010010", -- t[1490] = 0
      "0000000" when "00000010111010011", -- t[1491] = 0
      "0000000" when "00000010111010100", -- t[1492] = 0
      "0000000" when "00000010111010101", -- t[1493] = 0
      "0000000" when "00000010111010110", -- t[1494] = 0
      "0000000" when "00000010111010111", -- t[1495] = 0
      "0000000" when "00000010111011000", -- t[1496] = 0
      "0000000" when "00000010111011001", -- t[1497] = 0
      "0000000" when "00000010111011010", -- t[1498] = 0
      "0000000" when "00000010111011011", -- t[1499] = 0
      "0000000" when "00000010111011100", -- t[1500] = 0
      "0000000" when "00000010111011101", -- t[1501] = 0
      "0000000" when "00000010111011110", -- t[1502] = 0
      "0000000" when "00000010111011111", -- t[1503] = 0
      "0000000" when "00000010111100000", -- t[1504] = 0
      "0000000" when "00000010111100001", -- t[1505] = 0
      "0000000" when "00000010111100010", -- t[1506] = 0
      "0000000" when "00000010111100011", -- t[1507] = 0
      "0000000" when "00000010111100100", -- t[1508] = 0
      "0000000" when "00000010111100101", -- t[1509] = 0
      "0000000" when "00000010111100110", -- t[1510] = 0
      "0000000" when "00000010111100111", -- t[1511] = 0
      "0000000" when "00000010111101000", -- t[1512] = 0
      "0000000" when "00000010111101001", -- t[1513] = 0
      "0000000" when "00000010111101010", -- t[1514] = 0
      "0000000" when "00000010111101011", -- t[1515] = 0
      "0000000" when "00000010111101100", -- t[1516] = 0
      "0000000" when "00000010111101101", -- t[1517] = 0
      "0000000" when "00000010111101110", -- t[1518] = 0
      "0000000" when "00000010111101111", -- t[1519] = 0
      "0000000" when "00000010111110000", -- t[1520] = 0
      "0000000" when "00000010111110001", -- t[1521] = 0
      "0000000" when "00000010111110010", -- t[1522] = 0
      "0000000" when "00000010111110011", -- t[1523] = 0
      "0000000" when "00000010111110100", -- t[1524] = 0
      "0000000" when "00000010111110101", -- t[1525] = 0
      "0000000" when "00000010111110110", -- t[1526] = 0
      "0000000" when "00000010111110111", -- t[1527] = 0
      "0000000" when "00000010111111000", -- t[1528] = 0
      "0000000" when "00000010111111001", -- t[1529] = 0
      "0000000" when "00000010111111010", -- t[1530] = 0
      "0000000" when "00000010111111011", -- t[1531] = 0
      "0000000" when "00000010111111100", -- t[1532] = 0
      "0000000" when "00000010111111101", -- t[1533] = 0
      "0000000" when "00000010111111110", -- t[1534] = 0
      "0000000" when "00000010111111111", -- t[1535] = 0
      "0000000" when "00000011000000000", -- t[1536] = 0
      "0000000" when "00000011000000001", -- t[1537] = 0
      "0000000" when "00000011000000010", -- t[1538] = 0
      "0000000" when "00000011000000011", -- t[1539] = 0
      "0000000" when "00000011000000100", -- t[1540] = 0
      "0000000" when "00000011000000101", -- t[1541] = 0
      "0000000" when "00000011000000110", -- t[1542] = 0
      "0000000" when "00000011000000111", -- t[1543] = 0
      "0000000" when "00000011000001000", -- t[1544] = 0
      "0000000" when "00000011000001001", -- t[1545] = 0
      "0000000" when "00000011000001010", -- t[1546] = 0
      "0000000" when "00000011000001011", -- t[1547] = 0
      "0000000" when "00000011000001100", -- t[1548] = 0
      "0000000" when "00000011000001101", -- t[1549] = 0
      "0000000" when "00000011000001110", -- t[1550] = 0
      "0000000" when "00000011000001111", -- t[1551] = 0
      "0000000" when "00000011000010000", -- t[1552] = 0
      "0000000" when "00000011000010001", -- t[1553] = 0
      "0000000" when "00000011000010010", -- t[1554] = 0
      "0000000" when "00000011000010011", -- t[1555] = 0
      "0000000" when "00000011000010100", -- t[1556] = 0
      "0000000" when "00000011000010101", -- t[1557] = 0
      "0000000" when "00000011000010110", -- t[1558] = 0
      "0000000" when "00000011000010111", -- t[1559] = 0
      "0000000" when "00000011000011000", -- t[1560] = 0
      "0000000" when "00000011000011001", -- t[1561] = 0
      "0000000" when "00000011000011010", -- t[1562] = 0
      "0000000" when "00000011000011011", -- t[1563] = 0
      "0000000" when "00000011000011100", -- t[1564] = 0
      "0000000" when "00000011000011101", -- t[1565] = 0
      "0000000" when "00000011000011110", -- t[1566] = 0
      "0000000" when "00000011000011111", -- t[1567] = 0
      "0000000" when "00000011000100000", -- t[1568] = 0
      "0000000" when "00000011000100001", -- t[1569] = 0
      "0000000" when "00000011000100010", -- t[1570] = 0
      "0000000" when "00000011000100011", -- t[1571] = 0
      "0000000" when "00000011000100100", -- t[1572] = 0
      "0000000" when "00000011000100101", -- t[1573] = 0
      "0000000" when "00000011000100110", -- t[1574] = 0
      "0000000" when "00000011000100111", -- t[1575] = 0
      "0000000" when "00000011000101000", -- t[1576] = 0
      "0000000" when "00000011000101001", -- t[1577] = 0
      "0000000" when "00000011000101010", -- t[1578] = 0
      "0000000" when "00000011000101011", -- t[1579] = 0
      "0000000" when "00000011000101100", -- t[1580] = 0
      "0000000" when "00000011000101101", -- t[1581] = 0
      "0000000" when "00000011000101110", -- t[1582] = 0
      "0000000" when "00000011000101111", -- t[1583] = 0
      "0000000" when "00000011000110000", -- t[1584] = 0
      "0000000" when "00000011000110001", -- t[1585] = 0
      "0000000" when "00000011000110010", -- t[1586] = 0
      "0000000" when "00000011000110011", -- t[1587] = 0
      "0000000" when "00000011000110100", -- t[1588] = 0
      "0000000" when "00000011000110101", -- t[1589] = 0
      "0000000" when "00000011000110110", -- t[1590] = 0
      "0000000" when "00000011000110111", -- t[1591] = 0
      "0000000" when "00000011000111000", -- t[1592] = 0
      "0000000" when "00000011000111001", -- t[1593] = 0
      "0000000" when "00000011000111010", -- t[1594] = 0
      "0000000" when "00000011000111011", -- t[1595] = 0
      "0000000" when "00000011000111100", -- t[1596] = 0
      "0000000" when "00000011000111101", -- t[1597] = 0
      "0000000" when "00000011000111110", -- t[1598] = 0
      "0000000" when "00000011000111111", -- t[1599] = 0
      "0000000" when "00000011001000000", -- t[1600] = 0
      "0000000" when "00000011001000001", -- t[1601] = 0
      "0000000" when "00000011001000010", -- t[1602] = 0
      "0000000" when "00000011001000011", -- t[1603] = 0
      "0000000" when "00000011001000100", -- t[1604] = 0
      "0000000" when "00000011001000101", -- t[1605] = 0
      "0000000" when "00000011001000110", -- t[1606] = 0
      "0000000" when "00000011001000111", -- t[1607] = 0
      "0000000" when "00000011001001000", -- t[1608] = 0
      "0000000" when "00000011001001001", -- t[1609] = 0
      "0000000" when "00000011001001010", -- t[1610] = 0
      "0000000" when "00000011001001011", -- t[1611] = 0
      "0000000" when "00000011001001100", -- t[1612] = 0
      "0000000" when "00000011001001101", -- t[1613] = 0
      "0000000" when "00000011001001110", -- t[1614] = 0
      "0000000" when "00000011001001111", -- t[1615] = 0
      "0000000" when "00000011001010000", -- t[1616] = 0
      "0000000" when "00000011001010001", -- t[1617] = 0
      "0000000" when "00000011001010010", -- t[1618] = 0
      "0000000" when "00000011001010011", -- t[1619] = 0
      "0000000" when "00000011001010100", -- t[1620] = 0
      "0000000" when "00000011001010101", -- t[1621] = 0
      "0000000" when "00000011001010110", -- t[1622] = 0
      "0000000" when "00000011001010111", -- t[1623] = 0
      "0000000" when "00000011001011000", -- t[1624] = 0
      "0000000" when "00000011001011001", -- t[1625] = 0
      "0000000" when "00000011001011010", -- t[1626] = 0
      "0000000" when "00000011001011011", -- t[1627] = 0
      "0000000" when "00000011001011100", -- t[1628] = 0
      "0000000" when "00000011001011101", -- t[1629] = 0
      "0000000" when "00000011001011110", -- t[1630] = 0
      "0000000" when "00000011001011111", -- t[1631] = 0
      "0000000" when "00000011001100000", -- t[1632] = 0
      "0000000" when "00000011001100001", -- t[1633] = 0
      "0000000" when "00000011001100010", -- t[1634] = 0
      "0000000" when "00000011001100011", -- t[1635] = 0
      "0000000" when "00000011001100100", -- t[1636] = 0
      "0000000" when "00000011001100101", -- t[1637] = 0
      "0000000" when "00000011001100110", -- t[1638] = 0
      "0000000" when "00000011001100111", -- t[1639] = 0
      "0000000" when "00000011001101000", -- t[1640] = 0
      "0000000" when "00000011001101001", -- t[1641] = 0
      "0000000" when "00000011001101010", -- t[1642] = 0
      "0000000" when "00000011001101011", -- t[1643] = 0
      "0000000" when "00000011001101100", -- t[1644] = 0
      "0000000" when "00000011001101101", -- t[1645] = 0
      "0000000" when "00000011001101110", -- t[1646] = 0
      "0000000" when "00000011001101111", -- t[1647] = 0
      "0000000" when "00000011001110000", -- t[1648] = 0
      "0000000" when "00000011001110001", -- t[1649] = 0
      "0000000" when "00000011001110010", -- t[1650] = 0
      "0000000" when "00000011001110011", -- t[1651] = 0
      "0000000" when "00000011001110100", -- t[1652] = 0
      "0000000" when "00000011001110101", -- t[1653] = 0
      "0000000" when "00000011001110110", -- t[1654] = 0
      "0000000" when "00000011001110111", -- t[1655] = 0
      "0000000" when "00000011001111000", -- t[1656] = 0
      "0000000" when "00000011001111001", -- t[1657] = 0
      "0000000" when "00000011001111010", -- t[1658] = 0
      "0000000" when "00000011001111011", -- t[1659] = 0
      "0000000" when "00000011001111100", -- t[1660] = 0
      "0000000" when "00000011001111101", -- t[1661] = 0
      "0000000" when "00000011001111110", -- t[1662] = 0
      "0000000" when "00000011001111111", -- t[1663] = 0
      "0000000" when "00000011010000000", -- t[1664] = 0
      "0000000" when "00000011010000001", -- t[1665] = 0
      "0000000" when "00000011010000010", -- t[1666] = 0
      "0000000" when "00000011010000011", -- t[1667] = 0
      "0000000" when "00000011010000100", -- t[1668] = 0
      "0000000" when "00000011010000101", -- t[1669] = 0
      "0000000" when "00000011010000110", -- t[1670] = 0
      "0000000" when "00000011010000111", -- t[1671] = 0
      "0000000" when "00000011010001000", -- t[1672] = 0
      "0000000" when "00000011010001001", -- t[1673] = 0
      "0000000" when "00000011010001010", -- t[1674] = 0
      "0000000" when "00000011010001011", -- t[1675] = 0
      "0000000" when "00000011010001100", -- t[1676] = 0
      "0000000" when "00000011010001101", -- t[1677] = 0
      "0000000" when "00000011010001110", -- t[1678] = 0
      "0000000" when "00000011010001111", -- t[1679] = 0
      "0000000" when "00000011010010000", -- t[1680] = 0
      "0000000" when "00000011010010001", -- t[1681] = 0
      "0000000" when "00000011010010010", -- t[1682] = 0
      "0000000" when "00000011010010011", -- t[1683] = 0
      "0000000" when "00000011010010100", -- t[1684] = 0
      "0000000" when "00000011010010101", -- t[1685] = 0
      "0000000" when "00000011010010110", -- t[1686] = 0
      "0000000" when "00000011010010111", -- t[1687] = 0
      "0000000" when "00000011010011000", -- t[1688] = 0
      "0000000" when "00000011010011001", -- t[1689] = 0
      "0000000" when "00000011010011010", -- t[1690] = 0
      "0000000" when "00000011010011011", -- t[1691] = 0
      "0000000" when "00000011010011100", -- t[1692] = 0
      "0000000" when "00000011010011101", -- t[1693] = 0
      "0000000" when "00000011010011110", -- t[1694] = 0
      "0000000" when "00000011010011111", -- t[1695] = 0
      "0000000" when "00000011010100000", -- t[1696] = 0
      "0000000" when "00000011010100001", -- t[1697] = 0
      "0000000" when "00000011010100010", -- t[1698] = 0
      "0000000" when "00000011010100011", -- t[1699] = 0
      "0000000" when "00000011010100100", -- t[1700] = 0
      "0000000" when "00000011010100101", -- t[1701] = 0
      "0000000" when "00000011010100110", -- t[1702] = 0
      "0000000" when "00000011010100111", -- t[1703] = 0
      "0000000" when "00000011010101000", -- t[1704] = 0
      "0000000" when "00000011010101001", -- t[1705] = 0
      "0000000" when "00000011010101010", -- t[1706] = 0
      "0000000" when "00000011010101011", -- t[1707] = 0
      "0000000" when "00000011010101100", -- t[1708] = 0
      "0000000" when "00000011010101101", -- t[1709] = 0
      "0000000" when "00000011010101110", -- t[1710] = 0
      "0000000" when "00000011010101111", -- t[1711] = 0
      "0000000" when "00000011010110000", -- t[1712] = 0
      "0000000" when "00000011010110001", -- t[1713] = 0
      "0000000" when "00000011010110010", -- t[1714] = 0
      "0000000" when "00000011010110011", -- t[1715] = 0
      "0000000" when "00000011010110100", -- t[1716] = 0
      "0000000" when "00000011010110101", -- t[1717] = 0
      "0000000" when "00000011010110110", -- t[1718] = 0
      "0000000" when "00000011010110111", -- t[1719] = 0
      "0000000" when "00000011010111000", -- t[1720] = 0
      "0000000" when "00000011010111001", -- t[1721] = 0
      "0000000" when "00000011010111010", -- t[1722] = 0
      "0000000" when "00000011010111011", -- t[1723] = 0
      "0000000" when "00000011010111100", -- t[1724] = 0
      "0000000" when "00000011010111101", -- t[1725] = 0
      "0000000" when "00000011010111110", -- t[1726] = 0
      "0000000" when "00000011010111111", -- t[1727] = 0
      "0000000" when "00000011011000000", -- t[1728] = 0
      "0000000" when "00000011011000001", -- t[1729] = 0
      "0000000" when "00000011011000010", -- t[1730] = 0
      "0000000" when "00000011011000011", -- t[1731] = 0
      "0000000" when "00000011011000100", -- t[1732] = 0
      "0000000" when "00000011011000101", -- t[1733] = 0
      "0000000" when "00000011011000110", -- t[1734] = 0
      "0000000" when "00000011011000111", -- t[1735] = 0
      "0000000" when "00000011011001000", -- t[1736] = 0
      "0000000" when "00000011011001001", -- t[1737] = 0
      "0000000" when "00000011011001010", -- t[1738] = 0
      "0000000" when "00000011011001011", -- t[1739] = 0
      "0000000" when "00000011011001100", -- t[1740] = 0
      "0000000" when "00000011011001101", -- t[1741] = 0
      "0000000" when "00000011011001110", -- t[1742] = 0
      "0000000" when "00000011011001111", -- t[1743] = 0
      "0000000" when "00000011011010000", -- t[1744] = 0
      "0000000" when "00000011011010001", -- t[1745] = 0
      "0000000" when "00000011011010010", -- t[1746] = 0
      "0000000" when "00000011011010011", -- t[1747] = 0
      "0000000" when "00000011011010100", -- t[1748] = 0
      "0000000" when "00000011011010101", -- t[1749] = 0
      "0000000" when "00000011011010110", -- t[1750] = 0
      "0000000" when "00000011011010111", -- t[1751] = 0
      "0000000" when "00000011011011000", -- t[1752] = 0
      "0000000" when "00000011011011001", -- t[1753] = 0
      "0000000" when "00000011011011010", -- t[1754] = 0
      "0000000" when "00000011011011011", -- t[1755] = 0
      "0000000" when "00000011011011100", -- t[1756] = 0
      "0000000" when "00000011011011101", -- t[1757] = 0
      "0000000" when "00000011011011110", -- t[1758] = 0
      "0000000" when "00000011011011111", -- t[1759] = 0
      "0000000" when "00000011011100000", -- t[1760] = 0
      "0000000" when "00000011011100001", -- t[1761] = 0
      "0000000" when "00000011011100010", -- t[1762] = 0
      "0000000" when "00000011011100011", -- t[1763] = 0
      "0000000" when "00000011011100100", -- t[1764] = 0
      "0000000" when "00000011011100101", -- t[1765] = 0
      "0000000" when "00000011011100110", -- t[1766] = 0
      "0000000" when "00000011011100111", -- t[1767] = 0
      "0000000" when "00000011011101000", -- t[1768] = 0
      "0000000" when "00000011011101001", -- t[1769] = 0
      "0000000" when "00000011011101010", -- t[1770] = 0
      "0000000" when "00000011011101011", -- t[1771] = 0
      "0000000" when "00000011011101100", -- t[1772] = 0
      "0000000" when "00000011011101101", -- t[1773] = 0
      "0000000" when "00000011011101110", -- t[1774] = 0
      "0000000" when "00000011011101111", -- t[1775] = 0
      "0000000" when "00000011011110000", -- t[1776] = 0
      "0000000" when "00000011011110001", -- t[1777] = 0
      "0000000" when "00000011011110010", -- t[1778] = 0
      "0000000" when "00000011011110011", -- t[1779] = 0
      "0000000" when "00000011011110100", -- t[1780] = 0
      "0000000" when "00000011011110101", -- t[1781] = 0
      "0000000" when "00000011011110110", -- t[1782] = 0
      "0000000" when "00000011011110111", -- t[1783] = 0
      "0000000" when "00000011011111000", -- t[1784] = 0
      "0000000" when "00000011011111001", -- t[1785] = 0
      "0000000" when "00000011011111010", -- t[1786] = 0
      "0000000" when "00000011011111011", -- t[1787] = 0
      "0000000" when "00000011011111100", -- t[1788] = 0
      "0000000" when "00000011011111101", -- t[1789] = 0
      "0000000" when "00000011011111110", -- t[1790] = 0
      "0000000" when "00000011011111111", -- t[1791] = 0
      "0000000" when "00000011100000000", -- t[1792] = 0
      "0000000" when "00000011100000001", -- t[1793] = 0
      "0000000" when "00000011100000010", -- t[1794] = 0
      "0000000" when "00000011100000011", -- t[1795] = 0
      "0000000" when "00000011100000100", -- t[1796] = 0
      "0000000" when "00000011100000101", -- t[1797] = 0
      "0000000" when "00000011100000110", -- t[1798] = 0
      "0000000" when "00000011100000111", -- t[1799] = 0
      "0000000" when "00000011100001000", -- t[1800] = 0
      "0000000" when "00000011100001001", -- t[1801] = 0
      "0000000" when "00000011100001010", -- t[1802] = 0
      "0000000" when "00000011100001011", -- t[1803] = 0
      "0000000" when "00000011100001100", -- t[1804] = 0
      "0000000" when "00000011100001101", -- t[1805] = 0
      "0000000" when "00000011100001110", -- t[1806] = 0
      "0000000" when "00000011100001111", -- t[1807] = 0
      "0000000" when "00000011100010000", -- t[1808] = 0
      "0000000" when "00000011100010001", -- t[1809] = 0
      "0000000" when "00000011100010010", -- t[1810] = 0
      "0000000" when "00000011100010011", -- t[1811] = 0
      "0000000" when "00000011100010100", -- t[1812] = 0
      "0000000" when "00000011100010101", -- t[1813] = 0
      "0000000" when "00000011100010110", -- t[1814] = 0
      "0000000" when "00000011100010111", -- t[1815] = 0
      "0000000" when "00000011100011000", -- t[1816] = 0
      "0000000" when "00000011100011001", -- t[1817] = 0
      "0000000" when "00000011100011010", -- t[1818] = 0
      "0000000" when "00000011100011011", -- t[1819] = 0
      "0000000" when "00000011100011100", -- t[1820] = 0
      "0000000" when "00000011100011101", -- t[1821] = 0
      "0000000" when "00000011100011110", -- t[1822] = 0
      "0000000" when "00000011100011111", -- t[1823] = 0
      "0000000" when "00000011100100000", -- t[1824] = 0
      "0000000" when "00000011100100001", -- t[1825] = 0
      "0000000" when "00000011100100010", -- t[1826] = 0
      "0000000" when "00000011100100011", -- t[1827] = 0
      "0000000" when "00000011100100100", -- t[1828] = 0
      "0000000" when "00000011100100101", -- t[1829] = 0
      "0000000" when "00000011100100110", -- t[1830] = 0
      "0000000" when "00000011100100111", -- t[1831] = 0
      "0000000" when "00000011100101000", -- t[1832] = 0
      "0000000" when "00000011100101001", -- t[1833] = 0
      "0000000" when "00000011100101010", -- t[1834] = 0
      "0000000" when "00000011100101011", -- t[1835] = 0
      "0000000" when "00000011100101100", -- t[1836] = 0
      "0000000" when "00000011100101101", -- t[1837] = 0
      "0000000" when "00000011100101110", -- t[1838] = 0
      "0000000" when "00000011100101111", -- t[1839] = 0
      "0000000" when "00000011100110000", -- t[1840] = 0
      "0000000" when "00000011100110001", -- t[1841] = 0
      "0000000" when "00000011100110010", -- t[1842] = 0
      "0000000" when "00000011100110011", -- t[1843] = 0
      "0000000" when "00000011100110100", -- t[1844] = 0
      "0000000" when "00000011100110101", -- t[1845] = 0
      "0000000" when "00000011100110110", -- t[1846] = 0
      "0000000" when "00000011100110111", -- t[1847] = 0
      "0000000" when "00000011100111000", -- t[1848] = 0
      "0000000" when "00000011100111001", -- t[1849] = 0
      "0000000" when "00000011100111010", -- t[1850] = 0
      "0000000" when "00000011100111011", -- t[1851] = 0
      "0000000" when "00000011100111100", -- t[1852] = 0
      "0000000" when "00000011100111101", -- t[1853] = 0
      "0000000" when "00000011100111110", -- t[1854] = 0
      "0000000" when "00000011100111111", -- t[1855] = 0
      "0000000" when "00000011101000000", -- t[1856] = 0
      "0000000" when "00000011101000001", -- t[1857] = 0
      "0000000" when "00000011101000010", -- t[1858] = 0
      "0000000" when "00000011101000011", -- t[1859] = 0
      "0000000" when "00000011101000100", -- t[1860] = 0
      "0000000" when "00000011101000101", -- t[1861] = 0
      "0000000" when "00000011101000110", -- t[1862] = 0
      "0000000" when "00000011101000111", -- t[1863] = 0
      "0000000" when "00000011101001000", -- t[1864] = 0
      "0000000" when "00000011101001001", -- t[1865] = 0
      "0000000" when "00000011101001010", -- t[1866] = 0
      "0000000" when "00000011101001011", -- t[1867] = 0
      "0000000" when "00000011101001100", -- t[1868] = 0
      "0000000" when "00000011101001101", -- t[1869] = 0
      "0000000" when "00000011101001110", -- t[1870] = 0
      "0000000" when "00000011101001111", -- t[1871] = 0
      "0000000" when "00000011101010000", -- t[1872] = 0
      "0000000" when "00000011101010001", -- t[1873] = 0
      "0000000" when "00000011101010010", -- t[1874] = 0
      "0000000" when "00000011101010011", -- t[1875] = 0
      "0000000" when "00000011101010100", -- t[1876] = 0
      "0000000" when "00000011101010101", -- t[1877] = 0
      "0000000" when "00000011101010110", -- t[1878] = 0
      "0000000" when "00000011101010111", -- t[1879] = 0
      "0000000" when "00000011101011000", -- t[1880] = 0
      "0000000" when "00000011101011001", -- t[1881] = 0
      "0000000" when "00000011101011010", -- t[1882] = 0
      "0000000" when "00000011101011011", -- t[1883] = 0
      "0000000" when "00000011101011100", -- t[1884] = 0
      "0000000" when "00000011101011101", -- t[1885] = 0
      "0000000" when "00000011101011110", -- t[1886] = 0
      "0000000" when "00000011101011111", -- t[1887] = 0
      "0000000" when "00000011101100000", -- t[1888] = 0
      "0000000" when "00000011101100001", -- t[1889] = 0
      "0000000" when "00000011101100010", -- t[1890] = 0
      "0000000" when "00000011101100011", -- t[1891] = 0
      "0000000" when "00000011101100100", -- t[1892] = 0
      "0000000" when "00000011101100101", -- t[1893] = 0
      "0000000" when "00000011101100110", -- t[1894] = 0
      "0000000" when "00000011101100111", -- t[1895] = 0
      "0000000" when "00000011101101000", -- t[1896] = 0
      "0000000" when "00000011101101001", -- t[1897] = 0
      "0000000" when "00000011101101010", -- t[1898] = 0
      "0000000" when "00000011101101011", -- t[1899] = 0
      "0000000" when "00000011101101100", -- t[1900] = 0
      "0000000" when "00000011101101101", -- t[1901] = 0
      "0000000" when "00000011101101110", -- t[1902] = 0
      "0000000" when "00000011101101111", -- t[1903] = 0
      "0000000" when "00000011101110000", -- t[1904] = 0
      "0000000" when "00000011101110001", -- t[1905] = 0
      "0000000" when "00000011101110010", -- t[1906] = 0
      "0000000" when "00000011101110011", -- t[1907] = 0
      "0000000" when "00000011101110100", -- t[1908] = 0
      "0000000" when "00000011101110101", -- t[1909] = 0
      "0000000" when "00000011101110110", -- t[1910] = 0
      "0000000" when "00000011101110111", -- t[1911] = 0
      "0000000" when "00000011101111000", -- t[1912] = 0
      "0000000" when "00000011101111001", -- t[1913] = 0
      "0000000" when "00000011101111010", -- t[1914] = 0
      "0000000" when "00000011101111011", -- t[1915] = 0
      "0000000" when "00000011101111100", -- t[1916] = 0
      "0000000" when "00000011101111101", -- t[1917] = 0
      "0000000" when "00000011101111110", -- t[1918] = 0
      "0000000" when "00000011101111111", -- t[1919] = 0
      "0000000" when "00000011110000000", -- t[1920] = 0
      "0000000" when "00000011110000001", -- t[1921] = 0
      "0000000" when "00000011110000010", -- t[1922] = 0
      "0000000" when "00000011110000011", -- t[1923] = 0
      "0000000" when "00000011110000100", -- t[1924] = 0
      "0000000" when "00000011110000101", -- t[1925] = 0
      "0000000" when "00000011110000110", -- t[1926] = 0
      "0000000" when "00000011110000111", -- t[1927] = 0
      "0000000" when "00000011110001000", -- t[1928] = 0
      "0000000" when "00000011110001001", -- t[1929] = 0
      "0000000" when "00000011110001010", -- t[1930] = 0
      "0000000" when "00000011110001011", -- t[1931] = 0
      "0000000" when "00000011110001100", -- t[1932] = 0
      "0000000" when "00000011110001101", -- t[1933] = 0
      "0000000" when "00000011110001110", -- t[1934] = 0
      "0000000" when "00000011110001111", -- t[1935] = 0
      "0000000" when "00000011110010000", -- t[1936] = 0
      "0000000" when "00000011110010001", -- t[1937] = 0
      "0000000" when "00000011110010010", -- t[1938] = 0
      "0000000" when "00000011110010011", -- t[1939] = 0
      "0000000" when "00000011110010100", -- t[1940] = 0
      "0000000" when "00000011110010101", -- t[1941] = 0
      "0000000" when "00000011110010110", -- t[1942] = 0
      "0000000" when "00000011110010111", -- t[1943] = 0
      "0000000" when "00000011110011000", -- t[1944] = 0
      "0000000" when "00000011110011001", -- t[1945] = 0
      "0000000" when "00000011110011010", -- t[1946] = 0
      "0000000" when "00000011110011011", -- t[1947] = 0
      "0000000" when "00000011110011100", -- t[1948] = 0
      "0000000" when "00000011110011101", -- t[1949] = 0
      "0000000" when "00000011110011110", -- t[1950] = 0
      "0000000" when "00000011110011111", -- t[1951] = 0
      "0000000" when "00000011110100000", -- t[1952] = 0
      "0000000" when "00000011110100001", -- t[1953] = 0
      "0000000" when "00000011110100010", -- t[1954] = 0
      "0000000" when "00000011110100011", -- t[1955] = 0
      "0000000" when "00000011110100100", -- t[1956] = 0
      "0000000" when "00000011110100101", -- t[1957] = 0
      "0000000" when "00000011110100110", -- t[1958] = 0
      "0000000" when "00000011110100111", -- t[1959] = 0
      "0000000" when "00000011110101000", -- t[1960] = 0
      "0000000" when "00000011110101001", -- t[1961] = 0
      "0000000" when "00000011110101010", -- t[1962] = 0
      "0000000" when "00000011110101011", -- t[1963] = 0
      "0000000" when "00000011110101100", -- t[1964] = 0
      "0000000" when "00000011110101101", -- t[1965] = 0
      "0000000" when "00000011110101110", -- t[1966] = 0
      "0000000" when "00000011110101111", -- t[1967] = 0
      "0000000" when "00000011110110000", -- t[1968] = 0
      "0000000" when "00000011110110001", -- t[1969] = 0
      "0000000" when "00000011110110010", -- t[1970] = 0
      "0000000" when "00000011110110011", -- t[1971] = 0
      "0000000" when "00000011110110100", -- t[1972] = 0
      "0000000" when "00000011110110101", -- t[1973] = 0
      "0000000" when "00000011110110110", -- t[1974] = 0
      "0000000" when "00000011110110111", -- t[1975] = 0
      "0000000" when "00000011110111000", -- t[1976] = 0
      "0000000" when "00000011110111001", -- t[1977] = 0
      "0000000" when "00000011110111010", -- t[1978] = 0
      "0000000" when "00000011110111011", -- t[1979] = 0
      "0000000" when "00000011110111100", -- t[1980] = 0
      "0000000" when "00000011110111101", -- t[1981] = 0
      "0000000" when "00000011110111110", -- t[1982] = 0
      "0000000" when "00000011110111111", -- t[1983] = 0
      "0000000" when "00000011111000000", -- t[1984] = 0
      "0000000" when "00000011111000001", -- t[1985] = 0
      "0000000" when "00000011111000010", -- t[1986] = 0
      "0000000" when "00000011111000011", -- t[1987] = 0
      "0000000" when "00000011111000100", -- t[1988] = 0
      "0000000" when "00000011111000101", -- t[1989] = 0
      "0000000" when "00000011111000110", -- t[1990] = 0
      "0000000" when "00000011111000111", -- t[1991] = 0
      "0000000" when "00000011111001000", -- t[1992] = 0
      "0000000" when "00000011111001001", -- t[1993] = 0
      "0000000" when "00000011111001010", -- t[1994] = 0
      "0000000" when "00000011111001011", -- t[1995] = 0
      "0000000" when "00000011111001100", -- t[1996] = 0
      "0000000" when "00000011111001101", -- t[1997] = 0
      "0000000" when "00000011111001110", -- t[1998] = 0
      "0000000" when "00000011111001111", -- t[1999] = 0
      "0000000" when "00000011111010000", -- t[2000] = 0
      "0000000" when "00000011111010001", -- t[2001] = 0
      "0000000" when "00000011111010010", -- t[2002] = 0
      "0000000" when "00000011111010011", -- t[2003] = 0
      "0000000" when "00000011111010100", -- t[2004] = 0
      "0000000" when "00000011111010101", -- t[2005] = 0
      "0000000" when "00000011111010110", -- t[2006] = 0
      "0000000" when "00000011111010111", -- t[2007] = 0
      "0000000" when "00000011111011000", -- t[2008] = 0
      "0000000" when "00000011111011001", -- t[2009] = 0
      "0000000" when "00000011111011010", -- t[2010] = 0
      "0000000" when "00000011111011011", -- t[2011] = 0
      "0000000" when "00000011111011100", -- t[2012] = 0
      "0000000" when "00000011111011101", -- t[2013] = 0
      "0000000" when "00000011111011110", -- t[2014] = 0
      "0000000" when "00000011111011111", -- t[2015] = 0
      "0000000" when "00000011111100000", -- t[2016] = 0
      "0000000" when "00000011111100001", -- t[2017] = 0
      "0000000" when "00000011111100010", -- t[2018] = 0
      "0000000" when "00000011111100011", -- t[2019] = 0
      "0000000" when "00000011111100100", -- t[2020] = 0
      "0000000" when "00000011111100101", -- t[2021] = 0
      "0000000" when "00000011111100110", -- t[2022] = 0
      "0000000" when "00000011111100111", -- t[2023] = 0
      "0000000" when "00000011111101000", -- t[2024] = 0
      "0000000" when "00000011111101001", -- t[2025] = 0
      "0000000" when "00000011111101010", -- t[2026] = 0
      "0000000" when "00000011111101011", -- t[2027] = 0
      "0000000" when "00000011111101100", -- t[2028] = 0
      "0000000" when "00000011111101101", -- t[2029] = 0
      "0000000" when "00000011111101110", -- t[2030] = 0
      "0000000" when "00000011111101111", -- t[2031] = 0
      "0000000" when "00000011111110000", -- t[2032] = 0
      "0000000" when "00000011111110001", -- t[2033] = 0
      "0000000" when "00000011111110010", -- t[2034] = 0
      "0000000" when "00000011111110011", -- t[2035] = 0
      "0000000" when "00000011111110100", -- t[2036] = 0
      "0000000" when "00000011111110101", -- t[2037] = 0
      "0000000" when "00000011111110110", -- t[2038] = 0
      "0000000" when "00000011111110111", -- t[2039] = 0
      "0000000" when "00000011111111000", -- t[2040] = 0
      "0000000" when "00000011111111001", -- t[2041] = 0
      "0000000" when "00000011111111010", -- t[2042] = 0
      "0000000" when "00000011111111011", -- t[2043] = 0
      "0000000" when "00000011111111100", -- t[2044] = 0
      "0000000" when "00000011111111101", -- t[2045] = 0
      "0000000" when "00000011111111110", -- t[2046] = 0
      "0000000" when "00000011111111111", -- t[2047] = 0
      "0000000" when "00000100000000000", -- t[2048] = 0
      "0000000" when "00000100000000001", -- t[2049] = 0
      "0000000" when "00000100000000010", -- t[2050] = 0
      "0000000" when "00000100000000011", -- t[2051] = 0
      "0000000" when "00000100000000100", -- t[2052] = 0
      "0000000" when "00000100000000101", -- t[2053] = 0
      "0000000" when "00000100000000110", -- t[2054] = 0
      "0000000" when "00000100000000111", -- t[2055] = 0
      "0000000" when "00000100000001000", -- t[2056] = 0
      "0000000" when "00000100000001001", -- t[2057] = 0
      "0000000" when "00000100000001010", -- t[2058] = 0
      "0000000" when "00000100000001011", -- t[2059] = 0
      "0000000" when "00000100000001100", -- t[2060] = 0
      "0000000" when "00000100000001101", -- t[2061] = 0
      "0000000" when "00000100000001110", -- t[2062] = 0
      "0000000" when "00000100000001111", -- t[2063] = 0
      "0000000" when "00000100000010000", -- t[2064] = 0
      "0000000" when "00000100000010001", -- t[2065] = 0
      "0000000" when "00000100000010010", -- t[2066] = 0
      "0000000" when "00000100000010011", -- t[2067] = 0
      "0000000" when "00000100000010100", -- t[2068] = 0
      "0000000" when "00000100000010101", -- t[2069] = 0
      "0000000" when "00000100000010110", -- t[2070] = 0
      "0000000" when "00000100000010111", -- t[2071] = 0
      "0000000" when "00000100000011000", -- t[2072] = 0
      "0000000" when "00000100000011001", -- t[2073] = 0
      "0000000" when "00000100000011010", -- t[2074] = 0
      "0000000" when "00000100000011011", -- t[2075] = 0
      "0000000" when "00000100000011100", -- t[2076] = 0
      "0000000" when "00000100000011101", -- t[2077] = 0
      "0000000" when "00000100000011110", -- t[2078] = 0
      "0000000" when "00000100000011111", -- t[2079] = 0
      "0000000" when "00000100000100000", -- t[2080] = 0
      "0000000" when "00000100000100001", -- t[2081] = 0
      "0000000" when "00000100000100010", -- t[2082] = 0
      "0000000" when "00000100000100011", -- t[2083] = 0
      "0000000" when "00000100000100100", -- t[2084] = 0
      "0000000" when "00000100000100101", -- t[2085] = 0
      "0000000" when "00000100000100110", -- t[2086] = 0
      "0000000" when "00000100000100111", -- t[2087] = 0
      "0000000" when "00000100000101000", -- t[2088] = 0
      "0000000" when "00000100000101001", -- t[2089] = 0
      "0000000" when "00000100000101010", -- t[2090] = 0
      "0000000" when "00000100000101011", -- t[2091] = 0
      "0000000" when "00000100000101100", -- t[2092] = 0
      "0000000" when "00000100000101101", -- t[2093] = 0
      "0000000" when "00000100000101110", -- t[2094] = 0
      "0000000" when "00000100000101111", -- t[2095] = 0
      "0000000" when "00000100000110000", -- t[2096] = 0
      "0000000" when "00000100000110001", -- t[2097] = 0
      "0000000" when "00000100000110010", -- t[2098] = 0
      "0000000" when "00000100000110011", -- t[2099] = 0
      "0000000" when "00000100000110100", -- t[2100] = 0
      "0000000" when "00000100000110101", -- t[2101] = 0
      "0000000" when "00000100000110110", -- t[2102] = 0
      "0000000" when "00000100000110111", -- t[2103] = 0
      "0000000" when "00000100000111000", -- t[2104] = 0
      "0000000" when "00000100000111001", -- t[2105] = 0
      "0000000" when "00000100000111010", -- t[2106] = 0
      "0000000" when "00000100000111011", -- t[2107] = 0
      "0000000" when "00000100000111100", -- t[2108] = 0
      "0000000" when "00000100000111101", -- t[2109] = 0
      "0000000" when "00000100000111110", -- t[2110] = 0
      "0000000" when "00000100000111111", -- t[2111] = 0
      "0000000" when "00000100001000000", -- t[2112] = 0
      "0000000" when "00000100001000001", -- t[2113] = 0
      "0000000" when "00000100001000010", -- t[2114] = 0
      "0000000" when "00000100001000011", -- t[2115] = 0
      "0000000" when "00000100001000100", -- t[2116] = 0
      "0000000" when "00000100001000101", -- t[2117] = 0
      "0000000" when "00000100001000110", -- t[2118] = 0
      "0000000" when "00000100001000111", -- t[2119] = 0
      "0000000" when "00000100001001000", -- t[2120] = 0
      "0000000" when "00000100001001001", -- t[2121] = 0
      "0000000" when "00000100001001010", -- t[2122] = 0
      "0000000" when "00000100001001011", -- t[2123] = 0
      "0000000" when "00000100001001100", -- t[2124] = 0
      "0000000" when "00000100001001101", -- t[2125] = 0
      "0000000" when "00000100001001110", -- t[2126] = 0
      "0000000" when "00000100001001111", -- t[2127] = 0
      "0000000" when "00000100001010000", -- t[2128] = 0
      "0000000" when "00000100001010001", -- t[2129] = 0
      "0000000" when "00000100001010010", -- t[2130] = 0
      "0000000" when "00000100001010011", -- t[2131] = 0
      "0000000" when "00000100001010100", -- t[2132] = 0
      "0000000" when "00000100001010101", -- t[2133] = 0
      "0000000" when "00000100001010110", -- t[2134] = 0
      "0000000" when "00000100001010111", -- t[2135] = 0
      "0000000" when "00000100001011000", -- t[2136] = 0
      "0000000" when "00000100001011001", -- t[2137] = 0
      "0000000" when "00000100001011010", -- t[2138] = 0
      "0000000" when "00000100001011011", -- t[2139] = 0
      "0000000" when "00000100001011100", -- t[2140] = 0
      "0000000" when "00000100001011101", -- t[2141] = 0
      "0000000" when "00000100001011110", -- t[2142] = 0
      "0000000" when "00000100001011111", -- t[2143] = 0
      "0000000" when "00000100001100000", -- t[2144] = 0
      "0000000" when "00000100001100001", -- t[2145] = 0
      "0000000" when "00000100001100010", -- t[2146] = 0
      "0000000" when "00000100001100011", -- t[2147] = 0
      "0000000" when "00000100001100100", -- t[2148] = 0
      "0000000" when "00000100001100101", -- t[2149] = 0
      "0000000" when "00000100001100110", -- t[2150] = 0
      "0000000" when "00000100001100111", -- t[2151] = 0
      "0000000" when "00000100001101000", -- t[2152] = 0
      "0000000" when "00000100001101001", -- t[2153] = 0
      "0000000" when "00000100001101010", -- t[2154] = 0
      "0000000" when "00000100001101011", -- t[2155] = 0
      "0000000" when "00000100001101100", -- t[2156] = 0
      "0000000" when "00000100001101101", -- t[2157] = 0
      "0000000" when "00000100001101110", -- t[2158] = 0
      "0000000" when "00000100001101111", -- t[2159] = 0
      "0000000" when "00000100001110000", -- t[2160] = 0
      "0000000" when "00000100001110001", -- t[2161] = 0
      "0000000" when "00000100001110010", -- t[2162] = 0
      "0000000" when "00000100001110011", -- t[2163] = 0
      "0000000" when "00000100001110100", -- t[2164] = 0
      "0000000" when "00000100001110101", -- t[2165] = 0
      "0000000" when "00000100001110110", -- t[2166] = 0
      "0000000" when "00000100001110111", -- t[2167] = 0
      "0000000" when "00000100001111000", -- t[2168] = 0
      "0000000" when "00000100001111001", -- t[2169] = 0
      "0000000" when "00000100001111010", -- t[2170] = 0
      "0000000" when "00000100001111011", -- t[2171] = 0
      "0000000" when "00000100001111100", -- t[2172] = 0
      "0000000" when "00000100001111101", -- t[2173] = 0
      "0000000" when "00000100001111110", -- t[2174] = 0
      "0000000" when "00000100001111111", -- t[2175] = 0
      "0000000" when "00000100010000000", -- t[2176] = 0
      "0000000" when "00000100010000001", -- t[2177] = 0
      "0000000" when "00000100010000010", -- t[2178] = 0
      "0000000" when "00000100010000011", -- t[2179] = 0
      "0000000" when "00000100010000100", -- t[2180] = 0
      "0000000" when "00000100010000101", -- t[2181] = 0
      "0000000" when "00000100010000110", -- t[2182] = 0
      "0000000" when "00000100010000111", -- t[2183] = 0
      "0000000" when "00000100010001000", -- t[2184] = 0
      "0000000" when "00000100010001001", -- t[2185] = 0
      "0000000" when "00000100010001010", -- t[2186] = 0
      "0000000" when "00000100010001011", -- t[2187] = 0
      "0000000" when "00000100010001100", -- t[2188] = 0
      "0000000" when "00000100010001101", -- t[2189] = 0
      "0000000" when "00000100010001110", -- t[2190] = 0
      "0000000" when "00000100010001111", -- t[2191] = 0
      "0000000" when "00000100010010000", -- t[2192] = 0
      "0000000" when "00000100010010001", -- t[2193] = 0
      "0000000" when "00000100010010010", -- t[2194] = 0
      "0000000" when "00000100010010011", -- t[2195] = 0
      "0000000" when "00000100010010100", -- t[2196] = 0
      "0000000" when "00000100010010101", -- t[2197] = 0
      "0000000" when "00000100010010110", -- t[2198] = 0
      "0000000" when "00000100010010111", -- t[2199] = 0
      "0000000" when "00000100010011000", -- t[2200] = 0
      "0000000" when "00000100010011001", -- t[2201] = 0
      "0000000" when "00000100010011010", -- t[2202] = 0
      "0000000" when "00000100010011011", -- t[2203] = 0
      "0000000" when "00000100010011100", -- t[2204] = 0
      "0000000" when "00000100010011101", -- t[2205] = 0
      "0000000" when "00000100010011110", -- t[2206] = 0
      "0000000" when "00000100010011111", -- t[2207] = 0
      "0000000" when "00000100010100000", -- t[2208] = 0
      "0000000" when "00000100010100001", -- t[2209] = 0
      "0000000" when "00000100010100010", -- t[2210] = 0
      "0000000" when "00000100010100011", -- t[2211] = 0
      "0000000" when "00000100010100100", -- t[2212] = 0
      "0000000" when "00000100010100101", -- t[2213] = 0
      "0000000" when "00000100010100110", -- t[2214] = 0
      "0000000" when "00000100010100111", -- t[2215] = 0
      "0000000" when "00000100010101000", -- t[2216] = 0
      "0000000" when "00000100010101001", -- t[2217] = 0
      "0000000" when "00000100010101010", -- t[2218] = 0
      "0000000" when "00000100010101011", -- t[2219] = 0
      "0000000" when "00000100010101100", -- t[2220] = 0
      "0000000" when "00000100010101101", -- t[2221] = 0
      "0000000" when "00000100010101110", -- t[2222] = 0
      "0000000" when "00000100010101111", -- t[2223] = 0
      "0000000" when "00000100010110000", -- t[2224] = 0
      "0000000" when "00000100010110001", -- t[2225] = 0
      "0000000" when "00000100010110010", -- t[2226] = 0
      "0000000" when "00000100010110011", -- t[2227] = 0
      "0000000" when "00000100010110100", -- t[2228] = 0
      "0000000" when "00000100010110101", -- t[2229] = 0
      "0000000" when "00000100010110110", -- t[2230] = 0
      "0000000" when "00000100010110111", -- t[2231] = 0
      "0000000" when "00000100010111000", -- t[2232] = 0
      "0000000" when "00000100010111001", -- t[2233] = 0
      "0000000" when "00000100010111010", -- t[2234] = 0
      "0000000" when "00000100010111011", -- t[2235] = 0
      "0000000" when "00000100010111100", -- t[2236] = 0
      "0000000" when "00000100010111101", -- t[2237] = 0
      "0000000" when "00000100010111110", -- t[2238] = 0
      "0000000" when "00000100010111111", -- t[2239] = 0
      "0000000" when "00000100011000000", -- t[2240] = 0
      "0000000" when "00000100011000001", -- t[2241] = 0
      "0000000" when "00000100011000010", -- t[2242] = 0
      "0000000" when "00000100011000011", -- t[2243] = 0
      "0000000" when "00000100011000100", -- t[2244] = 0
      "0000000" when "00000100011000101", -- t[2245] = 0
      "0000000" when "00000100011000110", -- t[2246] = 0
      "0000000" when "00000100011000111", -- t[2247] = 0
      "0000000" when "00000100011001000", -- t[2248] = 0
      "0000000" when "00000100011001001", -- t[2249] = 0
      "0000000" when "00000100011001010", -- t[2250] = 0
      "0000000" when "00000100011001011", -- t[2251] = 0
      "0000000" when "00000100011001100", -- t[2252] = 0
      "0000000" when "00000100011001101", -- t[2253] = 0
      "0000000" when "00000100011001110", -- t[2254] = 0
      "0000000" when "00000100011001111", -- t[2255] = 0
      "0000000" when "00000100011010000", -- t[2256] = 0
      "0000000" when "00000100011010001", -- t[2257] = 0
      "0000000" when "00000100011010010", -- t[2258] = 0
      "0000000" when "00000100011010011", -- t[2259] = 0
      "0000000" when "00000100011010100", -- t[2260] = 0
      "0000000" when "00000100011010101", -- t[2261] = 0
      "0000000" when "00000100011010110", -- t[2262] = 0
      "0000000" when "00000100011010111", -- t[2263] = 0
      "0000000" when "00000100011011000", -- t[2264] = 0
      "0000000" when "00000100011011001", -- t[2265] = 0
      "0000000" when "00000100011011010", -- t[2266] = 0
      "0000000" when "00000100011011011", -- t[2267] = 0
      "0000000" when "00000100011011100", -- t[2268] = 0
      "0000000" when "00000100011011101", -- t[2269] = 0
      "0000000" when "00000100011011110", -- t[2270] = 0
      "0000000" when "00000100011011111", -- t[2271] = 0
      "0000000" when "00000100011100000", -- t[2272] = 0
      "0000000" when "00000100011100001", -- t[2273] = 0
      "0000000" when "00000100011100010", -- t[2274] = 0
      "0000000" when "00000100011100011", -- t[2275] = 0
      "0000000" when "00000100011100100", -- t[2276] = 0
      "0000000" when "00000100011100101", -- t[2277] = 0
      "0000000" when "00000100011100110", -- t[2278] = 0
      "0000000" when "00000100011100111", -- t[2279] = 0
      "0000000" when "00000100011101000", -- t[2280] = 0
      "0000000" when "00000100011101001", -- t[2281] = 0
      "0000000" when "00000100011101010", -- t[2282] = 0
      "0000000" when "00000100011101011", -- t[2283] = 0
      "0000000" when "00000100011101100", -- t[2284] = 0
      "0000000" when "00000100011101101", -- t[2285] = 0
      "0000000" when "00000100011101110", -- t[2286] = 0
      "0000000" when "00000100011101111", -- t[2287] = 0
      "0000000" when "00000100011110000", -- t[2288] = 0
      "0000000" when "00000100011110001", -- t[2289] = 0
      "0000000" when "00000100011110010", -- t[2290] = 0
      "0000000" when "00000100011110011", -- t[2291] = 0
      "0000000" when "00000100011110100", -- t[2292] = 0
      "0000000" when "00000100011110101", -- t[2293] = 0
      "0000000" when "00000100011110110", -- t[2294] = 0
      "0000000" when "00000100011110111", -- t[2295] = 0
      "0000000" when "00000100011111000", -- t[2296] = 0
      "0000000" when "00000100011111001", -- t[2297] = 0
      "0000000" when "00000100011111010", -- t[2298] = 0
      "0000000" when "00000100011111011", -- t[2299] = 0
      "0000000" when "00000100011111100", -- t[2300] = 0
      "0000000" when "00000100011111101", -- t[2301] = 0
      "0000000" when "00000100011111110", -- t[2302] = 0
      "0000000" when "00000100011111111", -- t[2303] = 0
      "0000000" when "00000100100000000", -- t[2304] = 0
      "0000000" when "00000100100000001", -- t[2305] = 0
      "0000000" when "00000100100000010", -- t[2306] = 0
      "0000000" when "00000100100000011", -- t[2307] = 0
      "0000000" when "00000100100000100", -- t[2308] = 0
      "0000000" when "00000100100000101", -- t[2309] = 0
      "0000000" when "00000100100000110", -- t[2310] = 0
      "0000000" when "00000100100000111", -- t[2311] = 0
      "0000000" when "00000100100001000", -- t[2312] = 0
      "0000000" when "00000100100001001", -- t[2313] = 0
      "0000000" when "00000100100001010", -- t[2314] = 0
      "0000000" when "00000100100001011", -- t[2315] = 0
      "0000000" when "00000100100001100", -- t[2316] = 0
      "0000000" when "00000100100001101", -- t[2317] = 0
      "0000000" when "00000100100001110", -- t[2318] = 0
      "0000000" when "00000100100001111", -- t[2319] = 0
      "0000000" when "00000100100010000", -- t[2320] = 0
      "0000000" when "00000100100010001", -- t[2321] = 0
      "0000000" when "00000100100010010", -- t[2322] = 0
      "0000000" when "00000100100010011", -- t[2323] = 0
      "0000000" when "00000100100010100", -- t[2324] = 0
      "0000000" when "00000100100010101", -- t[2325] = 0
      "0000000" when "00000100100010110", -- t[2326] = 0
      "0000000" when "00000100100010111", -- t[2327] = 0
      "0000000" when "00000100100011000", -- t[2328] = 0
      "0000000" when "00000100100011001", -- t[2329] = 0
      "0000000" when "00000100100011010", -- t[2330] = 0
      "0000000" when "00000100100011011", -- t[2331] = 0
      "0000000" when "00000100100011100", -- t[2332] = 0
      "0000000" when "00000100100011101", -- t[2333] = 0
      "0000000" when "00000100100011110", -- t[2334] = 0
      "0000000" when "00000100100011111", -- t[2335] = 0
      "0000000" when "00000100100100000", -- t[2336] = 0
      "0000000" when "00000100100100001", -- t[2337] = 0
      "0000000" when "00000100100100010", -- t[2338] = 0
      "0000000" when "00000100100100011", -- t[2339] = 0
      "0000000" when "00000100100100100", -- t[2340] = 0
      "0000000" when "00000100100100101", -- t[2341] = 0
      "0000000" when "00000100100100110", -- t[2342] = 0
      "0000000" when "00000100100100111", -- t[2343] = 0
      "0000000" when "00000100100101000", -- t[2344] = 0
      "0000000" when "00000100100101001", -- t[2345] = 0
      "0000000" when "00000100100101010", -- t[2346] = 0
      "0000000" when "00000100100101011", -- t[2347] = 0
      "0000000" when "00000100100101100", -- t[2348] = 0
      "0000000" when "00000100100101101", -- t[2349] = 0
      "0000000" when "00000100100101110", -- t[2350] = 0
      "0000000" when "00000100100101111", -- t[2351] = 0
      "0000000" when "00000100100110000", -- t[2352] = 0
      "0000000" when "00000100100110001", -- t[2353] = 0
      "0000000" when "00000100100110010", -- t[2354] = 0
      "0000000" when "00000100100110011", -- t[2355] = 0
      "0000000" when "00000100100110100", -- t[2356] = 0
      "0000000" when "00000100100110101", -- t[2357] = 0
      "0000000" when "00000100100110110", -- t[2358] = 0
      "0000000" when "00000100100110111", -- t[2359] = 0
      "0000000" when "00000100100111000", -- t[2360] = 0
      "0000000" when "00000100100111001", -- t[2361] = 0
      "0000000" when "00000100100111010", -- t[2362] = 0
      "0000000" when "00000100100111011", -- t[2363] = 0
      "0000000" when "00000100100111100", -- t[2364] = 0
      "0000000" when "00000100100111101", -- t[2365] = 0
      "0000000" when "00000100100111110", -- t[2366] = 0
      "0000000" when "00000100100111111", -- t[2367] = 0
      "0000000" when "00000100101000000", -- t[2368] = 0
      "0000000" when "00000100101000001", -- t[2369] = 0
      "0000000" when "00000100101000010", -- t[2370] = 0
      "0000000" when "00000100101000011", -- t[2371] = 0
      "0000000" when "00000100101000100", -- t[2372] = 0
      "0000000" when "00000100101000101", -- t[2373] = 0
      "0000000" when "00000100101000110", -- t[2374] = 0
      "0000000" when "00000100101000111", -- t[2375] = 0
      "0000000" when "00000100101001000", -- t[2376] = 0
      "0000000" when "00000100101001001", -- t[2377] = 0
      "0000000" when "00000100101001010", -- t[2378] = 0
      "0000000" when "00000100101001011", -- t[2379] = 0
      "0000000" when "00000100101001100", -- t[2380] = 0
      "0000000" when "00000100101001101", -- t[2381] = 0
      "0000000" when "00000100101001110", -- t[2382] = 0
      "0000000" when "00000100101001111", -- t[2383] = 0
      "0000000" when "00000100101010000", -- t[2384] = 0
      "0000000" when "00000100101010001", -- t[2385] = 0
      "0000000" when "00000100101010010", -- t[2386] = 0
      "0000000" when "00000100101010011", -- t[2387] = 0
      "0000000" when "00000100101010100", -- t[2388] = 0
      "0000000" when "00000100101010101", -- t[2389] = 0
      "0000000" when "00000100101010110", -- t[2390] = 0
      "0000000" when "00000100101010111", -- t[2391] = 0
      "0000000" when "00000100101011000", -- t[2392] = 0
      "0000000" when "00000100101011001", -- t[2393] = 0
      "0000000" when "00000100101011010", -- t[2394] = 0
      "0000000" when "00000100101011011", -- t[2395] = 0
      "0000000" when "00000100101011100", -- t[2396] = 0
      "0000000" when "00000100101011101", -- t[2397] = 0
      "0000000" when "00000100101011110", -- t[2398] = 0
      "0000000" when "00000100101011111", -- t[2399] = 0
      "0000000" when "00000100101100000", -- t[2400] = 0
      "0000000" when "00000100101100001", -- t[2401] = 0
      "0000000" when "00000100101100010", -- t[2402] = 0
      "0000000" when "00000100101100011", -- t[2403] = 0
      "0000000" when "00000100101100100", -- t[2404] = 0
      "0000000" when "00000100101100101", -- t[2405] = 0
      "0000000" when "00000100101100110", -- t[2406] = 0
      "0000000" when "00000100101100111", -- t[2407] = 0
      "0000000" when "00000100101101000", -- t[2408] = 0
      "0000000" when "00000100101101001", -- t[2409] = 0
      "0000000" when "00000100101101010", -- t[2410] = 0
      "0000000" when "00000100101101011", -- t[2411] = 0
      "0000000" when "00000100101101100", -- t[2412] = 0
      "0000000" when "00000100101101101", -- t[2413] = 0
      "0000000" when "00000100101101110", -- t[2414] = 0
      "0000000" when "00000100101101111", -- t[2415] = 0
      "0000000" when "00000100101110000", -- t[2416] = 0
      "0000000" when "00000100101110001", -- t[2417] = 0
      "0000000" when "00000100101110010", -- t[2418] = 0
      "0000000" when "00000100101110011", -- t[2419] = 0
      "0000000" when "00000100101110100", -- t[2420] = 0
      "0000000" when "00000100101110101", -- t[2421] = 0
      "0000000" when "00000100101110110", -- t[2422] = 0
      "0000000" when "00000100101110111", -- t[2423] = 0
      "0000000" when "00000100101111000", -- t[2424] = 0
      "0000000" when "00000100101111001", -- t[2425] = 0
      "0000000" when "00000100101111010", -- t[2426] = 0
      "0000000" when "00000100101111011", -- t[2427] = 0
      "0000000" when "00000100101111100", -- t[2428] = 0
      "0000000" when "00000100101111101", -- t[2429] = 0
      "0000000" when "00000100101111110", -- t[2430] = 0
      "0000000" when "00000100101111111", -- t[2431] = 0
      "0000000" when "00000100110000000", -- t[2432] = 0
      "0000000" when "00000100110000001", -- t[2433] = 0
      "0000000" when "00000100110000010", -- t[2434] = 0
      "0000000" when "00000100110000011", -- t[2435] = 0
      "0000000" when "00000100110000100", -- t[2436] = 0
      "0000000" when "00000100110000101", -- t[2437] = 0
      "0000000" when "00000100110000110", -- t[2438] = 0
      "0000000" when "00000100110000111", -- t[2439] = 0
      "0000000" when "00000100110001000", -- t[2440] = 0
      "0000000" when "00000100110001001", -- t[2441] = 0
      "0000000" when "00000100110001010", -- t[2442] = 0
      "0000000" when "00000100110001011", -- t[2443] = 0
      "0000000" when "00000100110001100", -- t[2444] = 0
      "0000000" when "00000100110001101", -- t[2445] = 0
      "0000000" when "00000100110001110", -- t[2446] = 0
      "0000000" when "00000100110001111", -- t[2447] = 0
      "0000000" when "00000100110010000", -- t[2448] = 0
      "0000000" when "00000100110010001", -- t[2449] = 0
      "0000000" when "00000100110010010", -- t[2450] = 0
      "0000000" when "00000100110010011", -- t[2451] = 0
      "0000000" when "00000100110010100", -- t[2452] = 0
      "0000000" when "00000100110010101", -- t[2453] = 0
      "0000000" when "00000100110010110", -- t[2454] = 0
      "0000000" when "00000100110010111", -- t[2455] = 0
      "0000000" when "00000100110011000", -- t[2456] = 0
      "0000000" when "00000100110011001", -- t[2457] = 0
      "0000000" when "00000100110011010", -- t[2458] = 0
      "0000000" when "00000100110011011", -- t[2459] = 0
      "0000000" when "00000100110011100", -- t[2460] = 0
      "0000000" when "00000100110011101", -- t[2461] = 0
      "0000000" when "00000100110011110", -- t[2462] = 0
      "0000000" when "00000100110011111", -- t[2463] = 0
      "0000000" when "00000100110100000", -- t[2464] = 0
      "0000000" when "00000100110100001", -- t[2465] = 0
      "0000000" when "00000100110100010", -- t[2466] = 0
      "0000000" when "00000100110100011", -- t[2467] = 0
      "0000000" when "00000100110100100", -- t[2468] = 0
      "0000000" when "00000100110100101", -- t[2469] = 0
      "0000000" when "00000100110100110", -- t[2470] = 0
      "0000000" when "00000100110100111", -- t[2471] = 0
      "0000000" when "00000100110101000", -- t[2472] = 0
      "0000000" when "00000100110101001", -- t[2473] = 0
      "0000000" when "00000100110101010", -- t[2474] = 0
      "0000000" when "00000100110101011", -- t[2475] = 0
      "0000000" when "00000100110101100", -- t[2476] = 0
      "0000000" when "00000100110101101", -- t[2477] = 0
      "0000000" when "00000100110101110", -- t[2478] = 0
      "0000000" when "00000100110101111", -- t[2479] = 0
      "0000000" when "00000100110110000", -- t[2480] = 0
      "0000000" when "00000100110110001", -- t[2481] = 0
      "0000000" when "00000100110110010", -- t[2482] = 0
      "0000000" when "00000100110110011", -- t[2483] = 0
      "0000000" when "00000100110110100", -- t[2484] = 0
      "0000000" when "00000100110110101", -- t[2485] = 0
      "0000000" when "00000100110110110", -- t[2486] = 0
      "0000000" when "00000100110110111", -- t[2487] = 0
      "0000000" when "00000100110111000", -- t[2488] = 0
      "0000000" when "00000100110111001", -- t[2489] = 0
      "0000000" when "00000100110111010", -- t[2490] = 0
      "0000000" when "00000100110111011", -- t[2491] = 0
      "0000000" when "00000100110111100", -- t[2492] = 0
      "0000000" when "00000100110111101", -- t[2493] = 0
      "0000000" when "00000100110111110", -- t[2494] = 0
      "0000000" when "00000100110111111", -- t[2495] = 0
      "0000000" when "00000100111000000", -- t[2496] = 0
      "0000000" when "00000100111000001", -- t[2497] = 0
      "0000000" when "00000100111000010", -- t[2498] = 0
      "0000000" when "00000100111000011", -- t[2499] = 0
      "0000000" when "00000100111000100", -- t[2500] = 0
      "0000000" when "00000100111000101", -- t[2501] = 0
      "0000000" when "00000100111000110", -- t[2502] = 0
      "0000000" when "00000100111000111", -- t[2503] = 0
      "0000000" when "00000100111001000", -- t[2504] = 0
      "0000000" when "00000100111001001", -- t[2505] = 0
      "0000000" when "00000100111001010", -- t[2506] = 0
      "0000000" when "00000100111001011", -- t[2507] = 0
      "0000000" when "00000100111001100", -- t[2508] = 0
      "0000000" when "00000100111001101", -- t[2509] = 0
      "0000000" when "00000100111001110", -- t[2510] = 0
      "0000000" when "00000100111001111", -- t[2511] = 0
      "0000000" when "00000100111010000", -- t[2512] = 0
      "0000000" when "00000100111010001", -- t[2513] = 0
      "0000000" when "00000100111010010", -- t[2514] = 0
      "0000000" when "00000100111010011", -- t[2515] = 0
      "0000000" when "00000100111010100", -- t[2516] = 0
      "0000000" when "00000100111010101", -- t[2517] = 0
      "0000000" when "00000100111010110", -- t[2518] = 0
      "0000000" when "00000100111010111", -- t[2519] = 0
      "0000000" when "00000100111011000", -- t[2520] = 0
      "0000000" when "00000100111011001", -- t[2521] = 0
      "0000000" when "00000100111011010", -- t[2522] = 0
      "0000000" when "00000100111011011", -- t[2523] = 0
      "0000000" when "00000100111011100", -- t[2524] = 0
      "0000000" when "00000100111011101", -- t[2525] = 0
      "0000000" when "00000100111011110", -- t[2526] = 0
      "0000000" when "00000100111011111", -- t[2527] = 0
      "0000000" when "00000100111100000", -- t[2528] = 0
      "0000000" when "00000100111100001", -- t[2529] = 0
      "0000000" when "00000100111100010", -- t[2530] = 0
      "0000000" when "00000100111100011", -- t[2531] = 0
      "0000000" when "00000100111100100", -- t[2532] = 0
      "0000000" when "00000100111100101", -- t[2533] = 0
      "0000000" when "00000100111100110", -- t[2534] = 0
      "0000000" when "00000100111100111", -- t[2535] = 0
      "0000000" when "00000100111101000", -- t[2536] = 0
      "0000000" when "00000100111101001", -- t[2537] = 0
      "0000000" when "00000100111101010", -- t[2538] = 0
      "0000000" when "00000100111101011", -- t[2539] = 0
      "0000000" when "00000100111101100", -- t[2540] = 0
      "0000000" when "00000100111101101", -- t[2541] = 0
      "0000000" when "00000100111101110", -- t[2542] = 0
      "0000000" when "00000100111101111", -- t[2543] = 0
      "0000000" when "00000100111110000", -- t[2544] = 0
      "0000000" when "00000100111110001", -- t[2545] = 0
      "0000000" when "00000100111110010", -- t[2546] = 0
      "0000000" when "00000100111110011", -- t[2547] = 0
      "0000000" when "00000100111110100", -- t[2548] = 0
      "0000000" when "00000100111110101", -- t[2549] = 0
      "0000000" when "00000100111110110", -- t[2550] = 0
      "0000000" when "00000100111110111", -- t[2551] = 0
      "0000000" when "00000100111111000", -- t[2552] = 0
      "0000000" when "00000100111111001", -- t[2553] = 0
      "0000000" when "00000100111111010", -- t[2554] = 0
      "0000000" when "00000100111111011", -- t[2555] = 0
      "0000000" when "00000100111111100", -- t[2556] = 0
      "0000000" when "00000100111111101", -- t[2557] = 0
      "0000000" when "00000100111111110", -- t[2558] = 0
      "0000000" when "00000100111111111", -- t[2559] = 0
      "0000000" when "00000101000000000", -- t[2560] = 0
      "0000000" when "00000101000000001", -- t[2561] = 0
      "0000000" when "00000101000000010", -- t[2562] = 0
      "0000000" when "00000101000000011", -- t[2563] = 0
      "0000000" when "00000101000000100", -- t[2564] = 0
      "0000000" when "00000101000000101", -- t[2565] = 0
      "0000000" when "00000101000000110", -- t[2566] = 0
      "0000000" when "00000101000000111", -- t[2567] = 0
      "0000000" when "00000101000001000", -- t[2568] = 0
      "0000000" when "00000101000001001", -- t[2569] = 0
      "0000000" when "00000101000001010", -- t[2570] = 0
      "0000000" when "00000101000001011", -- t[2571] = 0
      "0000000" when "00000101000001100", -- t[2572] = 0
      "0000000" when "00000101000001101", -- t[2573] = 0
      "0000000" when "00000101000001110", -- t[2574] = 0
      "0000000" when "00000101000001111", -- t[2575] = 0
      "0000000" when "00000101000010000", -- t[2576] = 0
      "0000000" when "00000101000010001", -- t[2577] = 0
      "0000000" when "00000101000010010", -- t[2578] = 0
      "0000000" when "00000101000010011", -- t[2579] = 0
      "0000000" when "00000101000010100", -- t[2580] = 0
      "0000000" when "00000101000010101", -- t[2581] = 0
      "0000000" when "00000101000010110", -- t[2582] = 0
      "0000000" when "00000101000010111", -- t[2583] = 0
      "0000000" when "00000101000011000", -- t[2584] = 0
      "0000000" when "00000101000011001", -- t[2585] = 0
      "0000000" when "00000101000011010", -- t[2586] = 0
      "0000000" when "00000101000011011", -- t[2587] = 0
      "0000000" when "00000101000011100", -- t[2588] = 0
      "0000000" when "00000101000011101", -- t[2589] = 0
      "0000000" when "00000101000011110", -- t[2590] = 0
      "0000000" when "00000101000011111", -- t[2591] = 0
      "0000000" when "00000101000100000", -- t[2592] = 0
      "0000000" when "00000101000100001", -- t[2593] = 0
      "0000000" when "00000101000100010", -- t[2594] = 0
      "0000000" when "00000101000100011", -- t[2595] = 0
      "0000000" when "00000101000100100", -- t[2596] = 0
      "0000000" when "00000101000100101", -- t[2597] = 0
      "0000000" when "00000101000100110", -- t[2598] = 0
      "0000000" when "00000101000100111", -- t[2599] = 0
      "0000000" when "00000101000101000", -- t[2600] = 0
      "0000000" when "00000101000101001", -- t[2601] = 0
      "0000000" when "00000101000101010", -- t[2602] = 0
      "0000000" when "00000101000101011", -- t[2603] = 0
      "0000000" when "00000101000101100", -- t[2604] = 0
      "0000000" when "00000101000101101", -- t[2605] = 0
      "0000000" when "00000101000101110", -- t[2606] = 0
      "0000000" when "00000101000101111", -- t[2607] = 0
      "0000000" when "00000101000110000", -- t[2608] = 0
      "0000000" when "00000101000110001", -- t[2609] = 0
      "0000000" when "00000101000110010", -- t[2610] = 0
      "0000000" when "00000101000110011", -- t[2611] = 0
      "0000000" when "00000101000110100", -- t[2612] = 0
      "0000000" when "00000101000110101", -- t[2613] = 0
      "0000000" when "00000101000110110", -- t[2614] = 0
      "0000000" when "00000101000110111", -- t[2615] = 0
      "0000000" when "00000101000111000", -- t[2616] = 0
      "0000000" when "00000101000111001", -- t[2617] = 0
      "0000000" when "00000101000111010", -- t[2618] = 0
      "0000000" when "00000101000111011", -- t[2619] = 0
      "0000000" when "00000101000111100", -- t[2620] = 0
      "0000000" when "00000101000111101", -- t[2621] = 0
      "0000000" when "00000101000111110", -- t[2622] = 0
      "0000000" when "00000101000111111", -- t[2623] = 0
      "0000000" when "00000101001000000", -- t[2624] = 0
      "0000000" when "00000101001000001", -- t[2625] = 0
      "0000000" when "00000101001000010", -- t[2626] = 0
      "0000000" when "00000101001000011", -- t[2627] = 0
      "0000000" when "00000101001000100", -- t[2628] = 0
      "0000000" when "00000101001000101", -- t[2629] = 0
      "0000000" when "00000101001000110", -- t[2630] = 0
      "0000000" when "00000101001000111", -- t[2631] = 0
      "0000000" when "00000101001001000", -- t[2632] = 0
      "0000000" when "00000101001001001", -- t[2633] = 0
      "0000000" when "00000101001001010", -- t[2634] = 0
      "0000000" when "00000101001001011", -- t[2635] = 0
      "0000000" when "00000101001001100", -- t[2636] = 0
      "0000000" when "00000101001001101", -- t[2637] = 0
      "0000000" when "00000101001001110", -- t[2638] = 0
      "0000000" when "00000101001001111", -- t[2639] = 0
      "0000000" when "00000101001010000", -- t[2640] = 0
      "0000000" when "00000101001010001", -- t[2641] = 0
      "0000000" when "00000101001010010", -- t[2642] = 0
      "0000000" when "00000101001010011", -- t[2643] = 0
      "0000000" when "00000101001010100", -- t[2644] = 0
      "0000000" when "00000101001010101", -- t[2645] = 0
      "0000000" when "00000101001010110", -- t[2646] = 0
      "0000000" when "00000101001010111", -- t[2647] = 0
      "0000000" when "00000101001011000", -- t[2648] = 0
      "0000000" when "00000101001011001", -- t[2649] = 0
      "0000000" when "00000101001011010", -- t[2650] = 0
      "0000000" when "00000101001011011", -- t[2651] = 0
      "0000000" when "00000101001011100", -- t[2652] = 0
      "0000000" when "00000101001011101", -- t[2653] = 0
      "0000000" when "00000101001011110", -- t[2654] = 0
      "0000000" when "00000101001011111", -- t[2655] = 0
      "0000000" when "00000101001100000", -- t[2656] = 0
      "0000000" when "00000101001100001", -- t[2657] = 0
      "0000000" when "00000101001100010", -- t[2658] = 0
      "0000000" when "00000101001100011", -- t[2659] = 0
      "0000000" when "00000101001100100", -- t[2660] = 0
      "0000000" when "00000101001100101", -- t[2661] = 0
      "0000000" when "00000101001100110", -- t[2662] = 0
      "0000000" when "00000101001100111", -- t[2663] = 0
      "0000000" when "00000101001101000", -- t[2664] = 0
      "0000000" when "00000101001101001", -- t[2665] = 0
      "0000000" when "00000101001101010", -- t[2666] = 0
      "0000000" when "00000101001101011", -- t[2667] = 0
      "0000000" when "00000101001101100", -- t[2668] = 0
      "0000000" when "00000101001101101", -- t[2669] = 0
      "0000000" when "00000101001101110", -- t[2670] = 0
      "0000000" when "00000101001101111", -- t[2671] = 0
      "0000000" when "00000101001110000", -- t[2672] = 0
      "0000000" when "00000101001110001", -- t[2673] = 0
      "0000000" when "00000101001110010", -- t[2674] = 0
      "0000000" when "00000101001110011", -- t[2675] = 0
      "0000000" when "00000101001110100", -- t[2676] = 0
      "0000000" when "00000101001110101", -- t[2677] = 0
      "0000000" when "00000101001110110", -- t[2678] = 0
      "0000000" when "00000101001110111", -- t[2679] = 0
      "0000000" when "00000101001111000", -- t[2680] = 0
      "0000000" when "00000101001111001", -- t[2681] = 0
      "0000000" when "00000101001111010", -- t[2682] = 0
      "0000000" when "00000101001111011", -- t[2683] = 0
      "0000000" when "00000101001111100", -- t[2684] = 0
      "0000000" when "00000101001111101", -- t[2685] = 0
      "0000000" when "00000101001111110", -- t[2686] = 0
      "0000000" when "00000101001111111", -- t[2687] = 0
      "0000000" when "00000101010000000", -- t[2688] = 0
      "0000000" when "00000101010000001", -- t[2689] = 0
      "0000000" when "00000101010000010", -- t[2690] = 0
      "0000000" when "00000101010000011", -- t[2691] = 0
      "0000000" when "00000101010000100", -- t[2692] = 0
      "0000000" when "00000101010000101", -- t[2693] = 0
      "0000000" when "00000101010000110", -- t[2694] = 0
      "0000000" when "00000101010000111", -- t[2695] = 0
      "0000000" when "00000101010001000", -- t[2696] = 0
      "0000000" when "00000101010001001", -- t[2697] = 0
      "0000000" when "00000101010001010", -- t[2698] = 0
      "0000000" when "00000101010001011", -- t[2699] = 0
      "0000000" when "00000101010001100", -- t[2700] = 0
      "0000000" when "00000101010001101", -- t[2701] = 0
      "0000000" when "00000101010001110", -- t[2702] = 0
      "0000000" when "00000101010001111", -- t[2703] = 0
      "0000000" when "00000101010010000", -- t[2704] = 0
      "0000000" when "00000101010010001", -- t[2705] = 0
      "0000000" when "00000101010010010", -- t[2706] = 0
      "0000000" when "00000101010010011", -- t[2707] = 0
      "0000000" when "00000101010010100", -- t[2708] = 0
      "0000000" when "00000101010010101", -- t[2709] = 0
      "0000000" when "00000101010010110", -- t[2710] = 0
      "0000000" when "00000101010010111", -- t[2711] = 0
      "0000000" when "00000101010011000", -- t[2712] = 0
      "0000000" when "00000101010011001", -- t[2713] = 0
      "0000000" when "00000101010011010", -- t[2714] = 0
      "0000000" when "00000101010011011", -- t[2715] = 0
      "0000000" when "00000101010011100", -- t[2716] = 0
      "0000000" when "00000101010011101", -- t[2717] = 0
      "0000000" when "00000101010011110", -- t[2718] = 0
      "0000000" when "00000101010011111", -- t[2719] = 0
      "0000000" when "00000101010100000", -- t[2720] = 0
      "0000000" when "00000101010100001", -- t[2721] = 0
      "0000000" when "00000101010100010", -- t[2722] = 0
      "0000000" when "00000101010100011", -- t[2723] = 0
      "0000000" when "00000101010100100", -- t[2724] = 0
      "0000000" when "00000101010100101", -- t[2725] = 0
      "0000000" when "00000101010100110", -- t[2726] = 0
      "0000000" when "00000101010100111", -- t[2727] = 0
      "0000000" when "00000101010101000", -- t[2728] = 0
      "0000000" when "00000101010101001", -- t[2729] = 0
      "0000000" when "00000101010101010", -- t[2730] = 0
      "0000000" when "00000101010101011", -- t[2731] = 0
      "0000000" when "00000101010101100", -- t[2732] = 0
      "0000000" when "00000101010101101", -- t[2733] = 0
      "0000000" when "00000101010101110", -- t[2734] = 0
      "0000000" when "00000101010101111", -- t[2735] = 0
      "0000000" when "00000101010110000", -- t[2736] = 0
      "0000000" when "00000101010110001", -- t[2737] = 0
      "0000000" when "00000101010110010", -- t[2738] = 0
      "0000000" when "00000101010110011", -- t[2739] = 0
      "0000000" when "00000101010110100", -- t[2740] = 0
      "0000000" when "00000101010110101", -- t[2741] = 0
      "0000000" when "00000101010110110", -- t[2742] = 0
      "0000000" when "00000101010110111", -- t[2743] = 0
      "0000000" when "00000101010111000", -- t[2744] = 0
      "0000000" when "00000101010111001", -- t[2745] = 0
      "0000000" when "00000101010111010", -- t[2746] = 0
      "0000000" when "00000101010111011", -- t[2747] = 0
      "0000000" when "00000101010111100", -- t[2748] = 0
      "0000000" when "00000101010111101", -- t[2749] = 0
      "0000000" when "00000101010111110", -- t[2750] = 0
      "0000000" when "00000101010111111", -- t[2751] = 0
      "0000000" when "00000101011000000", -- t[2752] = 0
      "0000000" when "00000101011000001", -- t[2753] = 0
      "0000000" when "00000101011000010", -- t[2754] = 0
      "0000000" when "00000101011000011", -- t[2755] = 0
      "0000000" when "00000101011000100", -- t[2756] = 0
      "0000000" when "00000101011000101", -- t[2757] = 0
      "0000000" when "00000101011000110", -- t[2758] = 0
      "0000000" when "00000101011000111", -- t[2759] = 0
      "0000000" when "00000101011001000", -- t[2760] = 0
      "0000000" when "00000101011001001", -- t[2761] = 0
      "0000000" when "00000101011001010", -- t[2762] = 0
      "0000000" when "00000101011001011", -- t[2763] = 0
      "0000000" when "00000101011001100", -- t[2764] = 0
      "0000000" when "00000101011001101", -- t[2765] = 0
      "0000000" when "00000101011001110", -- t[2766] = 0
      "0000000" when "00000101011001111", -- t[2767] = 0
      "0000000" when "00000101011010000", -- t[2768] = 0
      "0000000" when "00000101011010001", -- t[2769] = 0
      "0000000" when "00000101011010010", -- t[2770] = 0
      "0000000" when "00000101011010011", -- t[2771] = 0
      "0000000" when "00000101011010100", -- t[2772] = 0
      "0000000" when "00000101011010101", -- t[2773] = 0
      "0000000" when "00000101011010110", -- t[2774] = 0
      "0000000" when "00000101011010111", -- t[2775] = 0
      "0000000" when "00000101011011000", -- t[2776] = 0
      "0000000" when "00000101011011001", -- t[2777] = 0
      "0000000" when "00000101011011010", -- t[2778] = 0
      "0000000" when "00000101011011011", -- t[2779] = 0
      "0000000" when "00000101011011100", -- t[2780] = 0
      "0000000" when "00000101011011101", -- t[2781] = 0
      "0000000" when "00000101011011110", -- t[2782] = 0
      "0000000" when "00000101011011111", -- t[2783] = 0
      "0000000" when "00000101011100000", -- t[2784] = 0
      "0000000" when "00000101011100001", -- t[2785] = 0
      "0000000" when "00000101011100010", -- t[2786] = 0
      "0000000" when "00000101011100011", -- t[2787] = 0
      "0000000" when "00000101011100100", -- t[2788] = 0
      "0000000" when "00000101011100101", -- t[2789] = 0
      "0000000" when "00000101011100110", -- t[2790] = 0
      "0000000" when "00000101011100111", -- t[2791] = 0
      "0000000" when "00000101011101000", -- t[2792] = 0
      "0000000" when "00000101011101001", -- t[2793] = 0
      "0000000" when "00000101011101010", -- t[2794] = 0
      "0000000" when "00000101011101011", -- t[2795] = 0
      "0000000" when "00000101011101100", -- t[2796] = 0
      "0000000" when "00000101011101101", -- t[2797] = 0
      "0000000" when "00000101011101110", -- t[2798] = 0
      "0000000" when "00000101011101111", -- t[2799] = 0
      "0000000" when "00000101011110000", -- t[2800] = 0
      "0000000" when "00000101011110001", -- t[2801] = 0
      "0000000" when "00000101011110010", -- t[2802] = 0
      "0000000" when "00000101011110011", -- t[2803] = 0
      "0000000" when "00000101011110100", -- t[2804] = 0
      "0000000" when "00000101011110101", -- t[2805] = 0
      "0000000" when "00000101011110110", -- t[2806] = 0
      "0000000" when "00000101011110111", -- t[2807] = 0
      "0000000" when "00000101011111000", -- t[2808] = 0
      "0000000" when "00000101011111001", -- t[2809] = 0
      "0000000" when "00000101011111010", -- t[2810] = 0
      "0000000" when "00000101011111011", -- t[2811] = 0
      "0000000" when "00000101011111100", -- t[2812] = 0
      "0000000" when "00000101011111101", -- t[2813] = 0
      "0000000" when "00000101011111110", -- t[2814] = 0
      "0000000" when "00000101011111111", -- t[2815] = 0
      "0000000" when "00000101100000000", -- t[2816] = 0
      "0000000" when "00000101100000001", -- t[2817] = 0
      "0000000" when "00000101100000010", -- t[2818] = 0
      "0000000" when "00000101100000011", -- t[2819] = 0
      "0000000" when "00000101100000100", -- t[2820] = 0
      "0000000" when "00000101100000101", -- t[2821] = 0
      "0000000" when "00000101100000110", -- t[2822] = 0
      "0000000" when "00000101100000111", -- t[2823] = 0
      "0000000" when "00000101100001000", -- t[2824] = 0
      "0000000" when "00000101100001001", -- t[2825] = 0
      "0000000" when "00000101100001010", -- t[2826] = 0
      "0000000" when "00000101100001011", -- t[2827] = 0
      "0000000" when "00000101100001100", -- t[2828] = 0
      "0000000" when "00000101100001101", -- t[2829] = 0
      "0000000" when "00000101100001110", -- t[2830] = 0
      "0000000" when "00000101100001111", -- t[2831] = 0
      "0000000" when "00000101100010000", -- t[2832] = 0
      "0000000" when "00000101100010001", -- t[2833] = 0
      "0000000" when "00000101100010010", -- t[2834] = 0
      "0000000" when "00000101100010011", -- t[2835] = 0
      "0000000" when "00000101100010100", -- t[2836] = 0
      "0000000" when "00000101100010101", -- t[2837] = 0
      "0000000" when "00000101100010110", -- t[2838] = 0
      "0000000" when "00000101100010111", -- t[2839] = 0
      "0000000" when "00000101100011000", -- t[2840] = 0
      "0000000" when "00000101100011001", -- t[2841] = 0
      "0000000" when "00000101100011010", -- t[2842] = 0
      "0000000" when "00000101100011011", -- t[2843] = 0
      "0000000" when "00000101100011100", -- t[2844] = 0
      "0000000" when "00000101100011101", -- t[2845] = 0
      "0000000" when "00000101100011110", -- t[2846] = 0
      "0000000" when "00000101100011111", -- t[2847] = 0
      "0000000" when "00000101100100000", -- t[2848] = 0
      "0000000" when "00000101100100001", -- t[2849] = 0
      "0000000" when "00000101100100010", -- t[2850] = 0
      "0000000" when "00000101100100011", -- t[2851] = 0
      "0000000" when "00000101100100100", -- t[2852] = 0
      "0000000" when "00000101100100101", -- t[2853] = 0
      "0000000" when "00000101100100110", -- t[2854] = 0
      "0000000" when "00000101100100111", -- t[2855] = 0
      "0000000" when "00000101100101000", -- t[2856] = 0
      "0000000" when "00000101100101001", -- t[2857] = 0
      "0000000" when "00000101100101010", -- t[2858] = 0
      "0000000" when "00000101100101011", -- t[2859] = 0
      "0000000" when "00000101100101100", -- t[2860] = 0
      "0000000" when "00000101100101101", -- t[2861] = 0
      "0000000" when "00000101100101110", -- t[2862] = 0
      "0000000" when "00000101100101111", -- t[2863] = 0
      "0000000" when "00000101100110000", -- t[2864] = 0
      "0000000" when "00000101100110001", -- t[2865] = 0
      "0000000" when "00000101100110010", -- t[2866] = 0
      "0000000" when "00000101100110011", -- t[2867] = 0
      "0000000" when "00000101100110100", -- t[2868] = 0
      "0000000" when "00000101100110101", -- t[2869] = 0
      "0000000" when "00000101100110110", -- t[2870] = 0
      "0000000" when "00000101100110111", -- t[2871] = 0
      "0000000" when "00000101100111000", -- t[2872] = 0
      "0000000" when "00000101100111001", -- t[2873] = 0
      "0000000" when "00000101100111010", -- t[2874] = 0
      "0000000" when "00000101100111011", -- t[2875] = 0
      "0000000" when "00000101100111100", -- t[2876] = 0
      "0000000" when "00000101100111101", -- t[2877] = 0
      "0000000" when "00000101100111110", -- t[2878] = 0
      "0000000" when "00000101100111111", -- t[2879] = 0
      "0000000" when "00000101101000000", -- t[2880] = 0
      "0000000" when "00000101101000001", -- t[2881] = 0
      "0000000" when "00000101101000010", -- t[2882] = 0
      "0000000" when "00000101101000011", -- t[2883] = 0
      "0000000" when "00000101101000100", -- t[2884] = 0
      "0000000" when "00000101101000101", -- t[2885] = 0
      "0000000" when "00000101101000110", -- t[2886] = 0
      "0000000" when "00000101101000111", -- t[2887] = 0
      "0000000" when "00000101101001000", -- t[2888] = 0
      "0000000" when "00000101101001001", -- t[2889] = 0
      "0000000" when "00000101101001010", -- t[2890] = 0
      "0000000" when "00000101101001011", -- t[2891] = 0
      "0000000" when "00000101101001100", -- t[2892] = 0
      "0000000" when "00000101101001101", -- t[2893] = 0
      "0000000" when "00000101101001110", -- t[2894] = 0
      "0000000" when "00000101101001111", -- t[2895] = 0
      "0000000" when "00000101101010000", -- t[2896] = 0
      "0000000" when "00000101101010001", -- t[2897] = 0
      "0000000" when "00000101101010010", -- t[2898] = 0
      "0000000" when "00000101101010011", -- t[2899] = 0
      "0000000" when "00000101101010100", -- t[2900] = 0
      "0000000" when "00000101101010101", -- t[2901] = 0
      "0000000" when "00000101101010110", -- t[2902] = 0
      "0000000" when "00000101101010111", -- t[2903] = 0
      "0000000" when "00000101101011000", -- t[2904] = 0
      "0000000" when "00000101101011001", -- t[2905] = 0
      "0000000" when "00000101101011010", -- t[2906] = 0
      "0000000" when "00000101101011011", -- t[2907] = 0
      "0000000" when "00000101101011100", -- t[2908] = 0
      "0000000" when "00000101101011101", -- t[2909] = 0
      "0000000" when "00000101101011110", -- t[2910] = 0
      "0000000" when "00000101101011111", -- t[2911] = 0
      "0000000" when "00000101101100000", -- t[2912] = 0
      "0000000" when "00000101101100001", -- t[2913] = 0
      "0000000" when "00000101101100010", -- t[2914] = 0
      "0000000" when "00000101101100011", -- t[2915] = 0
      "0000000" when "00000101101100100", -- t[2916] = 0
      "0000000" when "00000101101100101", -- t[2917] = 0
      "0000000" when "00000101101100110", -- t[2918] = 0
      "0000000" when "00000101101100111", -- t[2919] = 0
      "0000000" when "00000101101101000", -- t[2920] = 0
      "0000000" when "00000101101101001", -- t[2921] = 0
      "0000000" when "00000101101101010", -- t[2922] = 0
      "0000000" when "00000101101101011", -- t[2923] = 0
      "0000000" when "00000101101101100", -- t[2924] = 0
      "0000000" when "00000101101101101", -- t[2925] = 0
      "0000000" when "00000101101101110", -- t[2926] = 0
      "0000000" when "00000101101101111", -- t[2927] = 0
      "0000000" when "00000101101110000", -- t[2928] = 0
      "0000000" when "00000101101110001", -- t[2929] = 0
      "0000000" when "00000101101110010", -- t[2930] = 0
      "0000000" when "00000101101110011", -- t[2931] = 0
      "0000000" when "00000101101110100", -- t[2932] = 0
      "0000000" when "00000101101110101", -- t[2933] = 0
      "0000000" when "00000101101110110", -- t[2934] = 0
      "0000000" when "00000101101110111", -- t[2935] = 0
      "0000000" when "00000101101111000", -- t[2936] = 0
      "0000000" when "00000101101111001", -- t[2937] = 0
      "0000000" when "00000101101111010", -- t[2938] = 0
      "0000000" when "00000101101111011", -- t[2939] = 0
      "0000000" when "00000101101111100", -- t[2940] = 0
      "0000000" when "00000101101111101", -- t[2941] = 0
      "0000000" when "00000101101111110", -- t[2942] = 0
      "0000000" when "00000101101111111", -- t[2943] = 0
      "0000000" when "00000101110000000", -- t[2944] = 0
      "0000000" when "00000101110000001", -- t[2945] = 0
      "0000000" when "00000101110000010", -- t[2946] = 0
      "0000000" when "00000101110000011", -- t[2947] = 0
      "0000000" when "00000101110000100", -- t[2948] = 0
      "0000000" when "00000101110000101", -- t[2949] = 0
      "0000000" when "00000101110000110", -- t[2950] = 0
      "0000000" when "00000101110000111", -- t[2951] = 0
      "0000000" when "00000101110001000", -- t[2952] = 0
      "0000000" when "00000101110001001", -- t[2953] = 0
      "0000000" when "00000101110001010", -- t[2954] = 0
      "0000000" when "00000101110001011", -- t[2955] = 0
      "0000000" when "00000101110001100", -- t[2956] = 0
      "0000000" when "00000101110001101", -- t[2957] = 0
      "0000000" when "00000101110001110", -- t[2958] = 0
      "0000000" when "00000101110001111", -- t[2959] = 0
      "0000000" when "00000101110010000", -- t[2960] = 0
      "0000000" when "00000101110010001", -- t[2961] = 0
      "0000000" when "00000101110010010", -- t[2962] = 0
      "0000000" when "00000101110010011", -- t[2963] = 0
      "0000000" when "00000101110010100", -- t[2964] = 0
      "0000000" when "00000101110010101", -- t[2965] = 0
      "0000000" when "00000101110010110", -- t[2966] = 0
      "0000000" when "00000101110010111", -- t[2967] = 0
      "0000000" when "00000101110011000", -- t[2968] = 0
      "0000000" when "00000101110011001", -- t[2969] = 0
      "0000000" when "00000101110011010", -- t[2970] = 0
      "0000000" when "00000101110011011", -- t[2971] = 0
      "0000000" when "00000101110011100", -- t[2972] = 0
      "0000000" when "00000101110011101", -- t[2973] = 0
      "0000000" when "00000101110011110", -- t[2974] = 0
      "0000000" when "00000101110011111", -- t[2975] = 0
      "0000000" when "00000101110100000", -- t[2976] = 0
      "0000000" when "00000101110100001", -- t[2977] = 0
      "0000000" when "00000101110100010", -- t[2978] = 0
      "0000000" when "00000101110100011", -- t[2979] = 0
      "0000000" when "00000101110100100", -- t[2980] = 0
      "0000000" when "00000101110100101", -- t[2981] = 0
      "0000000" when "00000101110100110", -- t[2982] = 0
      "0000000" when "00000101110100111", -- t[2983] = 0
      "0000000" when "00000101110101000", -- t[2984] = 0
      "0000000" when "00000101110101001", -- t[2985] = 0
      "0000000" when "00000101110101010", -- t[2986] = 0
      "0000000" when "00000101110101011", -- t[2987] = 0
      "0000000" when "00000101110101100", -- t[2988] = 0
      "0000000" when "00000101110101101", -- t[2989] = 0
      "0000000" when "00000101110101110", -- t[2990] = 0
      "0000000" when "00000101110101111", -- t[2991] = 0
      "0000000" when "00000101110110000", -- t[2992] = 0
      "0000000" when "00000101110110001", -- t[2993] = 0
      "0000000" when "00000101110110010", -- t[2994] = 0
      "0000000" when "00000101110110011", -- t[2995] = 0
      "0000000" when "00000101110110100", -- t[2996] = 0
      "0000000" when "00000101110110101", -- t[2997] = 0
      "0000000" when "00000101110110110", -- t[2998] = 0
      "0000000" when "00000101110110111", -- t[2999] = 0
      "0000000" when "00000101110111000", -- t[3000] = 0
      "0000000" when "00000101110111001", -- t[3001] = 0
      "0000000" when "00000101110111010", -- t[3002] = 0
      "0000000" when "00000101110111011", -- t[3003] = 0
      "0000000" when "00000101110111100", -- t[3004] = 0
      "0000000" when "00000101110111101", -- t[3005] = 0
      "0000000" when "00000101110111110", -- t[3006] = 0
      "0000000" when "00000101110111111", -- t[3007] = 0
      "0000000" when "00000101111000000", -- t[3008] = 0
      "0000000" when "00000101111000001", -- t[3009] = 0
      "0000000" when "00000101111000010", -- t[3010] = 0
      "0000000" when "00000101111000011", -- t[3011] = 0
      "0000000" when "00000101111000100", -- t[3012] = 0
      "0000000" when "00000101111000101", -- t[3013] = 0
      "0000000" when "00000101111000110", -- t[3014] = 0
      "0000000" when "00000101111000111", -- t[3015] = 0
      "0000000" when "00000101111001000", -- t[3016] = 0
      "0000000" when "00000101111001001", -- t[3017] = 0
      "0000000" when "00000101111001010", -- t[3018] = 0
      "0000000" when "00000101111001011", -- t[3019] = 0
      "0000000" when "00000101111001100", -- t[3020] = 0
      "0000000" when "00000101111001101", -- t[3021] = 0
      "0000000" when "00000101111001110", -- t[3022] = 0
      "0000000" when "00000101111001111", -- t[3023] = 0
      "0000000" when "00000101111010000", -- t[3024] = 0
      "0000000" when "00000101111010001", -- t[3025] = 0
      "0000000" when "00000101111010010", -- t[3026] = 0
      "0000000" when "00000101111010011", -- t[3027] = 0
      "0000000" when "00000101111010100", -- t[3028] = 0
      "0000000" when "00000101111010101", -- t[3029] = 0
      "0000000" when "00000101111010110", -- t[3030] = 0
      "0000000" when "00000101111010111", -- t[3031] = 0
      "0000000" when "00000101111011000", -- t[3032] = 0
      "0000000" when "00000101111011001", -- t[3033] = 0
      "0000000" when "00000101111011010", -- t[3034] = 0
      "0000000" when "00000101111011011", -- t[3035] = 0
      "0000000" when "00000101111011100", -- t[3036] = 0
      "0000000" when "00000101111011101", -- t[3037] = 0
      "0000000" when "00000101111011110", -- t[3038] = 0
      "0000000" when "00000101111011111", -- t[3039] = 0
      "0000000" when "00000101111100000", -- t[3040] = 0
      "0000000" when "00000101111100001", -- t[3041] = 0
      "0000000" when "00000101111100010", -- t[3042] = 0
      "0000000" when "00000101111100011", -- t[3043] = 0
      "0000000" when "00000101111100100", -- t[3044] = 0
      "0000000" when "00000101111100101", -- t[3045] = 0
      "0000000" when "00000101111100110", -- t[3046] = 0
      "0000000" when "00000101111100111", -- t[3047] = 0
      "0000000" when "00000101111101000", -- t[3048] = 0
      "0000000" when "00000101111101001", -- t[3049] = 0
      "0000000" when "00000101111101010", -- t[3050] = 0
      "0000000" when "00000101111101011", -- t[3051] = 0
      "0000000" when "00000101111101100", -- t[3052] = 0
      "0000000" when "00000101111101101", -- t[3053] = 0
      "0000000" when "00000101111101110", -- t[3054] = 0
      "0000000" when "00000101111101111", -- t[3055] = 0
      "0000000" when "00000101111110000", -- t[3056] = 0
      "0000000" when "00000101111110001", -- t[3057] = 0
      "0000000" when "00000101111110010", -- t[3058] = 0
      "0000000" when "00000101111110011", -- t[3059] = 0
      "0000000" when "00000101111110100", -- t[3060] = 0
      "0000000" when "00000101111110101", -- t[3061] = 0
      "0000000" when "00000101111110110", -- t[3062] = 0
      "0000000" when "00000101111110111", -- t[3063] = 0
      "0000000" when "00000101111111000", -- t[3064] = 0
      "0000000" when "00000101111111001", -- t[3065] = 0
      "0000000" when "00000101111111010", -- t[3066] = 0
      "0000000" when "00000101111111011", -- t[3067] = 0
      "0000000" when "00000101111111100", -- t[3068] = 0
      "0000000" when "00000101111111101", -- t[3069] = 0
      "0000000" when "00000101111111110", -- t[3070] = 0
      "0000000" when "00000101111111111", -- t[3071] = 0
      "0000000" when "00000110000000000", -- t[3072] = 0
      "0000000" when "00000110000000001", -- t[3073] = 0
      "0000000" when "00000110000000010", -- t[3074] = 0
      "0000000" when "00000110000000011", -- t[3075] = 0
      "0000000" when "00000110000000100", -- t[3076] = 0
      "0000000" when "00000110000000101", -- t[3077] = 0
      "0000000" when "00000110000000110", -- t[3078] = 0
      "0000000" when "00000110000000111", -- t[3079] = 0
      "0000000" when "00000110000001000", -- t[3080] = 0
      "0000000" when "00000110000001001", -- t[3081] = 0
      "0000000" when "00000110000001010", -- t[3082] = 0
      "0000000" when "00000110000001011", -- t[3083] = 0
      "0000000" when "00000110000001100", -- t[3084] = 0
      "0000000" when "00000110000001101", -- t[3085] = 0
      "0000000" when "00000110000001110", -- t[3086] = 0
      "0000000" when "00000110000001111", -- t[3087] = 0
      "0000000" when "00000110000010000", -- t[3088] = 0
      "0000000" when "00000110000010001", -- t[3089] = 0
      "0000000" when "00000110000010010", -- t[3090] = 0
      "0000000" when "00000110000010011", -- t[3091] = 0
      "0000000" when "00000110000010100", -- t[3092] = 0
      "0000000" when "00000110000010101", -- t[3093] = 0
      "0000000" when "00000110000010110", -- t[3094] = 0
      "0000000" when "00000110000010111", -- t[3095] = 0
      "0000000" when "00000110000011000", -- t[3096] = 0
      "0000000" when "00000110000011001", -- t[3097] = 0
      "0000000" when "00000110000011010", -- t[3098] = 0
      "0000000" when "00000110000011011", -- t[3099] = 0
      "0000000" when "00000110000011100", -- t[3100] = 0
      "0000000" when "00000110000011101", -- t[3101] = 0
      "0000000" when "00000110000011110", -- t[3102] = 0
      "0000000" when "00000110000011111", -- t[3103] = 0
      "0000000" when "00000110000100000", -- t[3104] = 0
      "0000000" when "00000110000100001", -- t[3105] = 0
      "0000000" when "00000110000100010", -- t[3106] = 0
      "0000000" when "00000110000100011", -- t[3107] = 0
      "0000000" when "00000110000100100", -- t[3108] = 0
      "0000000" when "00000110000100101", -- t[3109] = 0
      "0000000" when "00000110000100110", -- t[3110] = 0
      "0000000" when "00000110000100111", -- t[3111] = 0
      "0000000" when "00000110000101000", -- t[3112] = 0
      "0000000" when "00000110000101001", -- t[3113] = 0
      "0000000" when "00000110000101010", -- t[3114] = 0
      "0000000" when "00000110000101011", -- t[3115] = 0
      "0000000" when "00000110000101100", -- t[3116] = 0
      "0000000" when "00000110000101101", -- t[3117] = 0
      "0000000" when "00000110000101110", -- t[3118] = 0
      "0000000" when "00000110000101111", -- t[3119] = 0
      "0000000" when "00000110000110000", -- t[3120] = 0
      "0000000" when "00000110000110001", -- t[3121] = 0
      "0000000" when "00000110000110010", -- t[3122] = 0
      "0000000" when "00000110000110011", -- t[3123] = 0
      "0000000" when "00000110000110100", -- t[3124] = 0
      "0000000" when "00000110000110101", -- t[3125] = 0
      "0000000" when "00000110000110110", -- t[3126] = 0
      "0000000" when "00000110000110111", -- t[3127] = 0
      "0000000" when "00000110000111000", -- t[3128] = 0
      "0000000" when "00000110000111001", -- t[3129] = 0
      "0000000" when "00000110000111010", -- t[3130] = 0
      "0000000" when "00000110000111011", -- t[3131] = 0
      "0000000" when "00000110000111100", -- t[3132] = 0
      "0000000" when "00000110000111101", -- t[3133] = 0
      "0000000" when "00000110000111110", -- t[3134] = 0
      "0000000" when "00000110000111111", -- t[3135] = 0
      "0000000" when "00000110001000000", -- t[3136] = 0
      "0000000" when "00000110001000001", -- t[3137] = 0
      "0000000" when "00000110001000010", -- t[3138] = 0
      "0000000" when "00000110001000011", -- t[3139] = 0
      "0000000" when "00000110001000100", -- t[3140] = 0
      "0000000" when "00000110001000101", -- t[3141] = 0
      "0000000" when "00000110001000110", -- t[3142] = 0
      "0000000" when "00000110001000111", -- t[3143] = 0
      "0000000" when "00000110001001000", -- t[3144] = 0
      "0000000" when "00000110001001001", -- t[3145] = 0
      "0000000" when "00000110001001010", -- t[3146] = 0
      "0000000" when "00000110001001011", -- t[3147] = 0
      "0000000" when "00000110001001100", -- t[3148] = 0
      "0000000" when "00000110001001101", -- t[3149] = 0
      "0000000" when "00000110001001110", -- t[3150] = 0
      "0000000" when "00000110001001111", -- t[3151] = 0
      "0000000" when "00000110001010000", -- t[3152] = 0
      "0000000" when "00000110001010001", -- t[3153] = 0
      "0000000" when "00000110001010010", -- t[3154] = 0
      "0000000" when "00000110001010011", -- t[3155] = 0
      "0000000" when "00000110001010100", -- t[3156] = 0
      "0000000" when "00000110001010101", -- t[3157] = 0
      "0000000" when "00000110001010110", -- t[3158] = 0
      "0000000" when "00000110001010111", -- t[3159] = 0
      "0000000" when "00000110001011000", -- t[3160] = 0
      "0000000" when "00000110001011001", -- t[3161] = 0
      "0000000" when "00000110001011010", -- t[3162] = 0
      "0000000" when "00000110001011011", -- t[3163] = 0
      "0000000" when "00000110001011100", -- t[3164] = 0
      "0000000" when "00000110001011101", -- t[3165] = 0
      "0000000" when "00000110001011110", -- t[3166] = 0
      "0000000" when "00000110001011111", -- t[3167] = 0
      "0000000" when "00000110001100000", -- t[3168] = 0
      "0000000" when "00000110001100001", -- t[3169] = 0
      "0000000" when "00000110001100010", -- t[3170] = 0
      "0000000" when "00000110001100011", -- t[3171] = 0
      "0000000" when "00000110001100100", -- t[3172] = 0
      "0000000" when "00000110001100101", -- t[3173] = 0
      "0000000" when "00000110001100110", -- t[3174] = 0
      "0000000" when "00000110001100111", -- t[3175] = 0
      "0000000" when "00000110001101000", -- t[3176] = 0
      "0000000" when "00000110001101001", -- t[3177] = 0
      "0000000" when "00000110001101010", -- t[3178] = 0
      "0000000" when "00000110001101011", -- t[3179] = 0
      "0000000" when "00000110001101100", -- t[3180] = 0
      "0000000" when "00000110001101101", -- t[3181] = 0
      "0000000" when "00000110001101110", -- t[3182] = 0
      "0000000" when "00000110001101111", -- t[3183] = 0
      "0000000" when "00000110001110000", -- t[3184] = 0
      "0000000" when "00000110001110001", -- t[3185] = 0
      "0000000" when "00000110001110010", -- t[3186] = 0
      "0000000" when "00000110001110011", -- t[3187] = 0
      "0000000" when "00000110001110100", -- t[3188] = 0
      "0000000" when "00000110001110101", -- t[3189] = 0
      "0000000" when "00000110001110110", -- t[3190] = 0
      "0000000" when "00000110001110111", -- t[3191] = 0
      "0000000" when "00000110001111000", -- t[3192] = 0
      "0000000" when "00000110001111001", -- t[3193] = 0
      "0000000" when "00000110001111010", -- t[3194] = 0
      "0000000" when "00000110001111011", -- t[3195] = 0
      "0000000" when "00000110001111100", -- t[3196] = 0
      "0000000" when "00000110001111101", -- t[3197] = 0
      "0000000" when "00000110001111110", -- t[3198] = 0
      "0000000" when "00000110001111111", -- t[3199] = 0
      "0000000" when "00000110010000000", -- t[3200] = 0
      "0000000" when "00000110010000001", -- t[3201] = 0
      "0000000" when "00000110010000010", -- t[3202] = 0
      "0000000" when "00000110010000011", -- t[3203] = 0
      "0000000" when "00000110010000100", -- t[3204] = 0
      "0000000" when "00000110010000101", -- t[3205] = 0
      "0000000" when "00000110010000110", -- t[3206] = 0
      "0000000" when "00000110010000111", -- t[3207] = 0
      "0000000" when "00000110010001000", -- t[3208] = 0
      "0000000" when "00000110010001001", -- t[3209] = 0
      "0000000" when "00000110010001010", -- t[3210] = 0
      "0000000" when "00000110010001011", -- t[3211] = 0
      "0000000" when "00000110010001100", -- t[3212] = 0
      "0000000" when "00000110010001101", -- t[3213] = 0
      "0000000" when "00000110010001110", -- t[3214] = 0
      "0000000" when "00000110010001111", -- t[3215] = 0
      "0000000" when "00000110010010000", -- t[3216] = 0
      "0000000" when "00000110010010001", -- t[3217] = 0
      "0000000" when "00000110010010010", -- t[3218] = 0
      "0000000" when "00000110010010011", -- t[3219] = 0
      "0000000" when "00000110010010100", -- t[3220] = 0
      "0000000" when "00000110010010101", -- t[3221] = 0
      "0000000" when "00000110010010110", -- t[3222] = 0
      "0000000" when "00000110010010111", -- t[3223] = 0
      "0000000" when "00000110010011000", -- t[3224] = 0
      "0000000" when "00000110010011001", -- t[3225] = 0
      "0000000" when "00000110010011010", -- t[3226] = 0
      "0000000" when "00000110010011011", -- t[3227] = 0
      "0000000" when "00000110010011100", -- t[3228] = 0
      "0000000" when "00000110010011101", -- t[3229] = 0
      "0000000" when "00000110010011110", -- t[3230] = 0
      "0000000" when "00000110010011111", -- t[3231] = 0
      "0000000" when "00000110010100000", -- t[3232] = 0
      "0000000" when "00000110010100001", -- t[3233] = 0
      "0000000" when "00000110010100010", -- t[3234] = 0
      "0000000" when "00000110010100011", -- t[3235] = 0
      "0000000" when "00000110010100100", -- t[3236] = 0
      "0000000" when "00000110010100101", -- t[3237] = 0
      "0000000" when "00000110010100110", -- t[3238] = 0
      "0000000" when "00000110010100111", -- t[3239] = 0
      "0000000" when "00000110010101000", -- t[3240] = 0
      "0000000" when "00000110010101001", -- t[3241] = 0
      "0000000" when "00000110010101010", -- t[3242] = 0
      "0000000" when "00000110010101011", -- t[3243] = 0
      "0000000" when "00000110010101100", -- t[3244] = 0
      "0000000" when "00000110010101101", -- t[3245] = 0
      "0000000" when "00000110010101110", -- t[3246] = 0
      "0000000" when "00000110010101111", -- t[3247] = 0
      "0000000" when "00000110010110000", -- t[3248] = 0
      "0000000" when "00000110010110001", -- t[3249] = 0
      "0000000" when "00000110010110010", -- t[3250] = 0
      "0000000" when "00000110010110011", -- t[3251] = 0
      "0000000" when "00000110010110100", -- t[3252] = 0
      "0000000" when "00000110010110101", -- t[3253] = 0
      "0000000" when "00000110010110110", -- t[3254] = 0
      "0000000" when "00000110010110111", -- t[3255] = 0
      "0000000" when "00000110010111000", -- t[3256] = 0
      "0000000" when "00000110010111001", -- t[3257] = 0
      "0000000" when "00000110010111010", -- t[3258] = 0
      "0000000" when "00000110010111011", -- t[3259] = 0
      "0000000" when "00000110010111100", -- t[3260] = 0
      "0000000" when "00000110010111101", -- t[3261] = 0
      "0000000" when "00000110010111110", -- t[3262] = 0
      "0000000" when "00000110010111111", -- t[3263] = 0
      "0000000" when "00000110011000000", -- t[3264] = 0
      "0000000" when "00000110011000001", -- t[3265] = 0
      "0000000" when "00000110011000010", -- t[3266] = 0
      "0000000" when "00000110011000011", -- t[3267] = 0
      "0000000" when "00000110011000100", -- t[3268] = 0
      "0000000" when "00000110011000101", -- t[3269] = 0
      "0000000" when "00000110011000110", -- t[3270] = 0
      "0000000" when "00000110011000111", -- t[3271] = 0
      "0000000" when "00000110011001000", -- t[3272] = 0
      "0000000" when "00000110011001001", -- t[3273] = 0
      "0000000" when "00000110011001010", -- t[3274] = 0
      "0000000" when "00000110011001011", -- t[3275] = 0
      "0000000" when "00000110011001100", -- t[3276] = 0
      "0000000" when "00000110011001101", -- t[3277] = 0
      "0000000" when "00000110011001110", -- t[3278] = 0
      "0000000" when "00000110011001111", -- t[3279] = 0
      "0000000" when "00000110011010000", -- t[3280] = 0
      "0000000" when "00000110011010001", -- t[3281] = 0
      "0000000" when "00000110011010010", -- t[3282] = 0
      "0000000" when "00000110011010011", -- t[3283] = 0
      "0000000" when "00000110011010100", -- t[3284] = 0
      "0000000" when "00000110011010101", -- t[3285] = 0
      "0000000" when "00000110011010110", -- t[3286] = 0
      "0000000" when "00000110011010111", -- t[3287] = 0
      "0000000" when "00000110011011000", -- t[3288] = 0
      "0000000" when "00000110011011001", -- t[3289] = 0
      "0000000" when "00000110011011010", -- t[3290] = 0
      "0000000" when "00000110011011011", -- t[3291] = 0
      "0000000" when "00000110011011100", -- t[3292] = 0
      "0000000" when "00000110011011101", -- t[3293] = 0
      "0000000" when "00000110011011110", -- t[3294] = 0
      "0000000" when "00000110011011111", -- t[3295] = 0
      "0000000" when "00000110011100000", -- t[3296] = 0
      "0000000" when "00000110011100001", -- t[3297] = 0
      "0000000" when "00000110011100010", -- t[3298] = 0
      "0000000" when "00000110011100011", -- t[3299] = 0
      "0000000" when "00000110011100100", -- t[3300] = 0
      "0000000" when "00000110011100101", -- t[3301] = 0
      "0000000" when "00000110011100110", -- t[3302] = 0
      "0000000" when "00000110011100111", -- t[3303] = 0
      "0000000" when "00000110011101000", -- t[3304] = 0
      "0000000" when "00000110011101001", -- t[3305] = 0
      "0000000" when "00000110011101010", -- t[3306] = 0
      "0000000" when "00000110011101011", -- t[3307] = 0
      "0000000" when "00000110011101100", -- t[3308] = 0
      "0000000" when "00000110011101101", -- t[3309] = 0
      "0000000" when "00000110011101110", -- t[3310] = 0
      "0000000" when "00000110011101111", -- t[3311] = 0
      "0000000" when "00000110011110000", -- t[3312] = 0
      "0000000" when "00000110011110001", -- t[3313] = 0
      "0000000" when "00000110011110010", -- t[3314] = 0
      "0000000" when "00000110011110011", -- t[3315] = 0
      "0000000" when "00000110011110100", -- t[3316] = 0
      "0000000" when "00000110011110101", -- t[3317] = 0
      "0000000" when "00000110011110110", -- t[3318] = 0
      "0000000" when "00000110011110111", -- t[3319] = 0
      "0000000" when "00000110011111000", -- t[3320] = 0
      "0000000" when "00000110011111001", -- t[3321] = 0
      "0000000" when "00000110011111010", -- t[3322] = 0
      "0000000" when "00000110011111011", -- t[3323] = 0
      "0000000" when "00000110011111100", -- t[3324] = 0
      "0000000" when "00000110011111101", -- t[3325] = 0
      "0000000" when "00000110011111110", -- t[3326] = 0
      "0000000" when "00000110011111111", -- t[3327] = 0
      "0000000" when "00000110100000000", -- t[3328] = 0
      "0000000" when "00000110100000001", -- t[3329] = 0
      "0000000" when "00000110100000010", -- t[3330] = 0
      "0000000" when "00000110100000011", -- t[3331] = 0
      "0000000" when "00000110100000100", -- t[3332] = 0
      "0000000" when "00000110100000101", -- t[3333] = 0
      "0000000" when "00000110100000110", -- t[3334] = 0
      "0000000" when "00000110100000111", -- t[3335] = 0
      "0000000" when "00000110100001000", -- t[3336] = 0
      "0000000" when "00000110100001001", -- t[3337] = 0
      "0000000" when "00000110100001010", -- t[3338] = 0
      "0000000" when "00000110100001011", -- t[3339] = 0
      "0000000" when "00000110100001100", -- t[3340] = 0
      "0000000" when "00000110100001101", -- t[3341] = 0
      "0000000" when "00000110100001110", -- t[3342] = 0
      "0000000" when "00000110100001111", -- t[3343] = 0
      "0000000" when "00000110100010000", -- t[3344] = 0
      "0000000" when "00000110100010001", -- t[3345] = 0
      "0000000" when "00000110100010010", -- t[3346] = 0
      "0000000" when "00000110100010011", -- t[3347] = 0
      "0000000" when "00000110100010100", -- t[3348] = 0
      "0000000" when "00000110100010101", -- t[3349] = 0
      "0000000" when "00000110100010110", -- t[3350] = 0
      "0000000" when "00000110100010111", -- t[3351] = 0
      "0000000" when "00000110100011000", -- t[3352] = 0
      "0000000" when "00000110100011001", -- t[3353] = 0
      "0000000" when "00000110100011010", -- t[3354] = 0
      "0000000" when "00000110100011011", -- t[3355] = 0
      "0000000" when "00000110100011100", -- t[3356] = 0
      "0000000" when "00000110100011101", -- t[3357] = 0
      "0000000" when "00000110100011110", -- t[3358] = 0
      "0000000" when "00000110100011111", -- t[3359] = 0
      "0000000" when "00000110100100000", -- t[3360] = 0
      "0000000" when "00000110100100001", -- t[3361] = 0
      "0000000" when "00000110100100010", -- t[3362] = 0
      "0000000" when "00000110100100011", -- t[3363] = 0
      "0000000" when "00000110100100100", -- t[3364] = 0
      "0000000" when "00000110100100101", -- t[3365] = 0
      "0000000" when "00000110100100110", -- t[3366] = 0
      "0000000" when "00000110100100111", -- t[3367] = 0
      "0000000" when "00000110100101000", -- t[3368] = 0
      "0000000" when "00000110100101001", -- t[3369] = 0
      "0000000" when "00000110100101010", -- t[3370] = 0
      "0000000" when "00000110100101011", -- t[3371] = 0
      "0000000" when "00000110100101100", -- t[3372] = 0
      "0000000" when "00000110100101101", -- t[3373] = 0
      "0000000" when "00000110100101110", -- t[3374] = 0
      "0000000" when "00000110100101111", -- t[3375] = 0
      "0000000" when "00000110100110000", -- t[3376] = 0
      "0000000" when "00000110100110001", -- t[3377] = 0
      "0000000" when "00000110100110010", -- t[3378] = 0
      "0000000" when "00000110100110011", -- t[3379] = 0
      "0000000" when "00000110100110100", -- t[3380] = 0
      "0000000" when "00000110100110101", -- t[3381] = 0
      "0000000" when "00000110100110110", -- t[3382] = 0
      "0000000" when "00000110100110111", -- t[3383] = 0
      "0000000" when "00000110100111000", -- t[3384] = 0
      "0000000" when "00000110100111001", -- t[3385] = 0
      "0000000" when "00000110100111010", -- t[3386] = 0
      "0000000" when "00000110100111011", -- t[3387] = 0
      "0000000" when "00000110100111100", -- t[3388] = 0
      "0000000" when "00000110100111101", -- t[3389] = 0
      "0000000" when "00000110100111110", -- t[3390] = 0
      "0000000" when "00000110100111111", -- t[3391] = 0
      "0000000" when "00000110101000000", -- t[3392] = 0
      "0000000" when "00000110101000001", -- t[3393] = 0
      "0000000" when "00000110101000010", -- t[3394] = 0
      "0000000" when "00000110101000011", -- t[3395] = 0
      "0000000" when "00000110101000100", -- t[3396] = 0
      "0000000" when "00000110101000101", -- t[3397] = 0
      "0000000" when "00000110101000110", -- t[3398] = 0
      "0000000" when "00000110101000111", -- t[3399] = 0
      "0000000" when "00000110101001000", -- t[3400] = 0
      "0000000" when "00000110101001001", -- t[3401] = 0
      "0000000" when "00000110101001010", -- t[3402] = 0
      "0000000" when "00000110101001011", -- t[3403] = 0
      "0000000" when "00000110101001100", -- t[3404] = 0
      "0000000" when "00000110101001101", -- t[3405] = 0
      "0000000" when "00000110101001110", -- t[3406] = 0
      "0000000" when "00000110101001111", -- t[3407] = 0
      "0000000" when "00000110101010000", -- t[3408] = 0
      "0000000" when "00000110101010001", -- t[3409] = 0
      "0000000" when "00000110101010010", -- t[3410] = 0
      "0000000" when "00000110101010011", -- t[3411] = 0
      "0000000" when "00000110101010100", -- t[3412] = 0
      "0000000" when "00000110101010101", -- t[3413] = 0
      "0000000" when "00000110101010110", -- t[3414] = 0
      "0000000" when "00000110101010111", -- t[3415] = 0
      "0000000" when "00000110101011000", -- t[3416] = 0
      "0000000" when "00000110101011001", -- t[3417] = 0
      "0000000" when "00000110101011010", -- t[3418] = 0
      "0000000" when "00000110101011011", -- t[3419] = 0
      "0000000" when "00000110101011100", -- t[3420] = 0
      "0000000" when "00000110101011101", -- t[3421] = 0
      "0000000" when "00000110101011110", -- t[3422] = 0
      "0000000" when "00000110101011111", -- t[3423] = 0
      "0000000" when "00000110101100000", -- t[3424] = 0
      "0000000" when "00000110101100001", -- t[3425] = 0
      "0000000" when "00000110101100010", -- t[3426] = 0
      "0000000" when "00000110101100011", -- t[3427] = 0
      "0000000" when "00000110101100100", -- t[3428] = 0
      "0000000" when "00000110101100101", -- t[3429] = 0
      "0000000" when "00000110101100110", -- t[3430] = 0
      "0000000" when "00000110101100111", -- t[3431] = 0
      "0000000" when "00000110101101000", -- t[3432] = 0
      "0000000" when "00000110101101001", -- t[3433] = 0
      "0000000" when "00000110101101010", -- t[3434] = 0
      "0000000" when "00000110101101011", -- t[3435] = 0
      "0000000" when "00000110101101100", -- t[3436] = 0
      "0000000" when "00000110101101101", -- t[3437] = 0
      "0000000" when "00000110101101110", -- t[3438] = 0
      "0000000" when "00000110101101111", -- t[3439] = 0
      "0000000" when "00000110101110000", -- t[3440] = 0
      "0000000" when "00000110101110001", -- t[3441] = 0
      "0000000" when "00000110101110010", -- t[3442] = 0
      "0000000" when "00000110101110011", -- t[3443] = 0
      "0000000" when "00000110101110100", -- t[3444] = 0
      "0000000" when "00000110101110101", -- t[3445] = 0
      "0000000" when "00000110101110110", -- t[3446] = 0
      "0000000" when "00000110101110111", -- t[3447] = 0
      "0000000" when "00000110101111000", -- t[3448] = 0
      "0000000" when "00000110101111001", -- t[3449] = 0
      "0000000" when "00000110101111010", -- t[3450] = 0
      "0000000" when "00000110101111011", -- t[3451] = 0
      "0000000" when "00000110101111100", -- t[3452] = 0
      "0000000" when "00000110101111101", -- t[3453] = 0
      "0000000" when "00000110101111110", -- t[3454] = 0
      "0000000" when "00000110101111111", -- t[3455] = 0
      "0000000" when "00000110110000000", -- t[3456] = 0
      "0000000" when "00000110110000001", -- t[3457] = 0
      "0000000" when "00000110110000010", -- t[3458] = 0
      "0000000" when "00000110110000011", -- t[3459] = 0
      "0000000" when "00000110110000100", -- t[3460] = 0
      "0000000" when "00000110110000101", -- t[3461] = 0
      "0000000" when "00000110110000110", -- t[3462] = 0
      "0000000" when "00000110110000111", -- t[3463] = 0
      "0000000" when "00000110110001000", -- t[3464] = 0
      "0000000" when "00000110110001001", -- t[3465] = 0
      "0000000" when "00000110110001010", -- t[3466] = 0
      "0000000" when "00000110110001011", -- t[3467] = 0
      "0000000" when "00000110110001100", -- t[3468] = 0
      "0000000" when "00000110110001101", -- t[3469] = 0
      "0000000" when "00000110110001110", -- t[3470] = 0
      "0000000" when "00000110110001111", -- t[3471] = 0
      "0000000" when "00000110110010000", -- t[3472] = 0
      "0000000" when "00000110110010001", -- t[3473] = 0
      "0000000" when "00000110110010010", -- t[3474] = 0
      "0000000" when "00000110110010011", -- t[3475] = 0
      "0000000" when "00000110110010100", -- t[3476] = 0
      "0000000" when "00000110110010101", -- t[3477] = 0
      "0000000" when "00000110110010110", -- t[3478] = 0
      "0000000" when "00000110110010111", -- t[3479] = 0
      "0000000" when "00000110110011000", -- t[3480] = 0
      "0000000" when "00000110110011001", -- t[3481] = 0
      "0000000" when "00000110110011010", -- t[3482] = 0
      "0000000" when "00000110110011011", -- t[3483] = 0
      "0000000" when "00000110110011100", -- t[3484] = 0
      "0000000" when "00000110110011101", -- t[3485] = 0
      "0000000" when "00000110110011110", -- t[3486] = 0
      "0000000" when "00000110110011111", -- t[3487] = 0
      "0000000" when "00000110110100000", -- t[3488] = 0
      "0000000" when "00000110110100001", -- t[3489] = 0
      "0000000" when "00000110110100010", -- t[3490] = 0
      "0000000" when "00000110110100011", -- t[3491] = 0
      "0000000" when "00000110110100100", -- t[3492] = 0
      "0000000" when "00000110110100101", -- t[3493] = 0
      "0000000" when "00000110110100110", -- t[3494] = 0
      "0000000" when "00000110110100111", -- t[3495] = 0
      "0000000" when "00000110110101000", -- t[3496] = 0
      "0000000" when "00000110110101001", -- t[3497] = 0
      "0000000" when "00000110110101010", -- t[3498] = 0
      "0000000" when "00000110110101011", -- t[3499] = 0
      "0000000" when "00000110110101100", -- t[3500] = 0
      "0000000" when "00000110110101101", -- t[3501] = 0
      "0000000" when "00000110110101110", -- t[3502] = 0
      "0000000" when "00000110110101111", -- t[3503] = 0
      "0000000" when "00000110110110000", -- t[3504] = 0
      "0000000" when "00000110110110001", -- t[3505] = 0
      "0000000" when "00000110110110010", -- t[3506] = 0
      "0000000" when "00000110110110011", -- t[3507] = 0
      "0000000" when "00000110110110100", -- t[3508] = 0
      "0000000" when "00000110110110101", -- t[3509] = 0
      "0000000" when "00000110110110110", -- t[3510] = 0
      "0000000" when "00000110110110111", -- t[3511] = 0
      "0000000" when "00000110110111000", -- t[3512] = 0
      "0000000" when "00000110110111001", -- t[3513] = 0
      "0000000" when "00000110110111010", -- t[3514] = 0
      "0000000" when "00000110110111011", -- t[3515] = 0
      "0000000" when "00000110110111100", -- t[3516] = 0
      "0000000" when "00000110110111101", -- t[3517] = 0
      "0000000" when "00000110110111110", -- t[3518] = 0
      "0000000" when "00000110110111111", -- t[3519] = 0
      "0000000" when "00000110111000000", -- t[3520] = 0
      "0000000" when "00000110111000001", -- t[3521] = 0
      "0000000" when "00000110111000010", -- t[3522] = 0
      "0000000" when "00000110111000011", -- t[3523] = 0
      "0000000" when "00000110111000100", -- t[3524] = 0
      "0000000" when "00000110111000101", -- t[3525] = 0
      "0000000" when "00000110111000110", -- t[3526] = 0
      "0000000" when "00000110111000111", -- t[3527] = 0
      "0000000" when "00000110111001000", -- t[3528] = 0
      "0000000" when "00000110111001001", -- t[3529] = 0
      "0000000" when "00000110111001010", -- t[3530] = 0
      "0000000" when "00000110111001011", -- t[3531] = 0
      "0000000" when "00000110111001100", -- t[3532] = 0
      "0000000" when "00000110111001101", -- t[3533] = 0
      "0000000" when "00000110111001110", -- t[3534] = 0
      "0000000" when "00000110111001111", -- t[3535] = 0
      "0000000" when "00000110111010000", -- t[3536] = 0
      "0000000" when "00000110111010001", -- t[3537] = 0
      "0000000" when "00000110111010010", -- t[3538] = 0
      "0000000" when "00000110111010011", -- t[3539] = 0
      "0000000" when "00000110111010100", -- t[3540] = 0
      "0000000" when "00000110111010101", -- t[3541] = 0
      "0000000" when "00000110111010110", -- t[3542] = 0
      "0000000" when "00000110111010111", -- t[3543] = 0
      "0000000" when "00000110111011000", -- t[3544] = 0
      "0000000" when "00000110111011001", -- t[3545] = 0
      "0000000" when "00000110111011010", -- t[3546] = 0
      "0000000" when "00000110111011011", -- t[3547] = 0
      "0000000" when "00000110111011100", -- t[3548] = 0
      "0000000" when "00000110111011101", -- t[3549] = 0
      "0000000" when "00000110111011110", -- t[3550] = 0
      "0000000" when "00000110111011111", -- t[3551] = 0
      "0000000" when "00000110111100000", -- t[3552] = 0
      "0000000" when "00000110111100001", -- t[3553] = 0
      "0000000" when "00000110111100010", -- t[3554] = 0
      "0000000" when "00000110111100011", -- t[3555] = 0
      "0000000" when "00000110111100100", -- t[3556] = 0
      "0000000" when "00000110111100101", -- t[3557] = 0
      "0000000" when "00000110111100110", -- t[3558] = 0
      "0000000" when "00000110111100111", -- t[3559] = 0
      "0000000" when "00000110111101000", -- t[3560] = 0
      "0000000" when "00000110111101001", -- t[3561] = 0
      "0000000" when "00000110111101010", -- t[3562] = 0
      "0000000" when "00000110111101011", -- t[3563] = 0
      "0000000" when "00000110111101100", -- t[3564] = 0
      "0000000" when "00000110111101101", -- t[3565] = 0
      "0000000" when "00000110111101110", -- t[3566] = 0
      "0000000" when "00000110111101111", -- t[3567] = 0
      "0000000" when "00000110111110000", -- t[3568] = 0
      "0000000" when "00000110111110001", -- t[3569] = 0
      "0000000" when "00000110111110010", -- t[3570] = 0
      "0000000" when "00000110111110011", -- t[3571] = 0
      "0000000" when "00000110111110100", -- t[3572] = 0
      "0000000" when "00000110111110101", -- t[3573] = 0
      "0000000" when "00000110111110110", -- t[3574] = 0
      "0000000" when "00000110111110111", -- t[3575] = 0
      "0000000" when "00000110111111000", -- t[3576] = 0
      "0000000" when "00000110111111001", -- t[3577] = 0
      "0000000" when "00000110111111010", -- t[3578] = 0
      "0000000" when "00000110111111011", -- t[3579] = 0
      "0000000" when "00000110111111100", -- t[3580] = 0
      "0000000" when "00000110111111101", -- t[3581] = 0
      "0000000" when "00000110111111110", -- t[3582] = 0
      "0000000" when "00000110111111111", -- t[3583] = 0
      "0000000" when "00000111000000000", -- t[3584] = 0
      "0000000" when "00000111000000001", -- t[3585] = 0
      "0000000" when "00000111000000010", -- t[3586] = 0
      "0000000" when "00000111000000011", -- t[3587] = 0
      "0000000" when "00000111000000100", -- t[3588] = 0
      "0000000" when "00000111000000101", -- t[3589] = 0
      "0000000" when "00000111000000110", -- t[3590] = 0
      "0000000" when "00000111000000111", -- t[3591] = 0
      "0000000" when "00000111000001000", -- t[3592] = 0
      "0000000" when "00000111000001001", -- t[3593] = 0
      "0000000" when "00000111000001010", -- t[3594] = 0
      "0000000" when "00000111000001011", -- t[3595] = 0
      "0000000" when "00000111000001100", -- t[3596] = 0
      "0000000" when "00000111000001101", -- t[3597] = 0
      "0000000" when "00000111000001110", -- t[3598] = 0
      "0000000" when "00000111000001111", -- t[3599] = 0
      "0000000" when "00000111000010000", -- t[3600] = 0
      "0000000" when "00000111000010001", -- t[3601] = 0
      "0000000" when "00000111000010010", -- t[3602] = 0
      "0000000" when "00000111000010011", -- t[3603] = 0
      "0000000" when "00000111000010100", -- t[3604] = 0
      "0000000" when "00000111000010101", -- t[3605] = 0
      "0000000" when "00000111000010110", -- t[3606] = 0
      "0000000" when "00000111000010111", -- t[3607] = 0
      "0000000" when "00000111000011000", -- t[3608] = 0
      "0000000" when "00000111000011001", -- t[3609] = 0
      "0000000" when "00000111000011010", -- t[3610] = 0
      "0000000" when "00000111000011011", -- t[3611] = 0
      "0000000" when "00000111000011100", -- t[3612] = 0
      "0000000" when "00000111000011101", -- t[3613] = 0
      "0000000" when "00000111000011110", -- t[3614] = 0
      "0000000" when "00000111000011111", -- t[3615] = 0
      "0000000" when "00000111000100000", -- t[3616] = 0
      "0000000" when "00000111000100001", -- t[3617] = 0
      "0000000" when "00000111000100010", -- t[3618] = 0
      "0000000" when "00000111000100011", -- t[3619] = 0
      "0000000" when "00000111000100100", -- t[3620] = 0
      "0000000" when "00000111000100101", -- t[3621] = 0
      "0000000" when "00000111000100110", -- t[3622] = 0
      "0000000" when "00000111000100111", -- t[3623] = 0
      "0000000" when "00000111000101000", -- t[3624] = 0
      "0000000" when "00000111000101001", -- t[3625] = 0
      "0000000" when "00000111000101010", -- t[3626] = 0
      "0000000" when "00000111000101011", -- t[3627] = 0
      "0000000" when "00000111000101100", -- t[3628] = 0
      "0000000" when "00000111000101101", -- t[3629] = 0
      "0000000" when "00000111000101110", -- t[3630] = 0
      "0000000" when "00000111000101111", -- t[3631] = 0
      "0000000" when "00000111000110000", -- t[3632] = 0
      "0000000" when "00000111000110001", -- t[3633] = 0
      "0000000" when "00000111000110010", -- t[3634] = 0
      "0000000" when "00000111000110011", -- t[3635] = 0
      "0000000" when "00000111000110100", -- t[3636] = 0
      "0000000" when "00000111000110101", -- t[3637] = 0
      "0000000" when "00000111000110110", -- t[3638] = 0
      "0000000" when "00000111000110111", -- t[3639] = 0
      "0000000" when "00000111000111000", -- t[3640] = 0
      "0000000" when "00000111000111001", -- t[3641] = 0
      "0000000" when "00000111000111010", -- t[3642] = 0
      "0000000" when "00000111000111011", -- t[3643] = 0
      "0000000" when "00000111000111100", -- t[3644] = 0
      "0000000" when "00000111000111101", -- t[3645] = 0
      "0000000" when "00000111000111110", -- t[3646] = 0
      "0000000" when "00000111000111111", -- t[3647] = 0
      "0000000" when "00000111001000000", -- t[3648] = 0
      "0000000" when "00000111001000001", -- t[3649] = 0
      "0000000" when "00000111001000010", -- t[3650] = 0
      "0000000" when "00000111001000011", -- t[3651] = 0
      "0000000" when "00000111001000100", -- t[3652] = 0
      "0000000" when "00000111001000101", -- t[3653] = 0
      "0000000" when "00000111001000110", -- t[3654] = 0
      "0000000" when "00000111001000111", -- t[3655] = 0
      "0000000" when "00000111001001000", -- t[3656] = 0
      "0000000" when "00000111001001001", -- t[3657] = 0
      "0000000" when "00000111001001010", -- t[3658] = 0
      "0000000" when "00000111001001011", -- t[3659] = 0
      "0000000" when "00000111001001100", -- t[3660] = 0
      "0000000" when "00000111001001101", -- t[3661] = 0
      "0000000" when "00000111001001110", -- t[3662] = 0
      "0000000" when "00000111001001111", -- t[3663] = 0
      "0000000" when "00000111001010000", -- t[3664] = 0
      "0000000" when "00000111001010001", -- t[3665] = 0
      "0000000" when "00000111001010010", -- t[3666] = 0
      "0000000" when "00000111001010011", -- t[3667] = 0
      "0000000" when "00000111001010100", -- t[3668] = 0
      "0000000" when "00000111001010101", -- t[3669] = 0
      "0000000" when "00000111001010110", -- t[3670] = 0
      "0000000" when "00000111001010111", -- t[3671] = 0
      "0000000" when "00000111001011000", -- t[3672] = 0
      "0000000" when "00000111001011001", -- t[3673] = 0
      "0000000" when "00000111001011010", -- t[3674] = 0
      "0000000" when "00000111001011011", -- t[3675] = 0
      "0000000" when "00000111001011100", -- t[3676] = 0
      "0000000" when "00000111001011101", -- t[3677] = 0
      "0000000" when "00000111001011110", -- t[3678] = 0
      "0000000" when "00000111001011111", -- t[3679] = 0
      "0000000" when "00000111001100000", -- t[3680] = 0
      "0000000" when "00000111001100001", -- t[3681] = 0
      "0000000" when "00000111001100010", -- t[3682] = 0
      "0000000" when "00000111001100011", -- t[3683] = 0
      "0000000" when "00000111001100100", -- t[3684] = 0
      "0000000" when "00000111001100101", -- t[3685] = 0
      "0000000" when "00000111001100110", -- t[3686] = 0
      "0000000" when "00000111001100111", -- t[3687] = 0
      "0000000" when "00000111001101000", -- t[3688] = 0
      "0000000" when "00000111001101001", -- t[3689] = 0
      "0000000" when "00000111001101010", -- t[3690] = 0
      "0000000" when "00000111001101011", -- t[3691] = 0
      "0000000" when "00000111001101100", -- t[3692] = 0
      "0000000" when "00000111001101101", -- t[3693] = 0
      "0000000" when "00000111001101110", -- t[3694] = 0
      "0000000" when "00000111001101111", -- t[3695] = 0
      "0000000" when "00000111001110000", -- t[3696] = 0
      "0000000" when "00000111001110001", -- t[3697] = 0
      "0000000" when "00000111001110010", -- t[3698] = 0
      "0000000" when "00000111001110011", -- t[3699] = 0
      "0000000" when "00000111001110100", -- t[3700] = 0
      "0000000" when "00000111001110101", -- t[3701] = 0
      "0000000" when "00000111001110110", -- t[3702] = 0
      "0000000" when "00000111001110111", -- t[3703] = 0
      "0000000" when "00000111001111000", -- t[3704] = 0
      "0000000" when "00000111001111001", -- t[3705] = 0
      "0000000" when "00000111001111010", -- t[3706] = 0
      "0000000" when "00000111001111011", -- t[3707] = 0
      "0000000" when "00000111001111100", -- t[3708] = 0
      "0000000" when "00000111001111101", -- t[3709] = 0
      "0000000" when "00000111001111110", -- t[3710] = 0
      "0000000" when "00000111001111111", -- t[3711] = 0
      "0000000" when "00000111010000000", -- t[3712] = 0
      "0000000" when "00000111010000001", -- t[3713] = 0
      "0000000" when "00000111010000010", -- t[3714] = 0
      "0000000" when "00000111010000011", -- t[3715] = 0
      "0000000" when "00000111010000100", -- t[3716] = 0
      "0000000" when "00000111010000101", -- t[3717] = 0
      "0000000" when "00000111010000110", -- t[3718] = 0
      "0000000" when "00000111010000111", -- t[3719] = 0
      "0000000" when "00000111010001000", -- t[3720] = 0
      "0000000" when "00000111010001001", -- t[3721] = 0
      "0000000" when "00000111010001010", -- t[3722] = 0
      "0000000" when "00000111010001011", -- t[3723] = 0
      "0000000" when "00000111010001100", -- t[3724] = 0
      "0000000" when "00000111010001101", -- t[3725] = 0
      "0000000" when "00000111010001110", -- t[3726] = 0
      "0000000" when "00000111010001111", -- t[3727] = 0
      "0000000" when "00000111010010000", -- t[3728] = 0
      "0000000" when "00000111010010001", -- t[3729] = 0
      "0000000" when "00000111010010010", -- t[3730] = 0
      "0000000" when "00000111010010011", -- t[3731] = 0
      "0000000" when "00000111010010100", -- t[3732] = 0
      "0000000" when "00000111010010101", -- t[3733] = 0
      "0000000" when "00000111010010110", -- t[3734] = 0
      "0000000" when "00000111010010111", -- t[3735] = 0
      "0000000" when "00000111010011000", -- t[3736] = 0
      "0000000" when "00000111010011001", -- t[3737] = 0
      "0000000" when "00000111010011010", -- t[3738] = 0
      "0000000" when "00000111010011011", -- t[3739] = 0
      "0000000" when "00000111010011100", -- t[3740] = 0
      "0000000" when "00000111010011101", -- t[3741] = 0
      "0000000" when "00000111010011110", -- t[3742] = 0
      "0000000" when "00000111010011111", -- t[3743] = 0
      "0000000" when "00000111010100000", -- t[3744] = 0
      "0000000" when "00000111010100001", -- t[3745] = 0
      "0000000" when "00000111010100010", -- t[3746] = 0
      "0000000" when "00000111010100011", -- t[3747] = 0
      "0000000" when "00000111010100100", -- t[3748] = 0
      "0000000" when "00000111010100101", -- t[3749] = 0
      "0000000" when "00000111010100110", -- t[3750] = 0
      "0000000" when "00000111010100111", -- t[3751] = 0
      "0000000" when "00000111010101000", -- t[3752] = 0
      "0000000" when "00000111010101001", -- t[3753] = 0
      "0000000" when "00000111010101010", -- t[3754] = 0
      "0000000" when "00000111010101011", -- t[3755] = 0
      "0000000" when "00000111010101100", -- t[3756] = 0
      "0000000" when "00000111010101101", -- t[3757] = 0
      "0000000" when "00000111010101110", -- t[3758] = 0
      "0000000" when "00000111010101111", -- t[3759] = 0
      "0000000" when "00000111010110000", -- t[3760] = 0
      "0000000" when "00000111010110001", -- t[3761] = 0
      "0000000" when "00000111010110010", -- t[3762] = 0
      "0000000" when "00000111010110011", -- t[3763] = 0
      "0000000" when "00000111010110100", -- t[3764] = 0
      "0000000" when "00000111010110101", -- t[3765] = 0
      "0000000" when "00000111010110110", -- t[3766] = 0
      "0000000" when "00000111010110111", -- t[3767] = 0
      "0000000" when "00000111010111000", -- t[3768] = 0
      "0000000" when "00000111010111001", -- t[3769] = 0
      "0000000" when "00000111010111010", -- t[3770] = 0
      "0000000" when "00000111010111011", -- t[3771] = 0
      "0000000" when "00000111010111100", -- t[3772] = 0
      "0000000" when "00000111010111101", -- t[3773] = 0
      "0000000" when "00000111010111110", -- t[3774] = 0
      "0000000" when "00000111010111111", -- t[3775] = 0
      "0000000" when "00000111011000000", -- t[3776] = 0
      "0000000" when "00000111011000001", -- t[3777] = 0
      "0000000" when "00000111011000010", -- t[3778] = 0
      "0000000" when "00000111011000011", -- t[3779] = 0
      "0000000" when "00000111011000100", -- t[3780] = 0
      "0000000" when "00000111011000101", -- t[3781] = 0
      "0000000" when "00000111011000110", -- t[3782] = 0
      "0000000" when "00000111011000111", -- t[3783] = 0
      "0000000" when "00000111011001000", -- t[3784] = 0
      "0000000" when "00000111011001001", -- t[3785] = 0
      "0000000" when "00000111011001010", -- t[3786] = 0
      "0000000" when "00000111011001011", -- t[3787] = 0
      "0000000" when "00000111011001100", -- t[3788] = 0
      "0000000" when "00000111011001101", -- t[3789] = 0
      "0000000" when "00000111011001110", -- t[3790] = 0
      "0000000" when "00000111011001111", -- t[3791] = 0
      "0000000" when "00000111011010000", -- t[3792] = 0
      "0000000" when "00000111011010001", -- t[3793] = 0
      "0000000" when "00000111011010010", -- t[3794] = 0
      "0000000" when "00000111011010011", -- t[3795] = 0
      "0000000" when "00000111011010100", -- t[3796] = 0
      "0000000" when "00000111011010101", -- t[3797] = 0
      "0000000" when "00000111011010110", -- t[3798] = 0
      "0000000" when "00000111011010111", -- t[3799] = 0
      "0000000" when "00000111011011000", -- t[3800] = 0
      "0000000" when "00000111011011001", -- t[3801] = 0
      "0000000" when "00000111011011010", -- t[3802] = 0
      "0000000" when "00000111011011011", -- t[3803] = 0
      "0000000" when "00000111011011100", -- t[3804] = 0
      "0000000" when "00000111011011101", -- t[3805] = 0
      "0000000" when "00000111011011110", -- t[3806] = 0
      "0000000" when "00000111011011111", -- t[3807] = 0
      "0000000" when "00000111011100000", -- t[3808] = 0
      "0000000" when "00000111011100001", -- t[3809] = 0
      "0000000" when "00000111011100010", -- t[3810] = 0
      "0000000" when "00000111011100011", -- t[3811] = 0
      "0000000" when "00000111011100100", -- t[3812] = 0
      "0000000" when "00000111011100101", -- t[3813] = 0
      "0000000" when "00000111011100110", -- t[3814] = 0
      "0000000" when "00000111011100111", -- t[3815] = 0
      "0000000" when "00000111011101000", -- t[3816] = 0
      "0000000" when "00000111011101001", -- t[3817] = 0
      "0000000" when "00000111011101010", -- t[3818] = 0
      "0000000" when "00000111011101011", -- t[3819] = 0
      "0000000" when "00000111011101100", -- t[3820] = 0
      "0000000" when "00000111011101101", -- t[3821] = 0
      "0000000" when "00000111011101110", -- t[3822] = 0
      "0000000" when "00000111011101111", -- t[3823] = 0
      "0000000" when "00000111011110000", -- t[3824] = 0
      "0000000" when "00000111011110001", -- t[3825] = 0
      "0000000" when "00000111011110010", -- t[3826] = 0
      "0000000" when "00000111011110011", -- t[3827] = 0
      "0000000" when "00000111011110100", -- t[3828] = 0
      "0000000" when "00000111011110101", -- t[3829] = 0
      "0000000" when "00000111011110110", -- t[3830] = 0
      "0000000" when "00000111011110111", -- t[3831] = 0
      "0000000" when "00000111011111000", -- t[3832] = 0
      "0000000" when "00000111011111001", -- t[3833] = 0
      "0000000" when "00000111011111010", -- t[3834] = 0
      "0000000" when "00000111011111011", -- t[3835] = 0
      "0000000" when "00000111011111100", -- t[3836] = 0
      "0000000" when "00000111011111101", -- t[3837] = 0
      "0000000" when "00000111011111110", -- t[3838] = 0
      "0000000" when "00000111011111111", -- t[3839] = 0
      "0000000" when "00000111100000000", -- t[3840] = 0
      "0000000" when "00000111100000001", -- t[3841] = 0
      "0000000" when "00000111100000010", -- t[3842] = 0
      "0000000" when "00000111100000011", -- t[3843] = 0
      "0000000" when "00000111100000100", -- t[3844] = 0
      "0000000" when "00000111100000101", -- t[3845] = 0
      "0000000" when "00000111100000110", -- t[3846] = 0
      "0000000" when "00000111100000111", -- t[3847] = 0
      "0000000" when "00000111100001000", -- t[3848] = 0
      "0000000" when "00000111100001001", -- t[3849] = 0
      "0000000" when "00000111100001010", -- t[3850] = 0
      "0000000" when "00000111100001011", -- t[3851] = 0
      "0000000" when "00000111100001100", -- t[3852] = 0
      "0000000" when "00000111100001101", -- t[3853] = 0
      "0000000" when "00000111100001110", -- t[3854] = 0
      "0000000" when "00000111100001111", -- t[3855] = 0
      "0000000" when "00000111100010000", -- t[3856] = 0
      "0000000" when "00000111100010001", -- t[3857] = 0
      "0000000" when "00000111100010010", -- t[3858] = 0
      "0000000" when "00000111100010011", -- t[3859] = 0
      "0000000" when "00000111100010100", -- t[3860] = 0
      "0000000" when "00000111100010101", -- t[3861] = 0
      "0000000" when "00000111100010110", -- t[3862] = 0
      "0000000" when "00000111100010111", -- t[3863] = 0
      "0000000" when "00000111100011000", -- t[3864] = 0
      "0000000" when "00000111100011001", -- t[3865] = 0
      "0000000" when "00000111100011010", -- t[3866] = 0
      "0000000" when "00000111100011011", -- t[3867] = 0
      "0000000" when "00000111100011100", -- t[3868] = 0
      "0000000" when "00000111100011101", -- t[3869] = 0
      "0000000" when "00000111100011110", -- t[3870] = 0
      "0000000" when "00000111100011111", -- t[3871] = 0
      "0000000" when "00000111100100000", -- t[3872] = 0
      "0000000" when "00000111100100001", -- t[3873] = 0
      "0000000" when "00000111100100010", -- t[3874] = 0
      "0000000" when "00000111100100011", -- t[3875] = 0
      "0000000" when "00000111100100100", -- t[3876] = 0
      "0000000" when "00000111100100101", -- t[3877] = 0
      "0000000" when "00000111100100110", -- t[3878] = 0
      "0000000" when "00000111100100111", -- t[3879] = 0
      "0000000" when "00000111100101000", -- t[3880] = 0
      "0000000" when "00000111100101001", -- t[3881] = 0
      "0000000" when "00000111100101010", -- t[3882] = 0
      "0000000" when "00000111100101011", -- t[3883] = 0
      "0000000" when "00000111100101100", -- t[3884] = 0
      "0000000" when "00000111100101101", -- t[3885] = 0
      "0000000" when "00000111100101110", -- t[3886] = 0
      "0000000" when "00000111100101111", -- t[3887] = 0
      "0000000" when "00000111100110000", -- t[3888] = 0
      "0000000" when "00000111100110001", -- t[3889] = 0
      "0000000" when "00000111100110010", -- t[3890] = 0
      "0000000" when "00000111100110011", -- t[3891] = 0
      "0000000" when "00000111100110100", -- t[3892] = 0
      "0000000" when "00000111100110101", -- t[3893] = 0
      "0000000" when "00000111100110110", -- t[3894] = 0
      "0000000" when "00000111100110111", -- t[3895] = 0
      "0000000" when "00000111100111000", -- t[3896] = 0
      "0000000" when "00000111100111001", -- t[3897] = 0
      "0000000" when "00000111100111010", -- t[3898] = 0
      "0000000" when "00000111100111011", -- t[3899] = 0
      "0000000" when "00000111100111100", -- t[3900] = 0
      "0000000" when "00000111100111101", -- t[3901] = 0
      "0000000" when "00000111100111110", -- t[3902] = 0
      "0000000" when "00000111100111111", -- t[3903] = 0
      "0000000" when "00000111101000000", -- t[3904] = 0
      "0000000" when "00000111101000001", -- t[3905] = 0
      "0000000" when "00000111101000010", -- t[3906] = 0
      "0000000" when "00000111101000011", -- t[3907] = 0
      "0000000" when "00000111101000100", -- t[3908] = 0
      "0000000" when "00000111101000101", -- t[3909] = 0
      "0000000" when "00000111101000110", -- t[3910] = 0
      "0000000" when "00000111101000111", -- t[3911] = 0
      "0000000" when "00000111101001000", -- t[3912] = 0
      "0000000" when "00000111101001001", -- t[3913] = 0
      "0000000" when "00000111101001010", -- t[3914] = 0
      "0000000" when "00000111101001011", -- t[3915] = 0
      "0000000" when "00000111101001100", -- t[3916] = 0
      "0000000" when "00000111101001101", -- t[3917] = 0
      "0000000" when "00000111101001110", -- t[3918] = 0
      "0000000" when "00000111101001111", -- t[3919] = 0
      "0000000" when "00000111101010000", -- t[3920] = 0
      "0000000" when "00000111101010001", -- t[3921] = 0
      "0000000" when "00000111101010010", -- t[3922] = 0
      "0000000" when "00000111101010011", -- t[3923] = 0
      "0000000" when "00000111101010100", -- t[3924] = 0
      "0000000" when "00000111101010101", -- t[3925] = 0
      "0000000" when "00000111101010110", -- t[3926] = 0
      "0000000" when "00000111101010111", -- t[3927] = 0
      "0000000" when "00000111101011000", -- t[3928] = 0
      "0000000" when "00000111101011001", -- t[3929] = 0
      "0000000" when "00000111101011010", -- t[3930] = 0
      "0000000" when "00000111101011011", -- t[3931] = 0
      "0000000" when "00000111101011100", -- t[3932] = 0
      "0000000" when "00000111101011101", -- t[3933] = 0
      "0000000" when "00000111101011110", -- t[3934] = 0
      "0000000" when "00000111101011111", -- t[3935] = 0
      "0000000" when "00000111101100000", -- t[3936] = 0
      "0000000" when "00000111101100001", -- t[3937] = 0
      "0000000" when "00000111101100010", -- t[3938] = 0
      "0000000" when "00000111101100011", -- t[3939] = 0
      "0000000" when "00000111101100100", -- t[3940] = 0
      "0000000" when "00000111101100101", -- t[3941] = 0
      "0000000" when "00000111101100110", -- t[3942] = 0
      "0000000" when "00000111101100111", -- t[3943] = 0
      "0000000" when "00000111101101000", -- t[3944] = 0
      "0000000" when "00000111101101001", -- t[3945] = 0
      "0000000" when "00000111101101010", -- t[3946] = 0
      "0000000" when "00000111101101011", -- t[3947] = 0
      "0000000" when "00000111101101100", -- t[3948] = 0
      "0000000" when "00000111101101101", -- t[3949] = 0
      "0000000" when "00000111101101110", -- t[3950] = 0
      "0000000" when "00000111101101111", -- t[3951] = 0
      "0000000" when "00000111101110000", -- t[3952] = 0
      "0000000" when "00000111101110001", -- t[3953] = 0
      "0000000" when "00000111101110010", -- t[3954] = 0
      "0000000" when "00000111101110011", -- t[3955] = 0
      "0000000" when "00000111101110100", -- t[3956] = 0
      "0000000" when "00000111101110101", -- t[3957] = 0
      "0000000" when "00000111101110110", -- t[3958] = 0
      "0000000" when "00000111101110111", -- t[3959] = 0
      "0000000" when "00000111101111000", -- t[3960] = 0
      "0000000" when "00000111101111001", -- t[3961] = 0
      "0000000" when "00000111101111010", -- t[3962] = 0
      "0000000" when "00000111101111011", -- t[3963] = 0
      "0000000" when "00000111101111100", -- t[3964] = 0
      "0000000" when "00000111101111101", -- t[3965] = 0
      "0000000" when "00000111101111110", -- t[3966] = 0
      "0000000" when "00000111101111111", -- t[3967] = 0
      "0000000" when "00000111110000000", -- t[3968] = 0
      "0000000" when "00000111110000001", -- t[3969] = 0
      "0000000" when "00000111110000010", -- t[3970] = 0
      "0000000" when "00000111110000011", -- t[3971] = 0
      "0000000" when "00000111110000100", -- t[3972] = 0
      "0000000" when "00000111110000101", -- t[3973] = 0
      "0000000" when "00000111110000110", -- t[3974] = 0
      "0000000" when "00000111110000111", -- t[3975] = 0
      "0000000" when "00000111110001000", -- t[3976] = 0
      "0000000" when "00000111110001001", -- t[3977] = 0
      "0000000" when "00000111110001010", -- t[3978] = 0
      "0000000" when "00000111110001011", -- t[3979] = 0
      "0000000" when "00000111110001100", -- t[3980] = 0
      "0000000" when "00000111110001101", -- t[3981] = 0
      "0000000" when "00000111110001110", -- t[3982] = 0
      "0000000" when "00000111110001111", -- t[3983] = 0
      "0000000" when "00000111110010000", -- t[3984] = 0
      "0000000" when "00000111110010001", -- t[3985] = 0
      "0000000" when "00000111110010010", -- t[3986] = 0
      "0000000" when "00000111110010011", -- t[3987] = 0
      "0000000" when "00000111110010100", -- t[3988] = 0
      "0000000" when "00000111110010101", -- t[3989] = 0
      "0000000" when "00000111110010110", -- t[3990] = 0
      "0000000" when "00000111110010111", -- t[3991] = 0
      "0000000" when "00000111110011000", -- t[3992] = 0
      "0000000" when "00000111110011001", -- t[3993] = 0
      "0000000" when "00000111110011010", -- t[3994] = 0
      "0000000" when "00000111110011011", -- t[3995] = 0
      "0000000" when "00000111110011100", -- t[3996] = 0
      "0000000" when "00000111110011101", -- t[3997] = 0
      "0000000" when "00000111110011110", -- t[3998] = 0
      "0000000" when "00000111110011111", -- t[3999] = 0
      "0000000" when "00000111110100000", -- t[4000] = 0
      "0000000" when "00000111110100001", -- t[4001] = 0
      "0000000" when "00000111110100010", -- t[4002] = 0
      "0000000" when "00000111110100011", -- t[4003] = 0
      "0000000" when "00000111110100100", -- t[4004] = 0
      "0000000" when "00000111110100101", -- t[4005] = 0
      "0000000" when "00000111110100110", -- t[4006] = 0
      "0000000" when "00000111110100111", -- t[4007] = 0
      "0000000" when "00000111110101000", -- t[4008] = 0
      "0000000" when "00000111110101001", -- t[4009] = 0
      "0000000" when "00000111110101010", -- t[4010] = 0
      "0000000" when "00000111110101011", -- t[4011] = 0
      "0000000" when "00000111110101100", -- t[4012] = 0
      "0000000" when "00000111110101101", -- t[4013] = 0
      "0000000" when "00000111110101110", -- t[4014] = 0
      "0000000" when "00000111110101111", -- t[4015] = 0
      "0000000" when "00000111110110000", -- t[4016] = 0
      "0000000" when "00000111110110001", -- t[4017] = 0
      "0000000" when "00000111110110010", -- t[4018] = 0
      "0000000" when "00000111110110011", -- t[4019] = 0
      "0000000" when "00000111110110100", -- t[4020] = 0
      "0000000" when "00000111110110101", -- t[4021] = 0
      "0000000" when "00000111110110110", -- t[4022] = 0
      "0000000" when "00000111110110111", -- t[4023] = 0
      "0000000" when "00000111110111000", -- t[4024] = 0
      "0000000" when "00000111110111001", -- t[4025] = 0
      "0000000" when "00000111110111010", -- t[4026] = 0
      "0000000" when "00000111110111011", -- t[4027] = 0
      "0000000" when "00000111110111100", -- t[4028] = 0
      "0000000" when "00000111110111101", -- t[4029] = 0
      "0000000" when "00000111110111110", -- t[4030] = 0
      "0000000" when "00000111110111111", -- t[4031] = 0
      "0000000" when "00000111111000000", -- t[4032] = 0
      "0000000" when "00000111111000001", -- t[4033] = 0
      "0000000" when "00000111111000010", -- t[4034] = 0
      "0000000" when "00000111111000011", -- t[4035] = 0
      "0000000" when "00000111111000100", -- t[4036] = 0
      "0000000" when "00000111111000101", -- t[4037] = 0
      "0000000" when "00000111111000110", -- t[4038] = 0
      "0000000" when "00000111111000111", -- t[4039] = 0
      "0000000" when "00000111111001000", -- t[4040] = 0
      "0000000" when "00000111111001001", -- t[4041] = 0
      "0000000" when "00000111111001010", -- t[4042] = 0
      "0000000" when "00000111111001011", -- t[4043] = 0
      "0000000" when "00000111111001100", -- t[4044] = 0
      "0000000" when "00000111111001101", -- t[4045] = 0
      "0000000" when "00000111111001110", -- t[4046] = 0
      "0000000" when "00000111111001111", -- t[4047] = 0
      "0000000" when "00000111111010000", -- t[4048] = 0
      "0000000" when "00000111111010001", -- t[4049] = 0
      "0000000" when "00000111111010010", -- t[4050] = 0
      "0000000" when "00000111111010011", -- t[4051] = 0
      "0000000" when "00000111111010100", -- t[4052] = 0
      "0000000" when "00000111111010101", -- t[4053] = 0
      "0000000" when "00000111111010110", -- t[4054] = 0
      "0000000" when "00000111111010111", -- t[4055] = 0
      "0000000" when "00000111111011000", -- t[4056] = 0
      "0000000" when "00000111111011001", -- t[4057] = 0
      "0000000" when "00000111111011010", -- t[4058] = 0
      "0000000" when "00000111111011011", -- t[4059] = 0
      "0000000" when "00000111111011100", -- t[4060] = 0
      "0000000" when "00000111111011101", -- t[4061] = 0
      "0000000" when "00000111111011110", -- t[4062] = 0
      "0000000" when "00000111111011111", -- t[4063] = 0
      "0000000" when "00000111111100000", -- t[4064] = 0
      "0000000" when "00000111111100001", -- t[4065] = 0
      "0000000" when "00000111111100010", -- t[4066] = 0
      "0000000" when "00000111111100011", -- t[4067] = 0
      "0000000" when "00000111111100100", -- t[4068] = 0
      "0000000" when "00000111111100101", -- t[4069] = 0
      "0000000" when "00000111111100110", -- t[4070] = 0
      "0000000" when "00000111111100111", -- t[4071] = 0
      "0000000" when "00000111111101000", -- t[4072] = 0
      "0000000" when "00000111111101001", -- t[4073] = 0
      "0000000" when "00000111111101010", -- t[4074] = 0
      "0000000" when "00000111111101011", -- t[4075] = 0
      "0000000" when "00000111111101100", -- t[4076] = 0
      "0000000" when "00000111111101101", -- t[4077] = 0
      "0000000" when "00000111111101110", -- t[4078] = 0
      "0000000" when "00000111111101111", -- t[4079] = 0
      "0000000" when "00000111111110000", -- t[4080] = 0
      "0000000" when "00000111111110001", -- t[4081] = 0
      "0000000" when "00000111111110010", -- t[4082] = 0
      "0000000" when "00000111111110011", -- t[4083] = 0
      "0000000" when "00000111111110100", -- t[4084] = 0
      "0000000" when "00000111111110101", -- t[4085] = 0
      "0000000" when "00000111111110110", -- t[4086] = 0
      "0000000" when "00000111111110111", -- t[4087] = 0
      "0000000" when "00000111111111000", -- t[4088] = 0
      "0000000" when "00000111111111001", -- t[4089] = 0
      "0000000" when "00000111111111010", -- t[4090] = 0
      "0000000" when "00000111111111011", -- t[4091] = 0
      "0000000" when "00000111111111100", -- t[4092] = 0
      "0000000" when "00000111111111101", -- t[4093] = 0
      "0000000" when "00000111111111110", -- t[4094] = 0
      "0000000" when "00000111111111111", -- t[4095] = 0
      "0000000" when "00001000000000000", -- t[4096] = 0
      "0000000" when "00001000000000001", -- t[4097] = 0
      "0000000" when "00001000000000010", -- t[4098] = 0
      "0000000" when "00001000000000011", -- t[4099] = 0
      "0000000" when "00001000000000100", -- t[4100] = 0
      "0000000" when "00001000000000101", -- t[4101] = 0
      "0000000" when "00001000000000110", -- t[4102] = 0
      "0000000" when "00001000000000111", -- t[4103] = 0
      "0000000" when "00001000000001000", -- t[4104] = 0
      "0000000" when "00001000000001001", -- t[4105] = 0
      "0000000" when "00001000000001010", -- t[4106] = 0
      "0000000" when "00001000000001011", -- t[4107] = 0
      "0000000" when "00001000000001100", -- t[4108] = 0
      "0000000" when "00001000000001101", -- t[4109] = 0
      "0000000" when "00001000000001110", -- t[4110] = 0
      "0000000" when "00001000000001111", -- t[4111] = 0
      "0000000" when "00001000000010000", -- t[4112] = 0
      "0000000" when "00001000000010001", -- t[4113] = 0
      "0000000" when "00001000000010010", -- t[4114] = 0
      "0000000" when "00001000000010011", -- t[4115] = 0
      "0000000" when "00001000000010100", -- t[4116] = 0
      "0000000" when "00001000000010101", -- t[4117] = 0
      "0000000" when "00001000000010110", -- t[4118] = 0
      "0000000" when "00001000000010111", -- t[4119] = 0
      "0000000" when "00001000000011000", -- t[4120] = 0
      "0000000" when "00001000000011001", -- t[4121] = 0
      "0000000" when "00001000000011010", -- t[4122] = 0
      "0000000" when "00001000000011011", -- t[4123] = 0
      "0000000" when "00001000000011100", -- t[4124] = 0
      "0000000" when "00001000000011101", -- t[4125] = 0
      "0000000" when "00001000000011110", -- t[4126] = 0
      "0000000" when "00001000000011111", -- t[4127] = 0
      "0000000" when "00001000000100000", -- t[4128] = 0
      "0000000" when "00001000000100001", -- t[4129] = 0
      "0000000" when "00001000000100010", -- t[4130] = 0
      "0000000" when "00001000000100011", -- t[4131] = 0
      "0000000" when "00001000000100100", -- t[4132] = 0
      "0000000" when "00001000000100101", -- t[4133] = 0
      "0000000" when "00001000000100110", -- t[4134] = 0
      "0000000" when "00001000000100111", -- t[4135] = 0
      "0000000" when "00001000000101000", -- t[4136] = 0
      "0000000" when "00001000000101001", -- t[4137] = 0
      "0000000" when "00001000000101010", -- t[4138] = 0
      "0000000" when "00001000000101011", -- t[4139] = 0
      "0000000" when "00001000000101100", -- t[4140] = 0
      "0000000" when "00001000000101101", -- t[4141] = 0
      "0000000" when "00001000000101110", -- t[4142] = 0
      "0000000" when "00001000000101111", -- t[4143] = 0
      "0000000" when "00001000000110000", -- t[4144] = 0
      "0000000" when "00001000000110001", -- t[4145] = 0
      "0000000" when "00001000000110010", -- t[4146] = 0
      "0000000" when "00001000000110011", -- t[4147] = 0
      "0000000" when "00001000000110100", -- t[4148] = 0
      "0000000" when "00001000000110101", -- t[4149] = 0
      "0000000" when "00001000000110110", -- t[4150] = 0
      "0000000" when "00001000000110111", -- t[4151] = 0
      "0000000" when "00001000000111000", -- t[4152] = 0
      "0000000" when "00001000000111001", -- t[4153] = 0
      "0000000" when "00001000000111010", -- t[4154] = 0
      "0000000" when "00001000000111011", -- t[4155] = 0
      "0000000" when "00001000000111100", -- t[4156] = 0
      "0000000" when "00001000000111101", -- t[4157] = 0
      "0000000" when "00001000000111110", -- t[4158] = 0
      "0000000" when "00001000000111111", -- t[4159] = 0
      "0000000" when "00001000001000000", -- t[4160] = 0
      "0000000" when "00001000001000001", -- t[4161] = 0
      "0000000" when "00001000001000010", -- t[4162] = 0
      "0000000" when "00001000001000011", -- t[4163] = 0
      "0000000" when "00001000001000100", -- t[4164] = 0
      "0000000" when "00001000001000101", -- t[4165] = 0
      "0000000" when "00001000001000110", -- t[4166] = 0
      "0000000" when "00001000001000111", -- t[4167] = 0
      "0000000" when "00001000001001000", -- t[4168] = 0
      "0000000" when "00001000001001001", -- t[4169] = 0
      "0000000" when "00001000001001010", -- t[4170] = 0
      "0000000" when "00001000001001011", -- t[4171] = 0
      "0000000" when "00001000001001100", -- t[4172] = 0
      "0000000" when "00001000001001101", -- t[4173] = 0
      "0000000" when "00001000001001110", -- t[4174] = 0
      "0000000" when "00001000001001111", -- t[4175] = 0
      "0000000" when "00001000001010000", -- t[4176] = 0
      "0000000" when "00001000001010001", -- t[4177] = 0
      "0000000" when "00001000001010010", -- t[4178] = 0
      "0000000" when "00001000001010011", -- t[4179] = 0
      "0000000" when "00001000001010100", -- t[4180] = 0
      "0000000" when "00001000001010101", -- t[4181] = 0
      "0000000" when "00001000001010110", -- t[4182] = 0
      "0000000" when "00001000001010111", -- t[4183] = 0
      "0000000" when "00001000001011000", -- t[4184] = 0
      "0000000" when "00001000001011001", -- t[4185] = 0
      "0000000" when "00001000001011010", -- t[4186] = 0
      "0000000" when "00001000001011011", -- t[4187] = 0
      "0000000" when "00001000001011100", -- t[4188] = 0
      "0000000" when "00001000001011101", -- t[4189] = 0
      "0000000" when "00001000001011110", -- t[4190] = 0
      "0000000" when "00001000001011111", -- t[4191] = 0
      "0000000" when "00001000001100000", -- t[4192] = 0
      "0000000" when "00001000001100001", -- t[4193] = 0
      "0000000" when "00001000001100010", -- t[4194] = 0
      "0000000" when "00001000001100011", -- t[4195] = 0
      "0000000" when "00001000001100100", -- t[4196] = 0
      "0000000" when "00001000001100101", -- t[4197] = 0
      "0000000" when "00001000001100110", -- t[4198] = 0
      "0000000" when "00001000001100111", -- t[4199] = 0
      "0000000" when "00001000001101000", -- t[4200] = 0
      "0000000" when "00001000001101001", -- t[4201] = 0
      "0000000" when "00001000001101010", -- t[4202] = 0
      "0000000" when "00001000001101011", -- t[4203] = 0
      "0000000" when "00001000001101100", -- t[4204] = 0
      "0000000" when "00001000001101101", -- t[4205] = 0
      "0000000" when "00001000001101110", -- t[4206] = 0
      "0000000" when "00001000001101111", -- t[4207] = 0
      "0000000" when "00001000001110000", -- t[4208] = 0
      "0000000" when "00001000001110001", -- t[4209] = 0
      "0000000" when "00001000001110010", -- t[4210] = 0
      "0000000" when "00001000001110011", -- t[4211] = 0
      "0000000" when "00001000001110100", -- t[4212] = 0
      "0000000" when "00001000001110101", -- t[4213] = 0
      "0000000" when "00001000001110110", -- t[4214] = 0
      "0000000" when "00001000001110111", -- t[4215] = 0
      "0000000" when "00001000001111000", -- t[4216] = 0
      "0000000" when "00001000001111001", -- t[4217] = 0
      "0000000" when "00001000001111010", -- t[4218] = 0
      "0000000" when "00001000001111011", -- t[4219] = 0
      "0000000" when "00001000001111100", -- t[4220] = 0
      "0000000" when "00001000001111101", -- t[4221] = 0
      "0000000" when "00001000001111110", -- t[4222] = 0
      "0000000" when "00001000001111111", -- t[4223] = 0
      "0000000" when "00001000010000000", -- t[4224] = 0
      "0000000" when "00001000010000001", -- t[4225] = 0
      "0000000" when "00001000010000010", -- t[4226] = 0
      "0000000" when "00001000010000011", -- t[4227] = 0
      "0000000" when "00001000010000100", -- t[4228] = 0
      "0000000" when "00001000010000101", -- t[4229] = 0
      "0000000" when "00001000010000110", -- t[4230] = 0
      "0000000" when "00001000010000111", -- t[4231] = 0
      "0000000" when "00001000010001000", -- t[4232] = 0
      "0000000" when "00001000010001001", -- t[4233] = 0
      "0000000" when "00001000010001010", -- t[4234] = 0
      "0000000" when "00001000010001011", -- t[4235] = 0
      "0000000" when "00001000010001100", -- t[4236] = 0
      "0000000" when "00001000010001101", -- t[4237] = 0
      "0000000" when "00001000010001110", -- t[4238] = 0
      "0000000" when "00001000010001111", -- t[4239] = 0
      "0000000" when "00001000010010000", -- t[4240] = 0
      "0000000" when "00001000010010001", -- t[4241] = 0
      "0000000" when "00001000010010010", -- t[4242] = 0
      "0000000" when "00001000010010011", -- t[4243] = 0
      "0000000" when "00001000010010100", -- t[4244] = 0
      "0000000" when "00001000010010101", -- t[4245] = 0
      "0000000" when "00001000010010110", -- t[4246] = 0
      "0000000" when "00001000010010111", -- t[4247] = 0
      "0000000" when "00001000010011000", -- t[4248] = 0
      "0000000" when "00001000010011001", -- t[4249] = 0
      "0000000" when "00001000010011010", -- t[4250] = 0
      "0000000" when "00001000010011011", -- t[4251] = 0
      "0000000" when "00001000010011100", -- t[4252] = 0
      "0000000" when "00001000010011101", -- t[4253] = 0
      "0000000" when "00001000010011110", -- t[4254] = 0
      "0000000" when "00001000010011111", -- t[4255] = 0
      "0000000" when "00001000010100000", -- t[4256] = 0
      "0000000" when "00001000010100001", -- t[4257] = 0
      "0000000" when "00001000010100010", -- t[4258] = 0
      "0000000" when "00001000010100011", -- t[4259] = 0
      "0000000" when "00001000010100100", -- t[4260] = 0
      "0000000" when "00001000010100101", -- t[4261] = 0
      "0000000" when "00001000010100110", -- t[4262] = 0
      "0000000" when "00001000010100111", -- t[4263] = 0
      "0000000" when "00001000010101000", -- t[4264] = 0
      "0000000" when "00001000010101001", -- t[4265] = 0
      "0000000" when "00001000010101010", -- t[4266] = 0
      "0000000" when "00001000010101011", -- t[4267] = 0
      "0000000" when "00001000010101100", -- t[4268] = 0
      "0000000" when "00001000010101101", -- t[4269] = 0
      "0000000" when "00001000010101110", -- t[4270] = 0
      "0000000" when "00001000010101111", -- t[4271] = 0
      "0000000" when "00001000010110000", -- t[4272] = 0
      "0000000" when "00001000010110001", -- t[4273] = 0
      "0000000" when "00001000010110010", -- t[4274] = 0
      "0000000" when "00001000010110011", -- t[4275] = 0
      "0000000" when "00001000010110100", -- t[4276] = 0
      "0000000" when "00001000010110101", -- t[4277] = 0
      "0000000" when "00001000010110110", -- t[4278] = 0
      "0000000" when "00001000010110111", -- t[4279] = 0
      "0000000" when "00001000010111000", -- t[4280] = 0
      "0000000" when "00001000010111001", -- t[4281] = 0
      "0000000" when "00001000010111010", -- t[4282] = 0
      "0000000" when "00001000010111011", -- t[4283] = 0
      "0000000" when "00001000010111100", -- t[4284] = 0
      "0000000" when "00001000010111101", -- t[4285] = 0
      "0000000" when "00001000010111110", -- t[4286] = 0
      "0000000" when "00001000010111111", -- t[4287] = 0
      "0000000" when "00001000011000000", -- t[4288] = 0
      "0000000" when "00001000011000001", -- t[4289] = 0
      "0000000" when "00001000011000010", -- t[4290] = 0
      "0000000" when "00001000011000011", -- t[4291] = 0
      "0000000" when "00001000011000100", -- t[4292] = 0
      "0000000" when "00001000011000101", -- t[4293] = 0
      "0000000" when "00001000011000110", -- t[4294] = 0
      "0000000" when "00001000011000111", -- t[4295] = 0
      "0000000" when "00001000011001000", -- t[4296] = 0
      "0000000" when "00001000011001001", -- t[4297] = 0
      "0000000" when "00001000011001010", -- t[4298] = 0
      "0000000" when "00001000011001011", -- t[4299] = 0
      "0000000" when "00001000011001100", -- t[4300] = 0
      "0000000" when "00001000011001101", -- t[4301] = 0
      "0000000" when "00001000011001110", -- t[4302] = 0
      "0000000" when "00001000011001111", -- t[4303] = 0
      "0000000" when "00001000011010000", -- t[4304] = 0
      "0000000" when "00001000011010001", -- t[4305] = 0
      "0000000" when "00001000011010010", -- t[4306] = 0
      "0000000" when "00001000011010011", -- t[4307] = 0
      "0000000" when "00001000011010100", -- t[4308] = 0
      "0000000" when "00001000011010101", -- t[4309] = 0
      "0000000" when "00001000011010110", -- t[4310] = 0
      "0000000" when "00001000011010111", -- t[4311] = 0
      "0000000" when "00001000011011000", -- t[4312] = 0
      "0000000" when "00001000011011001", -- t[4313] = 0
      "0000000" when "00001000011011010", -- t[4314] = 0
      "0000000" when "00001000011011011", -- t[4315] = 0
      "0000000" when "00001000011011100", -- t[4316] = 0
      "0000000" when "00001000011011101", -- t[4317] = 0
      "0000000" when "00001000011011110", -- t[4318] = 0
      "0000000" when "00001000011011111", -- t[4319] = 0
      "0000000" when "00001000011100000", -- t[4320] = 0
      "0000000" when "00001000011100001", -- t[4321] = 0
      "0000000" when "00001000011100010", -- t[4322] = 0
      "0000000" when "00001000011100011", -- t[4323] = 0
      "0000000" when "00001000011100100", -- t[4324] = 0
      "0000000" when "00001000011100101", -- t[4325] = 0
      "0000000" when "00001000011100110", -- t[4326] = 0
      "0000000" when "00001000011100111", -- t[4327] = 0
      "0000000" when "00001000011101000", -- t[4328] = 0
      "0000000" when "00001000011101001", -- t[4329] = 0
      "0000000" when "00001000011101010", -- t[4330] = 0
      "0000000" when "00001000011101011", -- t[4331] = 0
      "0000000" when "00001000011101100", -- t[4332] = 0
      "0000000" when "00001000011101101", -- t[4333] = 0
      "0000000" when "00001000011101110", -- t[4334] = 0
      "0000000" when "00001000011101111", -- t[4335] = 0
      "0000000" when "00001000011110000", -- t[4336] = 0
      "0000000" when "00001000011110001", -- t[4337] = 0
      "0000000" when "00001000011110010", -- t[4338] = 0
      "0000000" when "00001000011110011", -- t[4339] = 0
      "0000000" when "00001000011110100", -- t[4340] = 0
      "0000000" when "00001000011110101", -- t[4341] = 0
      "0000000" when "00001000011110110", -- t[4342] = 0
      "0000000" when "00001000011110111", -- t[4343] = 0
      "0000000" when "00001000011111000", -- t[4344] = 0
      "0000000" when "00001000011111001", -- t[4345] = 0
      "0000000" when "00001000011111010", -- t[4346] = 0
      "0000000" when "00001000011111011", -- t[4347] = 0
      "0000000" when "00001000011111100", -- t[4348] = 0
      "0000000" when "00001000011111101", -- t[4349] = 0
      "0000000" when "00001000011111110", -- t[4350] = 0
      "0000000" when "00001000011111111", -- t[4351] = 0
      "0000000" when "00001000100000000", -- t[4352] = 0
      "0000000" when "00001000100000001", -- t[4353] = 0
      "0000000" when "00001000100000010", -- t[4354] = 0
      "0000000" when "00001000100000011", -- t[4355] = 0
      "0000000" when "00001000100000100", -- t[4356] = 0
      "0000000" when "00001000100000101", -- t[4357] = 0
      "0000000" when "00001000100000110", -- t[4358] = 0
      "0000000" when "00001000100000111", -- t[4359] = 0
      "0000000" when "00001000100001000", -- t[4360] = 0
      "0000000" when "00001000100001001", -- t[4361] = 0
      "0000000" when "00001000100001010", -- t[4362] = 0
      "0000000" when "00001000100001011", -- t[4363] = 0
      "0000000" when "00001000100001100", -- t[4364] = 0
      "0000000" when "00001000100001101", -- t[4365] = 0
      "0000000" when "00001000100001110", -- t[4366] = 0
      "0000000" when "00001000100001111", -- t[4367] = 0
      "0000000" when "00001000100010000", -- t[4368] = 0
      "0000000" when "00001000100010001", -- t[4369] = 0
      "0000000" when "00001000100010010", -- t[4370] = 0
      "0000000" when "00001000100010011", -- t[4371] = 0
      "0000000" when "00001000100010100", -- t[4372] = 0
      "0000000" when "00001000100010101", -- t[4373] = 0
      "0000000" when "00001000100010110", -- t[4374] = 0
      "0000000" when "00001000100010111", -- t[4375] = 0
      "0000000" when "00001000100011000", -- t[4376] = 0
      "0000000" when "00001000100011001", -- t[4377] = 0
      "0000000" when "00001000100011010", -- t[4378] = 0
      "0000000" when "00001000100011011", -- t[4379] = 0
      "0000000" when "00001000100011100", -- t[4380] = 0
      "0000000" when "00001000100011101", -- t[4381] = 0
      "0000000" when "00001000100011110", -- t[4382] = 0
      "0000000" when "00001000100011111", -- t[4383] = 0
      "0000000" when "00001000100100000", -- t[4384] = 0
      "0000000" when "00001000100100001", -- t[4385] = 0
      "0000000" when "00001000100100010", -- t[4386] = 0
      "0000000" when "00001000100100011", -- t[4387] = 0
      "0000000" when "00001000100100100", -- t[4388] = 0
      "0000000" when "00001000100100101", -- t[4389] = 0
      "0000000" when "00001000100100110", -- t[4390] = 0
      "0000000" when "00001000100100111", -- t[4391] = 0
      "0000000" when "00001000100101000", -- t[4392] = 0
      "0000000" when "00001000100101001", -- t[4393] = 0
      "0000000" when "00001000100101010", -- t[4394] = 0
      "0000000" when "00001000100101011", -- t[4395] = 0
      "0000000" when "00001000100101100", -- t[4396] = 0
      "0000000" when "00001000100101101", -- t[4397] = 0
      "0000000" when "00001000100101110", -- t[4398] = 0
      "0000000" when "00001000100101111", -- t[4399] = 0
      "0000000" when "00001000100110000", -- t[4400] = 0
      "0000000" when "00001000100110001", -- t[4401] = 0
      "0000000" when "00001000100110010", -- t[4402] = 0
      "0000000" when "00001000100110011", -- t[4403] = 0
      "0000000" when "00001000100110100", -- t[4404] = 0
      "0000000" when "00001000100110101", -- t[4405] = 0
      "0000000" when "00001000100110110", -- t[4406] = 0
      "0000000" when "00001000100110111", -- t[4407] = 0
      "0000000" when "00001000100111000", -- t[4408] = 0
      "0000000" when "00001000100111001", -- t[4409] = 0
      "0000000" when "00001000100111010", -- t[4410] = 0
      "0000000" when "00001000100111011", -- t[4411] = 0
      "0000000" when "00001000100111100", -- t[4412] = 0
      "0000000" when "00001000100111101", -- t[4413] = 0
      "0000000" when "00001000100111110", -- t[4414] = 0
      "0000000" when "00001000100111111", -- t[4415] = 0
      "0000000" when "00001000101000000", -- t[4416] = 0
      "0000000" when "00001000101000001", -- t[4417] = 0
      "0000000" when "00001000101000010", -- t[4418] = 0
      "0000000" when "00001000101000011", -- t[4419] = 0
      "0000000" when "00001000101000100", -- t[4420] = 0
      "0000000" when "00001000101000101", -- t[4421] = 0
      "0000000" when "00001000101000110", -- t[4422] = 0
      "0000000" when "00001000101000111", -- t[4423] = 0
      "0000000" when "00001000101001000", -- t[4424] = 0
      "0000000" when "00001000101001001", -- t[4425] = 0
      "0000000" when "00001000101001010", -- t[4426] = 0
      "0000000" when "00001000101001011", -- t[4427] = 0
      "0000000" when "00001000101001100", -- t[4428] = 0
      "0000000" when "00001000101001101", -- t[4429] = 0
      "0000000" when "00001000101001110", -- t[4430] = 0
      "0000000" when "00001000101001111", -- t[4431] = 0
      "0000000" when "00001000101010000", -- t[4432] = 0
      "0000000" when "00001000101010001", -- t[4433] = 0
      "0000000" when "00001000101010010", -- t[4434] = 0
      "0000000" when "00001000101010011", -- t[4435] = 0
      "0000000" when "00001000101010100", -- t[4436] = 0
      "0000000" when "00001000101010101", -- t[4437] = 0
      "0000000" when "00001000101010110", -- t[4438] = 0
      "0000000" when "00001000101010111", -- t[4439] = 0
      "0000000" when "00001000101011000", -- t[4440] = 0
      "0000000" when "00001000101011001", -- t[4441] = 0
      "0000000" when "00001000101011010", -- t[4442] = 0
      "0000000" when "00001000101011011", -- t[4443] = 0
      "0000000" when "00001000101011100", -- t[4444] = 0
      "0000000" when "00001000101011101", -- t[4445] = 0
      "0000000" when "00001000101011110", -- t[4446] = 0
      "0000000" when "00001000101011111", -- t[4447] = 0
      "0000000" when "00001000101100000", -- t[4448] = 0
      "0000000" when "00001000101100001", -- t[4449] = 0
      "0000000" when "00001000101100010", -- t[4450] = 0
      "0000000" when "00001000101100011", -- t[4451] = 0
      "0000000" when "00001000101100100", -- t[4452] = 0
      "0000000" when "00001000101100101", -- t[4453] = 0
      "0000000" when "00001000101100110", -- t[4454] = 0
      "0000000" when "00001000101100111", -- t[4455] = 0
      "0000000" when "00001000101101000", -- t[4456] = 0
      "0000000" when "00001000101101001", -- t[4457] = 0
      "0000000" when "00001000101101010", -- t[4458] = 0
      "0000000" when "00001000101101011", -- t[4459] = 0
      "0000000" when "00001000101101100", -- t[4460] = 0
      "0000000" when "00001000101101101", -- t[4461] = 0
      "0000000" when "00001000101101110", -- t[4462] = 0
      "0000000" when "00001000101101111", -- t[4463] = 0
      "0000000" when "00001000101110000", -- t[4464] = 0
      "0000000" when "00001000101110001", -- t[4465] = 0
      "0000000" when "00001000101110010", -- t[4466] = 0
      "0000000" when "00001000101110011", -- t[4467] = 0
      "0000000" when "00001000101110100", -- t[4468] = 0
      "0000000" when "00001000101110101", -- t[4469] = 0
      "0000000" when "00001000101110110", -- t[4470] = 0
      "0000000" when "00001000101110111", -- t[4471] = 0
      "0000000" when "00001000101111000", -- t[4472] = 0
      "0000000" when "00001000101111001", -- t[4473] = 0
      "0000000" when "00001000101111010", -- t[4474] = 0
      "0000000" when "00001000101111011", -- t[4475] = 0
      "0000000" when "00001000101111100", -- t[4476] = 0
      "0000000" when "00001000101111101", -- t[4477] = 0
      "0000000" when "00001000101111110", -- t[4478] = 0
      "0000000" when "00001000101111111", -- t[4479] = 0
      "0000000" when "00001000110000000", -- t[4480] = 0
      "0000000" when "00001000110000001", -- t[4481] = 0
      "0000000" when "00001000110000010", -- t[4482] = 0
      "0000000" when "00001000110000011", -- t[4483] = 0
      "0000000" when "00001000110000100", -- t[4484] = 0
      "0000000" when "00001000110000101", -- t[4485] = 0
      "0000000" when "00001000110000110", -- t[4486] = 0
      "0000000" when "00001000110000111", -- t[4487] = 0
      "0000000" when "00001000110001000", -- t[4488] = 0
      "0000000" when "00001000110001001", -- t[4489] = 0
      "0000000" when "00001000110001010", -- t[4490] = 0
      "0000000" when "00001000110001011", -- t[4491] = 0
      "0000000" when "00001000110001100", -- t[4492] = 0
      "0000000" when "00001000110001101", -- t[4493] = 0
      "0000000" when "00001000110001110", -- t[4494] = 0
      "0000000" when "00001000110001111", -- t[4495] = 0
      "0000000" when "00001000110010000", -- t[4496] = 0
      "0000000" when "00001000110010001", -- t[4497] = 0
      "0000000" when "00001000110010010", -- t[4498] = 0
      "0000000" when "00001000110010011", -- t[4499] = 0
      "0000000" when "00001000110010100", -- t[4500] = 0
      "0000000" when "00001000110010101", -- t[4501] = 0
      "0000000" when "00001000110010110", -- t[4502] = 0
      "0000000" when "00001000110010111", -- t[4503] = 0
      "0000000" when "00001000110011000", -- t[4504] = 0
      "0000000" when "00001000110011001", -- t[4505] = 0
      "0000000" when "00001000110011010", -- t[4506] = 0
      "0000000" when "00001000110011011", -- t[4507] = 0
      "0000000" when "00001000110011100", -- t[4508] = 0
      "0000000" when "00001000110011101", -- t[4509] = 0
      "0000000" when "00001000110011110", -- t[4510] = 0
      "0000000" when "00001000110011111", -- t[4511] = 0
      "0000000" when "00001000110100000", -- t[4512] = 0
      "0000000" when "00001000110100001", -- t[4513] = 0
      "0000000" when "00001000110100010", -- t[4514] = 0
      "0000000" when "00001000110100011", -- t[4515] = 0
      "0000000" when "00001000110100100", -- t[4516] = 0
      "0000000" when "00001000110100101", -- t[4517] = 0
      "0000000" when "00001000110100110", -- t[4518] = 0
      "0000000" when "00001000110100111", -- t[4519] = 0
      "0000000" when "00001000110101000", -- t[4520] = 0
      "0000000" when "00001000110101001", -- t[4521] = 0
      "0000000" when "00001000110101010", -- t[4522] = 0
      "0000000" when "00001000110101011", -- t[4523] = 0
      "0000000" when "00001000110101100", -- t[4524] = 0
      "0000000" when "00001000110101101", -- t[4525] = 0
      "0000000" when "00001000110101110", -- t[4526] = 0
      "0000000" when "00001000110101111", -- t[4527] = 0
      "0000000" when "00001000110110000", -- t[4528] = 0
      "0000000" when "00001000110110001", -- t[4529] = 0
      "0000000" when "00001000110110010", -- t[4530] = 0
      "0000000" when "00001000110110011", -- t[4531] = 0
      "0000000" when "00001000110110100", -- t[4532] = 0
      "0000000" when "00001000110110101", -- t[4533] = 0
      "0000000" when "00001000110110110", -- t[4534] = 0
      "0000000" when "00001000110110111", -- t[4535] = 0
      "0000000" when "00001000110111000", -- t[4536] = 0
      "0000000" when "00001000110111001", -- t[4537] = 0
      "0000000" when "00001000110111010", -- t[4538] = 0
      "0000000" when "00001000110111011", -- t[4539] = 0
      "0000000" when "00001000110111100", -- t[4540] = 0
      "0000000" when "00001000110111101", -- t[4541] = 0
      "0000000" when "00001000110111110", -- t[4542] = 0
      "0000000" when "00001000110111111", -- t[4543] = 0
      "0000000" when "00001000111000000", -- t[4544] = 0
      "0000000" when "00001000111000001", -- t[4545] = 0
      "0000000" when "00001000111000010", -- t[4546] = 0
      "0000000" when "00001000111000011", -- t[4547] = 0
      "0000000" when "00001000111000100", -- t[4548] = 0
      "0000000" when "00001000111000101", -- t[4549] = 0
      "0000000" when "00001000111000110", -- t[4550] = 0
      "0000000" when "00001000111000111", -- t[4551] = 0
      "0000000" when "00001000111001000", -- t[4552] = 0
      "0000000" when "00001000111001001", -- t[4553] = 0
      "0000000" when "00001000111001010", -- t[4554] = 0
      "0000000" when "00001000111001011", -- t[4555] = 0
      "0000000" when "00001000111001100", -- t[4556] = 0
      "0000000" when "00001000111001101", -- t[4557] = 0
      "0000000" when "00001000111001110", -- t[4558] = 0
      "0000000" when "00001000111001111", -- t[4559] = 0
      "0000000" when "00001000111010000", -- t[4560] = 0
      "0000000" when "00001000111010001", -- t[4561] = 0
      "0000000" when "00001000111010010", -- t[4562] = 0
      "0000000" when "00001000111010011", -- t[4563] = 0
      "0000000" when "00001000111010100", -- t[4564] = 0
      "0000000" when "00001000111010101", -- t[4565] = 0
      "0000000" when "00001000111010110", -- t[4566] = 0
      "0000000" when "00001000111010111", -- t[4567] = 0
      "0000000" when "00001000111011000", -- t[4568] = 0
      "0000000" when "00001000111011001", -- t[4569] = 0
      "0000000" when "00001000111011010", -- t[4570] = 0
      "0000000" when "00001000111011011", -- t[4571] = 0
      "0000000" when "00001000111011100", -- t[4572] = 0
      "0000000" when "00001000111011101", -- t[4573] = 0
      "0000000" when "00001000111011110", -- t[4574] = 0
      "0000000" when "00001000111011111", -- t[4575] = 0
      "0000000" when "00001000111100000", -- t[4576] = 0
      "0000000" when "00001000111100001", -- t[4577] = 0
      "0000000" when "00001000111100010", -- t[4578] = 0
      "0000000" when "00001000111100011", -- t[4579] = 0
      "0000000" when "00001000111100100", -- t[4580] = 0
      "0000000" when "00001000111100101", -- t[4581] = 0
      "0000000" when "00001000111100110", -- t[4582] = 0
      "0000000" when "00001000111100111", -- t[4583] = 0
      "0000000" when "00001000111101000", -- t[4584] = 0
      "0000000" when "00001000111101001", -- t[4585] = 0
      "0000000" when "00001000111101010", -- t[4586] = 0
      "0000000" when "00001000111101011", -- t[4587] = 0
      "0000000" when "00001000111101100", -- t[4588] = 0
      "0000000" when "00001000111101101", -- t[4589] = 0
      "0000000" when "00001000111101110", -- t[4590] = 0
      "0000000" when "00001000111101111", -- t[4591] = 0
      "0000000" when "00001000111110000", -- t[4592] = 0
      "0000000" when "00001000111110001", -- t[4593] = 0
      "0000000" when "00001000111110010", -- t[4594] = 0
      "0000000" when "00001000111110011", -- t[4595] = 0
      "0000000" when "00001000111110100", -- t[4596] = 0
      "0000000" when "00001000111110101", -- t[4597] = 0
      "0000000" when "00001000111110110", -- t[4598] = 0
      "0000000" when "00001000111110111", -- t[4599] = 0
      "0000000" when "00001000111111000", -- t[4600] = 0
      "0000000" when "00001000111111001", -- t[4601] = 0
      "0000000" when "00001000111111010", -- t[4602] = 0
      "0000000" when "00001000111111011", -- t[4603] = 0
      "0000000" when "00001000111111100", -- t[4604] = 0
      "0000000" when "00001000111111101", -- t[4605] = 0
      "0000000" when "00001000111111110", -- t[4606] = 0
      "0000000" when "00001000111111111", -- t[4607] = 0
      "0000000" when "00001001000000000", -- t[4608] = 0
      "0000000" when "00001001000000001", -- t[4609] = 0
      "0000000" when "00001001000000010", -- t[4610] = 0
      "0000000" when "00001001000000011", -- t[4611] = 0
      "0000000" when "00001001000000100", -- t[4612] = 0
      "0000000" when "00001001000000101", -- t[4613] = 0
      "0000000" when "00001001000000110", -- t[4614] = 0
      "0000000" when "00001001000000111", -- t[4615] = 0
      "0000000" when "00001001000001000", -- t[4616] = 0
      "0000000" when "00001001000001001", -- t[4617] = 0
      "0000000" when "00001001000001010", -- t[4618] = 0
      "0000000" when "00001001000001011", -- t[4619] = 0
      "0000000" when "00001001000001100", -- t[4620] = 0
      "0000000" when "00001001000001101", -- t[4621] = 0
      "0000000" when "00001001000001110", -- t[4622] = 0
      "0000000" when "00001001000001111", -- t[4623] = 0
      "0000000" when "00001001000010000", -- t[4624] = 0
      "0000000" when "00001001000010001", -- t[4625] = 0
      "0000000" when "00001001000010010", -- t[4626] = 0
      "0000000" when "00001001000010011", -- t[4627] = 0
      "0000000" when "00001001000010100", -- t[4628] = 0
      "0000000" when "00001001000010101", -- t[4629] = 0
      "0000000" when "00001001000010110", -- t[4630] = 0
      "0000000" when "00001001000010111", -- t[4631] = 0
      "0000000" when "00001001000011000", -- t[4632] = 0
      "0000000" when "00001001000011001", -- t[4633] = 0
      "0000000" when "00001001000011010", -- t[4634] = 0
      "0000000" when "00001001000011011", -- t[4635] = 0
      "0000000" when "00001001000011100", -- t[4636] = 0
      "0000000" when "00001001000011101", -- t[4637] = 0
      "0000000" when "00001001000011110", -- t[4638] = 0
      "0000000" when "00001001000011111", -- t[4639] = 0
      "0000000" when "00001001000100000", -- t[4640] = 0
      "0000000" when "00001001000100001", -- t[4641] = 0
      "0000000" when "00001001000100010", -- t[4642] = 0
      "0000000" when "00001001000100011", -- t[4643] = 0
      "0000000" when "00001001000100100", -- t[4644] = 0
      "0000000" when "00001001000100101", -- t[4645] = 0
      "0000000" when "00001001000100110", -- t[4646] = 0
      "0000000" when "00001001000100111", -- t[4647] = 0
      "0000000" when "00001001000101000", -- t[4648] = 0
      "0000000" when "00001001000101001", -- t[4649] = 0
      "0000000" when "00001001000101010", -- t[4650] = 0
      "0000000" when "00001001000101011", -- t[4651] = 0
      "0000000" when "00001001000101100", -- t[4652] = 0
      "0000000" when "00001001000101101", -- t[4653] = 0
      "0000000" when "00001001000101110", -- t[4654] = 0
      "0000000" when "00001001000101111", -- t[4655] = 0
      "0000000" when "00001001000110000", -- t[4656] = 0
      "0000000" when "00001001000110001", -- t[4657] = 0
      "0000000" when "00001001000110010", -- t[4658] = 0
      "0000000" when "00001001000110011", -- t[4659] = 0
      "0000000" when "00001001000110100", -- t[4660] = 0
      "0000000" when "00001001000110101", -- t[4661] = 0
      "0000000" when "00001001000110110", -- t[4662] = 0
      "0000000" when "00001001000110111", -- t[4663] = 0
      "0000000" when "00001001000111000", -- t[4664] = 0
      "0000000" when "00001001000111001", -- t[4665] = 0
      "0000000" when "00001001000111010", -- t[4666] = 0
      "0000000" when "00001001000111011", -- t[4667] = 0
      "0000000" when "00001001000111100", -- t[4668] = 0
      "0000000" when "00001001000111101", -- t[4669] = 0
      "0000000" when "00001001000111110", -- t[4670] = 0
      "0000000" when "00001001000111111", -- t[4671] = 0
      "0000000" when "00001001001000000", -- t[4672] = 0
      "0000000" when "00001001001000001", -- t[4673] = 0
      "0000000" when "00001001001000010", -- t[4674] = 0
      "0000000" when "00001001001000011", -- t[4675] = 0
      "0000000" when "00001001001000100", -- t[4676] = 0
      "0000000" when "00001001001000101", -- t[4677] = 0
      "0000000" when "00001001001000110", -- t[4678] = 0
      "0000000" when "00001001001000111", -- t[4679] = 0
      "0000000" when "00001001001001000", -- t[4680] = 0
      "0000000" when "00001001001001001", -- t[4681] = 0
      "0000000" when "00001001001001010", -- t[4682] = 0
      "0000000" when "00001001001001011", -- t[4683] = 0
      "0000000" when "00001001001001100", -- t[4684] = 0
      "0000000" when "00001001001001101", -- t[4685] = 0
      "0000000" when "00001001001001110", -- t[4686] = 0
      "0000000" when "00001001001001111", -- t[4687] = 0
      "0000000" when "00001001001010000", -- t[4688] = 0
      "0000000" when "00001001001010001", -- t[4689] = 0
      "0000000" when "00001001001010010", -- t[4690] = 0
      "0000000" when "00001001001010011", -- t[4691] = 0
      "0000000" when "00001001001010100", -- t[4692] = 0
      "0000000" when "00001001001010101", -- t[4693] = 0
      "0000000" when "00001001001010110", -- t[4694] = 0
      "0000000" when "00001001001010111", -- t[4695] = 0
      "0000000" when "00001001001011000", -- t[4696] = 0
      "0000000" when "00001001001011001", -- t[4697] = 0
      "0000000" when "00001001001011010", -- t[4698] = 0
      "0000000" when "00001001001011011", -- t[4699] = 0
      "0000000" when "00001001001011100", -- t[4700] = 0
      "0000000" when "00001001001011101", -- t[4701] = 0
      "0000000" when "00001001001011110", -- t[4702] = 0
      "0000000" when "00001001001011111", -- t[4703] = 0
      "0000000" when "00001001001100000", -- t[4704] = 0
      "0000000" when "00001001001100001", -- t[4705] = 0
      "0000000" when "00001001001100010", -- t[4706] = 0
      "0000000" when "00001001001100011", -- t[4707] = 0
      "0000000" when "00001001001100100", -- t[4708] = 0
      "0000000" when "00001001001100101", -- t[4709] = 0
      "0000000" when "00001001001100110", -- t[4710] = 0
      "0000000" when "00001001001100111", -- t[4711] = 0
      "0000000" when "00001001001101000", -- t[4712] = 0
      "0000000" when "00001001001101001", -- t[4713] = 0
      "0000000" when "00001001001101010", -- t[4714] = 0
      "0000000" when "00001001001101011", -- t[4715] = 0
      "0000000" when "00001001001101100", -- t[4716] = 0
      "0000000" when "00001001001101101", -- t[4717] = 0
      "0000000" when "00001001001101110", -- t[4718] = 0
      "0000000" when "00001001001101111", -- t[4719] = 0
      "0000000" when "00001001001110000", -- t[4720] = 0
      "0000000" when "00001001001110001", -- t[4721] = 0
      "0000000" when "00001001001110010", -- t[4722] = 0
      "0000000" when "00001001001110011", -- t[4723] = 0
      "0000000" when "00001001001110100", -- t[4724] = 0
      "0000000" when "00001001001110101", -- t[4725] = 0
      "0000000" when "00001001001110110", -- t[4726] = 0
      "0000000" when "00001001001110111", -- t[4727] = 0
      "0000000" when "00001001001111000", -- t[4728] = 0
      "0000000" when "00001001001111001", -- t[4729] = 0
      "0000000" when "00001001001111010", -- t[4730] = 0
      "0000000" when "00001001001111011", -- t[4731] = 0
      "0000000" when "00001001001111100", -- t[4732] = 0
      "0000000" when "00001001001111101", -- t[4733] = 0
      "0000000" when "00001001001111110", -- t[4734] = 0
      "0000000" when "00001001001111111", -- t[4735] = 0
      "0000000" when "00001001010000000", -- t[4736] = 0
      "0000000" when "00001001010000001", -- t[4737] = 0
      "0000000" when "00001001010000010", -- t[4738] = 0
      "0000000" when "00001001010000011", -- t[4739] = 0
      "0000000" when "00001001010000100", -- t[4740] = 0
      "0000000" when "00001001010000101", -- t[4741] = 0
      "0000000" when "00001001010000110", -- t[4742] = 0
      "0000000" when "00001001010000111", -- t[4743] = 0
      "0000000" when "00001001010001000", -- t[4744] = 0
      "0000000" when "00001001010001001", -- t[4745] = 0
      "0000000" when "00001001010001010", -- t[4746] = 0
      "0000000" when "00001001010001011", -- t[4747] = 0
      "0000000" when "00001001010001100", -- t[4748] = 0
      "0000000" when "00001001010001101", -- t[4749] = 0
      "0000000" when "00001001010001110", -- t[4750] = 0
      "0000000" when "00001001010001111", -- t[4751] = 0
      "0000000" when "00001001010010000", -- t[4752] = 0
      "0000000" when "00001001010010001", -- t[4753] = 0
      "0000000" when "00001001010010010", -- t[4754] = 0
      "0000000" when "00001001010010011", -- t[4755] = 0
      "0000000" when "00001001010010100", -- t[4756] = 0
      "0000000" when "00001001010010101", -- t[4757] = 0
      "0000000" when "00001001010010110", -- t[4758] = 0
      "0000000" when "00001001010010111", -- t[4759] = 0
      "0000000" when "00001001010011000", -- t[4760] = 0
      "0000000" when "00001001010011001", -- t[4761] = 0
      "0000000" when "00001001010011010", -- t[4762] = 0
      "0000000" when "00001001010011011", -- t[4763] = 0
      "0000000" when "00001001010011100", -- t[4764] = 0
      "0000000" when "00001001010011101", -- t[4765] = 0
      "0000000" when "00001001010011110", -- t[4766] = 0
      "0000000" when "00001001010011111", -- t[4767] = 0
      "0000000" when "00001001010100000", -- t[4768] = 0
      "0000000" when "00001001010100001", -- t[4769] = 0
      "0000000" when "00001001010100010", -- t[4770] = 0
      "0000000" when "00001001010100011", -- t[4771] = 0
      "0000000" when "00001001010100100", -- t[4772] = 0
      "0000000" when "00001001010100101", -- t[4773] = 0
      "0000000" when "00001001010100110", -- t[4774] = 0
      "0000000" when "00001001010100111", -- t[4775] = 0
      "0000000" when "00001001010101000", -- t[4776] = 0
      "0000000" when "00001001010101001", -- t[4777] = 0
      "0000000" when "00001001010101010", -- t[4778] = 0
      "0000000" when "00001001010101011", -- t[4779] = 0
      "0000000" when "00001001010101100", -- t[4780] = 0
      "0000000" when "00001001010101101", -- t[4781] = 0
      "0000000" when "00001001010101110", -- t[4782] = 0
      "0000000" when "00001001010101111", -- t[4783] = 0
      "0000000" when "00001001010110000", -- t[4784] = 0
      "0000000" when "00001001010110001", -- t[4785] = 0
      "0000000" when "00001001010110010", -- t[4786] = 0
      "0000000" when "00001001010110011", -- t[4787] = 0
      "0000000" when "00001001010110100", -- t[4788] = 0
      "0000000" when "00001001010110101", -- t[4789] = 0
      "0000000" when "00001001010110110", -- t[4790] = 0
      "0000000" when "00001001010110111", -- t[4791] = 0
      "0000000" when "00001001010111000", -- t[4792] = 0
      "0000000" when "00001001010111001", -- t[4793] = 0
      "0000000" when "00001001010111010", -- t[4794] = 0
      "0000000" when "00001001010111011", -- t[4795] = 0
      "0000000" when "00001001010111100", -- t[4796] = 0
      "0000000" when "00001001010111101", -- t[4797] = 0
      "0000000" when "00001001010111110", -- t[4798] = 0
      "0000000" when "00001001010111111", -- t[4799] = 0
      "0000000" when "00001001011000000", -- t[4800] = 0
      "0000000" when "00001001011000001", -- t[4801] = 0
      "0000000" when "00001001011000010", -- t[4802] = 0
      "0000000" when "00001001011000011", -- t[4803] = 0
      "0000000" when "00001001011000100", -- t[4804] = 0
      "0000000" when "00001001011000101", -- t[4805] = 0
      "0000000" when "00001001011000110", -- t[4806] = 0
      "0000000" when "00001001011000111", -- t[4807] = 0
      "0000000" when "00001001011001000", -- t[4808] = 0
      "0000000" when "00001001011001001", -- t[4809] = 0
      "0000000" when "00001001011001010", -- t[4810] = 0
      "0000000" when "00001001011001011", -- t[4811] = 0
      "0000000" when "00001001011001100", -- t[4812] = 0
      "0000000" when "00001001011001101", -- t[4813] = 0
      "0000000" when "00001001011001110", -- t[4814] = 0
      "0000000" when "00001001011001111", -- t[4815] = 0
      "0000000" when "00001001011010000", -- t[4816] = 0
      "0000000" when "00001001011010001", -- t[4817] = 0
      "0000000" when "00001001011010010", -- t[4818] = 0
      "0000000" when "00001001011010011", -- t[4819] = 0
      "0000000" when "00001001011010100", -- t[4820] = 0
      "0000000" when "00001001011010101", -- t[4821] = 0
      "0000000" when "00001001011010110", -- t[4822] = 0
      "0000000" when "00001001011010111", -- t[4823] = 0
      "0000000" when "00001001011011000", -- t[4824] = 0
      "0000000" when "00001001011011001", -- t[4825] = 0
      "0000000" when "00001001011011010", -- t[4826] = 0
      "0000000" when "00001001011011011", -- t[4827] = 0
      "0000000" when "00001001011011100", -- t[4828] = 0
      "0000000" when "00001001011011101", -- t[4829] = 0
      "0000000" when "00001001011011110", -- t[4830] = 0
      "0000000" when "00001001011011111", -- t[4831] = 0
      "0000000" when "00001001011100000", -- t[4832] = 0
      "0000000" when "00001001011100001", -- t[4833] = 0
      "0000000" when "00001001011100010", -- t[4834] = 0
      "0000000" when "00001001011100011", -- t[4835] = 0
      "0000000" when "00001001011100100", -- t[4836] = 0
      "0000000" when "00001001011100101", -- t[4837] = 0
      "0000000" when "00001001011100110", -- t[4838] = 0
      "0000000" when "00001001011100111", -- t[4839] = 0
      "0000000" when "00001001011101000", -- t[4840] = 0
      "0000000" when "00001001011101001", -- t[4841] = 0
      "0000000" when "00001001011101010", -- t[4842] = 0
      "0000000" when "00001001011101011", -- t[4843] = 0
      "0000000" when "00001001011101100", -- t[4844] = 0
      "0000000" when "00001001011101101", -- t[4845] = 0
      "0000000" when "00001001011101110", -- t[4846] = 0
      "0000000" when "00001001011101111", -- t[4847] = 0
      "0000000" when "00001001011110000", -- t[4848] = 0
      "0000000" when "00001001011110001", -- t[4849] = 0
      "0000000" when "00001001011110010", -- t[4850] = 0
      "0000000" when "00001001011110011", -- t[4851] = 0
      "0000000" when "00001001011110100", -- t[4852] = 0
      "0000000" when "00001001011110101", -- t[4853] = 0
      "0000000" when "00001001011110110", -- t[4854] = 0
      "0000000" when "00001001011110111", -- t[4855] = 0
      "0000000" when "00001001011111000", -- t[4856] = 0
      "0000000" when "00001001011111001", -- t[4857] = 0
      "0000000" when "00001001011111010", -- t[4858] = 0
      "0000000" when "00001001011111011", -- t[4859] = 0
      "0000000" when "00001001011111100", -- t[4860] = 0
      "0000000" when "00001001011111101", -- t[4861] = 0
      "0000000" when "00001001011111110", -- t[4862] = 0
      "0000000" when "00001001011111111", -- t[4863] = 0
      "0000000" when "00001001100000000", -- t[4864] = 0
      "0000000" when "00001001100000001", -- t[4865] = 0
      "0000000" when "00001001100000010", -- t[4866] = 0
      "0000000" when "00001001100000011", -- t[4867] = 0
      "0000000" when "00001001100000100", -- t[4868] = 0
      "0000000" when "00001001100000101", -- t[4869] = 0
      "0000000" when "00001001100000110", -- t[4870] = 0
      "0000000" when "00001001100000111", -- t[4871] = 0
      "0000000" when "00001001100001000", -- t[4872] = 0
      "0000000" when "00001001100001001", -- t[4873] = 0
      "0000000" when "00001001100001010", -- t[4874] = 0
      "0000000" when "00001001100001011", -- t[4875] = 0
      "0000000" when "00001001100001100", -- t[4876] = 0
      "0000000" when "00001001100001101", -- t[4877] = 0
      "0000000" when "00001001100001110", -- t[4878] = 0
      "0000000" when "00001001100001111", -- t[4879] = 0
      "0000000" when "00001001100010000", -- t[4880] = 0
      "0000000" when "00001001100010001", -- t[4881] = 0
      "0000000" when "00001001100010010", -- t[4882] = 0
      "0000000" when "00001001100010011", -- t[4883] = 0
      "0000000" when "00001001100010100", -- t[4884] = 0
      "0000000" when "00001001100010101", -- t[4885] = 0
      "0000000" when "00001001100010110", -- t[4886] = 0
      "0000000" when "00001001100010111", -- t[4887] = 0
      "0000000" when "00001001100011000", -- t[4888] = 0
      "0000000" when "00001001100011001", -- t[4889] = 0
      "0000000" when "00001001100011010", -- t[4890] = 0
      "0000000" when "00001001100011011", -- t[4891] = 0
      "0000000" when "00001001100011100", -- t[4892] = 0
      "0000000" when "00001001100011101", -- t[4893] = 0
      "0000000" when "00001001100011110", -- t[4894] = 0
      "0000000" when "00001001100011111", -- t[4895] = 0
      "0000000" when "00001001100100000", -- t[4896] = 0
      "0000000" when "00001001100100001", -- t[4897] = 0
      "0000000" when "00001001100100010", -- t[4898] = 0
      "0000000" when "00001001100100011", -- t[4899] = 0
      "0000000" when "00001001100100100", -- t[4900] = 0
      "0000000" when "00001001100100101", -- t[4901] = 0
      "0000000" when "00001001100100110", -- t[4902] = 0
      "0000000" when "00001001100100111", -- t[4903] = 0
      "0000000" when "00001001100101000", -- t[4904] = 0
      "0000000" when "00001001100101001", -- t[4905] = 0
      "0000000" when "00001001100101010", -- t[4906] = 0
      "0000000" when "00001001100101011", -- t[4907] = 0
      "0000000" when "00001001100101100", -- t[4908] = 0
      "0000000" when "00001001100101101", -- t[4909] = 0
      "0000000" when "00001001100101110", -- t[4910] = 0
      "0000000" when "00001001100101111", -- t[4911] = 0
      "0000000" when "00001001100110000", -- t[4912] = 0
      "0000000" when "00001001100110001", -- t[4913] = 0
      "0000000" when "00001001100110010", -- t[4914] = 0
      "0000000" when "00001001100110011", -- t[4915] = 0
      "0000000" when "00001001100110100", -- t[4916] = 0
      "0000000" when "00001001100110101", -- t[4917] = 0
      "0000000" when "00001001100110110", -- t[4918] = 0
      "0000000" when "00001001100110111", -- t[4919] = 0
      "0000000" when "00001001100111000", -- t[4920] = 0
      "0000000" when "00001001100111001", -- t[4921] = 0
      "0000000" when "00001001100111010", -- t[4922] = 0
      "0000000" when "00001001100111011", -- t[4923] = 0
      "0000000" when "00001001100111100", -- t[4924] = 0
      "0000000" when "00001001100111101", -- t[4925] = 0
      "0000000" when "00001001100111110", -- t[4926] = 0
      "0000000" when "00001001100111111", -- t[4927] = 0
      "0000000" when "00001001101000000", -- t[4928] = 0
      "0000000" when "00001001101000001", -- t[4929] = 0
      "0000000" when "00001001101000010", -- t[4930] = 0
      "0000000" when "00001001101000011", -- t[4931] = 0
      "0000000" when "00001001101000100", -- t[4932] = 0
      "0000000" when "00001001101000101", -- t[4933] = 0
      "0000000" when "00001001101000110", -- t[4934] = 0
      "0000000" when "00001001101000111", -- t[4935] = 0
      "0000000" when "00001001101001000", -- t[4936] = 0
      "0000000" when "00001001101001001", -- t[4937] = 0
      "0000000" when "00001001101001010", -- t[4938] = 0
      "0000000" when "00001001101001011", -- t[4939] = 0
      "0000000" when "00001001101001100", -- t[4940] = 0
      "0000000" when "00001001101001101", -- t[4941] = 0
      "0000000" when "00001001101001110", -- t[4942] = 0
      "0000000" when "00001001101001111", -- t[4943] = 0
      "0000000" when "00001001101010000", -- t[4944] = 0
      "0000000" when "00001001101010001", -- t[4945] = 0
      "0000000" when "00001001101010010", -- t[4946] = 0
      "0000000" when "00001001101010011", -- t[4947] = 0
      "0000000" when "00001001101010100", -- t[4948] = 0
      "0000000" when "00001001101010101", -- t[4949] = 0
      "0000000" when "00001001101010110", -- t[4950] = 0
      "0000000" when "00001001101010111", -- t[4951] = 0
      "0000000" when "00001001101011000", -- t[4952] = 0
      "0000000" when "00001001101011001", -- t[4953] = 0
      "0000000" when "00001001101011010", -- t[4954] = 0
      "0000000" when "00001001101011011", -- t[4955] = 0
      "0000000" when "00001001101011100", -- t[4956] = 0
      "0000000" when "00001001101011101", -- t[4957] = 0
      "0000000" when "00001001101011110", -- t[4958] = 0
      "0000000" when "00001001101011111", -- t[4959] = 0
      "0000000" when "00001001101100000", -- t[4960] = 0
      "0000000" when "00001001101100001", -- t[4961] = 0
      "0000000" when "00001001101100010", -- t[4962] = 0
      "0000000" when "00001001101100011", -- t[4963] = 0
      "0000000" when "00001001101100100", -- t[4964] = 0
      "0000000" when "00001001101100101", -- t[4965] = 0
      "0000000" when "00001001101100110", -- t[4966] = 0
      "0000000" when "00001001101100111", -- t[4967] = 0
      "0000000" when "00001001101101000", -- t[4968] = 0
      "0000000" when "00001001101101001", -- t[4969] = 0
      "0000000" when "00001001101101010", -- t[4970] = 0
      "0000000" when "00001001101101011", -- t[4971] = 0
      "0000000" when "00001001101101100", -- t[4972] = 0
      "0000000" when "00001001101101101", -- t[4973] = 0
      "0000000" when "00001001101101110", -- t[4974] = 0
      "0000000" when "00001001101101111", -- t[4975] = 0
      "0000000" when "00001001101110000", -- t[4976] = 0
      "0000000" when "00001001101110001", -- t[4977] = 0
      "0000000" when "00001001101110010", -- t[4978] = 0
      "0000000" when "00001001101110011", -- t[4979] = 0
      "0000000" when "00001001101110100", -- t[4980] = 0
      "0000000" when "00001001101110101", -- t[4981] = 0
      "0000000" when "00001001101110110", -- t[4982] = 0
      "0000000" when "00001001101110111", -- t[4983] = 0
      "0000000" when "00001001101111000", -- t[4984] = 0
      "0000000" when "00001001101111001", -- t[4985] = 0
      "0000000" when "00001001101111010", -- t[4986] = 0
      "0000000" when "00001001101111011", -- t[4987] = 0
      "0000000" when "00001001101111100", -- t[4988] = 0
      "0000000" when "00001001101111101", -- t[4989] = 0
      "0000000" when "00001001101111110", -- t[4990] = 0
      "0000000" when "00001001101111111", -- t[4991] = 0
      "0000000" when "00001001110000000", -- t[4992] = 0
      "0000000" when "00001001110000001", -- t[4993] = 0
      "0000000" when "00001001110000010", -- t[4994] = 0
      "0000000" when "00001001110000011", -- t[4995] = 0
      "0000000" when "00001001110000100", -- t[4996] = 0
      "0000000" when "00001001110000101", -- t[4997] = 0
      "0000000" when "00001001110000110", -- t[4998] = 0
      "0000000" when "00001001110000111", -- t[4999] = 0
      "0000000" when "00001001110001000", -- t[5000] = 0
      "0000000" when "00001001110001001", -- t[5001] = 0
      "0000000" when "00001001110001010", -- t[5002] = 0
      "0000000" when "00001001110001011", -- t[5003] = 0
      "0000000" when "00001001110001100", -- t[5004] = 0
      "0000000" when "00001001110001101", -- t[5005] = 0
      "0000000" when "00001001110001110", -- t[5006] = 0
      "0000000" when "00001001110001111", -- t[5007] = 0
      "0000000" when "00001001110010000", -- t[5008] = 0
      "0000000" when "00001001110010001", -- t[5009] = 0
      "0000000" when "00001001110010010", -- t[5010] = 0
      "0000000" when "00001001110010011", -- t[5011] = 0
      "0000000" when "00001001110010100", -- t[5012] = 0
      "0000000" when "00001001110010101", -- t[5013] = 0
      "0000000" when "00001001110010110", -- t[5014] = 0
      "0000000" when "00001001110010111", -- t[5015] = 0
      "0000000" when "00001001110011000", -- t[5016] = 0
      "0000000" when "00001001110011001", -- t[5017] = 0
      "0000000" when "00001001110011010", -- t[5018] = 0
      "0000000" when "00001001110011011", -- t[5019] = 0
      "0000000" when "00001001110011100", -- t[5020] = 0
      "0000000" when "00001001110011101", -- t[5021] = 0
      "0000000" when "00001001110011110", -- t[5022] = 0
      "0000000" when "00001001110011111", -- t[5023] = 0
      "0000000" when "00001001110100000", -- t[5024] = 0
      "0000000" when "00001001110100001", -- t[5025] = 0
      "0000000" when "00001001110100010", -- t[5026] = 0
      "0000000" when "00001001110100011", -- t[5027] = 0
      "0000000" when "00001001110100100", -- t[5028] = 0
      "0000000" when "00001001110100101", -- t[5029] = 0
      "0000000" when "00001001110100110", -- t[5030] = 0
      "0000000" when "00001001110100111", -- t[5031] = 0
      "0000000" when "00001001110101000", -- t[5032] = 0
      "0000000" when "00001001110101001", -- t[5033] = 0
      "0000000" when "00001001110101010", -- t[5034] = 0
      "0000000" when "00001001110101011", -- t[5035] = 0
      "0000000" when "00001001110101100", -- t[5036] = 0
      "0000000" when "00001001110101101", -- t[5037] = 0
      "0000000" when "00001001110101110", -- t[5038] = 0
      "0000000" when "00001001110101111", -- t[5039] = 0
      "0000000" when "00001001110110000", -- t[5040] = 0
      "0000000" when "00001001110110001", -- t[5041] = 0
      "0000000" when "00001001110110010", -- t[5042] = 0
      "0000000" when "00001001110110011", -- t[5043] = 0
      "0000000" when "00001001110110100", -- t[5044] = 0
      "0000000" when "00001001110110101", -- t[5045] = 0
      "0000000" when "00001001110110110", -- t[5046] = 0
      "0000000" when "00001001110110111", -- t[5047] = 0
      "0000000" when "00001001110111000", -- t[5048] = 0
      "0000000" when "00001001110111001", -- t[5049] = 0
      "0000000" when "00001001110111010", -- t[5050] = 0
      "0000000" when "00001001110111011", -- t[5051] = 0
      "0000000" when "00001001110111100", -- t[5052] = 0
      "0000000" when "00001001110111101", -- t[5053] = 0
      "0000000" when "00001001110111110", -- t[5054] = 0
      "0000000" when "00001001110111111", -- t[5055] = 0
      "0000000" when "00001001111000000", -- t[5056] = 0
      "0000000" when "00001001111000001", -- t[5057] = 0
      "0000000" when "00001001111000010", -- t[5058] = 0
      "0000000" when "00001001111000011", -- t[5059] = 0
      "0000000" when "00001001111000100", -- t[5060] = 0
      "0000000" when "00001001111000101", -- t[5061] = 0
      "0000000" when "00001001111000110", -- t[5062] = 0
      "0000000" when "00001001111000111", -- t[5063] = 0
      "0000000" when "00001001111001000", -- t[5064] = 0
      "0000000" when "00001001111001001", -- t[5065] = 0
      "0000000" when "00001001111001010", -- t[5066] = 0
      "0000000" when "00001001111001011", -- t[5067] = 0
      "0000000" when "00001001111001100", -- t[5068] = 0
      "0000000" when "00001001111001101", -- t[5069] = 0
      "0000000" when "00001001111001110", -- t[5070] = 0
      "0000000" when "00001001111001111", -- t[5071] = 0
      "0000000" when "00001001111010000", -- t[5072] = 0
      "0000000" when "00001001111010001", -- t[5073] = 0
      "0000000" when "00001001111010010", -- t[5074] = 0
      "0000000" when "00001001111010011", -- t[5075] = 0
      "0000000" when "00001001111010100", -- t[5076] = 0
      "0000000" when "00001001111010101", -- t[5077] = 0
      "0000000" when "00001001111010110", -- t[5078] = 0
      "0000000" when "00001001111010111", -- t[5079] = 0
      "0000000" when "00001001111011000", -- t[5080] = 0
      "0000000" when "00001001111011001", -- t[5081] = 0
      "0000000" when "00001001111011010", -- t[5082] = 0
      "0000000" when "00001001111011011", -- t[5083] = 0
      "0000000" when "00001001111011100", -- t[5084] = 0
      "0000000" when "00001001111011101", -- t[5085] = 0
      "0000000" when "00001001111011110", -- t[5086] = 0
      "0000000" when "00001001111011111", -- t[5087] = 0
      "0000000" when "00001001111100000", -- t[5088] = 0
      "0000000" when "00001001111100001", -- t[5089] = 0
      "0000000" when "00001001111100010", -- t[5090] = 0
      "0000000" when "00001001111100011", -- t[5091] = 0
      "0000000" when "00001001111100100", -- t[5092] = 0
      "0000000" when "00001001111100101", -- t[5093] = 0
      "0000000" when "00001001111100110", -- t[5094] = 0
      "0000000" when "00001001111100111", -- t[5095] = 0
      "0000000" when "00001001111101000", -- t[5096] = 0
      "0000000" when "00001001111101001", -- t[5097] = 0
      "0000000" when "00001001111101010", -- t[5098] = 0
      "0000000" when "00001001111101011", -- t[5099] = 0
      "0000000" when "00001001111101100", -- t[5100] = 0
      "0000000" when "00001001111101101", -- t[5101] = 0
      "0000000" when "00001001111101110", -- t[5102] = 0
      "0000000" when "00001001111101111", -- t[5103] = 0
      "0000000" when "00001001111110000", -- t[5104] = 0
      "0000000" when "00001001111110001", -- t[5105] = 0
      "0000000" when "00001001111110010", -- t[5106] = 0
      "0000000" when "00001001111110011", -- t[5107] = 0
      "0000000" when "00001001111110100", -- t[5108] = 0
      "0000000" when "00001001111110101", -- t[5109] = 0
      "0000000" when "00001001111110110", -- t[5110] = 0
      "0000000" when "00001001111110111", -- t[5111] = 0
      "0000000" when "00001001111111000", -- t[5112] = 0
      "0000000" when "00001001111111001", -- t[5113] = 0
      "0000000" when "00001001111111010", -- t[5114] = 0
      "0000000" when "00001001111111011", -- t[5115] = 0
      "0000000" when "00001001111111100", -- t[5116] = 0
      "0000000" when "00001001111111101", -- t[5117] = 0
      "0000000" when "00001001111111110", -- t[5118] = 0
      "0000000" when "00001001111111111", -- t[5119] = 0
      "0000000" when "00001010000000000", -- t[5120] = 0
      "0000000" when "00001010000000001", -- t[5121] = 0
      "0000000" when "00001010000000010", -- t[5122] = 0
      "0000000" when "00001010000000011", -- t[5123] = 0
      "0000000" when "00001010000000100", -- t[5124] = 0
      "0000000" when "00001010000000101", -- t[5125] = 0
      "0000000" when "00001010000000110", -- t[5126] = 0
      "0000000" when "00001010000000111", -- t[5127] = 0
      "0000000" when "00001010000001000", -- t[5128] = 0
      "0000000" when "00001010000001001", -- t[5129] = 0
      "0000000" when "00001010000001010", -- t[5130] = 0
      "0000000" when "00001010000001011", -- t[5131] = 0
      "0000000" when "00001010000001100", -- t[5132] = 0
      "0000000" when "00001010000001101", -- t[5133] = 0
      "0000000" when "00001010000001110", -- t[5134] = 0
      "0000000" when "00001010000001111", -- t[5135] = 0
      "0000000" when "00001010000010000", -- t[5136] = 0
      "0000000" when "00001010000010001", -- t[5137] = 0
      "0000000" when "00001010000010010", -- t[5138] = 0
      "0000000" when "00001010000010011", -- t[5139] = 0
      "0000000" when "00001010000010100", -- t[5140] = 0
      "0000000" when "00001010000010101", -- t[5141] = 0
      "0000000" when "00001010000010110", -- t[5142] = 0
      "0000000" when "00001010000010111", -- t[5143] = 0
      "0000000" when "00001010000011000", -- t[5144] = 0
      "0000000" when "00001010000011001", -- t[5145] = 0
      "0000000" when "00001010000011010", -- t[5146] = 0
      "0000000" when "00001010000011011", -- t[5147] = 0
      "0000000" when "00001010000011100", -- t[5148] = 0
      "0000000" when "00001010000011101", -- t[5149] = 0
      "0000000" when "00001010000011110", -- t[5150] = 0
      "0000000" when "00001010000011111", -- t[5151] = 0
      "0000000" when "00001010000100000", -- t[5152] = 0
      "0000000" when "00001010000100001", -- t[5153] = 0
      "0000000" when "00001010000100010", -- t[5154] = 0
      "0000000" when "00001010000100011", -- t[5155] = 0
      "0000000" when "00001010000100100", -- t[5156] = 0
      "0000000" when "00001010000100101", -- t[5157] = 0
      "0000000" when "00001010000100110", -- t[5158] = 0
      "0000000" when "00001010000100111", -- t[5159] = 0
      "0000000" when "00001010000101000", -- t[5160] = 0
      "0000000" when "00001010000101001", -- t[5161] = 0
      "0000000" when "00001010000101010", -- t[5162] = 0
      "0000000" when "00001010000101011", -- t[5163] = 0
      "0000000" when "00001010000101100", -- t[5164] = 0
      "0000000" when "00001010000101101", -- t[5165] = 0
      "0000000" when "00001010000101110", -- t[5166] = 0
      "0000000" when "00001010000101111", -- t[5167] = 0
      "0000000" when "00001010000110000", -- t[5168] = 0
      "0000000" when "00001010000110001", -- t[5169] = 0
      "0000000" when "00001010000110010", -- t[5170] = 0
      "0000000" when "00001010000110011", -- t[5171] = 0
      "0000000" when "00001010000110100", -- t[5172] = 0
      "0000000" when "00001010000110101", -- t[5173] = 0
      "0000000" when "00001010000110110", -- t[5174] = 0
      "0000000" when "00001010000110111", -- t[5175] = 0
      "0000000" when "00001010000111000", -- t[5176] = 0
      "0000000" when "00001010000111001", -- t[5177] = 0
      "0000000" when "00001010000111010", -- t[5178] = 0
      "0000000" when "00001010000111011", -- t[5179] = 0
      "0000000" when "00001010000111100", -- t[5180] = 0
      "0000000" when "00001010000111101", -- t[5181] = 0
      "0000000" when "00001010000111110", -- t[5182] = 0
      "0000000" when "00001010000111111", -- t[5183] = 0
      "0000000" when "00001010001000000", -- t[5184] = 0
      "0000000" when "00001010001000001", -- t[5185] = 0
      "0000000" when "00001010001000010", -- t[5186] = 0
      "0000000" when "00001010001000011", -- t[5187] = 0
      "0000000" when "00001010001000100", -- t[5188] = 0
      "0000000" when "00001010001000101", -- t[5189] = 0
      "0000000" when "00001010001000110", -- t[5190] = 0
      "0000000" when "00001010001000111", -- t[5191] = 0
      "0000000" when "00001010001001000", -- t[5192] = 0
      "0000000" when "00001010001001001", -- t[5193] = 0
      "0000000" when "00001010001001010", -- t[5194] = 0
      "0000000" when "00001010001001011", -- t[5195] = 0
      "0000000" when "00001010001001100", -- t[5196] = 0
      "0000000" when "00001010001001101", -- t[5197] = 0
      "0000000" when "00001010001001110", -- t[5198] = 0
      "0000000" when "00001010001001111", -- t[5199] = 0
      "0000000" when "00001010001010000", -- t[5200] = 0
      "0000000" when "00001010001010001", -- t[5201] = 0
      "0000000" when "00001010001010010", -- t[5202] = 0
      "0000000" when "00001010001010011", -- t[5203] = 0
      "0000000" when "00001010001010100", -- t[5204] = 0
      "0000000" when "00001010001010101", -- t[5205] = 0
      "0000000" when "00001010001010110", -- t[5206] = 0
      "0000000" when "00001010001010111", -- t[5207] = 0
      "0000000" when "00001010001011000", -- t[5208] = 0
      "0000000" when "00001010001011001", -- t[5209] = 0
      "0000000" when "00001010001011010", -- t[5210] = 0
      "0000000" when "00001010001011011", -- t[5211] = 0
      "0000000" when "00001010001011100", -- t[5212] = 0
      "0000000" when "00001010001011101", -- t[5213] = 0
      "0000000" when "00001010001011110", -- t[5214] = 0
      "0000000" when "00001010001011111", -- t[5215] = 0
      "0000000" when "00001010001100000", -- t[5216] = 0
      "0000000" when "00001010001100001", -- t[5217] = 0
      "0000000" when "00001010001100010", -- t[5218] = 0
      "0000000" when "00001010001100011", -- t[5219] = 0
      "0000000" when "00001010001100100", -- t[5220] = 0
      "0000000" when "00001010001100101", -- t[5221] = 0
      "0000000" when "00001010001100110", -- t[5222] = 0
      "0000000" when "00001010001100111", -- t[5223] = 0
      "0000000" when "00001010001101000", -- t[5224] = 0
      "0000000" when "00001010001101001", -- t[5225] = 0
      "0000000" when "00001010001101010", -- t[5226] = 0
      "0000000" when "00001010001101011", -- t[5227] = 0
      "0000000" when "00001010001101100", -- t[5228] = 0
      "0000000" when "00001010001101101", -- t[5229] = 0
      "0000000" when "00001010001101110", -- t[5230] = 0
      "0000000" when "00001010001101111", -- t[5231] = 0
      "0000000" when "00001010001110000", -- t[5232] = 0
      "0000000" when "00001010001110001", -- t[5233] = 0
      "0000000" when "00001010001110010", -- t[5234] = 0
      "0000000" when "00001010001110011", -- t[5235] = 0
      "0000000" when "00001010001110100", -- t[5236] = 0
      "0000000" when "00001010001110101", -- t[5237] = 0
      "0000000" when "00001010001110110", -- t[5238] = 0
      "0000000" when "00001010001110111", -- t[5239] = 0
      "0000000" when "00001010001111000", -- t[5240] = 0
      "0000000" when "00001010001111001", -- t[5241] = 0
      "0000000" when "00001010001111010", -- t[5242] = 0
      "0000000" when "00001010001111011", -- t[5243] = 0
      "0000000" when "00001010001111100", -- t[5244] = 0
      "0000000" when "00001010001111101", -- t[5245] = 0
      "0000000" when "00001010001111110", -- t[5246] = 0
      "0000000" when "00001010001111111", -- t[5247] = 0
      "0000000" when "00001010010000000", -- t[5248] = 0
      "0000000" when "00001010010000001", -- t[5249] = 0
      "0000000" when "00001010010000010", -- t[5250] = 0
      "0000000" when "00001010010000011", -- t[5251] = 0
      "0000000" when "00001010010000100", -- t[5252] = 0
      "0000000" when "00001010010000101", -- t[5253] = 0
      "0000000" when "00001010010000110", -- t[5254] = 0
      "0000000" when "00001010010000111", -- t[5255] = 0
      "0000000" when "00001010010001000", -- t[5256] = 0
      "0000000" when "00001010010001001", -- t[5257] = 0
      "0000000" when "00001010010001010", -- t[5258] = 0
      "0000000" when "00001010010001011", -- t[5259] = 0
      "0000000" when "00001010010001100", -- t[5260] = 0
      "0000000" when "00001010010001101", -- t[5261] = 0
      "0000000" when "00001010010001110", -- t[5262] = 0
      "0000000" when "00001010010001111", -- t[5263] = 0
      "0000000" when "00001010010010000", -- t[5264] = 0
      "0000000" when "00001010010010001", -- t[5265] = 0
      "0000000" when "00001010010010010", -- t[5266] = 0
      "0000000" when "00001010010010011", -- t[5267] = 0
      "0000000" when "00001010010010100", -- t[5268] = 0
      "0000000" when "00001010010010101", -- t[5269] = 0
      "0000000" when "00001010010010110", -- t[5270] = 0
      "0000000" when "00001010010010111", -- t[5271] = 0
      "0000000" when "00001010010011000", -- t[5272] = 0
      "0000000" when "00001010010011001", -- t[5273] = 0
      "0000000" when "00001010010011010", -- t[5274] = 0
      "0000000" when "00001010010011011", -- t[5275] = 0
      "0000000" when "00001010010011100", -- t[5276] = 0
      "0000000" when "00001010010011101", -- t[5277] = 0
      "0000000" when "00001010010011110", -- t[5278] = 0
      "0000000" when "00001010010011111", -- t[5279] = 0
      "0000000" when "00001010010100000", -- t[5280] = 0
      "0000000" when "00001010010100001", -- t[5281] = 0
      "0000000" when "00001010010100010", -- t[5282] = 0
      "0000000" when "00001010010100011", -- t[5283] = 0
      "0000000" when "00001010010100100", -- t[5284] = 0
      "0000000" when "00001010010100101", -- t[5285] = 0
      "0000000" when "00001010010100110", -- t[5286] = 0
      "0000000" when "00001010010100111", -- t[5287] = 0
      "0000000" when "00001010010101000", -- t[5288] = 0
      "0000000" when "00001010010101001", -- t[5289] = 0
      "0000000" when "00001010010101010", -- t[5290] = 0
      "0000000" when "00001010010101011", -- t[5291] = 0
      "0000000" when "00001010010101100", -- t[5292] = 0
      "0000000" when "00001010010101101", -- t[5293] = 0
      "0000000" when "00001010010101110", -- t[5294] = 0
      "0000000" when "00001010010101111", -- t[5295] = 0
      "0000000" when "00001010010110000", -- t[5296] = 0
      "0000000" when "00001010010110001", -- t[5297] = 0
      "0000000" when "00001010010110010", -- t[5298] = 0
      "0000000" when "00001010010110011", -- t[5299] = 0
      "0000000" when "00001010010110100", -- t[5300] = 0
      "0000000" when "00001010010110101", -- t[5301] = 0
      "0000000" when "00001010010110110", -- t[5302] = 0
      "0000000" when "00001010010110111", -- t[5303] = 0
      "0000000" when "00001010010111000", -- t[5304] = 0
      "0000000" when "00001010010111001", -- t[5305] = 0
      "0000000" when "00001010010111010", -- t[5306] = 0
      "0000000" when "00001010010111011", -- t[5307] = 0
      "0000000" when "00001010010111100", -- t[5308] = 0
      "0000000" when "00001010010111101", -- t[5309] = 0
      "0000000" when "00001010010111110", -- t[5310] = 0
      "0000000" when "00001010010111111", -- t[5311] = 0
      "0000000" when "00001010011000000", -- t[5312] = 0
      "0000000" when "00001010011000001", -- t[5313] = 0
      "0000000" when "00001010011000010", -- t[5314] = 0
      "0000000" when "00001010011000011", -- t[5315] = 0
      "0000000" when "00001010011000100", -- t[5316] = 0
      "0000000" when "00001010011000101", -- t[5317] = 0
      "0000000" when "00001010011000110", -- t[5318] = 0
      "0000000" when "00001010011000111", -- t[5319] = 0
      "0000000" when "00001010011001000", -- t[5320] = 0
      "0000000" when "00001010011001001", -- t[5321] = 0
      "0000000" when "00001010011001010", -- t[5322] = 0
      "0000000" when "00001010011001011", -- t[5323] = 0
      "0000000" when "00001010011001100", -- t[5324] = 0
      "0000000" when "00001010011001101", -- t[5325] = 0
      "0000000" when "00001010011001110", -- t[5326] = 0
      "0000000" when "00001010011001111", -- t[5327] = 0
      "0000000" when "00001010011010000", -- t[5328] = 0
      "0000000" when "00001010011010001", -- t[5329] = 0
      "0000000" when "00001010011010010", -- t[5330] = 0
      "0000000" when "00001010011010011", -- t[5331] = 0
      "0000000" when "00001010011010100", -- t[5332] = 0
      "0000000" when "00001010011010101", -- t[5333] = 0
      "0000000" when "00001010011010110", -- t[5334] = 0
      "0000000" when "00001010011010111", -- t[5335] = 0
      "0000000" when "00001010011011000", -- t[5336] = 0
      "0000000" when "00001010011011001", -- t[5337] = 0
      "0000000" when "00001010011011010", -- t[5338] = 0
      "0000000" when "00001010011011011", -- t[5339] = 0
      "0000000" when "00001010011011100", -- t[5340] = 0
      "0000000" when "00001010011011101", -- t[5341] = 0
      "0000000" when "00001010011011110", -- t[5342] = 0
      "0000000" when "00001010011011111", -- t[5343] = 0
      "0000000" when "00001010011100000", -- t[5344] = 0
      "0000000" when "00001010011100001", -- t[5345] = 0
      "0000000" when "00001010011100010", -- t[5346] = 0
      "0000000" when "00001010011100011", -- t[5347] = 0
      "0000000" when "00001010011100100", -- t[5348] = 0
      "0000000" when "00001010011100101", -- t[5349] = 0
      "0000000" when "00001010011100110", -- t[5350] = 0
      "0000000" when "00001010011100111", -- t[5351] = 0
      "0000000" when "00001010011101000", -- t[5352] = 0
      "0000000" when "00001010011101001", -- t[5353] = 0
      "0000000" when "00001010011101010", -- t[5354] = 0
      "0000000" when "00001010011101011", -- t[5355] = 0
      "0000000" when "00001010011101100", -- t[5356] = 0
      "0000000" when "00001010011101101", -- t[5357] = 0
      "0000000" when "00001010011101110", -- t[5358] = 0
      "0000000" when "00001010011101111", -- t[5359] = 0
      "0000000" when "00001010011110000", -- t[5360] = 0
      "0000000" when "00001010011110001", -- t[5361] = 0
      "0000000" when "00001010011110010", -- t[5362] = 0
      "0000000" when "00001010011110011", -- t[5363] = 0
      "0000000" when "00001010011110100", -- t[5364] = 0
      "0000000" when "00001010011110101", -- t[5365] = 0
      "0000000" when "00001010011110110", -- t[5366] = 0
      "0000000" when "00001010011110111", -- t[5367] = 0
      "0000000" when "00001010011111000", -- t[5368] = 0
      "0000000" when "00001010011111001", -- t[5369] = 0
      "0000000" when "00001010011111010", -- t[5370] = 0
      "0000000" when "00001010011111011", -- t[5371] = 0
      "0000000" when "00001010011111100", -- t[5372] = 0
      "0000000" when "00001010011111101", -- t[5373] = 0
      "0000000" when "00001010011111110", -- t[5374] = 0
      "0000000" when "00001010011111111", -- t[5375] = 0
      "0000000" when "00001010100000000", -- t[5376] = 0
      "0000000" when "00001010100000001", -- t[5377] = 0
      "0000000" when "00001010100000010", -- t[5378] = 0
      "0000000" when "00001010100000011", -- t[5379] = 0
      "0000000" when "00001010100000100", -- t[5380] = 0
      "0000000" when "00001010100000101", -- t[5381] = 0
      "0000000" when "00001010100000110", -- t[5382] = 0
      "0000000" when "00001010100000111", -- t[5383] = 0
      "0000000" when "00001010100001000", -- t[5384] = 0
      "0000000" when "00001010100001001", -- t[5385] = 0
      "0000000" when "00001010100001010", -- t[5386] = 0
      "0000000" when "00001010100001011", -- t[5387] = 0
      "0000000" when "00001010100001100", -- t[5388] = 0
      "0000000" when "00001010100001101", -- t[5389] = 0
      "0000000" when "00001010100001110", -- t[5390] = 0
      "0000000" when "00001010100001111", -- t[5391] = 0
      "0000000" when "00001010100010000", -- t[5392] = 0
      "0000000" when "00001010100010001", -- t[5393] = 0
      "0000000" when "00001010100010010", -- t[5394] = 0
      "0000000" when "00001010100010011", -- t[5395] = 0
      "0000000" when "00001010100010100", -- t[5396] = 0
      "0000000" when "00001010100010101", -- t[5397] = 0
      "0000000" when "00001010100010110", -- t[5398] = 0
      "0000000" when "00001010100010111", -- t[5399] = 0
      "0000000" when "00001010100011000", -- t[5400] = 0
      "0000000" when "00001010100011001", -- t[5401] = 0
      "0000000" when "00001010100011010", -- t[5402] = 0
      "0000000" when "00001010100011011", -- t[5403] = 0
      "0000000" when "00001010100011100", -- t[5404] = 0
      "0000000" when "00001010100011101", -- t[5405] = 0
      "0000000" when "00001010100011110", -- t[5406] = 0
      "0000000" when "00001010100011111", -- t[5407] = 0
      "0000000" when "00001010100100000", -- t[5408] = 0
      "0000000" when "00001010100100001", -- t[5409] = 0
      "0000000" when "00001010100100010", -- t[5410] = 0
      "0000000" when "00001010100100011", -- t[5411] = 0
      "0000000" when "00001010100100100", -- t[5412] = 0
      "0000000" when "00001010100100101", -- t[5413] = 0
      "0000000" when "00001010100100110", -- t[5414] = 0
      "0000000" when "00001010100100111", -- t[5415] = 0
      "0000000" when "00001010100101000", -- t[5416] = 0
      "0000000" when "00001010100101001", -- t[5417] = 0
      "0000000" when "00001010100101010", -- t[5418] = 0
      "0000000" when "00001010100101011", -- t[5419] = 0
      "0000000" when "00001010100101100", -- t[5420] = 0
      "0000000" when "00001010100101101", -- t[5421] = 0
      "0000000" when "00001010100101110", -- t[5422] = 0
      "0000000" when "00001010100101111", -- t[5423] = 0
      "0000000" when "00001010100110000", -- t[5424] = 0
      "0000000" when "00001010100110001", -- t[5425] = 0
      "0000000" when "00001010100110010", -- t[5426] = 0
      "0000000" when "00001010100110011", -- t[5427] = 0
      "0000000" when "00001010100110100", -- t[5428] = 0
      "0000000" when "00001010100110101", -- t[5429] = 0
      "0000000" when "00001010100110110", -- t[5430] = 0
      "0000000" when "00001010100110111", -- t[5431] = 0
      "0000000" when "00001010100111000", -- t[5432] = 0
      "0000000" when "00001010100111001", -- t[5433] = 0
      "0000000" when "00001010100111010", -- t[5434] = 0
      "0000000" when "00001010100111011", -- t[5435] = 0
      "0000000" when "00001010100111100", -- t[5436] = 0
      "0000000" when "00001010100111101", -- t[5437] = 0
      "0000000" when "00001010100111110", -- t[5438] = 0
      "0000000" when "00001010100111111", -- t[5439] = 0
      "0000000" when "00001010101000000", -- t[5440] = 0
      "0000000" when "00001010101000001", -- t[5441] = 0
      "0000000" when "00001010101000010", -- t[5442] = 0
      "0000000" when "00001010101000011", -- t[5443] = 0
      "0000000" when "00001010101000100", -- t[5444] = 0
      "0000000" when "00001010101000101", -- t[5445] = 0
      "0000000" when "00001010101000110", -- t[5446] = 0
      "0000000" when "00001010101000111", -- t[5447] = 0
      "0000000" when "00001010101001000", -- t[5448] = 0
      "0000000" when "00001010101001001", -- t[5449] = 0
      "0000000" when "00001010101001010", -- t[5450] = 0
      "0000000" when "00001010101001011", -- t[5451] = 0
      "0000000" when "00001010101001100", -- t[5452] = 0
      "0000000" when "00001010101001101", -- t[5453] = 0
      "0000000" when "00001010101001110", -- t[5454] = 0
      "0000000" when "00001010101001111", -- t[5455] = 0
      "0000000" when "00001010101010000", -- t[5456] = 0
      "0000000" when "00001010101010001", -- t[5457] = 0
      "0000000" when "00001010101010010", -- t[5458] = 0
      "0000000" when "00001010101010011", -- t[5459] = 0
      "0000000" when "00001010101010100", -- t[5460] = 0
      "0000000" when "00001010101010101", -- t[5461] = 0
      "0000000" when "00001010101010110", -- t[5462] = 0
      "0000000" when "00001010101010111", -- t[5463] = 0
      "0000000" when "00001010101011000", -- t[5464] = 0
      "0000000" when "00001010101011001", -- t[5465] = 0
      "0000000" when "00001010101011010", -- t[5466] = 0
      "0000000" when "00001010101011011", -- t[5467] = 0
      "0000000" when "00001010101011100", -- t[5468] = 0
      "0000000" when "00001010101011101", -- t[5469] = 0
      "0000000" when "00001010101011110", -- t[5470] = 0
      "0000000" when "00001010101011111", -- t[5471] = 0
      "0000000" when "00001010101100000", -- t[5472] = 0
      "0000000" when "00001010101100001", -- t[5473] = 0
      "0000000" when "00001010101100010", -- t[5474] = 0
      "0000000" when "00001010101100011", -- t[5475] = 0
      "0000000" when "00001010101100100", -- t[5476] = 0
      "0000000" when "00001010101100101", -- t[5477] = 0
      "0000000" when "00001010101100110", -- t[5478] = 0
      "0000000" when "00001010101100111", -- t[5479] = 0
      "0000000" when "00001010101101000", -- t[5480] = 0
      "0000000" when "00001010101101001", -- t[5481] = 0
      "0000000" when "00001010101101010", -- t[5482] = 0
      "0000000" when "00001010101101011", -- t[5483] = 0
      "0000000" when "00001010101101100", -- t[5484] = 0
      "0000000" when "00001010101101101", -- t[5485] = 0
      "0000000" when "00001010101101110", -- t[5486] = 0
      "0000000" when "00001010101101111", -- t[5487] = 0
      "0000000" when "00001010101110000", -- t[5488] = 0
      "0000000" when "00001010101110001", -- t[5489] = 0
      "0000000" when "00001010101110010", -- t[5490] = 0
      "0000000" when "00001010101110011", -- t[5491] = 0
      "0000000" when "00001010101110100", -- t[5492] = 0
      "0000000" when "00001010101110101", -- t[5493] = 0
      "0000000" when "00001010101110110", -- t[5494] = 0
      "0000000" when "00001010101110111", -- t[5495] = 0
      "0000000" when "00001010101111000", -- t[5496] = 0
      "0000000" when "00001010101111001", -- t[5497] = 0
      "0000000" when "00001010101111010", -- t[5498] = 0
      "0000000" when "00001010101111011", -- t[5499] = 0
      "0000000" when "00001010101111100", -- t[5500] = 0
      "0000000" when "00001010101111101", -- t[5501] = 0
      "0000000" when "00001010101111110", -- t[5502] = 0
      "0000000" when "00001010101111111", -- t[5503] = 0
      "0000000" when "00001010110000000", -- t[5504] = 0
      "0000000" when "00001010110000001", -- t[5505] = 0
      "0000000" when "00001010110000010", -- t[5506] = 0
      "0000000" when "00001010110000011", -- t[5507] = 0
      "0000000" when "00001010110000100", -- t[5508] = 0
      "0000000" when "00001010110000101", -- t[5509] = 0
      "0000000" when "00001010110000110", -- t[5510] = 0
      "0000000" when "00001010110000111", -- t[5511] = 0
      "0000000" when "00001010110001000", -- t[5512] = 0
      "0000000" when "00001010110001001", -- t[5513] = 0
      "0000000" when "00001010110001010", -- t[5514] = 0
      "0000000" when "00001010110001011", -- t[5515] = 0
      "0000000" when "00001010110001100", -- t[5516] = 0
      "0000000" when "00001010110001101", -- t[5517] = 0
      "0000000" when "00001010110001110", -- t[5518] = 0
      "0000000" when "00001010110001111", -- t[5519] = 0
      "0000000" when "00001010110010000", -- t[5520] = 0
      "0000000" when "00001010110010001", -- t[5521] = 0
      "0000000" when "00001010110010010", -- t[5522] = 0
      "0000000" when "00001010110010011", -- t[5523] = 0
      "0000000" when "00001010110010100", -- t[5524] = 0
      "0000000" when "00001010110010101", -- t[5525] = 0
      "0000000" when "00001010110010110", -- t[5526] = 0
      "0000000" when "00001010110010111", -- t[5527] = 0
      "0000000" when "00001010110011000", -- t[5528] = 0
      "0000000" when "00001010110011001", -- t[5529] = 0
      "0000000" when "00001010110011010", -- t[5530] = 0
      "0000000" when "00001010110011011", -- t[5531] = 0
      "0000000" when "00001010110011100", -- t[5532] = 0
      "0000000" when "00001010110011101", -- t[5533] = 0
      "0000000" when "00001010110011110", -- t[5534] = 0
      "0000000" when "00001010110011111", -- t[5535] = 0
      "0000000" when "00001010110100000", -- t[5536] = 0
      "0000000" when "00001010110100001", -- t[5537] = 0
      "0000000" when "00001010110100010", -- t[5538] = 0
      "0000000" when "00001010110100011", -- t[5539] = 0
      "0000000" when "00001010110100100", -- t[5540] = 0
      "0000000" when "00001010110100101", -- t[5541] = 0
      "0000000" when "00001010110100110", -- t[5542] = 0
      "0000000" when "00001010110100111", -- t[5543] = 0
      "0000000" when "00001010110101000", -- t[5544] = 0
      "0000000" when "00001010110101001", -- t[5545] = 0
      "0000000" when "00001010110101010", -- t[5546] = 0
      "0000000" when "00001010110101011", -- t[5547] = 0
      "0000000" when "00001010110101100", -- t[5548] = 0
      "0000000" when "00001010110101101", -- t[5549] = 0
      "0000000" when "00001010110101110", -- t[5550] = 0
      "0000000" when "00001010110101111", -- t[5551] = 0
      "0000000" when "00001010110110000", -- t[5552] = 0
      "0000000" when "00001010110110001", -- t[5553] = 0
      "0000000" when "00001010110110010", -- t[5554] = 0
      "0000000" when "00001010110110011", -- t[5555] = 0
      "0000000" when "00001010110110100", -- t[5556] = 0
      "0000000" when "00001010110110101", -- t[5557] = 0
      "0000000" when "00001010110110110", -- t[5558] = 0
      "0000000" when "00001010110110111", -- t[5559] = 0
      "0000000" when "00001010110111000", -- t[5560] = 0
      "0000000" when "00001010110111001", -- t[5561] = 0
      "0000000" when "00001010110111010", -- t[5562] = 0
      "0000000" when "00001010110111011", -- t[5563] = 0
      "0000000" when "00001010110111100", -- t[5564] = 0
      "0000000" when "00001010110111101", -- t[5565] = 0
      "0000000" when "00001010110111110", -- t[5566] = 0
      "0000000" when "00001010110111111", -- t[5567] = 0
      "0000000" when "00001010111000000", -- t[5568] = 0
      "0000000" when "00001010111000001", -- t[5569] = 0
      "0000000" when "00001010111000010", -- t[5570] = 0
      "0000000" when "00001010111000011", -- t[5571] = 0
      "0000000" when "00001010111000100", -- t[5572] = 0
      "0000000" when "00001010111000101", -- t[5573] = 0
      "0000000" when "00001010111000110", -- t[5574] = 0
      "0000000" when "00001010111000111", -- t[5575] = 0
      "0000000" when "00001010111001000", -- t[5576] = 0
      "0000000" when "00001010111001001", -- t[5577] = 0
      "0000000" when "00001010111001010", -- t[5578] = 0
      "0000000" when "00001010111001011", -- t[5579] = 0
      "0000000" when "00001010111001100", -- t[5580] = 0
      "0000000" when "00001010111001101", -- t[5581] = 0
      "0000000" when "00001010111001110", -- t[5582] = 0
      "0000000" when "00001010111001111", -- t[5583] = 0
      "0000000" when "00001010111010000", -- t[5584] = 0
      "0000000" when "00001010111010001", -- t[5585] = 0
      "0000000" when "00001010111010010", -- t[5586] = 0
      "0000000" when "00001010111010011", -- t[5587] = 0
      "0000000" when "00001010111010100", -- t[5588] = 0
      "0000000" when "00001010111010101", -- t[5589] = 0
      "0000000" when "00001010111010110", -- t[5590] = 0
      "0000000" when "00001010111010111", -- t[5591] = 0
      "0000000" when "00001010111011000", -- t[5592] = 0
      "0000000" when "00001010111011001", -- t[5593] = 0
      "0000000" when "00001010111011010", -- t[5594] = 0
      "0000000" when "00001010111011011", -- t[5595] = 0
      "0000000" when "00001010111011100", -- t[5596] = 0
      "0000000" when "00001010111011101", -- t[5597] = 0
      "0000000" when "00001010111011110", -- t[5598] = 0
      "0000000" when "00001010111011111", -- t[5599] = 0
      "0000000" when "00001010111100000", -- t[5600] = 0
      "0000000" when "00001010111100001", -- t[5601] = 0
      "0000000" when "00001010111100010", -- t[5602] = 0
      "0000000" when "00001010111100011", -- t[5603] = 0
      "0000000" when "00001010111100100", -- t[5604] = 0
      "0000000" when "00001010111100101", -- t[5605] = 0
      "0000000" when "00001010111100110", -- t[5606] = 0
      "0000000" when "00001010111100111", -- t[5607] = 0
      "0000000" when "00001010111101000", -- t[5608] = 0
      "0000000" when "00001010111101001", -- t[5609] = 0
      "0000000" when "00001010111101010", -- t[5610] = 0
      "0000000" when "00001010111101011", -- t[5611] = 0
      "0000000" when "00001010111101100", -- t[5612] = 0
      "0000000" when "00001010111101101", -- t[5613] = 0
      "0000000" when "00001010111101110", -- t[5614] = 0
      "0000000" when "00001010111101111", -- t[5615] = 0
      "0000000" when "00001010111110000", -- t[5616] = 0
      "0000000" when "00001010111110001", -- t[5617] = 0
      "0000000" when "00001010111110010", -- t[5618] = 0
      "0000000" when "00001010111110011", -- t[5619] = 0
      "0000000" when "00001010111110100", -- t[5620] = 0
      "0000000" when "00001010111110101", -- t[5621] = 0
      "0000000" when "00001010111110110", -- t[5622] = 0
      "0000000" when "00001010111110111", -- t[5623] = 0
      "0000000" when "00001010111111000", -- t[5624] = 0
      "0000000" when "00001010111111001", -- t[5625] = 0
      "0000000" when "00001010111111010", -- t[5626] = 0
      "0000000" when "00001010111111011", -- t[5627] = 0
      "0000000" when "00001010111111100", -- t[5628] = 0
      "0000000" when "00001010111111101", -- t[5629] = 0
      "0000000" when "00001010111111110", -- t[5630] = 0
      "0000000" when "00001010111111111", -- t[5631] = 0
      "0000000" when "00001011000000000", -- t[5632] = 0
      "0000000" when "00001011000000001", -- t[5633] = 0
      "0000000" when "00001011000000010", -- t[5634] = 0
      "0000000" when "00001011000000011", -- t[5635] = 0
      "0000000" when "00001011000000100", -- t[5636] = 0
      "0000000" when "00001011000000101", -- t[5637] = 0
      "0000000" when "00001011000000110", -- t[5638] = 0
      "0000000" when "00001011000000111", -- t[5639] = 0
      "0000000" when "00001011000001000", -- t[5640] = 0
      "0000000" when "00001011000001001", -- t[5641] = 0
      "0000000" when "00001011000001010", -- t[5642] = 0
      "0000000" when "00001011000001011", -- t[5643] = 0
      "0000000" when "00001011000001100", -- t[5644] = 0
      "0000000" when "00001011000001101", -- t[5645] = 0
      "0000000" when "00001011000001110", -- t[5646] = 0
      "0000000" when "00001011000001111", -- t[5647] = 0
      "0000000" when "00001011000010000", -- t[5648] = 0
      "0000000" when "00001011000010001", -- t[5649] = 0
      "0000000" when "00001011000010010", -- t[5650] = 0
      "0000000" when "00001011000010011", -- t[5651] = 0
      "0000000" when "00001011000010100", -- t[5652] = 0
      "0000000" when "00001011000010101", -- t[5653] = 0
      "0000000" when "00001011000010110", -- t[5654] = 0
      "0000000" when "00001011000010111", -- t[5655] = 0
      "0000000" when "00001011000011000", -- t[5656] = 0
      "0000000" when "00001011000011001", -- t[5657] = 0
      "0000000" when "00001011000011010", -- t[5658] = 0
      "0000000" when "00001011000011011", -- t[5659] = 0
      "0000000" when "00001011000011100", -- t[5660] = 0
      "0000000" when "00001011000011101", -- t[5661] = 0
      "0000000" when "00001011000011110", -- t[5662] = 0
      "0000000" when "00001011000011111", -- t[5663] = 0
      "0000000" when "00001011000100000", -- t[5664] = 0
      "0000000" when "00001011000100001", -- t[5665] = 0
      "0000000" when "00001011000100010", -- t[5666] = 0
      "0000000" when "00001011000100011", -- t[5667] = 0
      "0000000" when "00001011000100100", -- t[5668] = 0
      "0000000" when "00001011000100101", -- t[5669] = 0
      "0000000" when "00001011000100110", -- t[5670] = 0
      "0000000" when "00001011000100111", -- t[5671] = 0
      "0000000" when "00001011000101000", -- t[5672] = 0
      "0000000" when "00001011000101001", -- t[5673] = 0
      "0000000" when "00001011000101010", -- t[5674] = 0
      "0000000" when "00001011000101011", -- t[5675] = 0
      "0000000" when "00001011000101100", -- t[5676] = 0
      "0000000" when "00001011000101101", -- t[5677] = 0
      "0000000" when "00001011000101110", -- t[5678] = 0
      "0000000" when "00001011000101111", -- t[5679] = 0
      "0000000" when "00001011000110000", -- t[5680] = 0
      "0000000" when "00001011000110001", -- t[5681] = 0
      "0000000" when "00001011000110010", -- t[5682] = 0
      "0000000" when "00001011000110011", -- t[5683] = 0
      "0000000" when "00001011000110100", -- t[5684] = 0
      "0000000" when "00001011000110101", -- t[5685] = 0
      "0000000" when "00001011000110110", -- t[5686] = 0
      "0000000" when "00001011000110111", -- t[5687] = 0
      "0000000" when "00001011000111000", -- t[5688] = 0
      "0000000" when "00001011000111001", -- t[5689] = 0
      "0000000" when "00001011000111010", -- t[5690] = 0
      "0000000" when "00001011000111011", -- t[5691] = 0
      "0000000" when "00001011000111100", -- t[5692] = 0
      "0000000" when "00001011000111101", -- t[5693] = 0
      "0000000" when "00001011000111110", -- t[5694] = 0
      "0000000" when "00001011000111111", -- t[5695] = 0
      "0000000" when "00001011001000000", -- t[5696] = 0
      "0000000" when "00001011001000001", -- t[5697] = 0
      "0000000" when "00001011001000010", -- t[5698] = 0
      "0000000" when "00001011001000011", -- t[5699] = 0
      "0000000" when "00001011001000100", -- t[5700] = 0
      "0000000" when "00001011001000101", -- t[5701] = 0
      "0000000" when "00001011001000110", -- t[5702] = 0
      "0000000" when "00001011001000111", -- t[5703] = 0
      "0000000" when "00001011001001000", -- t[5704] = 0
      "0000000" when "00001011001001001", -- t[5705] = 0
      "0000000" when "00001011001001010", -- t[5706] = 0
      "0000000" when "00001011001001011", -- t[5707] = 0
      "0000000" when "00001011001001100", -- t[5708] = 0
      "0000000" when "00001011001001101", -- t[5709] = 0
      "0000000" when "00001011001001110", -- t[5710] = 0
      "0000000" when "00001011001001111", -- t[5711] = 0
      "0000000" when "00001011001010000", -- t[5712] = 0
      "0000000" when "00001011001010001", -- t[5713] = 0
      "0000000" when "00001011001010010", -- t[5714] = 0
      "0000000" when "00001011001010011", -- t[5715] = 0
      "0000000" when "00001011001010100", -- t[5716] = 0
      "0000000" when "00001011001010101", -- t[5717] = 0
      "0000000" when "00001011001010110", -- t[5718] = 0
      "0000000" when "00001011001010111", -- t[5719] = 0
      "0000000" when "00001011001011000", -- t[5720] = 0
      "0000000" when "00001011001011001", -- t[5721] = 0
      "0000000" when "00001011001011010", -- t[5722] = 0
      "0000000" when "00001011001011011", -- t[5723] = 0
      "0000000" when "00001011001011100", -- t[5724] = 0
      "0000000" when "00001011001011101", -- t[5725] = 0
      "0000000" when "00001011001011110", -- t[5726] = 0
      "0000000" when "00001011001011111", -- t[5727] = 0
      "0000000" when "00001011001100000", -- t[5728] = 0
      "0000000" when "00001011001100001", -- t[5729] = 0
      "0000000" when "00001011001100010", -- t[5730] = 0
      "0000000" when "00001011001100011", -- t[5731] = 0
      "0000000" when "00001011001100100", -- t[5732] = 0
      "0000000" when "00001011001100101", -- t[5733] = 0
      "0000000" when "00001011001100110", -- t[5734] = 0
      "0000000" when "00001011001100111", -- t[5735] = 0
      "0000000" when "00001011001101000", -- t[5736] = 0
      "0000000" when "00001011001101001", -- t[5737] = 0
      "0000000" when "00001011001101010", -- t[5738] = 0
      "0000000" when "00001011001101011", -- t[5739] = 0
      "0000000" when "00001011001101100", -- t[5740] = 0
      "0000000" when "00001011001101101", -- t[5741] = 0
      "0000000" when "00001011001101110", -- t[5742] = 0
      "0000000" when "00001011001101111", -- t[5743] = 0
      "0000000" when "00001011001110000", -- t[5744] = 0
      "0000000" when "00001011001110001", -- t[5745] = 0
      "0000000" when "00001011001110010", -- t[5746] = 0
      "0000000" when "00001011001110011", -- t[5747] = 0
      "0000000" when "00001011001110100", -- t[5748] = 0
      "0000000" when "00001011001110101", -- t[5749] = 0
      "0000000" when "00001011001110110", -- t[5750] = 0
      "0000000" when "00001011001110111", -- t[5751] = 0
      "0000000" when "00001011001111000", -- t[5752] = 0
      "0000000" when "00001011001111001", -- t[5753] = 0
      "0000000" when "00001011001111010", -- t[5754] = 0
      "0000000" when "00001011001111011", -- t[5755] = 0
      "0000000" when "00001011001111100", -- t[5756] = 0
      "0000000" when "00001011001111101", -- t[5757] = 0
      "0000000" when "00001011001111110", -- t[5758] = 0
      "0000000" when "00001011001111111", -- t[5759] = 0
      "0000000" when "00001011010000000", -- t[5760] = 0
      "0000000" when "00001011010000001", -- t[5761] = 0
      "0000000" when "00001011010000010", -- t[5762] = 0
      "0000000" when "00001011010000011", -- t[5763] = 0
      "0000000" when "00001011010000100", -- t[5764] = 0
      "0000000" when "00001011010000101", -- t[5765] = 0
      "0000000" when "00001011010000110", -- t[5766] = 0
      "0000000" when "00001011010000111", -- t[5767] = 0
      "0000000" when "00001011010001000", -- t[5768] = 0
      "0000000" when "00001011010001001", -- t[5769] = 0
      "0000000" when "00001011010001010", -- t[5770] = 0
      "0000000" when "00001011010001011", -- t[5771] = 0
      "0000000" when "00001011010001100", -- t[5772] = 0
      "0000000" when "00001011010001101", -- t[5773] = 0
      "0000000" when "00001011010001110", -- t[5774] = 0
      "0000000" when "00001011010001111", -- t[5775] = 0
      "0000000" when "00001011010010000", -- t[5776] = 0
      "0000000" when "00001011010010001", -- t[5777] = 0
      "0000000" when "00001011010010010", -- t[5778] = 0
      "0000000" when "00001011010010011", -- t[5779] = 0
      "0000000" when "00001011010010100", -- t[5780] = 0
      "0000000" when "00001011010010101", -- t[5781] = 0
      "0000000" when "00001011010010110", -- t[5782] = 0
      "0000000" when "00001011010010111", -- t[5783] = 0
      "0000000" when "00001011010011000", -- t[5784] = 0
      "0000000" when "00001011010011001", -- t[5785] = 0
      "0000000" when "00001011010011010", -- t[5786] = 0
      "0000000" when "00001011010011011", -- t[5787] = 0
      "0000000" when "00001011010011100", -- t[5788] = 0
      "0000000" when "00001011010011101", -- t[5789] = 0
      "0000000" when "00001011010011110", -- t[5790] = 0
      "0000000" when "00001011010011111", -- t[5791] = 0
      "0000000" when "00001011010100000", -- t[5792] = 0
      "0000000" when "00001011010100001", -- t[5793] = 0
      "0000000" when "00001011010100010", -- t[5794] = 0
      "0000000" when "00001011010100011", -- t[5795] = 0
      "0000000" when "00001011010100100", -- t[5796] = 0
      "0000000" when "00001011010100101", -- t[5797] = 0
      "0000000" when "00001011010100110", -- t[5798] = 0
      "0000000" when "00001011010100111", -- t[5799] = 0
      "0000000" when "00001011010101000", -- t[5800] = 0
      "0000000" when "00001011010101001", -- t[5801] = 0
      "0000000" when "00001011010101010", -- t[5802] = 0
      "0000000" when "00001011010101011", -- t[5803] = 0
      "0000000" when "00001011010101100", -- t[5804] = 0
      "0000000" when "00001011010101101", -- t[5805] = 0
      "0000000" when "00001011010101110", -- t[5806] = 0
      "0000000" when "00001011010101111", -- t[5807] = 0
      "0000000" when "00001011010110000", -- t[5808] = 0
      "0000000" when "00001011010110001", -- t[5809] = 0
      "0000000" when "00001011010110010", -- t[5810] = 0
      "0000000" when "00001011010110011", -- t[5811] = 0
      "0000000" when "00001011010110100", -- t[5812] = 0
      "0000000" when "00001011010110101", -- t[5813] = 0
      "0000000" when "00001011010110110", -- t[5814] = 0
      "0000000" when "00001011010110111", -- t[5815] = 0
      "0000000" when "00001011010111000", -- t[5816] = 0
      "0000000" when "00001011010111001", -- t[5817] = 0
      "0000000" when "00001011010111010", -- t[5818] = 0
      "0000000" when "00001011010111011", -- t[5819] = 0
      "0000000" when "00001011010111100", -- t[5820] = 0
      "0000000" when "00001011010111101", -- t[5821] = 0
      "0000000" when "00001011010111110", -- t[5822] = 0
      "0000000" when "00001011010111111", -- t[5823] = 0
      "0000000" when "00001011011000000", -- t[5824] = 0
      "0000000" when "00001011011000001", -- t[5825] = 0
      "0000000" when "00001011011000010", -- t[5826] = 0
      "0000000" when "00001011011000011", -- t[5827] = 0
      "0000000" when "00001011011000100", -- t[5828] = 0
      "0000000" when "00001011011000101", -- t[5829] = 0
      "0000000" when "00001011011000110", -- t[5830] = 0
      "0000000" when "00001011011000111", -- t[5831] = 0
      "0000000" when "00001011011001000", -- t[5832] = 0
      "0000000" when "00001011011001001", -- t[5833] = 0
      "0000000" when "00001011011001010", -- t[5834] = 0
      "0000000" when "00001011011001011", -- t[5835] = 0
      "0000000" when "00001011011001100", -- t[5836] = 0
      "0000000" when "00001011011001101", -- t[5837] = 0
      "0000000" when "00001011011001110", -- t[5838] = 0
      "0000000" when "00001011011001111", -- t[5839] = 0
      "0000000" when "00001011011010000", -- t[5840] = 0
      "0000000" when "00001011011010001", -- t[5841] = 0
      "0000000" when "00001011011010010", -- t[5842] = 0
      "0000000" when "00001011011010011", -- t[5843] = 0
      "0000000" when "00001011011010100", -- t[5844] = 0
      "0000000" when "00001011011010101", -- t[5845] = 0
      "0000000" when "00001011011010110", -- t[5846] = 0
      "0000000" when "00001011011010111", -- t[5847] = 0
      "0000000" when "00001011011011000", -- t[5848] = 0
      "0000000" when "00001011011011001", -- t[5849] = 0
      "0000000" when "00001011011011010", -- t[5850] = 0
      "0000000" when "00001011011011011", -- t[5851] = 0
      "0000000" when "00001011011011100", -- t[5852] = 0
      "0000000" when "00001011011011101", -- t[5853] = 0
      "0000000" when "00001011011011110", -- t[5854] = 0
      "0000000" when "00001011011011111", -- t[5855] = 0
      "0000000" when "00001011011100000", -- t[5856] = 0
      "0000000" when "00001011011100001", -- t[5857] = 0
      "0000000" when "00001011011100010", -- t[5858] = 0
      "0000000" when "00001011011100011", -- t[5859] = 0
      "0000000" when "00001011011100100", -- t[5860] = 0
      "0000000" when "00001011011100101", -- t[5861] = 0
      "0000000" when "00001011011100110", -- t[5862] = 0
      "0000000" when "00001011011100111", -- t[5863] = 0
      "0000000" when "00001011011101000", -- t[5864] = 0
      "0000000" when "00001011011101001", -- t[5865] = 0
      "0000000" when "00001011011101010", -- t[5866] = 0
      "0000000" when "00001011011101011", -- t[5867] = 0
      "0000000" when "00001011011101100", -- t[5868] = 0
      "0000000" when "00001011011101101", -- t[5869] = 0
      "0000000" when "00001011011101110", -- t[5870] = 0
      "0000000" when "00001011011101111", -- t[5871] = 0
      "0000000" when "00001011011110000", -- t[5872] = 0
      "0000000" when "00001011011110001", -- t[5873] = 0
      "0000000" when "00001011011110010", -- t[5874] = 0
      "0000000" when "00001011011110011", -- t[5875] = 0
      "0000000" when "00001011011110100", -- t[5876] = 0
      "0000000" when "00001011011110101", -- t[5877] = 0
      "0000000" when "00001011011110110", -- t[5878] = 0
      "0000000" when "00001011011110111", -- t[5879] = 0
      "0000000" when "00001011011111000", -- t[5880] = 0
      "0000000" when "00001011011111001", -- t[5881] = 0
      "0000000" when "00001011011111010", -- t[5882] = 0
      "0000000" when "00001011011111011", -- t[5883] = 0
      "0000000" when "00001011011111100", -- t[5884] = 0
      "0000000" when "00001011011111101", -- t[5885] = 0
      "0000000" when "00001011011111110", -- t[5886] = 0
      "0000000" when "00001011011111111", -- t[5887] = 0
      "0000000" when "00001011100000000", -- t[5888] = 0
      "0000000" when "00001011100000001", -- t[5889] = 0
      "0000000" when "00001011100000010", -- t[5890] = 0
      "0000000" when "00001011100000011", -- t[5891] = 0
      "0000000" when "00001011100000100", -- t[5892] = 0
      "0000000" when "00001011100000101", -- t[5893] = 0
      "0000000" when "00001011100000110", -- t[5894] = 0
      "0000000" when "00001011100000111", -- t[5895] = 0
      "0000000" when "00001011100001000", -- t[5896] = 0
      "0000000" when "00001011100001001", -- t[5897] = 0
      "0000000" when "00001011100001010", -- t[5898] = 0
      "0000000" when "00001011100001011", -- t[5899] = 0
      "0000000" when "00001011100001100", -- t[5900] = 0
      "0000000" when "00001011100001101", -- t[5901] = 0
      "0000000" when "00001011100001110", -- t[5902] = 0
      "0000000" when "00001011100001111", -- t[5903] = 0
      "0000000" when "00001011100010000", -- t[5904] = 0
      "0000000" when "00001011100010001", -- t[5905] = 0
      "0000000" when "00001011100010010", -- t[5906] = 0
      "0000000" when "00001011100010011", -- t[5907] = 0
      "0000000" when "00001011100010100", -- t[5908] = 0
      "0000000" when "00001011100010101", -- t[5909] = 0
      "0000000" when "00001011100010110", -- t[5910] = 0
      "0000000" when "00001011100010111", -- t[5911] = 0
      "0000000" when "00001011100011000", -- t[5912] = 0
      "0000000" when "00001011100011001", -- t[5913] = 0
      "0000000" when "00001011100011010", -- t[5914] = 0
      "0000000" when "00001011100011011", -- t[5915] = 0
      "0000000" when "00001011100011100", -- t[5916] = 0
      "0000000" when "00001011100011101", -- t[5917] = 0
      "0000000" when "00001011100011110", -- t[5918] = 0
      "0000000" when "00001011100011111", -- t[5919] = 0
      "0000000" when "00001011100100000", -- t[5920] = 0
      "0000000" when "00001011100100001", -- t[5921] = 0
      "0000000" when "00001011100100010", -- t[5922] = 0
      "0000000" when "00001011100100011", -- t[5923] = 0
      "0000000" when "00001011100100100", -- t[5924] = 0
      "0000000" when "00001011100100101", -- t[5925] = 0
      "0000000" when "00001011100100110", -- t[5926] = 0
      "0000000" when "00001011100100111", -- t[5927] = 0
      "0000000" when "00001011100101000", -- t[5928] = 0
      "0000000" when "00001011100101001", -- t[5929] = 0
      "0000000" when "00001011100101010", -- t[5930] = 0
      "0000000" when "00001011100101011", -- t[5931] = 0
      "0000000" when "00001011100101100", -- t[5932] = 0
      "0000000" when "00001011100101101", -- t[5933] = 0
      "0000000" when "00001011100101110", -- t[5934] = 0
      "0000000" when "00001011100101111", -- t[5935] = 0
      "0000000" when "00001011100110000", -- t[5936] = 0
      "0000000" when "00001011100110001", -- t[5937] = 0
      "0000000" when "00001011100110010", -- t[5938] = 0
      "0000000" when "00001011100110011", -- t[5939] = 0
      "0000000" when "00001011100110100", -- t[5940] = 0
      "0000000" when "00001011100110101", -- t[5941] = 0
      "0000000" when "00001011100110110", -- t[5942] = 0
      "0000000" when "00001011100110111", -- t[5943] = 0
      "0000000" when "00001011100111000", -- t[5944] = 0
      "0000000" when "00001011100111001", -- t[5945] = 0
      "0000000" when "00001011100111010", -- t[5946] = 0
      "0000000" when "00001011100111011", -- t[5947] = 0
      "0000000" when "00001011100111100", -- t[5948] = 0
      "0000000" when "00001011100111101", -- t[5949] = 0
      "0000000" when "00001011100111110", -- t[5950] = 0
      "0000000" when "00001011100111111", -- t[5951] = 0
      "0000000" when "00001011101000000", -- t[5952] = 0
      "0000000" when "00001011101000001", -- t[5953] = 0
      "0000000" when "00001011101000010", -- t[5954] = 0
      "0000000" when "00001011101000011", -- t[5955] = 0
      "0000000" when "00001011101000100", -- t[5956] = 0
      "0000000" when "00001011101000101", -- t[5957] = 0
      "0000000" when "00001011101000110", -- t[5958] = 0
      "0000000" when "00001011101000111", -- t[5959] = 0
      "0000000" when "00001011101001000", -- t[5960] = 0
      "0000000" when "00001011101001001", -- t[5961] = 0
      "0000000" when "00001011101001010", -- t[5962] = 0
      "0000000" when "00001011101001011", -- t[5963] = 0
      "0000000" when "00001011101001100", -- t[5964] = 0
      "0000000" when "00001011101001101", -- t[5965] = 0
      "0000000" when "00001011101001110", -- t[5966] = 0
      "0000000" when "00001011101001111", -- t[5967] = 0
      "0000000" when "00001011101010000", -- t[5968] = 0
      "0000000" when "00001011101010001", -- t[5969] = 0
      "0000000" when "00001011101010010", -- t[5970] = 0
      "0000000" when "00001011101010011", -- t[5971] = 0
      "0000000" when "00001011101010100", -- t[5972] = 0
      "0000000" when "00001011101010101", -- t[5973] = 0
      "0000000" when "00001011101010110", -- t[5974] = 0
      "0000000" when "00001011101010111", -- t[5975] = 0
      "0000000" when "00001011101011000", -- t[5976] = 0
      "0000000" when "00001011101011001", -- t[5977] = 0
      "0000000" when "00001011101011010", -- t[5978] = 0
      "0000000" when "00001011101011011", -- t[5979] = 0
      "0000000" when "00001011101011100", -- t[5980] = 0
      "0000000" when "00001011101011101", -- t[5981] = 0
      "0000000" when "00001011101011110", -- t[5982] = 0
      "0000000" when "00001011101011111", -- t[5983] = 0
      "0000000" when "00001011101100000", -- t[5984] = 0
      "0000000" when "00001011101100001", -- t[5985] = 0
      "0000000" when "00001011101100010", -- t[5986] = 0
      "0000000" when "00001011101100011", -- t[5987] = 0
      "0000000" when "00001011101100100", -- t[5988] = 0
      "0000000" when "00001011101100101", -- t[5989] = 0
      "0000000" when "00001011101100110", -- t[5990] = 0
      "0000000" when "00001011101100111", -- t[5991] = 0
      "0000000" when "00001011101101000", -- t[5992] = 0
      "0000000" when "00001011101101001", -- t[5993] = 0
      "0000000" when "00001011101101010", -- t[5994] = 0
      "0000000" when "00001011101101011", -- t[5995] = 0
      "0000000" when "00001011101101100", -- t[5996] = 0
      "0000000" when "00001011101101101", -- t[5997] = 0
      "0000000" when "00001011101101110", -- t[5998] = 0
      "0000000" when "00001011101101111", -- t[5999] = 0
      "0000000" when "00001011101110000", -- t[6000] = 0
      "0000000" when "00001011101110001", -- t[6001] = 0
      "0000000" when "00001011101110010", -- t[6002] = 0
      "0000000" when "00001011101110011", -- t[6003] = 0
      "0000000" when "00001011101110100", -- t[6004] = 0
      "0000000" when "00001011101110101", -- t[6005] = 0
      "0000000" when "00001011101110110", -- t[6006] = 0
      "0000000" when "00001011101110111", -- t[6007] = 0
      "0000000" when "00001011101111000", -- t[6008] = 0
      "0000000" when "00001011101111001", -- t[6009] = 0
      "0000000" when "00001011101111010", -- t[6010] = 0
      "0000000" when "00001011101111011", -- t[6011] = 0
      "0000000" when "00001011101111100", -- t[6012] = 0
      "0000000" when "00001011101111101", -- t[6013] = 0
      "0000000" when "00001011101111110", -- t[6014] = 0
      "0000000" when "00001011101111111", -- t[6015] = 0
      "0000000" when "00001011110000000", -- t[6016] = 0
      "0000000" when "00001011110000001", -- t[6017] = 0
      "0000000" when "00001011110000010", -- t[6018] = 0
      "0000000" when "00001011110000011", -- t[6019] = 0
      "0000000" when "00001011110000100", -- t[6020] = 0
      "0000000" when "00001011110000101", -- t[6021] = 0
      "0000000" when "00001011110000110", -- t[6022] = 0
      "0000000" when "00001011110000111", -- t[6023] = 0
      "0000000" when "00001011110001000", -- t[6024] = 0
      "0000000" when "00001011110001001", -- t[6025] = 0
      "0000000" when "00001011110001010", -- t[6026] = 0
      "0000000" when "00001011110001011", -- t[6027] = 0
      "0000000" when "00001011110001100", -- t[6028] = 0
      "0000000" when "00001011110001101", -- t[6029] = 0
      "0000000" when "00001011110001110", -- t[6030] = 0
      "0000000" when "00001011110001111", -- t[6031] = 0
      "0000000" when "00001011110010000", -- t[6032] = 0
      "0000000" when "00001011110010001", -- t[6033] = 0
      "0000000" when "00001011110010010", -- t[6034] = 0
      "0000000" when "00001011110010011", -- t[6035] = 0
      "0000000" when "00001011110010100", -- t[6036] = 0
      "0000000" when "00001011110010101", -- t[6037] = 0
      "0000000" when "00001011110010110", -- t[6038] = 0
      "0000000" when "00001011110010111", -- t[6039] = 0
      "0000000" when "00001011110011000", -- t[6040] = 0
      "0000000" when "00001011110011001", -- t[6041] = 0
      "0000000" when "00001011110011010", -- t[6042] = 0
      "0000000" when "00001011110011011", -- t[6043] = 0
      "0000000" when "00001011110011100", -- t[6044] = 0
      "0000000" when "00001011110011101", -- t[6045] = 0
      "0000000" when "00001011110011110", -- t[6046] = 0
      "0000000" when "00001011110011111", -- t[6047] = 0
      "0000000" when "00001011110100000", -- t[6048] = 0
      "0000000" when "00001011110100001", -- t[6049] = 0
      "0000000" when "00001011110100010", -- t[6050] = 0
      "0000000" when "00001011110100011", -- t[6051] = 0
      "0000000" when "00001011110100100", -- t[6052] = 0
      "0000000" when "00001011110100101", -- t[6053] = 0
      "0000000" when "00001011110100110", -- t[6054] = 0
      "0000000" when "00001011110100111", -- t[6055] = 0
      "0000000" when "00001011110101000", -- t[6056] = 0
      "0000000" when "00001011110101001", -- t[6057] = 0
      "0000000" when "00001011110101010", -- t[6058] = 0
      "0000000" when "00001011110101011", -- t[6059] = 0
      "0000000" when "00001011110101100", -- t[6060] = 0
      "0000000" when "00001011110101101", -- t[6061] = 0
      "0000000" when "00001011110101110", -- t[6062] = 0
      "0000000" when "00001011110101111", -- t[6063] = 0
      "0000000" when "00001011110110000", -- t[6064] = 0
      "0000000" when "00001011110110001", -- t[6065] = 0
      "0000000" when "00001011110110010", -- t[6066] = 0
      "0000000" when "00001011110110011", -- t[6067] = 0
      "0000000" when "00001011110110100", -- t[6068] = 0
      "0000000" when "00001011110110101", -- t[6069] = 0
      "0000000" when "00001011110110110", -- t[6070] = 0
      "0000000" when "00001011110110111", -- t[6071] = 0
      "0000000" when "00001011110111000", -- t[6072] = 0
      "0000000" when "00001011110111001", -- t[6073] = 0
      "0000000" when "00001011110111010", -- t[6074] = 0
      "0000000" when "00001011110111011", -- t[6075] = 0
      "0000000" when "00001011110111100", -- t[6076] = 0
      "0000000" when "00001011110111101", -- t[6077] = 0
      "0000000" when "00001011110111110", -- t[6078] = 0
      "0000000" when "00001011110111111", -- t[6079] = 0
      "0000000" when "00001011111000000", -- t[6080] = 0
      "0000000" when "00001011111000001", -- t[6081] = 0
      "0000000" when "00001011111000010", -- t[6082] = 0
      "0000000" when "00001011111000011", -- t[6083] = 0
      "0000000" when "00001011111000100", -- t[6084] = 0
      "0000000" when "00001011111000101", -- t[6085] = 0
      "0000000" when "00001011111000110", -- t[6086] = 0
      "0000000" when "00001011111000111", -- t[6087] = 0
      "0000000" when "00001011111001000", -- t[6088] = 0
      "0000000" when "00001011111001001", -- t[6089] = 0
      "0000000" when "00001011111001010", -- t[6090] = 0
      "0000000" when "00001011111001011", -- t[6091] = 0
      "0000000" when "00001011111001100", -- t[6092] = 0
      "0000000" when "00001011111001101", -- t[6093] = 0
      "0000000" when "00001011111001110", -- t[6094] = 0
      "0000000" when "00001011111001111", -- t[6095] = 0
      "0000000" when "00001011111010000", -- t[6096] = 0
      "0000000" when "00001011111010001", -- t[6097] = 0
      "0000000" when "00001011111010010", -- t[6098] = 0
      "0000000" when "00001011111010011", -- t[6099] = 0
      "0000000" when "00001011111010100", -- t[6100] = 0
      "0000000" when "00001011111010101", -- t[6101] = 0
      "0000000" when "00001011111010110", -- t[6102] = 0
      "0000000" when "00001011111010111", -- t[6103] = 0
      "0000000" when "00001011111011000", -- t[6104] = 0
      "0000000" when "00001011111011001", -- t[6105] = 0
      "0000000" when "00001011111011010", -- t[6106] = 0
      "0000000" when "00001011111011011", -- t[6107] = 0
      "0000000" when "00001011111011100", -- t[6108] = 0
      "0000000" when "00001011111011101", -- t[6109] = 0
      "0000000" when "00001011111011110", -- t[6110] = 0
      "0000000" when "00001011111011111", -- t[6111] = 0
      "0000000" when "00001011111100000", -- t[6112] = 0
      "0000000" when "00001011111100001", -- t[6113] = 0
      "0000000" when "00001011111100010", -- t[6114] = 0
      "0000000" when "00001011111100011", -- t[6115] = 0
      "0000000" when "00001011111100100", -- t[6116] = 0
      "0000000" when "00001011111100101", -- t[6117] = 0
      "0000000" when "00001011111100110", -- t[6118] = 0
      "0000000" when "00001011111100111", -- t[6119] = 0
      "0000000" when "00001011111101000", -- t[6120] = 0
      "0000000" when "00001011111101001", -- t[6121] = 0
      "0000000" when "00001011111101010", -- t[6122] = 0
      "0000000" when "00001011111101011", -- t[6123] = 0
      "0000000" when "00001011111101100", -- t[6124] = 0
      "0000000" when "00001011111101101", -- t[6125] = 0
      "0000000" when "00001011111101110", -- t[6126] = 0
      "0000000" when "00001011111101111", -- t[6127] = 0
      "0000000" when "00001011111110000", -- t[6128] = 0
      "0000000" when "00001011111110001", -- t[6129] = 0
      "0000000" when "00001011111110010", -- t[6130] = 0
      "0000000" when "00001011111110011", -- t[6131] = 0
      "0000000" when "00001011111110100", -- t[6132] = 0
      "0000000" when "00001011111110101", -- t[6133] = 0
      "0000000" when "00001011111110110", -- t[6134] = 0
      "0000000" when "00001011111110111", -- t[6135] = 0
      "0000000" when "00001011111111000", -- t[6136] = 0
      "0000000" when "00001011111111001", -- t[6137] = 0
      "0000000" when "00001011111111010", -- t[6138] = 0
      "0000000" when "00001011111111011", -- t[6139] = 0
      "0000000" when "00001011111111100", -- t[6140] = 0
      "0000000" when "00001011111111101", -- t[6141] = 0
      "0000000" when "00001011111111110", -- t[6142] = 0
      "0000000" when "00001011111111111", -- t[6143] = 0
      "0000000" when "00001100000000000", -- t[6144] = 0
      "0000000" when "00001100000000001", -- t[6145] = 0
      "0000000" when "00001100000000010", -- t[6146] = 0
      "0000000" when "00001100000000011", -- t[6147] = 0
      "0000000" when "00001100000000100", -- t[6148] = 0
      "0000000" when "00001100000000101", -- t[6149] = 0
      "0000000" when "00001100000000110", -- t[6150] = 0
      "0000000" when "00001100000000111", -- t[6151] = 0
      "0000000" when "00001100000001000", -- t[6152] = 0
      "0000000" when "00001100000001001", -- t[6153] = 0
      "0000000" when "00001100000001010", -- t[6154] = 0
      "0000000" when "00001100000001011", -- t[6155] = 0
      "0000000" when "00001100000001100", -- t[6156] = 0
      "0000000" when "00001100000001101", -- t[6157] = 0
      "0000000" when "00001100000001110", -- t[6158] = 0
      "0000000" when "00001100000001111", -- t[6159] = 0
      "0000000" when "00001100000010000", -- t[6160] = 0
      "0000000" when "00001100000010001", -- t[6161] = 0
      "0000000" when "00001100000010010", -- t[6162] = 0
      "0000000" when "00001100000010011", -- t[6163] = 0
      "0000000" when "00001100000010100", -- t[6164] = 0
      "0000000" when "00001100000010101", -- t[6165] = 0
      "0000000" when "00001100000010110", -- t[6166] = 0
      "0000000" when "00001100000010111", -- t[6167] = 0
      "0000000" when "00001100000011000", -- t[6168] = 0
      "0000000" when "00001100000011001", -- t[6169] = 0
      "0000000" when "00001100000011010", -- t[6170] = 0
      "0000000" when "00001100000011011", -- t[6171] = 0
      "0000000" when "00001100000011100", -- t[6172] = 0
      "0000000" when "00001100000011101", -- t[6173] = 0
      "0000000" when "00001100000011110", -- t[6174] = 0
      "0000000" when "00001100000011111", -- t[6175] = 0
      "0000000" when "00001100000100000", -- t[6176] = 0
      "0000000" when "00001100000100001", -- t[6177] = 0
      "0000000" when "00001100000100010", -- t[6178] = 0
      "0000000" when "00001100000100011", -- t[6179] = 0
      "0000000" when "00001100000100100", -- t[6180] = 0
      "0000000" when "00001100000100101", -- t[6181] = 0
      "0000000" when "00001100000100110", -- t[6182] = 0
      "0000000" when "00001100000100111", -- t[6183] = 0
      "0000000" when "00001100000101000", -- t[6184] = 0
      "0000000" when "00001100000101001", -- t[6185] = 0
      "0000000" when "00001100000101010", -- t[6186] = 0
      "0000000" when "00001100000101011", -- t[6187] = 0
      "0000000" when "00001100000101100", -- t[6188] = 0
      "0000000" when "00001100000101101", -- t[6189] = 0
      "0000000" when "00001100000101110", -- t[6190] = 0
      "0000000" when "00001100000101111", -- t[6191] = 0
      "0000000" when "00001100000110000", -- t[6192] = 0
      "0000000" when "00001100000110001", -- t[6193] = 0
      "0000000" when "00001100000110010", -- t[6194] = 0
      "0000000" when "00001100000110011", -- t[6195] = 0
      "0000000" when "00001100000110100", -- t[6196] = 0
      "0000000" when "00001100000110101", -- t[6197] = 0
      "0000000" when "00001100000110110", -- t[6198] = 0
      "0000000" when "00001100000110111", -- t[6199] = 0
      "0000000" when "00001100000111000", -- t[6200] = 0
      "0000000" when "00001100000111001", -- t[6201] = 0
      "0000000" when "00001100000111010", -- t[6202] = 0
      "0000000" when "00001100000111011", -- t[6203] = 0
      "0000000" when "00001100000111100", -- t[6204] = 0
      "0000000" when "00001100000111101", -- t[6205] = 0
      "0000000" when "00001100000111110", -- t[6206] = 0
      "0000000" when "00001100000111111", -- t[6207] = 0
      "0000000" when "00001100001000000", -- t[6208] = 0
      "0000000" when "00001100001000001", -- t[6209] = 0
      "0000000" when "00001100001000010", -- t[6210] = 0
      "0000000" when "00001100001000011", -- t[6211] = 0
      "0000000" when "00001100001000100", -- t[6212] = 0
      "0000000" when "00001100001000101", -- t[6213] = 0
      "0000000" when "00001100001000110", -- t[6214] = 0
      "0000000" when "00001100001000111", -- t[6215] = 0
      "0000000" when "00001100001001000", -- t[6216] = 0
      "0000000" when "00001100001001001", -- t[6217] = 0
      "0000000" when "00001100001001010", -- t[6218] = 0
      "0000000" when "00001100001001011", -- t[6219] = 0
      "0000000" when "00001100001001100", -- t[6220] = 0
      "0000000" when "00001100001001101", -- t[6221] = 0
      "0000000" when "00001100001001110", -- t[6222] = 0
      "0000000" when "00001100001001111", -- t[6223] = 0
      "0000000" when "00001100001010000", -- t[6224] = 0
      "0000000" when "00001100001010001", -- t[6225] = 0
      "0000000" when "00001100001010010", -- t[6226] = 0
      "0000000" when "00001100001010011", -- t[6227] = 0
      "0000000" when "00001100001010100", -- t[6228] = 0
      "0000000" when "00001100001010101", -- t[6229] = 0
      "0000000" when "00001100001010110", -- t[6230] = 0
      "0000000" when "00001100001010111", -- t[6231] = 0
      "0000000" when "00001100001011000", -- t[6232] = 0
      "0000000" when "00001100001011001", -- t[6233] = 0
      "0000000" when "00001100001011010", -- t[6234] = 0
      "0000000" when "00001100001011011", -- t[6235] = 0
      "0000000" when "00001100001011100", -- t[6236] = 0
      "0000000" when "00001100001011101", -- t[6237] = 0
      "0000000" when "00001100001011110", -- t[6238] = 0
      "0000000" when "00001100001011111", -- t[6239] = 0
      "0000000" when "00001100001100000", -- t[6240] = 0
      "0000000" when "00001100001100001", -- t[6241] = 0
      "0000000" when "00001100001100010", -- t[6242] = 0
      "0000000" when "00001100001100011", -- t[6243] = 0
      "0000000" when "00001100001100100", -- t[6244] = 0
      "0000000" when "00001100001100101", -- t[6245] = 0
      "0000000" when "00001100001100110", -- t[6246] = 0
      "0000000" when "00001100001100111", -- t[6247] = 0
      "0000000" when "00001100001101000", -- t[6248] = 0
      "0000000" when "00001100001101001", -- t[6249] = 0
      "0000000" when "00001100001101010", -- t[6250] = 0
      "0000000" when "00001100001101011", -- t[6251] = 0
      "0000000" when "00001100001101100", -- t[6252] = 0
      "0000000" when "00001100001101101", -- t[6253] = 0
      "0000000" when "00001100001101110", -- t[6254] = 0
      "0000000" when "00001100001101111", -- t[6255] = 0
      "0000000" when "00001100001110000", -- t[6256] = 0
      "0000000" when "00001100001110001", -- t[6257] = 0
      "0000000" when "00001100001110010", -- t[6258] = 0
      "0000000" when "00001100001110011", -- t[6259] = 0
      "0000000" when "00001100001110100", -- t[6260] = 0
      "0000000" when "00001100001110101", -- t[6261] = 0
      "0000000" when "00001100001110110", -- t[6262] = 0
      "0000000" when "00001100001110111", -- t[6263] = 0
      "0000000" when "00001100001111000", -- t[6264] = 0
      "0000000" when "00001100001111001", -- t[6265] = 0
      "0000000" when "00001100001111010", -- t[6266] = 0
      "0000000" when "00001100001111011", -- t[6267] = 0
      "0000000" when "00001100001111100", -- t[6268] = 0
      "0000000" when "00001100001111101", -- t[6269] = 0
      "0000000" when "00001100001111110", -- t[6270] = 0
      "0000000" when "00001100001111111", -- t[6271] = 0
      "0000000" when "00001100010000000", -- t[6272] = 0
      "0000000" when "00001100010000001", -- t[6273] = 0
      "0000000" when "00001100010000010", -- t[6274] = 0
      "0000000" when "00001100010000011", -- t[6275] = 0
      "0000000" when "00001100010000100", -- t[6276] = 0
      "0000000" when "00001100010000101", -- t[6277] = 0
      "0000000" when "00001100010000110", -- t[6278] = 0
      "0000000" when "00001100010000111", -- t[6279] = 0
      "0000000" when "00001100010001000", -- t[6280] = 0
      "0000000" when "00001100010001001", -- t[6281] = 0
      "0000000" when "00001100010001010", -- t[6282] = 0
      "0000000" when "00001100010001011", -- t[6283] = 0
      "0000000" when "00001100010001100", -- t[6284] = 0
      "0000000" when "00001100010001101", -- t[6285] = 0
      "0000000" when "00001100010001110", -- t[6286] = 0
      "0000000" when "00001100010001111", -- t[6287] = 0
      "0000000" when "00001100010010000", -- t[6288] = 0
      "0000000" when "00001100010010001", -- t[6289] = 0
      "0000000" when "00001100010010010", -- t[6290] = 0
      "0000000" when "00001100010010011", -- t[6291] = 0
      "0000000" when "00001100010010100", -- t[6292] = 0
      "0000000" when "00001100010010101", -- t[6293] = 0
      "0000000" when "00001100010010110", -- t[6294] = 0
      "0000000" when "00001100010010111", -- t[6295] = 0
      "0000000" when "00001100010011000", -- t[6296] = 0
      "0000000" when "00001100010011001", -- t[6297] = 0
      "0000000" when "00001100010011010", -- t[6298] = 0
      "0000000" when "00001100010011011", -- t[6299] = 0
      "0000000" when "00001100010011100", -- t[6300] = 0
      "0000000" when "00001100010011101", -- t[6301] = 0
      "0000000" when "00001100010011110", -- t[6302] = 0
      "0000000" when "00001100010011111", -- t[6303] = 0
      "0000000" when "00001100010100000", -- t[6304] = 0
      "0000000" when "00001100010100001", -- t[6305] = 0
      "0000000" when "00001100010100010", -- t[6306] = 0
      "0000000" when "00001100010100011", -- t[6307] = 0
      "0000000" when "00001100010100100", -- t[6308] = 0
      "0000000" when "00001100010100101", -- t[6309] = 0
      "0000000" when "00001100010100110", -- t[6310] = 0
      "0000000" when "00001100010100111", -- t[6311] = 0
      "0000000" when "00001100010101000", -- t[6312] = 0
      "0000000" when "00001100010101001", -- t[6313] = 0
      "0000000" when "00001100010101010", -- t[6314] = 0
      "0000000" when "00001100010101011", -- t[6315] = 0
      "0000000" when "00001100010101100", -- t[6316] = 0
      "0000000" when "00001100010101101", -- t[6317] = 0
      "0000000" when "00001100010101110", -- t[6318] = 0
      "0000000" when "00001100010101111", -- t[6319] = 0
      "0000000" when "00001100010110000", -- t[6320] = 0
      "0000000" when "00001100010110001", -- t[6321] = 0
      "0000000" when "00001100010110010", -- t[6322] = 0
      "0000000" when "00001100010110011", -- t[6323] = 0
      "0000000" when "00001100010110100", -- t[6324] = 0
      "0000000" when "00001100010110101", -- t[6325] = 0
      "0000000" when "00001100010110110", -- t[6326] = 0
      "0000000" when "00001100010110111", -- t[6327] = 0
      "0000000" when "00001100010111000", -- t[6328] = 0
      "0000000" when "00001100010111001", -- t[6329] = 0
      "0000000" when "00001100010111010", -- t[6330] = 0
      "0000000" when "00001100010111011", -- t[6331] = 0
      "0000000" when "00001100010111100", -- t[6332] = 0
      "0000000" when "00001100010111101", -- t[6333] = 0
      "0000000" when "00001100010111110", -- t[6334] = 0
      "0000000" when "00001100010111111", -- t[6335] = 0
      "0000000" when "00001100011000000", -- t[6336] = 0
      "0000000" when "00001100011000001", -- t[6337] = 0
      "0000000" when "00001100011000010", -- t[6338] = 0
      "0000000" when "00001100011000011", -- t[6339] = 0
      "0000000" when "00001100011000100", -- t[6340] = 0
      "0000000" when "00001100011000101", -- t[6341] = 0
      "0000000" when "00001100011000110", -- t[6342] = 0
      "0000000" when "00001100011000111", -- t[6343] = 0
      "0000000" when "00001100011001000", -- t[6344] = 0
      "0000000" when "00001100011001001", -- t[6345] = 0
      "0000000" when "00001100011001010", -- t[6346] = 0
      "0000000" when "00001100011001011", -- t[6347] = 0
      "0000000" when "00001100011001100", -- t[6348] = 0
      "0000000" when "00001100011001101", -- t[6349] = 0
      "0000000" when "00001100011001110", -- t[6350] = 0
      "0000000" when "00001100011001111", -- t[6351] = 0
      "0000000" when "00001100011010000", -- t[6352] = 0
      "0000000" when "00001100011010001", -- t[6353] = 0
      "0000000" when "00001100011010010", -- t[6354] = 0
      "0000000" when "00001100011010011", -- t[6355] = 0
      "0000000" when "00001100011010100", -- t[6356] = 0
      "0000000" when "00001100011010101", -- t[6357] = 0
      "0000000" when "00001100011010110", -- t[6358] = 0
      "0000000" when "00001100011010111", -- t[6359] = 0
      "0000000" when "00001100011011000", -- t[6360] = 0
      "0000000" when "00001100011011001", -- t[6361] = 0
      "0000000" when "00001100011011010", -- t[6362] = 0
      "0000000" when "00001100011011011", -- t[6363] = 0
      "0000000" when "00001100011011100", -- t[6364] = 0
      "0000000" when "00001100011011101", -- t[6365] = 0
      "0000000" when "00001100011011110", -- t[6366] = 0
      "0000000" when "00001100011011111", -- t[6367] = 0
      "0000000" when "00001100011100000", -- t[6368] = 0
      "0000000" when "00001100011100001", -- t[6369] = 0
      "0000000" when "00001100011100010", -- t[6370] = 0
      "0000000" when "00001100011100011", -- t[6371] = 0
      "0000000" when "00001100011100100", -- t[6372] = 0
      "0000000" when "00001100011100101", -- t[6373] = 0
      "0000000" when "00001100011100110", -- t[6374] = 0
      "0000000" when "00001100011100111", -- t[6375] = 0
      "0000000" when "00001100011101000", -- t[6376] = 0
      "0000000" when "00001100011101001", -- t[6377] = 0
      "0000000" when "00001100011101010", -- t[6378] = 0
      "0000000" when "00001100011101011", -- t[6379] = 0
      "0000000" when "00001100011101100", -- t[6380] = 0
      "0000000" when "00001100011101101", -- t[6381] = 0
      "0000000" when "00001100011101110", -- t[6382] = 0
      "0000000" when "00001100011101111", -- t[6383] = 0
      "0000000" when "00001100011110000", -- t[6384] = 0
      "0000000" when "00001100011110001", -- t[6385] = 0
      "0000000" when "00001100011110010", -- t[6386] = 0
      "0000000" when "00001100011110011", -- t[6387] = 0
      "0000000" when "00001100011110100", -- t[6388] = 0
      "0000000" when "00001100011110101", -- t[6389] = 0
      "0000000" when "00001100011110110", -- t[6390] = 0
      "0000000" when "00001100011110111", -- t[6391] = 0
      "0000000" when "00001100011111000", -- t[6392] = 0
      "0000000" when "00001100011111001", -- t[6393] = 0
      "0000000" when "00001100011111010", -- t[6394] = 0
      "0000000" when "00001100011111011", -- t[6395] = 0
      "0000000" when "00001100011111100", -- t[6396] = 0
      "0000000" when "00001100011111101", -- t[6397] = 0
      "0000000" when "00001100011111110", -- t[6398] = 0
      "0000000" when "00001100011111111", -- t[6399] = 0
      "0000000" when "00001100100000000", -- t[6400] = 0
      "0000000" when "00001100100000001", -- t[6401] = 0
      "0000000" when "00001100100000010", -- t[6402] = 0
      "0000000" when "00001100100000011", -- t[6403] = 0
      "0000000" when "00001100100000100", -- t[6404] = 0
      "0000000" when "00001100100000101", -- t[6405] = 0
      "0000000" when "00001100100000110", -- t[6406] = 0
      "0000000" when "00001100100000111", -- t[6407] = 0
      "0000000" when "00001100100001000", -- t[6408] = 0
      "0000000" when "00001100100001001", -- t[6409] = 0
      "0000000" when "00001100100001010", -- t[6410] = 0
      "0000000" when "00001100100001011", -- t[6411] = 0
      "0000000" when "00001100100001100", -- t[6412] = 0
      "0000000" when "00001100100001101", -- t[6413] = 0
      "0000000" when "00001100100001110", -- t[6414] = 0
      "0000000" when "00001100100001111", -- t[6415] = 0
      "0000000" when "00001100100010000", -- t[6416] = 0
      "0000000" when "00001100100010001", -- t[6417] = 0
      "0000000" when "00001100100010010", -- t[6418] = 0
      "0000000" when "00001100100010011", -- t[6419] = 0
      "0000000" when "00001100100010100", -- t[6420] = 0
      "0000000" when "00001100100010101", -- t[6421] = 0
      "0000000" when "00001100100010110", -- t[6422] = 0
      "0000000" when "00001100100010111", -- t[6423] = 0
      "0000000" when "00001100100011000", -- t[6424] = 0
      "0000000" when "00001100100011001", -- t[6425] = 0
      "0000000" when "00001100100011010", -- t[6426] = 0
      "0000000" when "00001100100011011", -- t[6427] = 0
      "0000000" when "00001100100011100", -- t[6428] = 0
      "0000000" when "00001100100011101", -- t[6429] = 0
      "0000000" when "00001100100011110", -- t[6430] = 0
      "0000000" when "00001100100011111", -- t[6431] = 0
      "0000000" when "00001100100100000", -- t[6432] = 0
      "0000000" when "00001100100100001", -- t[6433] = 0
      "0000000" when "00001100100100010", -- t[6434] = 0
      "0000000" when "00001100100100011", -- t[6435] = 0
      "0000000" when "00001100100100100", -- t[6436] = 0
      "0000000" when "00001100100100101", -- t[6437] = 0
      "0000000" when "00001100100100110", -- t[6438] = 0
      "0000000" when "00001100100100111", -- t[6439] = 0
      "0000000" when "00001100100101000", -- t[6440] = 0
      "0000000" when "00001100100101001", -- t[6441] = 0
      "0000000" when "00001100100101010", -- t[6442] = 0
      "0000000" when "00001100100101011", -- t[6443] = 0
      "0000000" when "00001100100101100", -- t[6444] = 0
      "0000000" when "00001100100101101", -- t[6445] = 0
      "0000000" when "00001100100101110", -- t[6446] = 0
      "0000000" when "00001100100101111", -- t[6447] = 0
      "0000000" when "00001100100110000", -- t[6448] = 0
      "0000000" when "00001100100110001", -- t[6449] = 0
      "0000000" when "00001100100110010", -- t[6450] = 0
      "0000000" when "00001100100110011", -- t[6451] = 0
      "0000000" when "00001100100110100", -- t[6452] = 0
      "0000000" when "00001100100110101", -- t[6453] = 0
      "0000000" when "00001100100110110", -- t[6454] = 0
      "0000000" when "00001100100110111", -- t[6455] = 0
      "0000000" when "00001100100111000", -- t[6456] = 0
      "0000000" when "00001100100111001", -- t[6457] = 0
      "0000000" when "00001100100111010", -- t[6458] = 0
      "0000000" when "00001100100111011", -- t[6459] = 0
      "0000000" when "00001100100111100", -- t[6460] = 0
      "0000000" when "00001100100111101", -- t[6461] = 0
      "0000000" when "00001100100111110", -- t[6462] = 0
      "0000000" when "00001100100111111", -- t[6463] = 0
      "0000000" when "00001100101000000", -- t[6464] = 0
      "0000000" when "00001100101000001", -- t[6465] = 0
      "0000000" when "00001100101000010", -- t[6466] = 0
      "0000000" when "00001100101000011", -- t[6467] = 0
      "0000000" when "00001100101000100", -- t[6468] = 0
      "0000000" when "00001100101000101", -- t[6469] = 0
      "0000000" when "00001100101000110", -- t[6470] = 0
      "0000000" when "00001100101000111", -- t[6471] = 0
      "0000000" when "00001100101001000", -- t[6472] = 0
      "0000000" when "00001100101001001", -- t[6473] = 0
      "0000000" when "00001100101001010", -- t[6474] = 0
      "0000000" when "00001100101001011", -- t[6475] = 0
      "0000000" when "00001100101001100", -- t[6476] = 0
      "0000000" when "00001100101001101", -- t[6477] = 0
      "0000000" when "00001100101001110", -- t[6478] = 0
      "0000000" when "00001100101001111", -- t[6479] = 0
      "0000000" when "00001100101010000", -- t[6480] = 0
      "0000000" when "00001100101010001", -- t[6481] = 0
      "0000000" when "00001100101010010", -- t[6482] = 0
      "0000000" when "00001100101010011", -- t[6483] = 0
      "0000000" when "00001100101010100", -- t[6484] = 0
      "0000000" when "00001100101010101", -- t[6485] = 0
      "0000000" when "00001100101010110", -- t[6486] = 0
      "0000000" when "00001100101010111", -- t[6487] = 0
      "0000000" when "00001100101011000", -- t[6488] = 0
      "0000000" when "00001100101011001", -- t[6489] = 0
      "0000000" when "00001100101011010", -- t[6490] = 0
      "0000000" when "00001100101011011", -- t[6491] = 0
      "0000000" when "00001100101011100", -- t[6492] = 0
      "0000000" when "00001100101011101", -- t[6493] = 0
      "0000000" when "00001100101011110", -- t[6494] = 0
      "0000000" when "00001100101011111", -- t[6495] = 0
      "0000000" when "00001100101100000", -- t[6496] = 0
      "0000000" when "00001100101100001", -- t[6497] = 0
      "0000000" when "00001100101100010", -- t[6498] = 0
      "0000000" when "00001100101100011", -- t[6499] = 0
      "0000000" when "00001100101100100", -- t[6500] = 0
      "0000000" when "00001100101100101", -- t[6501] = 0
      "0000000" when "00001100101100110", -- t[6502] = 0
      "0000000" when "00001100101100111", -- t[6503] = 0
      "0000000" when "00001100101101000", -- t[6504] = 0
      "0000000" when "00001100101101001", -- t[6505] = 0
      "0000000" when "00001100101101010", -- t[6506] = 0
      "0000000" when "00001100101101011", -- t[6507] = 0
      "0000000" when "00001100101101100", -- t[6508] = 0
      "0000000" when "00001100101101101", -- t[6509] = 0
      "0000000" when "00001100101101110", -- t[6510] = 0
      "0000000" when "00001100101101111", -- t[6511] = 0
      "0000000" when "00001100101110000", -- t[6512] = 0
      "0000000" when "00001100101110001", -- t[6513] = 0
      "0000000" when "00001100101110010", -- t[6514] = 0
      "0000000" when "00001100101110011", -- t[6515] = 0
      "0000000" when "00001100101110100", -- t[6516] = 0
      "0000000" when "00001100101110101", -- t[6517] = 0
      "0000000" when "00001100101110110", -- t[6518] = 0
      "0000000" when "00001100101110111", -- t[6519] = 0
      "0000000" when "00001100101111000", -- t[6520] = 0
      "0000000" when "00001100101111001", -- t[6521] = 0
      "0000000" when "00001100101111010", -- t[6522] = 0
      "0000000" when "00001100101111011", -- t[6523] = 0
      "0000000" when "00001100101111100", -- t[6524] = 0
      "0000000" when "00001100101111101", -- t[6525] = 0
      "0000000" when "00001100101111110", -- t[6526] = 0
      "0000000" when "00001100101111111", -- t[6527] = 0
      "0000000" when "00001100110000000", -- t[6528] = 0
      "0000000" when "00001100110000001", -- t[6529] = 0
      "0000000" when "00001100110000010", -- t[6530] = 0
      "0000000" when "00001100110000011", -- t[6531] = 0
      "0000000" when "00001100110000100", -- t[6532] = 0
      "0000000" when "00001100110000101", -- t[6533] = 0
      "0000000" when "00001100110000110", -- t[6534] = 0
      "0000000" when "00001100110000111", -- t[6535] = 0
      "0000000" when "00001100110001000", -- t[6536] = 0
      "0000000" when "00001100110001001", -- t[6537] = 0
      "0000000" when "00001100110001010", -- t[6538] = 0
      "0000000" when "00001100110001011", -- t[6539] = 0
      "0000000" when "00001100110001100", -- t[6540] = 0
      "0000000" when "00001100110001101", -- t[6541] = 0
      "0000000" when "00001100110001110", -- t[6542] = 0
      "0000000" when "00001100110001111", -- t[6543] = 0
      "0000000" when "00001100110010000", -- t[6544] = 0
      "0000000" when "00001100110010001", -- t[6545] = 0
      "0000000" when "00001100110010010", -- t[6546] = 0
      "0000000" when "00001100110010011", -- t[6547] = 0
      "0000000" when "00001100110010100", -- t[6548] = 0
      "0000000" when "00001100110010101", -- t[6549] = 0
      "0000000" when "00001100110010110", -- t[6550] = 0
      "0000000" when "00001100110010111", -- t[6551] = 0
      "0000000" when "00001100110011000", -- t[6552] = 0
      "0000000" when "00001100110011001", -- t[6553] = 0
      "0000000" when "00001100110011010", -- t[6554] = 0
      "0000000" when "00001100110011011", -- t[6555] = 0
      "0000000" when "00001100110011100", -- t[6556] = 0
      "0000000" when "00001100110011101", -- t[6557] = 0
      "0000000" when "00001100110011110", -- t[6558] = 0
      "0000000" when "00001100110011111", -- t[6559] = 0
      "0000000" when "00001100110100000", -- t[6560] = 0
      "0000000" when "00001100110100001", -- t[6561] = 0
      "0000000" when "00001100110100010", -- t[6562] = 0
      "0000000" when "00001100110100011", -- t[6563] = 0
      "0000000" when "00001100110100100", -- t[6564] = 0
      "0000000" when "00001100110100101", -- t[6565] = 0
      "0000000" when "00001100110100110", -- t[6566] = 0
      "0000000" when "00001100110100111", -- t[6567] = 0
      "0000000" when "00001100110101000", -- t[6568] = 0
      "0000000" when "00001100110101001", -- t[6569] = 0
      "0000000" when "00001100110101010", -- t[6570] = 0
      "0000000" when "00001100110101011", -- t[6571] = 0
      "0000000" when "00001100110101100", -- t[6572] = 0
      "0000000" when "00001100110101101", -- t[6573] = 0
      "0000000" when "00001100110101110", -- t[6574] = 0
      "0000000" when "00001100110101111", -- t[6575] = 0
      "0000000" when "00001100110110000", -- t[6576] = 0
      "0000000" when "00001100110110001", -- t[6577] = 0
      "0000000" when "00001100110110010", -- t[6578] = 0
      "0000000" when "00001100110110011", -- t[6579] = 0
      "0000000" when "00001100110110100", -- t[6580] = 0
      "0000000" when "00001100110110101", -- t[6581] = 0
      "0000000" when "00001100110110110", -- t[6582] = 0
      "0000000" when "00001100110110111", -- t[6583] = 0
      "0000000" when "00001100110111000", -- t[6584] = 0
      "0000000" when "00001100110111001", -- t[6585] = 0
      "0000000" when "00001100110111010", -- t[6586] = 0
      "0000000" when "00001100110111011", -- t[6587] = 0
      "0000000" when "00001100110111100", -- t[6588] = 0
      "0000000" when "00001100110111101", -- t[6589] = 0
      "0000000" when "00001100110111110", -- t[6590] = 0
      "0000000" when "00001100110111111", -- t[6591] = 0
      "0000000" when "00001100111000000", -- t[6592] = 0
      "0000000" when "00001100111000001", -- t[6593] = 0
      "0000000" when "00001100111000010", -- t[6594] = 0
      "0000000" when "00001100111000011", -- t[6595] = 0
      "0000000" when "00001100111000100", -- t[6596] = 0
      "0000000" when "00001100111000101", -- t[6597] = 0
      "0000000" when "00001100111000110", -- t[6598] = 0
      "0000000" when "00001100111000111", -- t[6599] = 0
      "0000000" when "00001100111001000", -- t[6600] = 0
      "0000000" when "00001100111001001", -- t[6601] = 0
      "0000000" when "00001100111001010", -- t[6602] = 0
      "0000000" when "00001100111001011", -- t[6603] = 0
      "0000000" when "00001100111001100", -- t[6604] = 0
      "0000000" when "00001100111001101", -- t[6605] = 0
      "0000000" when "00001100111001110", -- t[6606] = 0
      "0000000" when "00001100111001111", -- t[6607] = 0
      "0000000" when "00001100111010000", -- t[6608] = 0
      "0000000" when "00001100111010001", -- t[6609] = 0
      "0000000" when "00001100111010010", -- t[6610] = 0
      "0000000" when "00001100111010011", -- t[6611] = 0
      "0000000" when "00001100111010100", -- t[6612] = 0
      "0000000" when "00001100111010101", -- t[6613] = 0
      "0000000" when "00001100111010110", -- t[6614] = 0
      "0000000" when "00001100111010111", -- t[6615] = 0
      "0000000" when "00001100111011000", -- t[6616] = 0
      "0000000" when "00001100111011001", -- t[6617] = 0
      "0000000" when "00001100111011010", -- t[6618] = 0
      "0000000" when "00001100111011011", -- t[6619] = 0
      "0000000" when "00001100111011100", -- t[6620] = 0
      "0000000" when "00001100111011101", -- t[6621] = 0
      "0000000" when "00001100111011110", -- t[6622] = 0
      "0000000" when "00001100111011111", -- t[6623] = 0
      "0000000" when "00001100111100000", -- t[6624] = 0
      "0000000" when "00001100111100001", -- t[6625] = 0
      "0000000" when "00001100111100010", -- t[6626] = 0
      "0000000" when "00001100111100011", -- t[6627] = 0
      "0000000" when "00001100111100100", -- t[6628] = 0
      "0000000" when "00001100111100101", -- t[6629] = 0
      "0000000" when "00001100111100110", -- t[6630] = 0
      "0000000" when "00001100111100111", -- t[6631] = 0
      "0000000" when "00001100111101000", -- t[6632] = 0
      "0000000" when "00001100111101001", -- t[6633] = 0
      "0000000" when "00001100111101010", -- t[6634] = 0
      "0000000" when "00001100111101011", -- t[6635] = 0
      "0000000" when "00001100111101100", -- t[6636] = 0
      "0000000" when "00001100111101101", -- t[6637] = 0
      "0000000" when "00001100111101110", -- t[6638] = 0
      "0000000" when "00001100111101111", -- t[6639] = 0
      "0000000" when "00001100111110000", -- t[6640] = 0
      "0000000" when "00001100111110001", -- t[6641] = 0
      "0000000" when "00001100111110010", -- t[6642] = 0
      "0000000" when "00001100111110011", -- t[6643] = 0
      "0000000" when "00001100111110100", -- t[6644] = 0
      "0000000" when "00001100111110101", -- t[6645] = 0
      "0000000" when "00001100111110110", -- t[6646] = 0
      "0000000" when "00001100111110111", -- t[6647] = 0
      "0000000" when "00001100111111000", -- t[6648] = 0
      "0000000" when "00001100111111001", -- t[6649] = 0
      "0000000" when "00001100111111010", -- t[6650] = 0
      "0000000" when "00001100111111011", -- t[6651] = 0
      "0000000" when "00001100111111100", -- t[6652] = 0
      "0000000" when "00001100111111101", -- t[6653] = 0
      "0000000" when "00001100111111110", -- t[6654] = 0
      "0000000" when "00001100111111111", -- t[6655] = 0
      "0000000" when "00001101000000000", -- t[6656] = 0
      "0000000" when "00001101000000001", -- t[6657] = 0
      "0000000" when "00001101000000010", -- t[6658] = 0
      "0000000" when "00001101000000011", -- t[6659] = 0
      "0000000" when "00001101000000100", -- t[6660] = 0
      "0000000" when "00001101000000101", -- t[6661] = 0
      "0000000" when "00001101000000110", -- t[6662] = 0
      "0000000" when "00001101000000111", -- t[6663] = 0
      "0000000" when "00001101000001000", -- t[6664] = 0
      "0000000" when "00001101000001001", -- t[6665] = 0
      "0000000" when "00001101000001010", -- t[6666] = 0
      "0000000" when "00001101000001011", -- t[6667] = 0
      "0000000" when "00001101000001100", -- t[6668] = 0
      "0000000" when "00001101000001101", -- t[6669] = 0
      "0000000" when "00001101000001110", -- t[6670] = 0
      "0000000" when "00001101000001111", -- t[6671] = 0
      "0000000" when "00001101000010000", -- t[6672] = 0
      "0000000" when "00001101000010001", -- t[6673] = 0
      "0000000" when "00001101000010010", -- t[6674] = 0
      "0000000" when "00001101000010011", -- t[6675] = 0
      "0000000" when "00001101000010100", -- t[6676] = 0
      "0000000" when "00001101000010101", -- t[6677] = 0
      "0000000" when "00001101000010110", -- t[6678] = 0
      "0000000" when "00001101000010111", -- t[6679] = 0
      "0000000" when "00001101000011000", -- t[6680] = 0
      "0000000" when "00001101000011001", -- t[6681] = 0
      "0000000" when "00001101000011010", -- t[6682] = 0
      "0000000" when "00001101000011011", -- t[6683] = 0
      "0000000" when "00001101000011100", -- t[6684] = 0
      "0000000" when "00001101000011101", -- t[6685] = 0
      "0000000" when "00001101000011110", -- t[6686] = 0
      "0000000" when "00001101000011111", -- t[6687] = 0
      "0000000" when "00001101000100000", -- t[6688] = 0
      "0000000" when "00001101000100001", -- t[6689] = 0
      "0000000" when "00001101000100010", -- t[6690] = 0
      "0000000" when "00001101000100011", -- t[6691] = 0
      "0000000" when "00001101000100100", -- t[6692] = 0
      "0000000" when "00001101000100101", -- t[6693] = 0
      "0000000" when "00001101000100110", -- t[6694] = 0
      "0000000" when "00001101000100111", -- t[6695] = 0
      "0000000" when "00001101000101000", -- t[6696] = 0
      "0000000" when "00001101000101001", -- t[6697] = 0
      "0000000" when "00001101000101010", -- t[6698] = 0
      "0000000" when "00001101000101011", -- t[6699] = 0
      "0000000" when "00001101000101100", -- t[6700] = 0
      "0000000" when "00001101000101101", -- t[6701] = 0
      "0000000" when "00001101000101110", -- t[6702] = 0
      "0000000" when "00001101000101111", -- t[6703] = 0
      "0000000" when "00001101000110000", -- t[6704] = 0
      "0000000" when "00001101000110001", -- t[6705] = 0
      "0000000" when "00001101000110010", -- t[6706] = 0
      "0000000" when "00001101000110011", -- t[6707] = 0
      "0000000" when "00001101000110100", -- t[6708] = 0
      "0000000" when "00001101000110101", -- t[6709] = 0
      "0000000" when "00001101000110110", -- t[6710] = 0
      "0000000" when "00001101000110111", -- t[6711] = 0
      "0000000" when "00001101000111000", -- t[6712] = 0
      "0000000" when "00001101000111001", -- t[6713] = 0
      "0000000" when "00001101000111010", -- t[6714] = 0
      "0000000" when "00001101000111011", -- t[6715] = 0
      "0000000" when "00001101000111100", -- t[6716] = 0
      "0000000" when "00001101000111101", -- t[6717] = 0
      "0000000" when "00001101000111110", -- t[6718] = 0
      "0000000" when "00001101000111111", -- t[6719] = 0
      "0000000" when "00001101001000000", -- t[6720] = 0
      "0000000" when "00001101001000001", -- t[6721] = 0
      "0000000" when "00001101001000010", -- t[6722] = 0
      "0000000" when "00001101001000011", -- t[6723] = 0
      "0000000" when "00001101001000100", -- t[6724] = 0
      "0000000" when "00001101001000101", -- t[6725] = 0
      "0000000" when "00001101001000110", -- t[6726] = 0
      "0000000" when "00001101001000111", -- t[6727] = 0
      "0000000" when "00001101001001000", -- t[6728] = 0
      "0000000" when "00001101001001001", -- t[6729] = 0
      "0000000" when "00001101001001010", -- t[6730] = 0
      "0000000" when "00001101001001011", -- t[6731] = 0
      "0000000" when "00001101001001100", -- t[6732] = 0
      "0000000" when "00001101001001101", -- t[6733] = 0
      "0000000" when "00001101001001110", -- t[6734] = 0
      "0000000" when "00001101001001111", -- t[6735] = 0
      "0000000" when "00001101001010000", -- t[6736] = 0
      "0000000" when "00001101001010001", -- t[6737] = 0
      "0000000" when "00001101001010010", -- t[6738] = 0
      "0000000" when "00001101001010011", -- t[6739] = 0
      "0000000" when "00001101001010100", -- t[6740] = 0
      "0000000" when "00001101001010101", -- t[6741] = 0
      "0000000" when "00001101001010110", -- t[6742] = 0
      "0000000" when "00001101001010111", -- t[6743] = 0
      "0000000" when "00001101001011000", -- t[6744] = 0
      "0000000" when "00001101001011001", -- t[6745] = 0
      "0000000" when "00001101001011010", -- t[6746] = 0
      "0000000" when "00001101001011011", -- t[6747] = 0
      "0000000" when "00001101001011100", -- t[6748] = 0
      "0000000" when "00001101001011101", -- t[6749] = 0
      "0000000" when "00001101001011110", -- t[6750] = 0
      "0000000" when "00001101001011111", -- t[6751] = 0
      "0000000" when "00001101001100000", -- t[6752] = 0
      "0000000" when "00001101001100001", -- t[6753] = 0
      "0000000" when "00001101001100010", -- t[6754] = 0
      "0000000" when "00001101001100011", -- t[6755] = 0
      "0000000" when "00001101001100100", -- t[6756] = 0
      "0000000" when "00001101001100101", -- t[6757] = 0
      "0000000" when "00001101001100110", -- t[6758] = 0
      "0000000" when "00001101001100111", -- t[6759] = 0
      "0000000" when "00001101001101000", -- t[6760] = 0
      "0000000" when "00001101001101001", -- t[6761] = 0
      "0000000" when "00001101001101010", -- t[6762] = 0
      "0000000" when "00001101001101011", -- t[6763] = 0
      "0000000" when "00001101001101100", -- t[6764] = 0
      "0000000" when "00001101001101101", -- t[6765] = 0
      "0000000" when "00001101001101110", -- t[6766] = 0
      "0000000" when "00001101001101111", -- t[6767] = 0
      "0000000" when "00001101001110000", -- t[6768] = 0
      "0000000" when "00001101001110001", -- t[6769] = 0
      "0000000" when "00001101001110010", -- t[6770] = 0
      "0000000" when "00001101001110011", -- t[6771] = 0
      "0000000" when "00001101001110100", -- t[6772] = 0
      "0000000" when "00001101001110101", -- t[6773] = 0
      "0000000" when "00001101001110110", -- t[6774] = 0
      "0000000" when "00001101001110111", -- t[6775] = 0
      "0000000" when "00001101001111000", -- t[6776] = 0
      "0000000" when "00001101001111001", -- t[6777] = 0
      "0000000" when "00001101001111010", -- t[6778] = 0
      "0000000" when "00001101001111011", -- t[6779] = 0
      "0000000" when "00001101001111100", -- t[6780] = 0
      "0000000" when "00001101001111101", -- t[6781] = 0
      "0000000" when "00001101001111110", -- t[6782] = 0
      "0000000" when "00001101001111111", -- t[6783] = 0
      "0000000" when "00001101010000000", -- t[6784] = 0
      "0000000" when "00001101010000001", -- t[6785] = 0
      "0000000" when "00001101010000010", -- t[6786] = 0
      "0000000" when "00001101010000011", -- t[6787] = 0
      "0000000" when "00001101010000100", -- t[6788] = 0
      "0000000" when "00001101010000101", -- t[6789] = 0
      "0000000" when "00001101010000110", -- t[6790] = 0
      "0000000" when "00001101010000111", -- t[6791] = 0
      "0000000" when "00001101010001000", -- t[6792] = 0
      "0000000" when "00001101010001001", -- t[6793] = 0
      "0000000" when "00001101010001010", -- t[6794] = 0
      "0000000" when "00001101010001011", -- t[6795] = 0
      "0000000" when "00001101010001100", -- t[6796] = 0
      "0000000" when "00001101010001101", -- t[6797] = 0
      "0000000" when "00001101010001110", -- t[6798] = 0
      "0000000" when "00001101010001111", -- t[6799] = 0
      "0000000" when "00001101010010000", -- t[6800] = 0
      "0000000" when "00001101010010001", -- t[6801] = 0
      "0000000" when "00001101010010010", -- t[6802] = 0
      "0000000" when "00001101010010011", -- t[6803] = 0
      "0000000" when "00001101010010100", -- t[6804] = 0
      "0000000" when "00001101010010101", -- t[6805] = 0
      "0000000" when "00001101010010110", -- t[6806] = 0
      "0000000" when "00001101010010111", -- t[6807] = 0
      "0000000" when "00001101010011000", -- t[6808] = 0
      "0000000" when "00001101010011001", -- t[6809] = 0
      "0000000" when "00001101010011010", -- t[6810] = 0
      "0000000" when "00001101010011011", -- t[6811] = 0
      "0000000" when "00001101010011100", -- t[6812] = 0
      "0000000" when "00001101010011101", -- t[6813] = 0
      "0000000" when "00001101010011110", -- t[6814] = 0
      "0000000" when "00001101010011111", -- t[6815] = 0
      "0000000" when "00001101010100000", -- t[6816] = 0
      "0000000" when "00001101010100001", -- t[6817] = 0
      "0000000" when "00001101010100010", -- t[6818] = 0
      "0000000" when "00001101010100011", -- t[6819] = 0
      "0000000" when "00001101010100100", -- t[6820] = 0
      "0000000" when "00001101010100101", -- t[6821] = 0
      "0000000" when "00001101010100110", -- t[6822] = 0
      "0000000" when "00001101010100111", -- t[6823] = 0
      "0000000" when "00001101010101000", -- t[6824] = 0
      "0000000" when "00001101010101001", -- t[6825] = 0
      "0000000" when "00001101010101010", -- t[6826] = 0
      "0000000" when "00001101010101011", -- t[6827] = 0
      "0000000" when "00001101010101100", -- t[6828] = 0
      "0000000" when "00001101010101101", -- t[6829] = 0
      "0000000" when "00001101010101110", -- t[6830] = 0
      "0000000" when "00001101010101111", -- t[6831] = 0
      "0000000" when "00001101010110000", -- t[6832] = 0
      "0000000" when "00001101010110001", -- t[6833] = 0
      "0000000" when "00001101010110010", -- t[6834] = 0
      "0000000" when "00001101010110011", -- t[6835] = 0
      "0000000" when "00001101010110100", -- t[6836] = 0
      "0000000" when "00001101010110101", -- t[6837] = 0
      "0000000" when "00001101010110110", -- t[6838] = 0
      "0000000" when "00001101010110111", -- t[6839] = 0
      "0000000" when "00001101010111000", -- t[6840] = 0
      "0000000" when "00001101010111001", -- t[6841] = 0
      "0000000" when "00001101010111010", -- t[6842] = 0
      "0000000" when "00001101010111011", -- t[6843] = 0
      "0000000" when "00001101010111100", -- t[6844] = 0
      "0000000" when "00001101010111101", -- t[6845] = 0
      "0000000" when "00001101010111110", -- t[6846] = 0
      "0000000" when "00001101010111111", -- t[6847] = 0
      "0000000" when "00001101011000000", -- t[6848] = 0
      "0000000" when "00001101011000001", -- t[6849] = 0
      "0000000" when "00001101011000010", -- t[6850] = 0
      "0000000" when "00001101011000011", -- t[6851] = 0
      "0000000" when "00001101011000100", -- t[6852] = 0
      "0000000" when "00001101011000101", -- t[6853] = 0
      "0000000" when "00001101011000110", -- t[6854] = 0
      "0000000" when "00001101011000111", -- t[6855] = 0
      "0000000" when "00001101011001000", -- t[6856] = 0
      "0000000" when "00001101011001001", -- t[6857] = 0
      "0000000" when "00001101011001010", -- t[6858] = 0
      "0000000" when "00001101011001011", -- t[6859] = 0
      "0000000" when "00001101011001100", -- t[6860] = 0
      "0000000" when "00001101011001101", -- t[6861] = 0
      "0000000" when "00001101011001110", -- t[6862] = 0
      "0000000" when "00001101011001111", -- t[6863] = 0
      "0000000" when "00001101011010000", -- t[6864] = 0
      "0000000" when "00001101011010001", -- t[6865] = 0
      "0000000" when "00001101011010010", -- t[6866] = 0
      "0000000" when "00001101011010011", -- t[6867] = 0
      "0000000" when "00001101011010100", -- t[6868] = 0
      "0000000" when "00001101011010101", -- t[6869] = 0
      "0000000" when "00001101011010110", -- t[6870] = 0
      "0000000" when "00001101011010111", -- t[6871] = 0
      "0000000" when "00001101011011000", -- t[6872] = 0
      "0000000" when "00001101011011001", -- t[6873] = 0
      "0000000" when "00001101011011010", -- t[6874] = 0
      "0000000" when "00001101011011011", -- t[6875] = 0
      "0000000" when "00001101011011100", -- t[6876] = 0
      "0000000" when "00001101011011101", -- t[6877] = 0
      "0000000" when "00001101011011110", -- t[6878] = 0
      "0000000" when "00001101011011111", -- t[6879] = 0
      "0000000" when "00001101011100000", -- t[6880] = 0
      "0000000" when "00001101011100001", -- t[6881] = 0
      "0000000" when "00001101011100010", -- t[6882] = 0
      "0000000" when "00001101011100011", -- t[6883] = 0
      "0000000" when "00001101011100100", -- t[6884] = 0
      "0000000" when "00001101011100101", -- t[6885] = 0
      "0000000" when "00001101011100110", -- t[6886] = 0
      "0000000" when "00001101011100111", -- t[6887] = 0
      "0000000" when "00001101011101000", -- t[6888] = 0
      "0000000" when "00001101011101001", -- t[6889] = 0
      "0000000" when "00001101011101010", -- t[6890] = 0
      "0000000" when "00001101011101011", -- t[6891] = 0
      "0000000" when "00001101011101100", -- t[6892] = 0
      "0000000" when "00001101011101101", -- t[6893] = 0
      "0000000" when "00001101011101110", -- t[6894] = 0
      "0000000" when "00001101011101111", -- t[6895] = 0
      "0000000" when "00001101011110000", -- t[6896] = 0
      "0000000" when "00001101011110001", -- t[6897] = 0
      "0000000" when "00001101011110010", -- t[6898] = 0
      "0000000" when "00001101011110011", -- t[6899] = 0
      "0000000" when "00001101011110100", -- t[6900] = 0
      "0000000" when "00001101011110101", -- t[6901] = 0
      "0000000" when "00001101011110110", -- t[6902] = 0
      "0000000" when "00001101011110111", -- t[6903] = 0
      "0000000" when "00001101011111000", -- t[6904] = 0
      "0000000" when "00001101011111001", -- t[6905] = 0
      "0000000" when "00001101011111010", -- t[6906] = 0
      "0000000" when "00001101011111011", -- t[6907] = 0
      "0000000" when "00001101011111100", -- t[6908] = 0
      "0000000" when "00001101011111101", -- t[6909] = 0
      "0000000" when "00001101011111110", -- t[6910] = 0
      "0000000" when "00001101011111111", -- t[6911] = 0
      "0000000" when "00001101100000000", -- t[6912] = 0
      "0000000" when "00001101100000001", -- t[6913] = 0
      "0000000" when "00001101100000010", -- t[6914] = 0
      "0000000" when "00001101100000011", -- t[6915] = 0
      "0000000" when "00001101100000100", -- t[6916] = 0
      "0000000" when "00001101100000101", -- t[6917] = 0
      "0000000" when "00001101100000110", -- t[6918] = 0
      "0000000" when "00001101100000111", -- t[6919] = 0
      "0000000" when "00001101100001000", -- t[6920] = 0
      "0000000" when "00001101100001001", -- t[6921] = 0
      "0000000" when "00001101100001010", -- t[6922] = 0
      "0000000" when "00001101100001011", -- t[6923] = 0
      "0000000" when "00001101100001100", -- t[6924] = 0
      "0000000" when "00001101100001101", -- t[6925] = 0
      "0000000" when "00001101100001110", -- t[6926] = 0
      "0000000" when "00001101100001111", -- t[6927] = 0
      "0000000" when "00001101100010000", -- t[6928] = 0
      "0000000" when "00001101100010001", -- t[6929] = 0
      "0000000" when "00001101100010010", -- t[6930] = 0
      "0000000" when "00001101100010011", -- t[6931] = 0
      "0000000" when "00001101100010100", -- t[6932] = 0
      "0000000" when "00001101100010101", -- t[6933] = 0
      "0000000" when "00001101100010110", -- t[6934] = 0
      "0000000" when "00001101100010111", -- t[6935] = 0
      "0000000" when "00001101100011000", -- t[6936] = 0
      "0000000" when "00001101100011001", -- t[6937] = 0
      "0000000" when "00001101100011010", -- t[6938] = 0
      "0000000" when "00001101100011011", -- t[6939] = 0
      "0000000" when "00001101100011100", -- t[6940] = 0
      "0000000" when "00001101100011101", -- t[6941] = 0
      "0000000" when "00001101100011110", -- t[6942] = 0
      "0000000" when "00001101100011111", -- t[6943] = 0
      "0000000" when "00001101100100000", -- t[6944] = 0
      "0000000" when "00001101100100001", -- t[6945] = 0
      "0000000" when "00001101100100010", -- t[6946] = 0
      "0000000" when "00001101100100011", -- t[6947] = 0
      "0000000" when "00001101100100100", -- t[6948] = 0
      "0000000" when "00001101100100101", -- t[6949] = 0
      "0000000" when "00001101100100110", -- t[6950] = 0
      "0000000" when "00001101100100111", -- t[6951] = 0
      "0000000" when "00001101100101000", -- t[6952] = 0
      "0000000" when "00001101100101001", -- t[6953] = 0
      "0000000" when "00001101100101010", -- t[6954] = 0
      "0000000" when "00001101100101011", -- t[6955] = 0
      "0000000" when "00001101100101100", -- t[6956] = 0
      "0000000" when "00001101100101101", -- t[6957] = 0
      "0000000" when "00001101100101110", -- t[6958] = 0
      "0000000" when "00001101100101111", -- t[6959] = 0
      "0000000" when "00001101100110000", -- t[6960] = 0
      "0000000" when "00001101100110001", -- t[6961] = 0
      "0000000" when "00001101100110010", -- t[6962] = 0
      "0000000" when "00001101100110011", -- t[6963] = 0
      "0000000" when "00001101100110100", -- t[6964] = 0
      "0000000" when "00001101100110101", -- t[6965] = 0
      "0000000" when "00001101100110110", -- t[6966] = 0
      "0000000" when "00001101100110111", -- t[6967] = 0
      "0000000" when "00001101100111000", -- t[6968] = 0
      "0000000" when "00001101100111001", -- t[6969] = 0
      "0000000" when "00001101100111010", -- t[6970] = 0
      "0000000" when "00001101100111011", -- t[6971] = 0
      "0000000" when "00001101100111100", -- t[6972] = 0
      "0000000" when "00001101100111101", -- t[6973] = 0
      "0000000" when "00001101100111110", -- t[6974] = 0
      "0000000" when "00001101100111111", -- t[6975] = 0
      "0000000" when "00001101101000000", -- t[6976] = 0
      "0000000" when "00001101101000001", -- t[6977] = 0
      "0000000" when "00001101101000010", -- t[6978] = 0
      "0000000" when "00001101101000011", -- t[6979] = 0
      "0000000" when "00001101101000100", -- t[6980] = 0
      "0000000" when "00001101101000101", -- t[6981] = 0
      "0000000" when "00001101101000110", -- t[6982] = 0
      "0000000" when "00001101101000111", -- t[6983] = 0
      "0000000" when "00001101101001000", -- t[6984] = 0
      "0000000" when "00001101101001001", -- t[6985] = 0
      "0000000" when "00001101101001010", -- t[6986] = 0
      "0000000" when "00001101101001011", -- t[6987] = 0
      "0000000" when "00001101101001100", -- t[6988] = 0
      "0000000" when "00001101101001101", -- t[6989] = 0
      "0000000" when "00001101101001110", -- t[6990] = 0
      "0000000" when "00001101101001111", -- t[6991] = 0
      "0000000" when "00001101101010000", -- t[6992] = 0
      "0000000" when "00001101101010001", -- t[6993] = 0
      "0000000" when "00001101101010010", -- t[6994] = 0
      "0000000" when "00001101101010011", -- t[6995] = 0
      "0000000" when "00001101101010100", -- t[6996] = 0
      "0000000" when "00001101101010101", -- t[6997] = 0
      "0000000" when "00001101101010110", -- t[6998] = 0
      "0000000" when "00001101101010111", -- t[6999] = 0
      "0000000" when "00001101101011000", -- t[7000] = 0
      "0000000" when "00001101101011001", -- t[7001] = 0
      "0000000" when "00001101101011010", -- t[7002] = 0
      "0000000" when "00001101101011011", -- t[7003] = 0
      "0000000" when "00001101101011100", -- t[7004] = 0
      "0000000" when "00001101101011101", -- t[7005] = 0
      "0000000" when "00001101101011110", -- t[7006] = 0
      "0000000" when "00001101101011111", -- t[7007] = 0
      "0000000" when "00001101101100000", -- t[7008] = 0
      "0000000" when "00001101101100001", -- t[7009] = 0
      "0000000" when "00001101101100010", -- t[7010] = 0
      "0000000" when "00001101101100011", -- t[7011] = 0
      "0000000" when "00001101101100100", -- t[7012] = 0
      "0000000" when "00001101101100101", -- t[7013] = 0
      "0000000" when "00001101101100110", -- t[7014] = 0
      "0000000" when "00001101101100111", -- t[7015] = 0
      "0000000" when "00001101101101000", -- t[7016] = 0
      "0000000" when "00001101101101001", -- t[7017] = 0
      "0000000" when "00001101101101010", -- t[7018] = 0
      "0000000" when "00001101101101011", -- t[7019] = 0
      "0000000" when "00001101101101100", -- t[7020] = 0
      "0000000" when "00001101101101101", -- t[7021] = 0
      "0000000" when "00001101101101110", -- t[7022] = 0
      "0000000" when "00001101101101111", -- t[7023] = 0
      "0000000" when "00001101101110000", -- t[7024] = 0
      "0000000" when "00001101101110001", -- t[7025] = 0
      "0000000" when "00001101101110010", -- t[7026] = 0
      "0000000" when "00001101101110011", -- t[7027] = 0
      "0000000" when "00001101101110100", -- t[7028] = 0
      "0000000" when "00001101101110101", -- t[7029] = 0
      "0000000" when "00001101101110110", -- t[7030] = 0
      "0000000" when "00001101101110111", -- t[7031] = 0
      "0000000" when "00001101101111000", -- t[7032] = 0
      "0000000" when "00001101101111001", -- t[7033] = 0
      "0000000" when "00001101101111010", -- t[7034] = 0
      "0000000" when "00001101101111011", -- t[7035] = 0
      "0000000" when "00001101101111100", -- t[7036] = 0
      "0000000" when "00001101101111101", -- t[7037] = 0
      "0000000" when "00001101101111110", -- t[7038] = 0
      "0000000" when "00001101101111111", -- t[7039] = 0
      "0000000" when "00001101110000000", -- t[7040] = 0
      "0000000" when "00001101110000001", -- t[7041] = 0
      "0000000" when "00001101110000010", -- t[7042] = 0
      "0000000" when "00001101110000011", -- t[7043] = 0
      "0000000" when "00001101110000100", -- t[7044] = 0
      "0000000" when "00001101110000101", -- t[7045] = 0
      "0000000" when "00001101110000110", -- t[7046] = 0
      "0000000" when "00001101110000111", -- t[7047] = 0
      "0000000" when "00001101110001000", -- t[7048] = 0
      "0000000" when "00001101110001001", -- t[7049] = 0
      "0000000" when "00001101110001010", -- t[7050] = 0
      "0000000" when "00001101110001011", -- t[7051] = 0
      "0000000" when "00001101110001100", -- t[7052] = 0
      "0000000" when "00001101110001101", -- t[7053] = 0
      "0000000" when "00001101110001110", -- t[7054] = 0
      "0000000" when "00001101110001111", -- t[7055] = 0
      "0000000" when "00001101110010000", -- t[7056] = 0
      "0000000" when "00001101110010001", -- t[7057] = 0
      "0000000" when "00001101110010010", -- t[7058] = 0
      "0000000" when "00001101110010011", -- t[7059] = 0
      "0000000" when "00001101110010100", -- t[7060] = 0
      "0000000" when "00001101110010101", -- t[7061] = 0
      "0000000" when "00001101110010110", -- t[7062] = 0
      "0000000" when "00001101110010111", -- t[7063] = 0
      "0000000" when "00001101110011000", -- t[7064] = 0
      "0000000" when "00001101110011001", -- t[7065] = 0
      "0000000" when "00001101110011010", -- t[7066] = 0
      "0000000" when "00001101110011011", -- t[7067] = 0
      "0000000" when "00001101110011100", -- t[7068] = 0
      "0000000" when "00001101110011101", -- t[7069] = 0
      "0000000" when "00001101110011110", -- t[7070] = 0
      "0000000" when "00001101110011111", -- t[7071] = 0
      "0000000" when "00001101110100000", -- t[7072] = 0
      "0000000" when "00001101110100001", -- t[7073] = 0
      "0000000" when "00001101110100010", -- t[7074] = 0
      "0000000" when "00001101110100011", -- t[7075] = 0
      "0000000" when "00001101110100100", -- t[7076] = 0
      "0000000" when "00001101110100101", -- t[7077] = 0
      "0000000" when "00001101110100110", -- t[7078] = 0
      "0000000" when "00001101110100111", -- t[7079] = 0
      "0000000" when "00001101110101000", -- t[7080] = 0
      "0000000" when "00001101110101001", -- t[7081] = 0
      "0000000" when "00001101110101010", -- t[7082] = 0
      "0000000" when "00001101110101011", -- t[7083] = 0
      "0000000" when "00001101110101100", -- t[7084] = 0
      "0000000" when "00001101110101101", -- t[7085] = 0
      "0000000" when "00001101110101110", -- t[7086] = 0
      "0000000" when "00001101110101111", -- t[7087] = 0
      "0000000" when "00001101110110000", -- t[7088] = 0
      "0000000" when "00001101110110001", -- t[7089] = 0
      "0000000" when "00001101110110010", -- t[7090] = 0
      "0000000" when "00001101110110011", -- t[7091] = 0
      "0000000" when "00001101110110100", -- t[7092] = 0
      "0000000" when "00001101110110101", -- t[7093] = 0
      "0000000" when "00001101110110110", -- t[7094] = 0
      "0000000" when "00001101110110111", -- t[7095] = 0
      "0000000" when "00001101110111000", -- t[7096] = 0
      "0000000" when "00001101110111001", -- t[7097] = 0
      "0000000" when "00001101110111010", -- t[7098] = 0
      "0000000" when "00001101110111011", -- t[7099] = 0
      "0000000" when "00001101110111100", -- t[7100] = 0
      "0000000" when "00001101110111101", -- t[7101] = 0
      "0000000" when "00001101110111110", -- t[7102] = 0
      "0000000" when "00001101110111111", -- t[7103] = 0
      "0000000" when "00001101111000000", -- t[7104] = 0
      "0000000" when "00001101111000001", -- t[7105] = 0
      "0000000" when "00001101111000010", -- t[7106] = 0
      "0000000" when "00001101111000011", -- t[7107] = 0
      "0000000" when "00001101111000100", -- t[7108] = 0
      "0000000" when "00001101111000101", -- t[7109] = 0
      "0000000" when "00001101111000110", -- t[7110] = 0
      "0000000" when "00001101111000111", -- t[7111] = 0
      "0000000" when "00001101111001000", -- t[7112] = 0
      "0000000" when "00001101111001001", -- t[7113] = 0
      "0000000" when "00001101111001010", -- t[7114] = 0
      "0000000" when "00001101111001011", -- t[7115] = 0
      "0000000" when "00001101111001100", -- t[7116] = 0
      "0000000" when "00001101111001101", -- t[7117] = 0
      "0000000" when "00001101111001110", -- t[7118] = 0
      "0000000" when "00001101111001111", -- t[7119] = 0
      "0000000" when "00001101111010000", -- t[7120] = 0
      "0000000" when "00001101111010001", -- t[7121] = 0
      "0000000" when "00001101111010010", -- t[7122] = 0
      "0000000" when "00001101111010011", -- t[7123] = 0
      "0000000" when "00001101111010100", -- t[7124] = 0
      "0000000" when "00001101111010101", -- t[7125] = 0
      "0000000" when "00001101111010110", -- t[7126] = 0
      "0000000" when "00001101111010111", -- t[7127] = 0
      "0000000" when "00001101111011000", -- t[7128] = 0
      "0000000" when "00001101111011001", -- t[7129] = 0
      "0000000" when "00001101111011010", -- t[7130] = 0
      "0000000" when "00001101111011011", -- t[7131] = 0
      "0000000" when "00001101111011100", -- t[7132] = 0
      "0000000" when "00001101111011101", -- t[7133] = 0
      "0000000" when "00001101111011110", -- t[7134] = 0
      "0000000" when "00001101111011111", -- t[7135] = 0
      "0000000" when "00001101111100000", -- t[7136] = 0
      "0000000" when "00001101111100001", -- t[7137] = 0
      "0000000" when "00001101111100010", -- t[7138] = 0
      "0000000" when "00001101111100011", -- t[7139] = 0
      "0000000" when "00001101111100100", -- t[7140] = 0
      "0000000" when "00001101111100101", -- t[7141] = 0
      "0000000" when "00001101111100110", -- t[7142] = 0
      "0000000" when "00001101111100111", -- t[7143] = 0
      "0000000" when "00001101111101000", -- t[7144] = 0
      "0000000" when "00001101111101001", -- t[7145] = 0
      "0000000" when "00001101111101010", -- t[7146] = 0
      "0000000" when "00001101111101011", -- t[7147] = 0
      "0000000" when "00001101111101100", -- t[7148] = 0
      "0000000" when "00001101111101101", -- t[7149] = 0
      "0000000" when "00001101111101110", -- t[7150] = 0
      "0000000" when "00001101111101111", -- t[7151] = 0
      "0000000" when "00001101111110000", -- t[7152] = 0
      "0000000" when "00001101111110001", -- t[7153] = 0
      "0000000" when "00001101111110010", -- t[7154] = 0
      "0000000" when "00001101111110011", -- t[7155] = 0
      "0000000" when "00001101111110100", -- t[7156] = 0
      "0000000" when "00001101111110101", -- t[7157] = 0
      "0000000" when "00001101111110110", -- t[7158] = 0
      "0000000" when "00001101111110111", -- t[7159] = 0
      "0000000" when "00001101111111000", -- t[7160] = 0
      "0000000" when "00001101111111001", -- t[7161] = 0
      "0000000" when "00001101111111010", -- t[7162] = 0
      "0000000" when "00001101111111011", -- t[7163] = 0
      "0000000" when "00001101111111100", -- t[7164] = 0
      "0000000" when "00001101111111101", -- t[7165] = 0
      "0000000" when "00001101111111110", -- t[7166] = 0
      "0000000" when "00001101111111111", -- t[7167] = 0
      "0000000" when "00001110000000000", -- t[7168] = 0
      "0000000" when "00001110000000001", -- t[7169] = 0
      "0000000" when "00001110000000010", -- t[7170] = 0
      "0000000" when "00001110000000011", -- t[7171] = 0
      "0000000" when "00001110000000100", -- t[7172] = 0
      "0000000" when "00001110000000101", -- t[7173] = 0
      "0000000" when "00001110000000110", -- t[7174] = 0
      "0000000" when "00001110000000111", -- t[7175] = 0
      "0000000" when "00001110000001000", -- t[7176] = 0
      "0000000" when "00001110000001001", -- t[7177] = 0
      "0000000" when "00001110000001010", -- t[7178] = 0
      "0000000" when "00001110000001011", -- t[7179] = 0
      "0000000" when "00001110000001100", -- t[7180] = 0
      "0000000" when "00001110000001101", -- t[7181] = 0
      "0000000" when "00001110000001110", -- t[7182] = 0
      "0000000" when "00001110000001111", -- t[7183] = 0
      "0000000" when "00001110000010000", -- t[7184] = 0
      "0000000" when "00001110000010001", -- t[7185] = 0
      "0000000" when "00001110000010010", -- t[7186] = 0
      "0000000" when "00001110000010011", -- t[7187] = 0
      "0000000" when "00001110000010100", -- t[7188] = 0
      "0000000" when "00001110000010101", -- t[7189] = 0
      "0000000" when "00001110000010110", -- t[7190] = 0
      "0000000" when "00001110000010111", -- t[7191] = 0
      "0000000" when "00001110000011000", -- t[7192] = 0
      "0000000" when "00001110000011001", -- t[7193] = 0
      "0000000" when "00001110000011010", -- t[7194] = 0
      "0000000" when "00001110000011011", -- t[7195] = 0
      "0000000" when "00001110000011100", -- t[7196] = 0
      "0000000" when "00001110000011101", -- t[7197] = 0
      "0000000" when "00001110000011110", -- t[7198] = 0
      "0000000" when "00001110000011111", -- t[7199] = 0
      "0000000" when "00001110000100000", -- t[7200] = 0
      "0000000" when "00001110000100001", -- t[7201] = 0
      "0000000" when "00001110000100010", -- t[7202] = 0
      "0000000" when "00001110000100011", -- t[7203] = 0
      "0000000" when "00001110000100100", -- t[7204] = 0
      "0000000" when "00001110000100101", -- t[7205] = 0
      "0000000" when "00001110000100110", -- t[7206] = 0
      "0000000" when "00001110000100111", -- t[7207] = 0
      "0000000" when "00001110000101000", -- t[7208] = 0
      "0000000" when "00001110000101001", -- t[7209] = 0
      "0000000" when "00001110000101010", -- t[7210] = 0
      "0000000" when "00001110000101011", -- t[7211] = 0
      "0000000" when "00001110000101100", -- t[7212] = 0
      "0000000" when "00001110000101101", -- t[7213] = 0
      "0000000" when "00001110000101110", -- t[7214] = 0
      "0000000" when "00001110000101111", -- t[7215] = 0
      "0000000" when "00001110000110000", -- t[7216] = 0
      "0000000" when "00001110000110001", -- t[7217] = 0
      "0000000" when "00001110000110010", -- t[7218] = 0
      "0000000" when "00001110000110011", -- t[7219] = 0
      "0000000" when "00001110000110100", -- t[7220] = 0
      "0000000" when "00001110000110101", -- t[7221] = 0
      "0000000" when "00001110000110110", -- t[7222] = 0
      "0000000" when "00001110000110111", -- t[7223] = 0
      "0000000" when "00001110000111000", -- t[7224] = 0
      "0000000" when "00001110000111001", -- t[7225] = 0
      "0000000" when "00001110000111010", -- t[7226] = 0
      "0000000" when "00001110000111011", -- t[7227] = 0
      "0000000" when "00001110000111100", -- t[7228] = 0
      "0000000" when "00001110000111101", -- t[7229] = 0
      "0000000" when "00001110000111110", -- t[7230] = 0
      "0000000" when "00001110000111111", -- t[7231] = 0
      "0000000" when "00001110001000000", -- t[7232] = 0
      "0000000" when "00001110001000001", -- t[7233] = 0
      "0000000" when "00001110001000010", -- t[7234] = 0
      "0000000" when "00001110001000011", -- t[7235] = 0
      "0000000" when "00001110001000100", -- t[7236] = 0
      "0000000" when "00001110001000101", -- t[7237] = 0
      "0000000" when "00001110001000110", -- t[7238] = 0
      "0000000" when "00001110001000111", -- t[7239] = 0
      "0000000" when "00001110001001000", -- t[7240] = 0
      "0000000" when "00001110001001001", -- t[7241] = 0
      "0000000" when "00001110001001010", -- t[7242] = 0
      "0000000" when "00001110001001011", -- t[7243] = 0
      "0000000" when "00001110001001100", -- t[7244] = 0
      "0000000" when "00001110001001101", -- t[7245] = 0
      "0000000" when "00001110001001110", -- t[7246] = 0
      "0000000" when "00001110001001111", -- t[7247] = 0
      "0000000" when "00001110001010000", -- t[7248] = 0
      "0000000" when "00001110001010001", -- t[7249] = 0
      "0000000" when "00001110001010010", -- t[7250] = 0
      "0000000" when "00001110001010011", -- t[7251] = 0
      "0000000" when "00001110001010100", -- t[7252] = 0
      "0000000" when "00001110001010101", -- t[7253] = 0
      "0000000" when "00001110001010110", -- t[7254] = 0
      "0000000" when "00001110001010111", -- t[7255] = 0
      "0000000" when "00001110001011000", -- t[7256] = 0
      "0000000" when "00001110001011001", -- t[7257] = 0
      "0000000" when "00001110001011010", -- t[7258] = 0
      "0000000" when "00001110001011011", -- t[7259] = 0
      "0000000" when "00001110001011100", -- t[7260] = 0
      "0000000" when "00001110001011101", -- t[7261] = 0
      "0000000" when "00001110001011110", -- t[7262] = 0
      "0000000" when "00001110001011111", -- t[7263] = 0
      "0000000" when "00001110001100000", -- t[7264] = 0
      "0000000" when "00001110001100001", -- t[7265] = 0
      "0000000" when "00001110001100010", -- t[7266] = 0
      "0000000" when "00001110001100011", -- t[7267] = 0
      "0000000" when "00001110001100100", -- t[7268] = 0
      "0000000" when "00001110001100101", -- t[7269] = 0
      "0000000" when "00001110001100110", -- t[7270] = 0
      "0000000" when "00001110001100111", -- t[7271] = 0
      "0000000" when "00001110001101000", -- t[7272] = 0
      "0000000" when "00001110001101001", -- t[7273] = 0
      "0000000" when "00001110001101010", -- t[7274] = 0
      "0000000" when "00001110001101011", -- t[7275] = 0
      "0000000" when "00001110001101100", -- t[7276] = 0
      "0000000" when "00001110001101101", -- t[7277] = 0
      "0000000" when "00001110001101110", -- t[7278] = 0
      "0000000" when "00001110001101111", -- t[7279] = 0
      "0000000" when "00001110001110000", -- t[7280] = 0
      "0000000" when "00001110001110001", -- t[7281] = 0
      "0000000" when "00001110001110010", -- t[7282] = 0
      "0000000" when "00001110001110011", -- t[7283] = 0
      "0000000" when "00001110001110100", -- t[7284] = 0
      "0000000" when "00001110001110101", -- t[7285] = 0
      "0000000" when "00001110001110110", -- t[7286] = 0
      "0000000" when "00001110001110111", -- t[7287] = 0
      "0000000" when "00001110001111000", -- t[7288] = 0
      "0000000" when "00001110001111001", -- t[7289] = 0
      "0000000" when "00001110001111010", -- t[7290] = 0
      "0000000" when "00001110001111011", -- t[7291] = 0
      "0000000" when "00001110001111100", -- t[7292] = 0
      "0000000" when "00001110001111101", -- t[7293] = 0
      "0000000" when "00001110001111110", -- t[7294] = 0
      "0000000" when "00001110001111111", -- t[7295] = 0
      "0000000" when "00001110010000000", -- t[7296] = 0
      "0000000" when "00001110010000001", -- t[7297] = 0
      "0000000" when "00001110010000010", -- t[7298] = 0
      "0000000" when "00001110010000011", -- t[7299] = 0
      "0000000" when "00001110010000100", -- t[7300] = 0
      "0000000" when "00001110010000101", -- t[7301] = 0
      "0000000" when "00001110010000110", -- t[7302] = 0
      "0000000" when "00001110010000111", -- t[7303] = 0
      "0000000" when "00001110010001000", -- t[7304] = 0
      "0000000" when "00001110010001001", -- t[7305] = 0
      "0000000" when "00001110010001010", -- t[7306] = 0
      "0000000" when "00001110010001011", -- t[7307] = 0
      "0000000" when "00001110010001100", -- t[7308] = 0
      "0000000" when "00001110010001101", -- t[7309] = 0
      "0000000" when "00001110010001110", -- t[7310] = 0
      "0000000" when "00001110010001111", -- t[7311] = 0
      "0000000" when "00001110010010000", -- t[7312] = 0
      "0000000" when "00001110010010001", -- t[7313] = 0
      "0000000" when "00001110010010010", -- t[7314] = 0
      "0000000" when "00001110010010011", -- t[7315] = 0
      "0000000" when "00001110010010100", -- t[7316] = 0
      "0000000" when "00001110010010101", -- t[7317] = 0
      "0000000" when "00001110010010110", -- t[7318] = 0
      "0000000" when "00001110010010111", -- t[7319] = 0
      "0000000" when "00001110010011000", -- t[7320] = 0
      "0000000" when "00001110010011001", -- t[7321] = 0
      "0000000" when "00001110010011010", -- t[7322] = 0
      "0000000" when "00001110010011011", -- t[7323] = 0
      "0000000" when "00001110010011100", -- t[7324] = 0
      "0000000" when "00001110010011101", -- t[7325] = 0
      "0000000" when "00001110010011110", -- t[7326] = 0
      "0000000" when "00001110010011111", -- t[7327] = 0
      "0000000" when "00001110010100000", -- t[7328] = 0
      "0000000" when "00001110010100001", -- t[7329] = 0
      "0000000" when "00001110010100010", -- t[7330] = 0
      "0000000" when "00001110010100011", -- t[7331] = 0
      "0000000" when "00001110010100100", -- t[7332] = 0
      "0000000" when "00001110010100101", -- t[7333] = 0
      "0000000" when "00001110010100110", -- t[7334] = 0
      "0000000" when "00001110010100111", -- t[7335] = 0
      "0000000" when "00001110010101000", -- t[7336] = 0
      "0000000" when "00001110010101001", -- t[7337] = 0
      "0000000" when "00001110010101010", -- t[7338] = 0
      "0000000" when "00001110010101011", -- t[7339] = 0
      "0000000" when "00001110010101100", -- t[7340] = 0
      "0000000" when "00001110010101101", -- t[7341] = 0
      "0000000" when "00001110010101110", -- t[7342] = 0
      "0000000" when "00001110010101111", -- t[7343] = 0
      "0000000" when "00001110010110000", -- t[7344] = 0
      "0000000" when "00001110010110001", -- t[7345] = 0
      "0000000" when "00001110010110010", -- t[7346] = 0
      "0000000" when "00001110010110011", -- t[7347] = 0
      "0000000" when "00001110010110100", -- t[7348] = 0
      "0000000" when "00001110010110101", -- t[7349] = 0
      "0000000" when "00001110010110110", -- t[7350] = 0
      "0000000" when "00001110010110111", -- t[7351] = 0
      "0000000" when "00001110010111000", -- t[7352] = 0
      "0000000" when "00001110010111001", -- t[7353] = 0
      "0000000" when "00001110010111010", -- t[7354] = 0
      "0000000" when "00001110010111011", -- t[7355] = 0
      "0000000" when "00001110010111100", -- t[7356] = 0
      "0000000" when "00001110010111101", -- t[7357] = 0
      "0000000" when "00001110010111110", -- t[7358] = 0
      "0000000" when "00001110010111111", -- t[7359] = 0
      "0000000" when "00001110011000000", -- t[7360] = 0
      "0000000" when "00001110011000001", -- t[7361] = 0
      "0000000" when "00001110011000010", -- t[7362] = 0
      "0000000" when "00001110011000011", -- t[7363] = 0
      "0000000" when "00001110011000100", -- t[7364] = 0
      "0000000" when "00001110011000101", -- t[7365] = 0
      "0000000" when "00001110011000110", -- t[7366] = 0
      "0000000" when "00001110011000111", -- t[7367] = 0
      "0000000" when "00001110011001000", -- t[7368] = 0
      "0000000" when "00001110011001001", -- t[7369] = 0
      "0000000" when "00001110011001010", -- t[7370] = 0
      "0000000" when "00001110011001011", -- t[7371] = 0
      "0000000" when "00001110011001100", -- t[7372] = 0
      "0000000" when "00001110011001101", -- t[7373] = 0
      "0000000" when "00001110011001110", -- t[7374] = 0
      "0000000" when "00001110011001111", -- t[7375] = 0
      "0000000" when "00001110011010000", -- t[7376] = 0
      "0000000" when "00001110011010001", -- t[7377] = 0
      "0000000" when "00001110011010010", -- t[7378] = 0
      "0000000" when "00001110011010011", -- t[7379] = 0
      "0000000" when "00001110011010100", -- t[7380] = 0
      "0000000" when "00001110011010101", -- t[7381] = 0
      "0000000" when "00001110011010110", -- t[7382] = 0
      "0000000" when "00001110011010111", -- t[7383] = 0
      "0000000" when "00001110011011000", -- t[7384] = 0
      "0000000" when "00001110011011001", -- t[7385] = 0
      "0000000" when "00001110011011010", -- t[7386] = 0
      "0000000" when "00001110011011011", -- t[7387] = 0
      "0000000" when "00001110011011100", -- t[7388] = 0
      "0000000" when "00001110011011101", -- t[7389] = 0
      "0000000" when "00001110011011110", -- t[7390] = 0
      "0000000" when "00001110011011111", -- t[7391] = 0
      "0000000" when "00001110011100000", -- t[7392] = 0
      "0000000" when "00001110011100001", -- t[7393] = 0
      "0000000" when "00001110011100010", -- t[7394] = 0
      "0000000" when "00001110011100011", -- t[7395] = 0
      "0000000" when "00001110011100100", -- t[7396] = 0
      "0000000" when "00001110011100101", -- t[7397] = 0
      "0000000" when "00001110011100110", -- t[7398] = 0
      "0000000" when "00001110011100111", -- t[7399] = 0
      "0000000" when "00001110011101000", -- t[7400] = 0
      "0000000" when "00001110011101001", -- t[7401] = 0
      "0000000" when "00001110011101010", -- t[7402] = 0
      "0000000" when "00001110011101011", -- t[7403] = 0
      "0000000" when "00001110011101100", -- t[7404] = 0
      "0000000" when "00001110011101101", -- t[7405] = 0
      "0000000" when "00001110011101110", -- t[7406] = 0
      "0000000" when "00001110011101111", -- t[7407] = 0
      "0000000" when "00001110011110000", -- t[7408] = 0
      "0000000" when "00001110011110001", -- t[7409] = 0
      "0000000" when "00001110011110010", -- t[7410] = 0
      "0000000" when "00001110011110011", -- t[7411] = 0
      "0000000" when "00001110011110100", -- t[7412] = 0
      "0000000" when "00001110011110101", -- t[7413] = 0
      "0000000" when "00001110011110110", -- t[7414] = 0
      "0000000" when "00001110011110111", -- t[7415] = 0
      "0000000" when "00001110011111000", -- t[7416] = 0
      "0000000" when "00001110011111001", -- t[7417] = 0
      "0000000" when "00001110011111010", -- t[7418] = 0
      "0000000" when "00001110011111011", -- t[7419] = 0
      "0000000" when "00001110011111100", -- t[7420] = 0
      "0000000" when "00001110011111101", -- t[7421] = 0
      "0000000" when "00001110011111110", -- t[7422] = 0
      "0000000" when "00001110011111111", -- t[7423] = 0
      "0000000" when "00001110100000000", -- t[7424] = 0
      "0000000" when "00001110100000001", -- t[7425] = 0
      "0000000" when "00001110100000010", -- t[7426] = 0
      "0000000" when "00001110100000011", -- t[7427] = 0
      "0000000" when "00001110100000100", -- t[7428] = 0
      "0000000" when "00001110100000101", -- t[7429] = 0
      "0000000" when "00001110100000110", -- t[7430] = 0
      "0000000" when "00001110100000111", -- t[7431] = 0
      "0000000" when "00001110100001000", -- t[7432] = 0
      "0000000" when "00001110100001001", -- t[7433] = 0
      "0000000" when "00001110100001010", -- t[7434] = 0
      "0000000" when "00001110100001011", -- t[7435] = 0
      "0000000" when "00001110100001100", -- t[7436] = 0
      "0000000" when "00001110100001101", -- t[7437] = 0
      "0000000" when "00001110100001110", -- t[7438] = 0
      "0000000" when "00001110100001111", -- t[7439] = 0
      "0000000" when "00001110100010000", -- t[7440] = 0
      "0000000" when "00001110100010001", -- t[7441] = 0
      "0000000" when "00001110100010010", -- t[7442] = 0
      "0000000" when "00001110100010011", -- t[7443] = 0
      "0000000" when "00001110100010100", -- t[7444] = 0
      "0000000" when "00001110100010101", -- t[7445] = 0
      "0000000" when "00001110100010110", -- t[7446] = 0
      "0000000" when "00001110100010111", -- t[7447] = 0
      "0000000" when "00001110100011000", -- t[7448] = 0
      "0000000" when "00001110100011001", -- t[7449] = 0
      "0000000" when "00001110100011010", -- t[7450] = 0
      "0000000" when "00001110100011011", -- t[7451] = 0
      "0000000" when "00001110100011100", -- t[7452] = 0
      "0000000" when "00001110100011101", -- t[7453] = 0
      "0000000" when "00001110100011110", -- t[7454] = 0
      "0000000" when "00001110100011111", -- t[7455] = 0
      "0000000" when "00001110100100000", -- t[7456] = 0
      "0000000" when "00001110100100001", -- t[7457] = 0
      "0000000" when "00001110100100010", -- t[7458] = 0
      "0000000" when "00001110100100011", -- t[7459] = 0
      "0000000" when "00001110100100100", -- t[7460] = 0
      "0000000" when "00001110100100101", -- t[7461] = 0
      "0000000" when "00001110100100110", -- t[7462] = 0
      "0000000" when "00001110100100111", -- t[7463] = 0
      "0000000" when "00001110100101000", -- t[7464] = 0
      "0000000" when "00001110100101001", -- t[7465] = 0
      "0000000" when "00001110100101010", -- t[7466] = 0
      "0000000" when "00001110100101011", -- t[7467] = 0
      "0000000" when "00001110100101100", -- t[7468] = 0
      "0000000" when "00001110100101101", -- t[7469] = 0
      "0000000" when "00001110100101110", -- t[7470] = 0
      "0000000" when "00001110100101111", -- t[7471] = 0
      "0000000" when "00001110100110000", -- t[7472] = 0
      "0000000" when "00001110100110001", -- t[7473] = 0
      "0000000" when "00001110100110010", -- t[7474] = 0
      "0000000" when "00001110100110011", -- t[7475] = 0
      "0000000" when "00001110100110100", -- t[7476] = 0
      "0000000" when "00001110100110101", -- t[7477] = 0
      "0000000" when "00001110100110110", -- t[7478] = 0
      "0000000" when "00001110100110111", -- t[7479] = 0
      "0000000" when "00001110100111000", -- t[7480] = 0
      "0000000" when "00001110100111001", -- t[7481] = 0
      "0000000" when "00001110100111010", -- t[7482] = 0
      "0000000" when "00001110100111011", -- t[7483] = 0
      "0000000" when "00001110100111100", -- t[7484] = 0
      "0000000" when "00001110100111101", -- t[7485] = 0
      "0000000" when "00001110100111110", -- t[7486] = 0
      "0000000" when "00001110100111111", -- t[7487] = 0
      "0000000" when "00001110101000000", -- t[7488] = 0
      "0000000" when "00001110101000001", -- t[7489] = 0
      "0000000" when "00001110101000010", -- t[7490] = 0
      "0000000" when "00001110101000011", -- t[7491] = 0
      "0000000" when "00001110101000100", -- t[7492] = 0
      "0000000" when "00001110101000101", -- t[7493] = 0
      "0000000" when "00001110101000110", -- t[7494] = 0
      "0000000" when "00001110101000111", -- t[7495] = 0
      "0000000" when "00001110101001000", -- t[7496] = 0
      "0000000" when "00001110101001001", -- t[7497] = 0
      "0000000" when "00001110101001010", -- t[7498] = 0
      "0000000" when "00001110101001011", -- t[7499] = 0
      "0000000" when "00001110101001100", -- t[7500] = 0
      "0000000" when "00001110101001101", -- t[7501] = 0
      "0000000" when "00001110101001110", -- t[7502] = 0
      "0000000" when "00001110101001111", -- t[7503] = 0
      "0000000" when "00001110101010000", -- t[7504] = 0
      "0000000" when "00001110101010001", -- t[7505] = 0
      "0000000" when "00001110101010010", -- t[7506] = 0
      "0000000" when "00001110101010011", -- t[7507] = 0
      "0000000" when "00001110101010100", -- t[7508] = 0
      "0000000" when "00001110101010101", -- t[7509] = 0
      "0000000" when "00001110101010110", -- t[7510] = 0
      "0000000" when "00001110101010111", -- t[7511] = 0
      "0000000" when "00001110101011000", -- t[7512] = 0
      "0000000" when "00001110101011001", -- t[7513] = 0
      "0000000" when "00001110101011010", -- t[7514] = 0
      "0000000" when "00001110101011011", -- t[7515] = 0
      "0000000" when "00001110101011100", -- t[7516] = 0
      "0000000" when "00001110101011101", -- t[7517] = 0
      "0000000" when "00001110101011110", -- t[7518] = 0
      "0000000" when "00001110101011111", -- t[7519] = 0
      "0000000" when "00001110101100000", -- t[7520] = 0
      "0000000" when "00001110101100001", -- t[7521] = 0
      "0000000" when "00001110101100010", -- t[7522] = 0
      "0000000" when "00001110101100011", -- t[7523] = 0
      "0000000" when "00001110101100100", -- t[7524] = 0
      "0000000" when "00001110101100101", -- t[7525] = 0
      "0000000" when "00001110101100110", -- t[7526] = 0
      "0000000" when "00001110101100111", -- t[7527] = 0
      "0000000" when "00001110101101000", -- t[7528] = 0
      "0000000" when "00001110101101001", -- t[7529] = 0
      "0000000" when "00001110101101010", -- t[7530] = 0
      "0000000" when "00001110101101011", -- t[7531] = 0
      "0000000" when "00001110101101100", -- t[7532] = 0
      "0000000" when "00001110101101101", -- t[7533] = 0
      "0000000" when "00001110101101110", -- t[7534] = 0
      "0000000" when "00001110101101111", -- t[7535] = 0
      "0000000" when "00001110101110000", -- t[7536] = 0
      "0000000" when "00001110101110001", -- t[7537] = 0
      "0000000" when "00001110101110010", -- t[7538] = 0
      "0000000" when "00001110101110011", -- t[7539] = 0
      "0000000" when "00001110101110100", -- t[7540] = 0
      "0000000" when "00001110101110101", -- t[7541] = 0
      "0000000" when "00001110101110110", -- t[7542] = 0
      "0000000" when "00001110101110111", -- t[7543] = 0
      "0000000" when "00001110101111000", -- t[7544] = 0
      "0000000" when "00001110101111001", -- t[7545] = 0
      "0000000" when "00001110101111010", -- t[7546] = 0
      "0000000" when "00001110101111011", -- t[7547] = 0
      "0000000" when "00001110101111100", -- t[7548] = 0
      "0000000" when "00001110101111101", -- t[7549] = 0
      "0000000" when "00001110101111110", -- t[7550] = 0
      "0000000" when "00001110101111111", -- t[7551] = 0
      "0000000" when "00001110110000000", -- t[7552] = 0
      "0000000" when "00001110110000001", -- t[7553] = 0
      "0000000" when "00001110110000010", -- t[7554] = 0
      "0000000" when "00001110110000011", -- t[7555] = 0
      "0000000" when "00001110110000100", -- t[7556] = 0
      "0000000" when "00001110110000101", -- t[7557] = 0
      "0000000" when "00001110110000110", -- t[7558] = 0
      "0000000" when "00001110110000111", -- t[7559] = 0
      "0000000" when "00001110110001000", -- t[7560] = 0
      "0000000" when "00001110110001001", -- t[7561] = 0
      "0000000" when "00001110110001010", -- t[7562] = 0
      "0000000" when "00001110110001011", -- t[7563] = 0
      "0000000" when "00001110110001100", -- t[7564] = 0
      "0000000" when "00001110110001101", -- t[7565] = 0
      "0000000" when "00001110110001110", -- t[7566] = 0
      "0000000" when "00001110110001111", -- t[7567] = 0
      "0000000" when "00001110110010000", -- t[7568] = 0
      "0000000" when "00001110110010001", -- t[7569] = 0
      "0000000" when "00001110110010010", -- t[7570] = 0
      "0000000" when "00001110110010011", -- t[7571] = 0
      "0000000" when "00001110110010100", -- t[7572] = 0
      "0000000" when "00001110110010101", -- t[7573] = 0
      "0000000" when "00001110110010110", -- t[7574] = 0
      "0000000" when "00001110110010111", -- t[7575] = 0
      "0000000" when "00001110110011000", -- t[7576] = 0
      "0000000" when "00001110110011001", -- t[7577] = 0
      "0000000" when "00001110110011010", -- t[7578] = 0
      "0000000" when "00001110110011011", -- t[7579] = 0
      "0000000" when "00001110110011100", -- t[7580] = 0
      "0000000" when "00001110110011101", -- t[7581] = 0
      "0000000" when "00001110110011110", -- t[7582] = 0
      "0000000" when "00001110110011111", -- t[7583] = 0
      "0000000" when "00001110110100000", -- t[7584] = 0
      "0000000" when "00001110110100001", -- t[7585] = 0
      "0000000" when "00001110110100010", -- t[7586] = 0
      "0000000" when "00001110110100011", -- t[7587] = 0
      "0000000" when "00001110110100100", -- t[7588] = 0
      "0000000" when "00001110110100101", -- t[7589] = 0
      "0000000" when "00001110110100110", -- t[7590] = 0
      "0000000" when "00001110110100111", -- t[7591] = 0
      "0000000" when "00001110110101000", -- t[7592] = 0
      "0000000" when "00001110110101001", -- t[7593] = 0
      "0000000" when "00001110110101010", -- t[7594] = 0
      "0000000" when "00001110110101011", -- t[7595] = 0
      "0000000" when "00001110110101100", -- t[7596] = 0
      "0000000" when "00001110110101101", -- t[7597] = 0
      "0000000" when "00001110110101110", -- t[7598] = 0
      "0000000" when "00001110110101111", -- t[7599] = 0
      "0000000" when "00001110110110000", -- t[7600] = 0
      "0000000" when "00001110110110001", -- t[7601] = 0
      "0000000" when "00001110110110010", -- t[7602] = 0
      "0000000" when "00001110110110011", -- t[7603] = 0
      "0000000" when "00001110110110100", -- t[7604] = 0
      "0000000" when "00001110110110101", -- t[7605] = 0
      "0000000" when "00001110110110110", -- t[7606] = 0
      "0000000" when "00001110110110111", -- t[7607] = 0
      "0000000" when "00001110110111000", -- t[7608] = 0
      "0000000" when "00001110110111001", -- t[7609] = 0
      "0000000" when "00001110110111010", -- t[7610] = 0
      "0000000" when "00001110110111011", -- t[7611] = 0
      "0000000" when "00001110110111100", -- t[7612] = 0
      "0000000" when "00001110110111101", -- t[7613] = 0
      "0000000" when "00001110110111110", -- t[7614] = 0
      "0000000" when "00001110110111111", -- t[7615] = 0
      "0000000" when "00001110111000000", -- t[7616] = 0
      "0000000" when "00001110111000001", -- t[7617] = 0
      "0000000" when "00001110111000010", -- t[7618] = 0
      "0000000" when "00001110111000011", -- t[7619] = 0
      "0000000" when "00001110111000100", -- t[7620] = 0
      "0000000" when "00001110111000101", -- t[7621] = 0
      "0000000" when "00001110111000110", -- t[7622] = 0
      "0000000" when "00001110111000111", -- t[7623] = 0
      "0000000" when "00001110111001000", -- t[7624] = 0
      "0000000" when "00001110111001001", -- t[7625] = 0
      "0000000" when "00001110111001010", -- t[7626] = 0
      "0000000" when "00001110111001011", -- t[7627] = 0
      "0000000" when "00001110111001100", -- t[7628] = 0
      "0000000" when "00001110111001101", -- t[7629] = 0
      "0000000" when "00001110111001110", -- t[7630] = 0
      "0000000" when "00001110111001111", -- t[7631] = 0
      "0000000" when "00001110111010000", -- t[7632] = 0
      "0000000" when "00001110111010001", -- t[7633] = 0
      "0000000" when "00001110111010010", -- t[7634] = 0
      "0000000" when "00001110111010011", -- t[7635] = 0
      "0000000" when "00001110111010100", -- t[7636] = 0
      "0000000" when "00001110111010101", -- t[7637] = 0
      "0000000" when "00001110111010110", -- t[7638] = 0
      "0000000" when "00001110111010111", -- t[7639] = 0
      "0000000" when "00001110111011000", -- t[7640] = 0
      "0000000" when "00001110111011001", -- t[7641] = 0
      "0000000" when "00001110111011010", -- t[7642] = 0
      "0000000" when "00001110111011011", -- t[7643] = 0
      "0000000" when "00001110111011100", -- t[7644] = 0
      "0000000" when "00001110111011101", -- t[7645] = 0
      "0000000" when "00001110111011110", -- t[7646] = 0
      "0000000" when "00001110111011111", -- t[7647] = 0
      "0000000" when "00001110111100000", -- t[7648] = 0
      "0000000" when "00001110111100001", -- t[7649] = 0
      "0000000" when "00001110111100010", -- t[7650] = 0
      "0000000" when "00001110111100011", -- t[7651] = 0
      "0000000" when "00001110111100100", -- t[7652] = 0
      "0000000" when "00001110111100101", -- t[7653] = 0
      "0000000" when "00001110111100110", -- t[7654] = 0
      "0000000" when "00001110111100111", -- t[7655] = 0
      "0000000" when "00001110111101000", -- t[7656] = 0
      "0000000" when "00001110111101001", -- t[7657] = 0
      "0000000" when "00001110111101010", -- t[7658] = 0
      "0000000" when "00001110111101011", -- t[7659] = 0
      "0000000" when "00001110111101100", -- t[7660] = 0
      "0000000" when "00001110111101101", -- t[7661] = 0
      "0000000" when "00001110111101110", -- t[7662] = 0
      "0000000" when "00001110111101111", -- t[7663] = 0
      "0000000" when "00001110111110000", -- t[7664] = 0
      "0000000" when "00001110111110001", -- t[7665] = 0
      "0000000" when "00001110111110010", -- t[7666] = 0
      "0000000" when "00001110111110011", -- t[7667] = 0
      "0000000" when "00001110111110100", -- t[7668] = 0
      "0000000" when "00001110111110101", -- t[7669] = 0
      "0000000" when "00001110111110110", -- t[7670] = 0
      "0000000" when "00001110111110111", -- t[7671] = 0
      "0000000" when "00001110111111000", -- t[7672] = 0
      "0000000" when "00001110111111001", -- t[7673] = 0
      "0000000" when "00001110111111010", -- t[7674] = 0
      "0000000" when "00001110111111011", -- t[7675] = 0
      "0000000" when "00001110111111100", -- t[7676] = 0
      "0000000" when "00001110111111101", -- t[7677] = 0
      "0000000" when "00001110111111110", -- t[7678] = 0
      "0000000" when "00001110111111111", -- t[7679] = 0
      "0000000" when "00001111000000000", -- t[7680] = 0
      "0000000" when "00001111000000001", -- t[7681] = 0
      "0000000" when "00001111000000010", -- t[7682] = 0
      "0000000" when "00001111000000011", -- t[7683] = 0
      "0000000" when "00001111000000100", -- t[7684] = 0
      "0000000" when "00001111000000101", -- t[7685] = 0
      "0000000" when "00001111000000110", -- t[7686] = 0
      "0000000" when "00001111000000111", -- t[7687] = 0
      "0000000" when "00001111000001000", -- t[7688] = 0
      "0000000" when "00001111000001001", -- t[7689] = 0
      "0000000" when "00001111000001010", -- t[7690] = 0
      "0000000" when "00001111000001011", -- t[7691] = 0
      "0000000" when "00001111000001100", -- t[7692] = 0
      "0000000" when "00001111000001101", -- t[7693] = 0
      "0000000" when "00001111000001110", -- t[7694] = 0
      "0000000" when "00001111000001111", -- t[7695] = 0
      "0000000" when "00001111000010000", -- t[7696] = 0
      "0000000" when "00001111000010001", -- t[7697] = 0
      "0000000" when "00001111000010010", -- t[7698] = 0
      "0000000" when "00001111000010011", -- t[7699] = 0
      "0000000" when "00001111000010100", -- t[7700] = 0
      "0000000" when "00001111000010101", -- t[7701] = 0
      "0000000" when "00001111000010110", -- t[7702] = 0
      "0000000" when "00001111000010111", -- t[7703] = 0
      "0000000" when "00001111000011000", -- t[7704] = 0
      "0000000" when "00001111000011001", -- t[7705] = 0
      "0000000" when "00001111000011010", -- t[7706] = 0
      "0000000" when "00001111000011011", -- t[7707] = 0
      "0000000" when "00001111000011100", -- t[7708] = 0
      "0000000" when "00001111000011101", -- t[7709] = 0
      "0000000" when "00001111000011110", -- t[7710] = 0
      "0000000" when "00001111000011111", -- t[7711] = 0
      "0000000" when "00001111000100000", -- t[7712] = 0
      "0000000" when "00001111000100001", -- t[7713] = 0
      "0000000" when "00001111000100010", -- t[7714] = 0
      "0000000" when "00001111000100011", -- t[7715] = 0
      "0000000" when "00001111000100100", -- t[7716] = 0
      "0000000" when "00001111000100101", -- t[7717] = 0
      "0000000" when "00001111000100110", -- t[7718] = 0
      "0000000" when "00001111000100111", -- t[7719] = 0
      "0000000" when "00001111000101000", -- t[7720] = 0
      "0000000" when "00001111000101001", -- t[7721] = 0
      "0000000" when "00001111000101010", -- t[7722] = 0
      "0000000" when "00001111000101011", -- t[7723] = 0
      "0000000" when "00001111000101100", -- t[7724] = 0
      "0000000" when "00001111000101101", -- t[7725] = 0
      "0000000" when "00001111000101110", -- t[7726] = 0
      "0000000" when "00001111000101111", -- t[7727] = 0
      "0000000" when "00001111000110000", -- t[7728] = 0
      "0000000" when "00001111000110001", -- t[7729] = 0
      "0000000" when "00001111000110010", -- t[7730] = 0
      "0000000" when "00001111000110011", -- t[7731] = 0
      "0000000" when "00001111000110100", -- t[7732] = 0
      "0000000" when "00001111000110101", -- t[7733] = 0
      "0000000" when "00001111000110110", -- t[7734] = 0
      "0000000" when "00001111000110111", -- t[7735] = 0
      "0000000" when "00001111000111000", -- t[7736] = 0
      "0000000" when "00001111000111001", -- t[7737] = 0
      "0000000" when "00001111000111010", -- t[7738] = 0
      "0000000" when "00001111000111011", -- t[7739] = 0
      "0000000" when "00001111000111100", -- t[7740] = 0
      "0000000" when "00001111000111101", -- t[7741] = 0
      "0000000" when "00001111000111110", -- t[7742] = 0
      "0000000" when "00001111000111111", -- t[7743] = 0
      "0000000" when "00001111001000000", -- t[7744] = 0
      "0000000" when "00001111001000001", -- t[7745] = 0
      "0000000" when "00001111001000010", -- t[7746] = 0
      "0000000" when "00001111001000011", -- t[7747] = 0
      "0000000" when "00001111001000100", -- t[7748] = 0
      "0000000" when "00001111001000101", -- t[7749] = 0
      "0000000" when "00001111001000110", -- t[7750] = 0
      "0000000" when "00001111001000111", -- t[7751] = 0
      "0000000" when "00001111001001000", -- t[7752] = 0
      "0000000" when "00001111001001001", -- t[7753] = 0
      "0000000" when "00001111001001010", -- t[7754] = 0
      "0000000" when "00001111001001011", -- t[7755] = 0
      "0000000" when "00001111001001100", -- t[7756] = 0
      "0000000" when "00001111001001101", -- t[7757] = 0
      "0000000" when "00001111001001110", -- t[7758] = 0
      "0000000" when "00001111001001111", -- t[7759] = 0
      "0000000" when "00001111001010000", -- t[7760] = 0
      "0000000" when "00001111001010001", -- t[7761] = 0
      "0000000" when "00001111001010010", -- t[7762] = 0
      "0000000" when "00001111001010011", -- t[7763] = 0
      "0000000" when "00001111001010100", -- t[7764] = 0
      "0000000" when "00001111001010101", -- t[7765] = 0
      "0000000" when "00001111001010110", -- t[7766] = 0
      "0000000" when "00001111001010111", -- t[7767] = 0
      "0000000" when "00001111001011000", -- t[7768] = 0
      "0000000" when "00001111001011001", -- t[7769] = 0
      "0000000" when "00001111001011010", -- t[7770] = 0
      "0000000" when "00001111001011011", -- t[7771] = 0
      "0000000" when "00001111001011100", -- t[7772] = 0
      "0000000" when "00001111001011101", -- t[7773] = 0
      "0000000" when "00001111001011110", -- t[7774] = 0
      "0000000" when "00001111001011111", -- t[7775] = 0
      "0000000" when "00001111001100000", -- t[7776] = 0
      "0000000" when "00001111001100001", -- t[7777] = 0
      "0000000" when "00001111001100010", -- t[7778] = 0
      "0000000" when "00001111001100011", -- t[7779] = 0
      "0000000" when "00001111001100100", -- t[7780] = 0
      "0000000" when "00001111001100101", -- t[7781] = 0
      "0000000" when "00001111001100110", -- t[7782] = 0
      "0000000" when "00001111001100111", -- t[7783] = 0
      "0000000" when "00001111001101000", -- t[7784] = 0
      "0000000" when "00001111001101001", -- t[7785] = 0
      "0000000" when "00001111001101010", -- t[7786] = 0
      "0000000" when "00001111001101011", -- t[7787] = 0
      "0000000" when "00001111001101100", -- t[7788] = 0
      "0000000" when "00001111001101101", -- t[7789] = 0
      "0000000" when "00001111001101110", -- t[7790] = 0
      "0000000" when "00001111001101111", -- t[7791] = 0
      "0000000" when "00001111001110000", -- t[7792] = 0
      "0000000" when "00001111001110001", -- t[7793] = 0
      "0000000" when "00001111001110010", -- t[7794] = 0
      "0000000" when "00001111001110011", -- t[7795] = 0
      "0000000" when "00001111001110100", -- t[7796] = 0
      "0000000" when "00001111001110101", -- t[7797] = 0
      "0000000" when "00001111001110110", -- t[7798] = 0
      "0000000" when "00001111001110111", -- t[7799] = 0
      "0000000" when "00001111001111000", -- t[7800] = 0
      "0000000" when "00001111001111001", -- t[7801] = 0
      "0000000" when "00001111001111010", -- t[7802] = 0
      "0000000" when "00001111001111011", -- t[7803] = 0
      "0000000" when "00001111001111100", -- t[7804] = 0
      "0000000" when "00001111001111101", -- t[7805] = 0
      "0000000" when "00001111001111110", -- t[7806] = 0
      "0000000" when "00001111001111111", -- t[7807] = 0
      "0000000" when "00001111010000000", -- t[7808] = 0
      "0000000" when "00001111010000001", -- t[7809] = 0
      "0000000" when "00001111010000010", -- t[7810] = 0
      "0000000" when "00001111010000011", -- t[7811] = 0
      "0000000" when "00001111010000100", -- t[7812] = 0
      "0000000" when "00001111010000101", -- t[7813] = 0
      "0000000" when "00001111010000110", -- t[7814] = 0
      "0000000" when "00001111010000111", -- t[7815] = 0
      "0000000" when "00001111010001000", -- t[7816] = 0
      "0000000" when "00001111010001001", -- t[7817] = 0
      "0000000" when "00001111010001010", -- t[7818] = 0
      "0000000" when "00001111010001011", -- t[7819] = 0
      "0000000" when "00001111010001100", -- t[7820] = 0
      "0000000" when "00001111010001101", -- t[7821] = 0
      "0000000" when "00001111010001110", -- t[7822] = 0
      "0000000" when "00001111010001111", -- t[7823] = 0
      "0000000" when "00001111010010000", -- t[7824] = 0
      "0000000" when "00001111010010001", -- t[7825] = 0
      "0000000" when "00001111010010010", -- t[7826] = 0
      "0000000" when "00001111010010011", -- t[7827] = 0
      "0000000" when "00001111010010100", -- t[7828] = 0
      "0000000" when "00001111010010101", -- t[7829] = 0
      "0000000" when "00001111010010110", -- t[7830] = 0
      "0000000" when "00001111010010111", -- t[7831] = 0
      "0000000" when "00001111010011000", -- t[7832] = 0
      "0000000" when "00001111010011001", -- t[7833] = 0
      "0000000" when "00001111010011010", -- t[7834] = 0
      "0000000" when "00001111010011011", -- t[7835] = 0
      "0000000" when "00001111010011100", -- t[7836] = 0
      "0000000" when "00001111010011101", -- t[7837] = 0
      "0000000" when "00001111010011110", -- t[7838] = 0
      "0000000" when "00001111010011111", -- t[7839] = 0
      "0000000" when "00001111010100000", -- t[7840] = 0
      "0000000" when "00001111010100001", -- t[7841] = 0
      "0000000" when "00001111010100010", -- t[7842] = 0
      "0000000" when "00001111010100011", -- t[7843] = 0
      "0000000" when "00001111010100100", -- t[7844] = 0
      "0000000" when "00001111010100101", -- t[7845] = 0
      "0000000" when "00001111010100110", -- t[7846] = 0
      "0000000" when "00001111010100111", -- t[7847] = 0
      "0000000" when "00001111010101000", -- t[7848] = 0
      "0000000" when "00001111010101001", -- t[7849] = 0
      "0000000" when "00001111010101010", -- t[7850] = 0
      "0000000" when "00001111010101011", -- t[7851] = 0
      "0000000" when "00001111010101100", -- t[7852] = 0
      "0000000" when "00001111010101101", -- t[7853] = 0
      "0000000" when "00001111010101110", -- t[7854] = 0
      "0000000" when "00001111010101111", -- t[7855] = 0
      "0000000" when "00001111010110000", -- t[7856] = 0
      "0000000" when "00001111010110001", -- t[7857] = 0
      "0000000" when "00001111010110010", -- t[7858] = 0
      "0000000" when "00001111010110011", -- t[7859] = 0
      "0000000" when "00001111010110100", -- t[7860] = 0
      "0000000" when "00001111010110101", -- t[7861] = 0
      "0000000" when "00001111010110110", -- t[7862] = 0
      "0000000" when "00001111010110111", -- t[7863] = 0
      "0000000" when "00001111010111000", -- t[7864] = 0
      "0000000" when "00001111010111001", -- t[7865] = 0
      "0000000" when "00001111010111010", -- t[7866] = 0
      "0000000" when "00001111010111011", -- t[7867] = 0
      "0000000" when "00001111010111100", -- t[7868] = 0
      "0000000" when "00001111010111101", -- t[7869] = 0
      "0000000" when "00001111010111110", -- t[7870] = 0
      "0000000" when "00001111010111111", -- t[7871] = 0
      "0000000" when "00001111011000000", -- t[7872] = 0
      "0000000" when "00001111011000001", -- t[7873] = 0
      "0000000" when "00001111011000010", -- t[7874] = 0
      "0000000" when "00001111011000011", -- t[7875] = 0
      "0000000" when "00001111011000100", -- t[7876] = 0
      "0000000" when "00001111011000101", -- t[7877] = 0
      "0000000" when "00001111011000110", -- t[7878] = 0
      "0000000" when "00001111011000111", -- t[7879] = 0
      "0000000" when "00001111011001000", -- t[7880] = 0
      "0000000" when "00001111011001001", -- t[7881] = 0
      "0000000" when "00001111011001010", -- t[7882] = 0
      "0000000" when "00001111011001011", -- t[7883] = 0
      "0000000" when "00001111011001100", -- t[7884] = 0
      "0000000" when "00001111011001101", -- t[7885] = 0
      "0000000" when "00001111011001110", -- t[7886] = 0
      "0000000" when "00001111011001111", -- t[7887] = 0
      "0000000" when "00001111011010000", -- t[7888] = 0
      "0000000" when "00001111011010001", -- t[7889] = 0
      "0000000" when "00001111011010010", -- t[7890] = 0
      "0000000" when "00001111011010011", -- t[7891] = 0
      "0000000" when "00001111011010100", -- t[7892] = 0
      "0000000" when "00001111011010101", -- t[7893] = 0
      "0000000" when "00001111011010110", -- t[7894] = 0
      "0000000" when "00001111011010111", -- t[7895] = 0
      "0000000" when "00001111011011000", -- t[7896] = 0
      "0000000" when "00001111011011001", -- t[7897] = 0
      "0000000" when "00001111011011010", -- t[7898] = 0
      "0000000" when "00001111011011011", -- t[7899] = 0
      "0000000" when "00001111011011100", -- t[7900] = 0
      "0000000" when "00001111011011101", -- t[7901] = 0
      "0000000" when "00001111011011110", -- t[7902] = 0
      "0000000" when "00001111011011111", -- t[7903] = 0
      "0000000" when "00001111011100000", -- t[7904] = 0
      "0000000" when "00001111011100001", -- t[7905] = 0
      "0000000" when "00001111011100010", -- t[7906] = 0
      "0000000" when "00001111011100011", -- t[7907] = 0
      "0000000" when "00001111011100100", -- t[7908] = 0
      "0000000" when "00001111011100101", -- t[7909] = 0
      "0000000" when "00001111011100110", -- t[7910] = 0
      "0000000" when "00001111011100111", -- t[7911] = 0
      "0000000" when "00001111011101000", -- t[7912] = 0
      "0000000" when "00001111011101001", -- t[7913] = 0
      "0000000" when "00001111011101010", -- t[7914] = 0
      "0000000" when "00001111011101011", -- t[7915] = 0
      "0000000" when "00001111011101100", -- t[7916] = 0
      "0000000" when "00001111011101101", -- t[7917] = 0
      "0000000" when "00001111011101110", -- t[7918] = 0
      "0000000" when "00001111011101111", -- t[7919] = 0
      "0000000" when "00001111011110000", -- t[7920] = 0
      "0000000" when "00001111011110001", -- t[7921] = 0
      "0000000" when "00001111011110010", -- t[7922] = 0
      "0000000" when "00001111011110011", -- t[7923] = 0
      "0000000" when "00001111011110100", -- t[7924] = 0
      "0000000" when "00001111011110101", -- t[7925] = 0
      "0000000" when "00001111011110110", -- t[7926] = 0
      "0000000" when "00001111011110111", -- t[7927] = 0
      "0000000" when "00001111011111000", -- t[7928] = 0
      "0000000" when "00001111011111001", -- t[7929] = 0
      "0000000" when "00001111011111010", -- t[7930] = 0
      "0000000" when "00001111011111011", -- t[7931] = 0
      "0000000" when "00001111011111100", -- t[7932] = 0
      "0000000" when "00001111011111101", -- t[7933] = 0
      "0000000" when "00001111011111110", -- t[7934] = 0
      "0000000" when "00001111011111111", -- t[7935] = 0
      "0000000" when "00001111100000000", -- t[7936] = 0
      "0000000" when "00001111100000001", -- t[7937] = 0
      "0000000" when "00001111100000010", -- t[7938] = 0
      "0000000" when "00001111100000011", -- t[7939] = 0
      "0000000" when "00001111100000100", -- t[7940] = 0
      "0000000" when "00001111100000101", -- t[7941] = 0
      "0000000" when "00001111100000110", -- t[7942] = 0
      "0000000" when "00001111100000111", -- t[7943] = 0
      "0000000" when "00001111100001000", -- t[7944] = 0
      "0000000" when "00001111100001001", -- t[7945] = 0
      "0000000" when "00001111100001010", -- t[7946] = 0
      "0000000" when "00001111100001011", -- t[7947] = 0
      "0000000" when "00001111100001100", -- t[7948] = 0
      "0000000" when "00001111100001101", -- t[7949] = 0
      "0000000" when "00001111100001110", -- t[7950] = 0
      "0000000" when "00001111100001111", -- t[7951] = 0
      "0000000" when "00001111100010000", -- t[7952] = 0
      "0000000" when "00001111100010001", -- t[7953] = 0
      "0000000" when "00001111100010010", -- t[7954] = 0
      "0000000" when "00001111100010011", -- t[7955] = 0
      "0000000" when "00001111100010100", -- t[7956] = 0
      "0000000" when "00001111100010101", -- t[7957] = 0
      "0000000" when "00001111100010110", -- t[7958] = 0
      "0000000" when "00001111100010111", -- t[7959] = 0
      "0000000" when "00001111100011000", -- t[7960] = 0
      "0000000" when "00001111100011001", -- t[7961] = 0
      "0000000" when "00001111100011010", -- t[7962] = 0
      "0000000" when "00001111100011011", -- t[7963] = 0
      "0000000" when "00001111100011100", -- t[7964] = 0
      "0000000" when "00001111100011101", -- t[7965] = 0
      "0000000" when "00001111100011110", -- t[7966] = 0
      "0000000" when "00001111100011111", -- t[7967] = 0
      "0000000" when "00001111100100000", -- t[7968] = 0
      "0000000" when "00001111100100001", -- t[7969] = 0
      "0000000" when "00001111100100010", -- t[7970] = 0
      "0000000" when "00001111100100011", -- t[7971] = 0
      "0000000" when "00001111100100100", -- t[7972] = 0
      "0000000" when "00001111100100101", -- t[7973] = 0
      "0000000" when "00001111100100110", -- t[7974] = 0
      "0000000" when "00001111100100111", -- t[7975] = 0
      "0000000" when "00001111100101000", -- t[7976] = 0
      "0000000" when "00001111100101001", -- t[7977] = 0
      "0000000" when "00001111100101010", -- t[7978] = 0
      "0000000" when "00001111100101011", -- t[7979] = 0
      "0000000" when "00001111100101100", -- t[7980] = 0
      "0000000" when "00001111100101101", -- t[7981] = 0
      "0000000" when "00001111100101110", -- t[7982] = 0
      "0000000" when "00001111100101111", -- t[7983] = 0
      "0000000" when "00001111100110000", -- t[7984] = 0
      "0000000" when "00001111100110001", -- t[7985] = 0
      "0000000" when "00001111100110010", -- t[7986] = 0
      "0000000" when "00001111100110011", -- t[7987] = 0
      "0000000" when "00001111100110100", -- t[7988] = 0
      "0000000" when "00001111100110101", -- t[7989] = 0
      "0000000" when "00001111100110110", -- t[7990] = 0
      "0000000" when "00001111100110111", -- t[7991] = 0
      "0000000" when "00001111100111000", -- t[7992] = 0
      "0000000" when "00001111100111001", -- t[7993] = 0
      "0000000" when "00001111100111010", -- t[7994] = 0
      "0000000" when "00001111100111011", -- t[7995] = 0
      "0000000" when "00001111100111100", -- t[7996] = 0
      "0000000" when "00001111100111101", -- t[7997] = 0
      "0000000" when "00001111100111110", -- t[7998] = 0
      "0000000" when "00001111100111111", -- t[7999] = 0
      "0000000" when "00001111101000000", -- t[8000] = 0
      "0000000" when "00001111101000001", -- t[8001] = 0
      "0000000" when "00001111101000010", -- t[8002] = 0
      "0000000" when "00001111101000011", -- t[8003] = 0
      "0000000" when "00001111101000100", -- t[8004] = 0
      "0000000" when "00001111101000101", -- t[8005] = 0
      "0000000" when "00001111101000110", -- t[8006] = 0
      "0000000" when "00001111101000111", -- t[8007] = 0
      "0000000" when "00001111101001000", -- t[8008] = 0
      "0000000" when "00001111101001001", -- t[8009] = 0
      "0000000" when "00001111101001010", -- t[8010] = 0
      "0000000" when "00001111101001011", -- t[8011] = 0
      "0000000" when "00001111101001100", -- t[8012] = 0
      "0000000" when "00001111101001101", -- t[8013] = 0
      "0000000" when "00001111101001110", -- t[8014] = 0
      "0000000" when "00001111101001111", -- t[8015] = 0
      "0000000" when "00001111101010000", -- t[8016] = 0
      "0000000" when "00001111101010001", -- t[8017] = 0
      "0000000" when "00001111101010010", -- t[8018] = 0
      "0000000" when "00001111101010011", -- t[8019] = 0
      "0000000" when "00001111101010100", -- t[8020] = 0
      "0000000" when "00001111101010101", -- t[8021] = 0
      "0000000" when "00001111101010110", -- t[8022] = 0
      "0000000" when "00001111101010111", -- t[8023] = 0
      "0000000" when "00001111101011000", -- t[8024] = 0
      "0000000" when "00001111101011001", -- t[8025] = 0
      "0000000" when "00001111101011010", -- t[8026] = 0
      "0000000" when "00001111101011011", -- t[8027] = 0
      "0000000" when "00001111101011100", -- t[8028] = 0
      "0000000" when "00001111101011101", -- t[8029] = 0
      "0000000" when "00001111101011110", -- t[8030] = 0
      "0000000" when "00001111101011111", -- t[8031] = 0
      "0000000" when "00001111101100000", -- t[8032] = 0
      "0000000" when "00001111101100001", -- t[8033] = 0
      "0000000" when "00001111101100010", -- t[8034] = 0
      "0000000" when "00001111101100011", -- t[8035] = 0
      "0000000" when "00001111101100100", -- t[8036] = 0
      "0000000" when "00001111101100101", -- t[8037] = 0
      "0000000" when "00001111101100110", -- t[8038] = 0
      "0000000" when "00001111101100111", -- t[8039] = 0
      "0000000" when "00001111101101000", -- t[8040] = 0
      "0000000" when "00001111101101001", -- t[8041] = 0
      "0000000" when "00001111101101010", -- t[8042] = 0
      "0000000" when "00001111101101011", -- t[8043] = 0
      "0000000" when "00001111101101100", -- t[8044] = 0
      "0000000" when "00001111101101101", -- t[8045] = 0
      "0000000" when "00001111101101110", -- t[8046] = 0
      "0000000" when "00001111101101111", -- t[8047] = 0
      "0000000" when "00001111101110000", -- t[8048] = 0
      "0000000" when "00001111101110001", -- t[8049] = 0
      "0000000" when "00001111101110010", -- t[8050] = 0
      "0000000" when "00001111101110011", -- t[8051] = 0
      "0000000" when "00001111101110100", -- t[8052] = 0
      "0000000" when "00001111101110101", -- t[8053] = 0
      "0000000" when "00001111101110110", -- t[8054] = 0
      "0000000" when "00001111101110111", -- t[8055] = 0
      "0000000" when "00001111101111000", -- t[8056] = 0
      "0000000" when "00001111101111001", -- t[8057] = 0
      "0000000" when "00001111101111010", -- t[8058] = 0
      "0000000" when "00001111101111011", -- t[8059] = 0
      "0000000" when "00001111101111100", -- t[8060] = 0
      "0000000" when "00001111101111101", -- t[8061] = 0
      "0000000" when "00001111101111110", -- t[8062] = 0
      "0000000" when "00001111101111111", -- t[8063] = 0
      "0000000" when "00001111110000000", -- t[8064] = 0
      "0000000" when "00001111110000001", -- t[8065] = 0
      "0000000" when "00001111110000010", -- t[8066] = 0
      "0000000" when "00001111110000011", -- t[8067] = 0
      "0000000" when "00001111110000100", -- t[8068] = 0
      "0000000" when "00001111110000101", -- t[8069] = 0
      "0000000" when "00001111110000110", -- t[8070] = 0
      "0000000" when "00001111110000111", -- t[8071] = 0
      "0000000" when "00001111110001000", -- t[8072] = 0
      "0000000" when "00001111110001001", -- t[8073] = 0
      "0000000" when "00001111110001010", -- t[8074] = 0
      "0000000" when "00001111110001011", -- t[8075] = 0
      "0000000" when "00001111110001100", -- t[8076] = 0
      "0000000" when "00001111110001101", -- t[8077] = 0
      "0000000" when "00001111110001110", -- t[8078] = 0
      "0000000" when "00001111110001111", -- t[8079] = 0
      "0000000" when "00001111110010000", -- t[8080] = 0
      "0000000" when "00001111110010001", -- t[8081] = 0
      "0000000" when "00001111110010010", -- t[8082] = 0
      "0000000" when "00001111110010011", -- t[8083] = 0
      "0000000" when "00001111110010100", -- t[8084] = 0
      "0000000" when "00001111110010101", -- t[8085] = 0
      "0000000" when "00001111110010110", -- t[8086] = 0
      "0000000" when "00001111110010111", -- t[8087] = 0
      "0000000" when "00001111110011000", -- t[8088] = 0
      "0000000" when "00001111110011001", -- t[8089] = 0
      "0000000" when "00001111110011010", -- t[8090] = 0
      "0000000" when "00001111110011011", -- t[8091] = 0
      "0000000" when "00001111110011100", -- t[8092] = 0
      "0000000" when "00001111110011101", -- t[8093] = 0
      "0000000" when "00001111110011110", -- t[8094] = 0
      "0000000" when "00001111110011111", -- t[8095] = 0
      "0000000" when "00001111110100000", -- t[8096] = 0
      "0000000" when "00001111110100001", -- t[8097] = 0
      "0000000" when "00001111110100010", -- t[8098] = 0
      "0000000" when "00001111110100011", -- t[8099] = 0
      "0000000" when "00001111110100100", -- t[8100] = 0
      "0000000" when "00001111110100101", -- t[8101] = 0
      "0000000" when "00001111110100110", -- t[8102] = 0
      "0000000" when "00001111110100111", -- t[8103] = 0
      "0000000" when "00001111110101000", -- t[8104] = 0
      "0000000" when "00001111110101001", -- t[8105] = 0
      "0000000" when "00001111110101010", -- t[8106] = 0
      "0000000" when "00001111110101011", -- t[8107] = 0
      "0000000" when "00001111110101100", -- t[8108] = 0
      "0000000" when "00001111110101101", -- t[8109] = 0
      "0000000" when "00001111110101110", -- t[8110] = 0
      "0000000" when "00001111110101111", -- t[8111] = 0
      "0000000" when "00001111110110000", -- t[8112] = 0
      "0000000" when "00001111110110001", -- t[8113] = 0
      "0000000" when "00001111110110010", -- t[8114] = 0
      "0000000" when "00001111110110011", -- t[8115] = 0
      "0000000" when "00001111110110100", -- t[8116] = 0
      "0000000" when "00001111110110101", -- t[8117] = 0
      "0000000" when "00001111110110110", -- t[8118] = 0
      "0000000" when "00001111110110111", -- t[8119] = 0
      "0000000" when "00001111110111000", -- t[8120] = 0
      "0000000" when "00001111110111001", -- t[8121] = 0
      "0000000" when "00001111110111010", -- t[8122] = 0
      "0000000" when "00001111110111011", -- t[8123] = 0
      "0000000" when "00001111110111100", -- t[8124] = 0
      "0000000" when "00001111110111101", -- t[8125] = 0
      "0000000" when "00001111110111110", -- t[8126] = 0
      "0000000" when "00001111110111111", -- t[8127] = 0
      "0000000" when "00001111111000000", -- t[8128] = 0
      "0000000" when "00001111111000001", -- t[8129] = 0
      "0000000" when "00001111111000010", -- t[8130] = 0
      "0000000" when "00001111111000011", -- t[8131] = 0
      "0000000" when "00001111111000100", -- t[8132] = 0
      "0000000" when "00001111111000101", -- t[8133] = 0
      "0000000" when "00001111111000110", -- t[8134] = 0
      "0000000" when "00001111111000111", -- t[8135] = 0
      "0000000" when "00001111111001000", -- t[8136] = 0
      "0000000" when "00001111111001001", -- t[8137] = 0
      "0000000" when "00001111111001010", -- t[8138] = 0
      "0000000" when "00001111111001011", -- t[8139] = 0
      "0000000" when "00001111111001100", -- t[8140] = 0
      "0000000" when "00001111111001101", -- t[8141] = 0
      "0000000" when "00001111111001110", -- t[8142] = 0
      "0000000" when "00001111111001111", -- t[8143] = 0
      "0000000" when "00001111111010000", -- t[8144] = 0
      "0000000" when "00001111111010001", -- t[8145] = 0
      "0000000" when "00001111111010010", -- t[8146] = 0
      "0000000" when "00001111111010011", -- t[8147] = 0
      "0000000" when "00001111111010100", -- t[8148] = 0
      "0000000" when "00001111111010101", -- t[8149] = 0
      "0000000" when "00001111111010110", -- t[8150] = 0
      "0000000" when "00001111111010111", -- t[8151] = 0
      "0000000" when "00001111111011000", -- t[8152] = 0
      "0000000" when "00001111111011001", -- t[8153] = 0
      "0000000" when "00001111111011010", -- t[8154] = 0
      "0000000" when "00001111111011011", -- t[8155] = 0
      "0000000" when "00001111111011100", -- t[8156] = 0
      "0000000" when "00001111111011101", -- t[8157] = 0
      "0000000" when "00001111111011110", -- t[8158] = 0
      "0000000" when "00001111111011111", -- t[8159] = 0
      "0000000" when "00001111111100000", -- t[8160] = 0
      "0000000" when "00001111111100001", -- t[8161] = 0
      "0000000" when "00001111111100010", -- t[8162] = 0
      "0000000" when "00001111111100011", -- t[8163] = 0
      "0000000" when "00001111111100100", -- t[8164] = 0
      "0000000" when "00001111111100101", -- t[8165] = 0
      "0000000" when "00001111111100110", -- t[8166] = 0
      "0000000" when "00001111111100111", -- t[8167] = 0
      "0000000" when "00001111111101000", -- t[8168] = 0
      "0000000" when "00001111111101001", -- t[8169] = 0
      "0000000" when "00001111111101010", -- t[8170] = 0
      "0000000" when "00001111111101011", -- t[8171] = 0
      "0000000" when "00001111111101100", -- t[8172] = 0
      "0000000" when "00001111111101101", -- t[8173] = 0
      "0000000" when "00001111111101110", -- t[8174] = 0
      "0000000" when "00001111111101111", -- t[8175] = 0
      "0000000" when "00001111111110000", -- t[8176] = 0
      "0000000" when "00001111111110001", -- t[8177] = 0
      "0000000" when "00001111111110010", -- t[8178] = 0
      "0000000" when "00001111111110011", -- t[8179] = 0
      "0000000" when "00001111111110100", -- t[8180] = 0
      "0000000" when "00001111111110101", -- t[8181] = 0
      "0000000" when "00001111111110110", -- t[8182] = 0
      "0000000" when "00001111111110111", -- t[8183] = 0
      "0000000" when "00001111111111000", -- t[8184] = 0
      "0000000" when "00001111111111001", -- t[8185] = 0
      "0000000" when "00001111111111010", -- t[8186] = 0
      "0000000" when "00001111111111011", -- t[8187] = 0
      "0000000" when "00001111111111100", -- t[8188] = 0
      "0000000" when "00001111111111101", -- t[8189] = 0
      "0000000" when "00001111111111110", -- t[8190] = 0
      "0000000" when "00001111111111111", -- t[8191] = 0
      "0000000" when "00010000000000000", -- t[8192] = 0
      "0000000" when "00010000000000001", -- t[8193] = 0
      "0000000" when "00010000000000010", -- t[8194] = 0
      "0000000" when "00010000000000011", -- t[8195] = 0
      "0000000" when "00010000000000100", -- t[8196] = 0
      "0000000" when "00010000000000101", -- t[8197] = 0
      "0000000" when "00010000000000110", -- t[8198] = 0
      "0000000" when "00010000000000111", -- t[8199] = 0
      "0000000" when "00010000000001000", -- t[8200] = 0
      "0000000" when "00010000000001001", -- t[8201] = 0
      "0000000" when "00010000000001010", -- t[8202] = 0
      "0000000" when "00010000000001011", -- t[8203] = 0
      "0000000" when "00010000000001100", -- t[8204] = 0
      "0000000" when "00010000000001101", -- t[8205] = 0
      "0000000" when "00010000000001110", -- t[8206] = 0
      "0000000" when "00010000000001111", -- t[8207] = 0
      "0000000" when "00010000000010000", -- t[8208] = 0
      "0000000" when "00010000000010001", -- t[8209] = 0
      "0000000" when "00010000000010010", -- t[8210] = 0
      "0000000" when "00010000000010011", -- t[8211] = 0
      "0000000" when "00010000000010100", -- t[8212] = 0
      "0000000" when "00010000000010101", -- t[8213] = 0
      "0000000" when "00010000000010110", -- t[8214] = 0
      "0000000" when "00010000000010111", -- t[8215] = 0
      "0000000" when "00010000000011000", -- t[8216] = 0
      "0000000" when "00010000000011001", -- t[8217] = 0
      "0000000" when "00010000000011010", -- t[8218] = 0
      "0000000" when "00010000000011011", -- t[8219] = 0
      "0000000" when "00010000000011100", -- t[8220] = 0
      "0000000" when "00010000000011101", -- t[8221] = 0
      "0000000" when "00010000000011110", -- t[8222] = 0
      "0000000" when "00010000000011111", -- t[8223] = 0
      "0000000" when "00010000000100000", -- t[8224] = 0
      "0000000" when "00010000000100001", -- t[8225] = 0
      "0000000" when "00010000000100010", -- t[8226] = 0
      "0000000" when "00010000000100011", -- t[8227] = 0
      "0000000" when "00010000000100100", -- t[8228] = 0
      "0000000" when "00010000000100101", -- t[8229] = 0
      "0000000" when "00010000000100110", -- t[8230] = 0
      "0000000" when "00010000000100111", -- t[8231] = 0
      "0000000" when "00010000000101000", -- t[8232] = 0
      "0000000" when "00010000000101001", -- t[8233] = 0
      "0000000" when "00010000000101010", -- t[8234] = 0
      "0000000" when "00010000000101011", -- t[8235] = 0
      "0000000" when "00010000000101100", -- t[8236] = 0
      "0000000" when "00010000000101101", -- t[8237] = 0
      "0000000" when "00010000000101110", -- t[8238] = 0
      "0000000" when "00010000000101111", -- t[8239] = 0
      "0000000" when "00010000000110000", -- t[8240] = 0
      "0000000" when "00010000000110001", -- t[8241] = 0
      "0000000" when "00010000000110010", -- t[8242] = 0
      "0000000" when "00010000000110011", -- t[8243] = 0
      "0000000" when "00010000000110100", -- t[8244] = 0
      "0000000" when "00010000000110101", -- t[8245] = 0
      "0000000" when "00010000000110110", -- t[8246] = 0
      "0000000" when "00010000000110111", -- t[8247] = 0
      "0000000" when "00010000000111000", -- t[8248] = 0
      "0000000" when "00010000000111001", -- t[8249] = 0
      "0000000" when "00010000000111010", -- t[8250] = 0
      "0000000" when "00010000000111011", -- t[8251] = 0
      "0000000" when "00010000000111100", -- t[8252] = 0
      "0000000" when "00010000000111101", -- t[8253] = 0
      "0000000" when "00010000000111110", -- t[8254] = 0
      "0000000" when "00010000000111111", -- t[8255] = 0
      "0000000" when "00010000001000000", -- t[8256] = 0
      "0000000" when "00010000001000001", -- t[8257] = 0
      "0000000" when "00010000001000010", -- t[8258] = 0
      "0000000" when "00010000001000011", -- t[8259] = 0
      "0000000" when "00010000001000100", -- t[8260] = 0
      "0000000" when "00010000001000101", -- t[8261] = 0
      "0000000" when "00010000001000110", -- t[8262] = 0
      "0000000" when "00010000001000111", -- t[8263] = 0
      "0000000" when "00010000001001000", -- t[8264] = 0
      "0000000" when "00010000001001001", -- t[8265] = 0
      "0000000" when "00010000001001010", -- t[8266] = 0
      "0000000" when "00010000001001011", -- t[8267] = 0
      "0000000" when "00010000001001100", -- t[8268] = 0
      "0000000" when "00010000001001101", -- t[8269] = 0
      "0000000" when "00010000001001110", -- t[8270] = 0
      "0000000" when "00010000001001111", -- t[8271] = 0
      "0000000" when "00010000001010000", -- t[8272] = 0
      "0000000" when "00010000001010001", -- t[8273] = 0
      "0000000" when "00010000001010010", -- t[8274] = 0
      "0000000" when "00010000001010011", -- t[8275] = 0
      "0000000" when "00010000001010100", -- t[8276] = 0
      "0000000" when "00010000001010101", -- t[8277] = 0
      "0000000" when "00010000001010110", -- t[8278] = 0
      "0000000" when "00010000001010111", -- t[8279] = 0
      "0000000" when "00010000001011000", -- t[8280] = 0
      "0000000" when "00010000001011001", -- t[8281] = 0
      "0000000" when "00010000001011010", -- t[8282] = 0
      "0000000" when "00010000001011011", -- t[8283] = 0
      "0000000" when "00010000001011100", -- t[8284] = 0
      "0000000" when "00010000001011101", -- t[8285] = 0
      "0000000" when "00010000001011110", -- t[8286] = 0
      "0000000" when "00010000001011111", -- t[8287] = 0
      "0000000" when "00010000001100000", -- t[8288] = 0
      "0000000" when "00010000001100001", -- t[8289] = 0
      "0000000" when "00010000001100010", -- t[8290] = 0
      "0000000" when "00010000001100011", -- t[8291] = 0
      "0000000" when "00010000001100100", -- t[8292] = 0
      "0000000" when "00010000001100101", -- t[8293] = 0
      "0000000" when "00010000001100110", -- t[8294] = 0
      "0000000" when "00010000001100111", -- t[8295] = 0
      "0000000" when "00010000001101000", -- t[8296] = 0
      "0000000" when "00010000001101001", -- t[8297] = 0
      "0000000" when "00010000001101010", -- t[8298] = 0
      "0000000" when "00010000001101011", -- t[8299] = 0
      "0000000" when "00010000001101100", -- t[8300] = 0
      "0000000" when "00010000001101101", -- t[8301] = 0
      "0000000" when "00010000001101110", -- t[8302] = 0
      "0000000" when "00010000001101111", -- t[8303] = 0
      "0000000" when "00010000001110000", -- t[8304] = 0
      "0000000" when "00010000001110001", -- t[8305] = 0
      "0000000" when "00010000001110010", -- t[8306] = 0
      "0000000" when "00010000001110011", -- t[8307] = 0
      "0000000" when "00010000001110100", -- t[8308] = 0
      "0000000" when "00010000001110101", -- t[8309] = 0
      "0000000" when "00010000001110110", -- t[8310] = 0
      "0000000" when "00010000001110111", -- t[8311] = 0
      "0000000" when "00010000001111000", -- t[8312] = 0
      "0000000" when "00010000001111001", -- t[8313] = 0
      "0000000" when "00010000001111010", -- t[8314] = 0
      "0000000" when "00010000001111011", -- t[8315] = 0
      "0000000" when "00010000001111100", -- t[8316] = 0
      "0000000" when "00010000001111101", -- t[8317] = 0
      "0000000" when "00010000001111110", -- t[8318] = 0
      "0000000" when "00010000001111111", -- t[8319] = 0
      "0000000" when "00010000010000000", -- t[8320] = 0
      "0000000" when "00010000010000001", -- t[8321] = 0
      "0000000" when "00010000010000010", -- t[8322] = 0
      "0000000" when "00010000010000011", -- t[8323] = 0
      "0000000" when "00010000010000100", -- t[8324] = 0
      "0000000" when "00010000010000101", -- t[8325] = 0
      "0000000" when "00010000010000110", -- t[8326] = 0
      "0000000" when "00010000010000111", -- t[8327] = 0
      "0000000" when "00010000010001000", -- t[8328] = 0
      "0000000" when "00010000010001001", -- t[8329] = 0
      "0000000" when "00010000010001010", -- t[8330] = 0
      "0000000" when "00010000010001011", -- t[8331] = 0
      "0000000" when "00010000010001100", -- t[8332] = 0
      "0000000" when "00010000010001101", -- t[8333] = 0
      "0000000" when "00010000010001110", -- t[8334] = 0
      "0000000" when "00010000010001111", -- t[8335] = 0
      "0000000" when "00010000010010000", -- t[8336] = 0
      "0000000" when "00010000010010001", -- t[8337] = 0
      "0000000" when "00010000010010010", -- t[8338] = 0
      "0000000" when "00010000010010011", -- t[8339] = 0
      "0000000" when "00010000010010100", -- t[8340] = 0
      "0000000" when "00010000010010101", -- t[8341] = 0
      "0000000" when "00010000010010110", -- t[8342] = 0
      "0000000" when "00010000010010111", -- t[8343] = 0
      "0000000" when "00010000010011000", -- t[8344] = 0
      "0000000" when "00010000010011001", -- t[8345] = 0
      "0000000" when "00010000010011010", -- t[8346] = 0
      "0000000" when "00010000010011011", -- t[8347] = 0
      "0000000" when "00010000010011100", -- t[8348] = 0
      "0000000" when "00010000010011101", -- t[8349] = 0
      "0000000" when "00010000010011110", -- t[8350] = 0
      "0000000" when "00010000010011111", -- t[8351] = 0
      "0000000" when "00010000010100000", -- t[8352] = 0
      "0000000" when "00010000010100001", -- t[8353] = 0
      "0000000" when "00010000010100010", -- t[8354] = 0
      "0000000" when "00010000010100011", -- t[8355] = 0
      "0000000" when "00010000010100100", -- t[8356] = 0
      "0000000" when "00010000010100101", -- t[8357] = 0
      "0000000" when "00010000010100110", -- t[8358] = 0
      "0000000" when "00010000010100111", -- t[8359] = 0
      "0000000" when "00010000010101000", -- t[8360] = 0
      "0000000" when "00010000010101001", -- t[8361] = 0
      "0000000" when "00010000010101010", -- t[8362] = 0
      "0000000" when "00010000010101011", -- t[8363] = 0
      "0000000" when "00010000010101100", -- t[8364] = 0
      "0000000" when "00010000010101101", -- t[8365] = 0
      "0000000" when "00010000010101110", -- t[8366] = 0
      "0000000" when "00010000010101111", -- t[8367] = 0
      "0000000" when "00010000010110000", -- t[8368] = 0
      "0000000" when "00010000010110001", -- t[8369] = 0
      "0000000" when "00010000010110010", -- t[8370] = 0
      "0000000" when "00010000010110011", -- t[8371] = 0
      "0000000" when "00010000010110100", -- t[8372] = 0
      "0000000" when "00010000010110101", -- t[8373] = 0
      "0000000" when "00010000010110110", -- t[8374] = 0
      "0000000" when "00010000010110111", -- t[8375] = 0
      "0000000" when "00010000010111000", -- t[8376] = 0
      "0000000" when "00010000010111001", -- t[8377] = 0
      "0000000" when "00010000010111010", -- t[8378] = 0
      "0000000" when "00010000010111011", -- t[8379] = 0
      "0000000" when "00010000010111100", -- t[8380] = 0
      "0000000" when "00010000010111101", -- t[8381] = 0
      "0000000" when "00010000010111110", -- t[8382] = 0
      "0000000" when "00010000010111111", -- t[8383] = 0
      "0000000" when "00010000011000000", -- t[8384] = 0
      "0000000" when "00010000011000001", -- t[8385] = 0
      "0000000" when "00010000011000010", -- t[8386] = 0
      "0000000" when "00010000011000011", -- t[8387] = 0
      "0000000" when "00010000011000100", -- t[8388] = 0
      "0000000" when "00010000011000101", -- t[8389] = 0
      "0000000" when "00010000011000110", -- t[8390] = 0
      "0000000" when "00010000011000111", -- t[8391] = 0
      "0000000" when "00010000011001000", -- t[8392] = 0
      "0000000" when "00010000011001001", -- t[8393] = 0
      "0000000" when "00010000011001010", -- t[8394] = 0
      "0000000" when "00010000011001011", -- t[8395] = 0
      "0000000" when "00010000011001100", -- t[8396] = 0
      "0000000" when "00010000011001101", -- t[8397] = 0
      "0000000" when "00010000011001110", -- t[8398] = 0
      "0000000" when "00010000011001111", -- t[8399] = 0
      "0000000" when "00010000011010000", -- t[8400] = 0
      "0000000" when "00010000011010001", -- t[8401] = 0
      "0000000" when "00010000011010010", -- t[8402] = 0
      "0000000" when "00010000011010011", -- t[8403] = 0
      "0000000" when "00010000011010100", -- t[8404] = 0
      "0000000" when "00010000011010101", -- t[8405] = 0
      "0000000" when "00010000011010110", -- t[8406] = 0
      "0000000" when "00010000011010111", -- t[8407] = 0
      "0000000" when "00010000011011000", -- t[8408] = 0
      "0000000" when "00010000011011001", -- t[8409] = 0
      "0000000" when "00010000011011010", -- t[8410] = 0
      "0000000" when "00010000011011011", -- t[8411] = 0
      "0000000" when "00010000011011100", -- t[8412] = 0
      "0000000" when "00010000011011101", -- t[8413] = 0
      "0000000" when "00010000011011110", -- t[8414] = 0
      "0000000" when "00010000011011111", -- t[8415] = 0
      "0000000" when "00010000011100000", -- t[8416] = 0
      "0000000" when "00010000011100001", -- t[8417] = 0
      "0000000" when "00010000011100010", -- t[8418] = 0
      "0000000" when "00010000011100011", -- t[8419] = 0
      "0000000" when "00010000011100100", -- t[8420] = 0
      "0000000" when "00010000011100101", -- t[8421] = 0
      "0000000" when "00010000011100110", -- t[8422] = 0
      "0000000" when "00010000011100111", -- t[8423] = 0
      "0000000" when "00010000011101000", -- t[8424] = 0
      "0000000" when "00010000011101001", -- t[8425] = 0
      "0000000" when "00010000011101010", -- t[8426] = 0
      "0000000" when "00010000011101011", -- t[8427] = 0
      "0000000" when "00010000011101100", -- t[8428] = 0
      "0000000" when "00010000011101101", -- t[8429] = 0
      "0000000" when "00010000011101110", -- t[8430] = 0
      "0000000" when "00010000011101111", -- t[8431] = 0
      "0000000" when "00010000011110000", -- t[8432] = 0
      "0000000" when "00010000011110001", -- t[8433] = 0
      "0000000" when "00010000011110010", -- t[8434] = 0
      "0000000" when "00010000011110011", -- t[8435] = 0
      "0000000" when "00010000011110100", -- t[8436] = 0
      "0000000" when "00010000011110101", -- t[8437] = 0
      "0000000" when "00010000011110110", -- t[8438] = 0
      "0000000" when "00010000011110111", -- t[8439] = 0
      "0000000" when "00010000011111000", -- t[8440] = 0
      "0000000" when "00010000011111001", -- t[8441] = 0
      "0000000" when "00010000011111010", -- t[8442] = 0
      "0000000" when "00010000011111011", -- t[8443] = 0
      "0000000" when "00010000011111100", -- t[8444] = 0
      "0000000" when "00010000011111101", -- t[8445] = 0
      "0000000" when "00010000011111110", -- t[8446] = 0
      "0000000" when "00010000011111111", -- t[8447] = 0
      "0000000" when "00010000100000000", -- t[8448] = 0
      "0000000" when "00010000100000001", -- t[8449] = 0
      "0000000" when "00010000100000010", -- t[8450] = 0
      "0000000" when "00010000100000011", -- t[8451] = 0
      "0000000" when "00010000100000100", -- t[8452] = 0
      "0000000" when "00010000100000101", -- t[8453] = 0
      "0000000" when "00010000100000110", -- t[8454] = 0
      "0000000" when "00010000100000111", -- t[8455] = 0
      "0000000" when "00010000100001000", -- t[8456] = 0
      "0000000" when "00010000100001001", -- t[8457] = 0
      "0000000" when "00010000100001010", -- t[8458] = 0
      "0000000" when "00010000100001011", -- t[8459] = 0
      "0000000" when "00010000100001100", -- t[8460] = 0
      "0000000" when "00010000100001101", -- t[8461] = 0
      "0000000" when "00010000100001110", -- t[8462] = 0
      "0000000" when "00010000100001111", -- t[8463] = 0
      "0000000" when "00010000100010000", -- t[8464] = 0
      "0000000" when "00010000100010001", -- t[8465] = 0
      "0000000" when "00010000100010010", -- t[8466] = 0
      "0000000" when "00010000100010011", -- t[8467] = 0
      "0000000" when "00010000100010100", -- t[8468] = 0
      "0000000" when "00010000100010101", -- t[8469] = 0
      "0000000" when "00010000100010110", -- t[8470] = 0
      "0000000" when "00010000100010111", -- t[8471] = 0
      "0000000" when "00010000100011000", -- t[8472] = 0
      "0000000" when "00010000100011001", -- t[8473] = 0
      "0000000" when "00010000100011010", -- t[8474] = 0
      "0000000" when "00010000100011011", -- t[8475] = 0
      "0000000" when "00010000100011100", -- t[8476] = 0
      "0000000" when "00010000100011101", -- t[8477] = 0
      "0000000" when "00010000100011110", -- t[8478] = 0
      "0000000" when "00010000100011111", -- t[8479] = 0
      "0000000" when "00010000100100000", -- t[8480] = 0
      "0000000" when "00010000100100001", -- t[8481] = 0
      "0000000" when "00010000100100010", -- t[8482] = 0
      "0000000" when "00010000100100011", -- t[8483] = 0
      "0000000" when "00010000100100100", -- t[8484] = 0
      "0000000" when "00010000100100101", -- t[8485] = 0
      "0000000" when "00010000100100110", -- t[8486] = 0
      "0000000" when "00010000100100111", -- t[8487] = 0
      "0000000" when "00010000100101000", -- t[8488] = 0
      "0000000" when "00010000100101001", -- t[8489] = 0
      "0000000" when "00010000100101010", -- t[8490] = 0
      "0000000" when "00010000100101011", -- t[8491] = 0
      "0000000" when "00010000100101100", -- t[8492] = 0
      "0000000" when "00010000100101101", -- t[8493] = 0
      "0000000" when "00010000100101110", -- t[8494] = 0
      "0000000" when "00010000100101111", -- t[8495] = 0
      "0000000" when "00010000100110000", -- t[8496] = 0
      "0000000" when "00010000100110001", -- t[8497] = 0
      "0000000" when "00010000100110010", -- t[8498] = 0
      "0000000" when "00010000100110011", -- t[8499] = 0
      "0000000" when "00010000100110100", -- t[8500] = 0
      "0000000" when "00010000100110101", -- t[8501] = 0
      "0000000" when "00010000100110110", -- t[8502] = 0
      "0000000" when "00010000100110111", -- t[8503] = 0
      "0000000" when "00010000100111000", -- t[8504] = 0
      "0000000" when "00010000100111001", -- t[8505] = 0
      "0000000" when "00010000100111010", -- t[8506] = 0
      "0000000" when "00010000100111011", -- t[8507] = 0
      "0000000" when "00010000100111100", -- t[8508] = 0
      "0000000" when "00010000100111101", -- t[8509] = 0
      "0000000" when "00010000100111110", -- t[8510] = 0
      "0000000" when "00010000100111111", -- t[8511] = 0
      "0000000" when "00010000101000000", -- t[8512] = 0
      "0000000" when "00010000101000001", -- t[8513] = 0
      "0000000" when "00010000101000010", -- t[8514] = 0
      "0000000" when "00010000101000011", -- t[8515] = 0
      "0000000" when "00010000101000100", -- t[8516] = 0
      "0000000" when "00010000101000101", -- t[8517] = 0
      "0000000" when "00010000101000110", -- t[8518] = 0
      "0000000" when "00010000101000111", -- t[8519] = 0
      "0000000" when "00010000101001000", -- t[8520] = 0
      "0000000" when "00010000101001001", -- t[8521] = 0
      "0000000" when "00010000101001010", -- t[8522] = 0
      "0000000" when "00010000101001011", -- t[8523] = 0
      "0000000" when "00010000101001100", -- t[8524] = 0
      "0000000" when "00010000101001101", -- t[8525] = 0
      "0000000" when "00010000101001110", -- t[8526] = 0
      "0000000" when "00010000101001111", -- t[8527] = 0
      "0000000" when "00010000101010000", -- t[8528] = 0
      "0000000" when "00010000101010001", -- t[8529] = 0
      "0000000" when "00010000101010010", -- t[8530] = 0
      "0000000" when "00010000101010011", -- t[8531] = 0
      "0000000" when "00010000101010100", -- t[8532] = 0
      "0000000" when "00010000101010101", -- t[8533] = 0
      "0000000" when "00010000101010110", -- t[8534] = 0
      "0000000" when "00010000101010111", -- t[8535] = 0
      "0000000" when "00010000101011000", -- t[8536] = 0
      "0000000" when "00010000101011001", -- t[8537] = 0
      "0000000" when "00010000101011010", -- t[8538] = 0
      "0000000" when "00010000101011011", -- t[8539] = 0
      "0000000" when "00010000101011100", -- t[8540] = 0
      "0000000" when "00010000101011101", -- t[8541] = 0
      "0000000" when "00010000101011110", -- t[8542] = 0
      "0000000" when "00010000101011111", -- t[8543] = 0
      "0000000" when "00010000101100000", -- t[8544] = 0
      "0000000" when "00010000101100001", -- t[8545] = 0
      "0000000" when "00010000101100010", -- t[8546] = 0
      "0000000" when "00010000101100011", -- t[8547] = 0
      "0000000" when "00010000101100100", -- t[8548] = 0
      "0000000" when "00010000101100101", -- t[8549] = 0
      "0000000" when "00010000101100110", -- t[8550] = 0
      "0000000" when "00010000101100111", -- t[8551] = 0
      "0000000" when "00010000101101000", -- t[8552] = 0
      "0000000" when "00010000101101001", -- t[8553] = 0
      "0000000" when "00010000101101010", -- t[8554] = 0
      "0000000" when "00010000101101011", -- t[8555] = 0
      "0000000" when "00010000101101100", -- t[8556] = 0
      "0000000" when "00010000101101101", -- t[8557] = 0
      "0000000" when "00010000101101110", -- t[8558] = 0
      "0000000" when "00010000101101111", -- t[8559] = 0
      "0000000" when "00010000101110000", -- t[8560] = 0
      "0000000" when "00010000101110001", -- t[8561] = 0
      "0000000" when "00010000101110010", -- t[8562] = 0
      "0000000" when "00010000101110011", -- t[8563] = 0
      "0000000" when "00010000101110100", -- t[8564] = 0
      "0000000" when "00010000101110101", -- t[8565] = 0
      "0000000" when "00010000101110110", -- t[8566] = 0
      "0000000" when "00010000101110111", -- t[8567] = 0
      "0000000" when "00010000101111000", -- t[8568] = 0
      "0000000" when "00010000101111001", -- t[8569] = 0
      "0000000" when "00010000101111010", -- t[8570] = 0
      "0000000" when "00010000101111011", -- t[8571] = 0
      "0000000" when "00010000101111100", -- t[8572] = 0
      "0000000" when "00010000101111101", -- t[8573] = 0
      "0000000" when "00010000101111110", -- t[8574] = 0
      "0000000" when "00010000101111111", -- t[8575] = 0
      "0000000" when "00010000110000000", -- t[8576] = 0
      "0000000" when "00010000110000001", -- t[8577] = 0
      "0000000" when "00010000110000010", -- t[8578] = 0
      "0000000" when "00010000110000011", -- t[8579] = 0
      "0000000" when "00010000110000100", -- t[8580] = 0
      "0000000" when "00010000110000101", -- t[8581] = 0
      "0000000" when "00010000110000110", -- t[8582] = 0
      "0000000" when "00010000110000111", -- t[8583] = 0
      "0000000" when "00010000110001000", -- t[8584] = 0
      "0000000" when "00010000110001001", -- t[8585] = 0
      "0000000" when "00010000110001010", -- t[8586] = 0
      "0000000" when "00010000110001011", -- t[8587] = 0
      "0000000" when "00010000110001100", -- t[8588] = 0
      "0000000" when "00010000110001101", -- t[8589] = 0
      "0000000" when "00010000110001110", -- t[8590] = 0
      "0000000" when "00010000110001111", -- t[8591] = 0
      "0000000" when "00010000110010000", -- t[8592] = 0
      "0000000" when "00010000110010001", -- t[8593] = 0
      "0000000" when "00010000110010010", -- t[8594] = 0
      "0000000" when "00010000110010011", -- t[8595] = 0
      "0000000" when "00010000110010100", -- t[8596] = 0
      "0000000" when "00010000110010101", -- t[8597] = 0
      "0000000" when "00010000110010110", -- t[8598] = 0
      "0000000" when "00010000110010111", -- t[8599] = 0
      "0000000" when "00010000110011000", -- t[8600] = 0
      "0000000" when "00010000110011001", -- t[8601] = 0
      "0000000" when "00010000110011010", -- t[8602] = 0
      "0000000" when "00010000110011011", -- t[8603] = 0
      "0000000" when "00010000110011100", -- t[8604] = 0
      "0000000" when "00010000110011101", -- t[8605] = 0
      "0000000" when "00010000110011110", -- t[8606] = 0
      "0000000" when "00010000110011111", -- t[8607] = 0
      "0000000" when "00010000110100000", -- t[8608] = 0
      "0000000" when "00010000110100001", -- t[8609] = 0
      "0000000" when "00010000110100010", -- t[8610] = 0
      "0000000" when "00010000110100011", -- t[8611] = 0
      "0000000" when "00010000110100100", -- t[8612] = 0
      "0000000" when "00010000110100101", -- t[8613] = 0
      "0000000" when "00010000110100110", -- t[8614] = 0
      "0000000" when "00010000110100111", -- t[8615] = 0
      "0000000" when "00010000110101000", -- t[8616] = 0
      "0000000" when "00010000110101001", -- t[8617] = 0
      "0000000" when "00010000110101010", -- t[8618] = 0
      "0000000" when "00010000110101011", -- t[8619] = 0
      "0000000" when "00010000110101100", -- t[8620] = 0
      "0000000" when "00010000110101101", -- t[8621] = 0
      "0000000" when "00010000110101110", -- t[8622] = 0
      "0000000" when "00010000110101111", -- t[8623] = 0
      "0000000" when "00010000110110000", -- t[8624] = 0
      "0000000" when "00010000110110001", -- t[8625] = 0
      "0000000" when "00010000110110010", -- t[8626] = 0
      "0000000" when "00010000110110011", -- t[8627] = 0
      "0000000" when "00010000110110100", -- t[8628] = 0
      "0000000" when "00010000110110101", -- t[8629] = 0
      "0000000" when "00010000110110110", -- t[8630] = 0
      "0000000" when "00010000110110111", -- t[8631] = 0
      "0000000" when "00010000110111000", -- t[8632] = 0
      "0000000" when "00010000110111001", -- t[8633] = 0
      "0000000" when "00010000110111010", -- t[8634] = 0
      "0000000" when "00010000110111011", -- t[8635] = 0
      "0000000" when "00010000110111100", -- t[8636] = 0
      "0000000" when "00010000110111101", -- t[8637] = 0
      "0000000" when "00010000110111110", -- t[8638] = 0
      "0000000" when "00010000110111111", -- t[8639] = 0
      "0000000" when "00010000111000000", -- t[8640] = 0
      "0000000" when "00010000111000001", -- t[8641] = 0
      "0000000" when "00010000111000010", -- t[8642] = 0
      "0000000" when "00010000111000011", -- t[8643] = 0
      "0000000" when "00010000111000100", -- t[8644] = 0
      "0000000" when "00010000111000101", -- t[8645] = 0
      "0000000" when "00010000111000110", -- t[8646] = 0
      "0000000" when "00010000111000111", -- t[8647] = 0
      "0000000" when "00010000111001000", -- t[8648] = 0
      "0000000" when "00010000111001001", -- t[8649] = 0
      "0000000" when "00010000111001010", -- t[8650] = 0
      "0000000" when "00010000111001011", -- t[8651] = 0
      "0000000" when "00010000111001100", -- t[8652] = 0
      "0000000" when "00010000111001101", -- t[8653] = 0
      "0000000" when "00010000111001110", -- t[8654] = 0
      "0000000" when "00010000111001111", -- t[8655] = 0
      "0000000" when "00010000111010000", -- t[8656] = 0
      "0000000" when "00010000111010001", -- t[8657] = 0
      "0000000" when "00010000111010010", -- t[8658] = 0
      "0000000" when "00010000111010011", -- t[8659] = 0
      "0000000" when "00010000111010100", -- t[8660] = 0
      "0000000" when "00010000111010101", -- t[8661] = 0
      "0000000" when "00010000111010110", -- t[8662] = 0
      "0000000" when "00010000111010111", -- t[8663] = 0
      "0000000" when "00010000111011000", -- t[8664] = 0
      "0000000" when "00010000111011001", -- t[8665] = 0
      "0000000" when "00010000111011010", -- t[8666] = 0
      "0000000" when "00010000111011011", -- t[8667] = 0
      "0000000" when "00010000111011100", -- t[8668] = 0
      "0000000" when "00010000111011101", -- t[8669] = 0
      "0000000" when "00010000111011110", -- t[8670] = 0
      "0000000" when "00010000111011111", -- t[8671] = 0
      "0000000" when "00010000111100000", -- t[8672] = 0
      "0000000" when "00010000111100001", -- t[8673] = 0
      "0000000" when "00010000111100010", -- t[8674] = 0
      "0000000" when "00010000111100011", -- t[8675] = 0
      "0000000" when "00010000111100100", -- t[8676] = 0
      "0000000" when "00010000111100101", -- t[8677] = 0
      "0000000" when "00010000111100110", -- t[8678] = 0
      "0000000" when "00010000111100111", -- t[8679] = 0
      "0000000" when "00010000111101000", -- t[8680] = 0
      "0000000" when "00010000111101001", -- t[8681] = 0
      "0000000" when "00010000111101010", -- t[8682] = 0
      "0000000" when "00010000111101011", -- t[8683] = 0
      "0000000" when "00010000111101100", -- t[8684] = 0
      "0000000" when "00010000111101101", -- t[8685] = 0
      "0000000" when "00010000111101110", -- t[8686] = 0
      "0000000" when "00010000111101111", -- t[8687] = 0
      "0000000" when "00010000111110000", -- t[8688] = 0
      "0000000" when "00010000111110001", -- t[8689] = 0
      "0000000" when "00010000111110010", -- t[8690] = 0
      "0000000" when "00010000111110011", -- t[8691] = 0
      "0000000" when "00010000111110100", -- t[8692] = 0
      "0000000" when "00010000111110101", -- t[8693] = 0
      "0000000" when "00010000111110110", -- t[8694] = 0
      "0000000" when "00010000111110111", -- t[8695] = 0
      "0000000" when "00010000111111000", -- t[8696] = 0
      "0000000" when "00010000111111001", -- t[8697] = 0
      "0000000" when "00010000111111010", -- t[8698] = 0
      "0000000" when "00010000111111011", -- t[8699] = 0
      "0000000" when "00010000111111100", -- t[8700] = 0
      "0000000" when "00010000111111101", -- t[8701] = 0
      "0000000" when "00010000111111110", -- t[8702] = 0
      "0000000" when "00010000111111111", -- t[8703] = 0
      "0000000" when "00010001000000000", -- t[8704] = 0
      "0000000" when "00010001000000001", -- t[8705] = 0
      "0000000" when "00010001000000010", -- t[8706] = 0
      "0000000" when "00010001000000011", -- t[8707] = 0
      "0000000" when "00010001000000100", -- t[8708] = 0
      "0000000" when "00010001000000101", -- t[8709] = 0
      "0000000" when "00010001000000110", -- t[8710] = 0
      "0000000" when "00010001000000111", -- t[8711] = 0
      "0000000" when "00010001000001000", -- t[8712] = 0
      "0000000" when "00010001000001001", -- t[8713] = 0
      "0000000" when "00010001000001010", -- t[8714] = 0
      "0000000" when "00010001000001011", -- t[8715] = 0
      "0000000" when "00010001000001100", -- t[8716] = 0
      "0000000" when "00010001000001101", -- t[8717] = 0
      "0000000" when "00010001000001110", -- t[8718] = 0
      "0000000" when "00010001000001111", -- t[8719] = 0
      "0000000" when "00010001000010000", -- t[8720] = 0
      "0000000" when "00010001000010001", -- t[8721] = 0
      "0000000" when "00010001000010010", -- t[8722] = 0
      "0000000" when "00010001000010011", -- t[8723] = 0
      "0000000" when "00010001000010100", -- t[8724] = 0
      "0000000" when "00010001000010101", -- t[8725] = 0
      "0000000" when "00010001000010110", -- t[8726] = 0
      "0000000" when "00010001000010111", -- t[8727] = 0
      "0000000" when "00010001000011000", -- t[8728] = 0
      "0000000" when "00010001000011001", -- t[8729] = 0
      "0000000" when "00010001000011010", -- t[8730] = 0
      "0000000" when "00010001000011011", -- t[8731] = 0
      "0000000" when "00010001000011100", -- t[8732] = 0
      "0000000" when "00010001000011101", -- t[8733] = 0
      "0000000" when "00010001000011110", -- t[8734] = 0
      "0000000" when "00010001000011111", -- t[8735] = 0
      "0000000" when "00010001000100000", -- t[8736] = 0
      "0000000" when "00010001000100001", -- t[8737] = 0
      "0000000" when "00010001000100010", -- t[8738] = 0
      "0000000" when "00010001000100011", -- t[8739] = 0
      "0000000" when "00010001000100100", -- t[8740] = 0
      "0000000" when "00010001000100101", -- t[8741] = 0
      "0000000" when "00010001000100110", -- t[8742] = 0
      "0000000" when "00010001000100111", -- t[8743] = 0
      "0000000" when "00010001000101000", -- t[8744] = 0
      "0000000" when "00010001000101001", -- t[8745] = 0
      "0000000" when "00010001000101010", -- t[8746] = 0
      "0000000" when "00010001000101011", -- t[8747] = 0
      "0000000" when "00010001000101100", -- t[8748] = 0
      "0000000" when "00010001000101101", -- t[8749] = 0
      "0000000" when "00010001000101110", -- t[8750] = 0
      "0000000" when "00010001000101111", -- t[8751] = 0
      "0000000" when "00010001000110000", -- t[8752] = 0
      "0000000" when "00010001000110001", -- t[8753] = 0
      "0000000" when "00010001000110010", -- t[8754] = 0
      "0000000" when "00010001000110011", -- t[8755] = 0
      "0000000" when "00010001000110100", -- t[8756] = 0
      "0000000" when "00010001000110101", -- t[8757] = 0
      "0000000" when "00010001000110110", -- t[8758] = 0
      "0000000" when "00010001000110111", -- t[8759] = 0
      "0000000" when "00010001000111000", -- t[8760] = 0
      "0000000" when "00010001000111001", -- t[8761] = 0
      "0000000" when "00010001000111010", -- t[8762] = 0
      "0000000" when "00010001000111011", -- t[8763] = 0
      "0000000" when "00010001000111100", -- t[8764] = 0
      "0000000" when "00010001000111101", -- t[8765] = 0
      "0000000" when "00010001000111110", -- t[8766] = 0
      "0000000" when "00010001000111111", -- t[8767] = 0
      "0000000" when "00010001001000000", -- t[8768] = 0
      "0000000" when "00010001001000001", -- t[8769] = 0
      "0000000" when "00010001001000010", -- t[8770] = 0
      "0000000" when "00010001001000011", -- t[8771] = 0
      "0000000" when "00010001001000100", -- t[8772] = 0
      "0000000" when "00010001001000101", -- t[8773] = 0
      "0000000" when "00010001001000110", -- t[8774] = 0
      "0000000" when "00010001001000111", -- t[8775] = 0
      "0000000" when "00010001001001000", -- t[8776] = 0
      "0000000" when "00010001001001001", -- t[8777] = 0
      "0000000" when "00010001001001010", -- t[8778] = 0
      "0000000" when "00010001001001011", -- t[8779] = 0
      "0000000" when "00010001001001100", -- t[8780] = 0
      "0000000" when "00010001001001101", -- t[8781] = 0
      "0000000" when "00010001001001110", -- t[8782] = 0
      "0000000" when "00010001001001111", -- t[8783] = 0
      "0000000" when "00010001001010000", -- t[8784] = 0
      "0000000" when "00010001001010001", -- t[8785] = 0
      "0000000" when "00010001001010010", -- t[8786] = 0
      "0000000" when "00010001001010011", -- t[8787] = 0
      "0000000" when "00010001001010100", -- t[8788] = 0
      "0000000" when "00010001001010101", -- t[8789] = 0
      "0000000" when "00010001001010110", -- t[8790] = 0
      "0000000" when "00010001001010111", -- t[8791] = 0
      "0000000" when "00010001001011000", -- t[8792] = 0
      "0000000" when "00010001001011001", -- t[8793] = 0
      "0000000" when "00010001001011010", -- t[8794] = 0
      "0000000" when "00010001001011011", -- t[8795] = 0
      "0000000" when "00010001001011100", -- t[8796] = 0
      "0000000" when "00010001001011101", -- t[8797] = 0
      "0000000" when "00010001001011110", -- t[8798] = 0
      "0000000" when "00010001001011111", -- t[8799] = 0
      "0000000" when "00010001001100000", -- t[8800] = 0
      "0000000" when "00010001001100001", -- t[8801] = 0
      "0000000" when "00010001001100010", -- t[8802] = 0
      "0000000" when "00010001001100011", -- t[8803] = 0
      "0000000" when "00010001001100100", -- t[8804] = 0
      "0000000" when "00010001001100101", -- t[8805] = 0
      "0000000" when "00010001001100110", -- t[8806] = 0
      "0000000" when "00010001001100111", -- t[8807] = 0
      "0000000" when "00010001001101000", -- t[8808] = 0
      "0000000" when "00010001001101001", -- t[8809] = 0
      "0000000" when "00010001001101010", -- t[8810] = 0
      "0000000" when "00010001001101011", -- t[8811] = 0
      "0000000" when "00010001001101100", -- t[8812] = 0
      "0000000" when "00010001001101101", -- t[8813] = 0
      "0000000" when "00010001001101110", -- t[8814] = 0
      "0000000" when "00010001001101111", -- t[8815] = 0
      "0000000" when "00010001001110000", -- t[8816] = 0
      "0000000" when "00010001001110001", -- t[8817] = 0
      "0000000" when "00010001001110010", -- t[8818] = 0
      "0000000" when "00010001001110011", -- t[8819] = 0
      "0000000" when "00010001001110100", -- t[8820] = 0
      "0000000" when "00010001001110101", -- t[8821] = 0
      "0000000" when "00010001001110110", -- t[8822] = 0
      "0000000" when "00010001001110111", -- t[8823] = 0
      "0000000" when "00010001001111000", -- t[8824] = 0
      "0000000" when "00010001001111001", -- t[8825] = 0
      "0000000" when "00010001001111010", -- t[8826] = 0
      "0000000" when "00010001001111011", -- t[8827] = 0
      "0000000" when "00010001001111100", -- t[8828] = 0
      "0000000" when "00010001001111101", -- t[8829] = 0
      "0000000" when "00010001001111110", -- t[8830] = 0
      "0000000" when "00010001001111111", -- t[8831] = 0
      "0000000" when "00010001010000000", -- t[8832] = 0
      "0000000" when "00010001010000001", -- t[8833] = 0
      "0000000" when "00010001010000010", -- t[8834] = 0
      "0000000" when "00010001010000011", -- t[8835] = 0
      "0000000" when "00010001010000100", -- t[8836] = 0
      "0000000" when "00010001010000101", -- t[8837] = 0
      "0000000" when "00010001010000110", -- t[8838] = 0
      "0000000" when "00010001010000111", -- t[8839] = 0
      "0000000" when "00010001010001000", -- t[8840] = 0
      "0000000" when "00010001010001001", -- t[8841] = 0
      "0000000" when "00010001010001010", -- t[8842] = 0
      "0000000" when "00010001010001011", -- t[8843] = 0
      "0000000" when "00010001010001100", -- t[8844] = 0
      "0000000" when "00010001010001101", -- t[8845] = 0
      "0000000" when "00010001010001110", -- t[8846] = 0
      "0000000" when "00010001010001111", -- t[8847] = 0
      "0000000" when "00010001010010000", -- t[8848] = 0
      "0000000" when "00010001010010001", -- t[8849] = 0
      "0000000" when "00010001010010010", -- t[8850] = 0
      "0000000" when "00010001010010011", -- t[8851] = 0
      "0000000" when "00010001010010100", -- t[8852] = 0
      "0000000" when "00010001010010101", -- t[8853] = 0
      "0000000" when "00010001010010110", -- t[8854] = 0
      "0000000" when "00010001010010111", -- t[8855] = 0
      "0000000" when "00010001010011000", -- t[8856] = 0
      "0000000" when "00010001010011001", -- t[8857] = 0
      "0000000" when "00010001010011010", -- t[8858] = 0
      "0000000" when "00010001010011011", -- t[8859] = 0
      "0000000" when "00010001010011100", -- t[8860] = 0
      "0000000" when "00010001010011101", -- t[8861] = 0
      "0000000" when "00010001010011110", -- t[8862] = 0
      "0000000" when "00010001010011111", -- t[8863] = 0
      "0000000" when "00010001010100000", -- t[8864] = 0
      "0000000" when "00010001010100001", -- t[8865] = 0
      "0000000" when "00010001010100010", -- t[8866] = 0
      "0000000" when "00010001010100011", -- t[8867] = 0
      "0000000" when "00010001010100100", -- t[8868] = 0
      "0000000" when "00010001010100101", -- t[8869] = 0
      "0000000" when "00010001010100110", -- t[8870] = 0
      "0000000" when "00010001010100111", -- t[8871] = 0
      "0000000" when "00010001010101000", -- t[8872] = 0
      "0000000" when "00010001010101001", -- t[8873] = 0
      "0000000" when "00010001010101010", -- t[8874] = 0
      "0000000" when "00010001010101011", -- t[8875] = 0
      "0000000" when "00010001010101100", -- t[8876] = 0
      "0000000" when "00010001010101101", -- t[8877] = 0
      "0000000" when "00010001010101110", -- t[8878] = 0
      "0000000" when "00010001010101111", -- t[8879] = 0
      "0000000" when "00010001010110000", -- t[8880] = 0
      "0000000" when "00010001010110001", -- t[8881] = 0
      "0000000" when "00010001010110010", -- t[8882] = 0
      "0000000" when "00010001010110011", -- t[8883] = 0
      "0000000" when "00010001010110100", -- t[8884] = 0
      "0000000" when "00010001010110101", -- t[8885] = 0
      "0000000" when "00010001010110110", -- t[8886] = 0
      "0000000" when "00010001010110111", -- t[8887] = 0
      "0000000" when "00010001010111000", -- t[8888] = 0
      "0000000" when "00010001010111001", -- t[8889] = 0
      "0000000" when "00010001010111010", -- t[8890] = 0
      "0000000" when "00010001010111011", -- t[8891] = 0
      "0000000" when "00010001010111100", -- t[8892] = 0
      "0000000" when "00010001010111101", -- t[8893] = 0
      "0000000" when "00010001010111110", -- t[8894] = 0
      "0000000" when "00010001010111111", -- t[8895] = 0
      "0000000" when "00010001011000000", -- t[8896] = 0
      "0000000" when "00010001011000001", -- t[8897] = 0
      "0000000" when "00010001011000010", -- t[8898] = 0
      "0000000" when "00010001011000011", -- t[8899] = 0
      "0000000" when "00010001011000100", -- t[8900] = 0
      "0000000" when "00010001011000101", -- t[8901] = 0
      "0000000" when "00010001011000110", -- t[8902] = 0
      "0000000" when "00010001011000111", -- t[8903] = 0
      "0000000" when "00010001011001000", -- t[8904] = 0
      "0000000" when "00010001011001001", -- t[8905] = 0
      "0000000" when "00010001011001010", -- t[8906] = 0
      "0000000" when "00010001011001011", -- t[8907] = 0
      "0000000" when "00010001011001100", -- t[8908] = 0
      "0000000" when "00010001011001101", -- t[8909] = 0
      "0000000" when "00010001011001110", -- t[8910] = 0
      "0000000" when "00010001011001111", -- t[8911] = 0
      "0000000" when "00010001011010000", -- t[8912] = 0
      "0000000" when "00010001011010001", -- t[8913] = 0
      "0000000" when "00010001011010010", -- t[8914] = 0
      "0000000" when "00010001011010011", -- t[8915] = 0
      "0000000" when "00010001011010100", -- t[8916] = 0
      "0000000" when "00010001011010101", -- t[8917] = 0
      "0000000" when "00010001011010110", -- t[8918] = 0
      "0000000" when "00010001011010111", -- t[8919] = 0
      "0000000" when "00010001011011000", -- t[8920] = 0
      "0000000" when "00010001011011001", -- t[8921] = 0
      "0000000" when "00010001011011010", -- t[8922] = 0
      "0000000" when "00010001011011011", -- t[8923] = 0
      "0000000" when "00010001011011100", -- t[8924] = 0
      "0000000" when "00010001011011101", -- t[8925] = 0
      "0000000" when "00010001011011110", -- t[8926] = 0
      "0000000" when "00010001011011111", -- t[8927] = 0
      "0000000" when "00010001011100000", -- t[8928] = 0
      "0000000" when "00010001011100001", -- t[8929] = 0
      "0000000" when "00010001011100010", -- t[8930] = 0
      "0000000" when "00010001011100011", -- t[8931] = 0
      "0000000" when "00010001011100100", -- t[8932] = 0
      "0000000" when "00010001011100101", -- t[8933] = 0
      "0000000" when "00010001011100110", -- t[8934] = 0
      "0000000" when "00010001011100111", -- t[8935] = 0
      "0000000" when "00010001011101000", -- t[8936] = 0
      "0000000" when "00010001011101001", -- t[8937] = 0
      "0000000" when "00010001011101010", -- t[8938] = 0
      "0000000" when "00010001011101011", -- t[8939] = 0
      "0000000" when "00010001011101100", -- t[8940] = 0
      "0000000" when "00010001011101101", -- t[8941] = 0
      "0000000" when "00010001011101110", -- t[8942] = 0
      "0000000" when "00010001011101111", -- t[8943] = 0
      "0000000" when "00010001011110000", -- t[8944] = 0
      "0000000" when "00010001011110001", -- t[8945] = 0
      "0000000" when "00010001011110010", -- t[8946] = 0
      "0000000" when "00010001011110011", -- t[8947] = 0
      "0000000" when "00010001011110100", -- t[8948] = 0
      "0000000" when "00010001011110101", -- t[8949] = 0
      "0000000" when "00010001011110110", -- t[8950] = 0
      "0000000" when "00010001011110111", -- t[8951] = 0
      "0000000" when "00010001011111000", -- t[8952] = 0
      "0000000" when "00010001011111001", -- t[8953] = 0
      "0000000" when "00010001011111010", -- t[8954] = 0
      "0000000" when "00010001011111011", -- t[8955] = 0
      "0000000" when "00010001011111100", -- t[8956] = 0
      "0000000" when "00010001011111101", -- t[8957] = 0
      "0000000" when "00010001011111110", -- t[8958] = 0
      "0000000" when "00010001011111111", -- t[8959] = 0
      "0000000" when "00010001100000000", -- t[8960] = 0
      "0000000" when "00010001100000001", -- t[8961] = 0
      "0000000" when "00010001100000010", -- t[8962] = 0
      "0000000" when "00010001100000011", -- t[8963] = 0
      "0000000" when "00010001100000100", -- t[8964] = 0
      "0000000" when "00010001100000101", -- t[8965] = 0
      "0000000" when "00010001100000110", -- t[8966] = 0
      "0000000" when "00010001100000111", -- t[8967] = 0
      "0000000" when "00010001100001000", -- t[8968] = 0
      "0000000" when "00010001100001001", -- t[8969] = 0
      "0000000" when "00010001100001010", -- t[8970] = 0
      "0000000" when "00010001100001011", -- t[8971] = 0
      "0000000" when "00010001100001100", -- t[8972] = 0
      "0000000" when "00010001100001101", -- t[8973] = 0
      "0000000" when "00010001100001110", -- t[8974] = 0
      "0000000" when "00010001100001111", -- t[8975] = 0
      "0000000" when "00010001100010000", -- t[8976] = 0
      "0000000" when "00010001100010001", -- t[8977] = 0
      "0000000" when "00010001100010010", -- t[8978] = 0
      "0000000" when "00010001100010011", -- t[8979] = 0
      "0000000" when "00010001100010100", -- t[8980] = 0
      "0000000" when "00010001100010101", -- t[8981] = 0
      "0000000" when "00010001100010110", -- t[8982] = 0
      "0000000" when "00010001100010111", -- t[8983] = 0
      "0000000" when "00010001100011000", -- t[8984] = 0
      "0000000" when "00010001100011001", -- t[8985] = 0
      "0000000" when "00010001100011010", -- t[8986] = 0
      "0000000" when "00010001100011011", -- t[8987] = 0
      "0000000" when "00010001100011100", -- t[8988] = 0
      "0000000" when "00010001100011101", -- t[8989] = 0
      "0000000" when "00010001100011110", -- t[8990] = 0
      "0000000" when "00010001100011111", -- t[8991] = 0
      "0000000" when "00010001100100000", -- t[8992] = 0
      "0000000" when "00010001100100001", -- t[8993] = 0
      "0000000" when "00010001100100010", -- t[8994] = 0
      "0000000" when "00010001100100011", -- t[8995] = 0
      "0000000" when "00010001100100100", -- t[8996] = 0
      "0000000" when "00010001100100101", -- t[8997] = 0
      "0000000" when "00010001100100110", -- t[8998] = 0
      "0000000" when "00010001100100111", -- t[8999] = 0
      "0000000" when "00010001100101000", -- t[9000] = 0
      "0000000" when "00010001100101001", -- t[9001] = 0
      "0000000" when "00010001100101010", -- t[9002] = 0
      "0000000" when "00010001100101011", -- t[9003] = 0
      "0000000" when "00010001100101100", -- t[9004] = 0
      "0000000" when "00010001100101101", -- t[9005] = 0
      "0000000" when "00010001100101110", -- t[9006] = 0
      "0000000" when "00010001100101111", -- t[9007] = 0
      "0000000" when "00010001100110000", -- t[9008] = 0
      "0000000" when "00010001100110001", -- t[9009] = 0
      "0000000" when "00010001100110010", -- t[9010] = 0
      "0000000" when "00010001100110011", -- t[9011] = 0
      "0000000" when "00010001100110100", -- t[9012] = 0
      "0000000" when "00010001100110101", -- t[9013] = 0
      "0000000" when "00010001100110110", -- t[9014] = 0
      "0000000" when "00010001100110111", -- t[9015] = 0
      "0000000" when "00010001100111000", -- t[9016] = 0
      "0000000" when "00010001100111001", -- t[9017] = 0
      "0000000" when "00010001100111010", -- t[9018] = 0
      "0000000" when "00010001100111011", -- t[9019] = 0
      "0000000" when "00010001100111100", -- t[9020] = 0
      "0000000" when "00010001100111101", -- t[9021] = 0
      "0000000" when "00010001100111110", -- t[9022] = 0
      "0000000" when "00010001100111111", -- t[9023] = 0
      "0000000" when "00010001101000000", -- t[9024] = 0
      "0000000" when "00010001101000001", -- t[9025] = 0
      "0000000" when "00010001101000010", -- t[9026] = 0
      "0000000" when "00010001101000011", -- t[9027] = 0
      "0000000" when "00010001101000100", -- t[9028] = 0
      "0000000" when "00010001101000101", -- t[9029] = 0
      "0000000" when "00010001101000110", -- t[9030] = 0
      "0000000" when "00010001101000111", -- t[9031] = 0
      "0000000" when "00010001101001000", -- t[9032] = 0
      "0000000" when "00010001101001001", -- t[9033] = 0
      "0000000" when "00010001101001010", -- t[9034] = 0
      "0000000" when "00010001101001011", -- t[9035] = 0
      "0000000" when "00010001101001100", -- t[9036] = 0
      "0000000" when "00010001101001101", -- t[9037] = 0
      "0000000" when "00010001101001110", -- t[9038] = 0
      "0000000" when "00010001101001111", -- t[9039] = 0
      "0000000" when "00010001101010000", -- t[9040] = 0
      "0000000" when "00010001101010001", -- t[9041] = 0
      "0000000" when "00010001101010010", -- t[9042] = 0
      "0000000" when "00010001101010011", -- t[9043] = 0
      "0000000" when "00010001101010100", -- t[9044] = 0
      "0000000" when "00010001101010101", -- t[9045] = 0
      "0000000" when "00010001101010110", -- t[9046] = 0
      "0000000" when "00010001101010111", -- t[9047] = 0
      "0000000" when "00010001101011000", -- t[9048] = 0
      "0000000" when "00010001101011001", -- t[9049] = 0
      "0000000" when "00010001101011010", -- t[9050] = 0
      "0000000" when "00010001101011011", -- t[9051] = 0
      "0000000" when "00010001101011100", -- t[9052] = 0
      "0000000" when "00010001101011101", -- t[9053] = 0
      "0000000" when "00010001101011110", -- t[9054] = 0
      "0000000" when "00010001101011111", -- t[9055] = 0
      "0000000" when "00010001101100000", -- t[9056] = 0
      "0000000" when "00010001101100001", -- t[9057] = 0
      "0000000" when "00010001101100010", -- t[9058] = 0
      "0000000" when "00010001101100011", -- t[9059] = 0
      "0000000" when "00010001101100100", -- t[9060] = 0
      "0000000" when "00010001101100101", -- t[9061] = 0
      "0000000" when "00010001101100110", -- t[9062] = 0
      "0000000" when "00010001101100111", -- t[9063] = 0
      "0000000" when "00010001101101000", -- t[9064] = 0
      "0000000" when "00010001101101001", -- t[9065] = 0
      "0000000" when "00010001101101010", -- t[9066] = 0
      "0000000" when "00010001101101011", -- t[9067] = 0
      "0000000" when "00010001101101100", -- t[9068] = 0
      "0000000" when "00010001101101101", -- t[9069] = 0
      "0000000" when "00010001101101110", -- t[9070] = 0
      "0000000" when "00010001101101111", -- t[9071] = 0
      "0000000" when "00010001101110000", -- t[9072] = 0
      "0000000" when "00010001101110001", -- t[9073] = 0
      "0000000" when "00010001101110010", -- t[9074] = 0
      "0000000" when "00010001101110011", -- t[9075] = 0
      "0000000" when "00010001101110100", -- t[9076] = 0
      "0000000" when "00010001101110101", -- t[9077] = 0
      "0000000" when "00010001101110110", -- t[9078] = 0
      "0000000" when "00010001101110111", -- t[9079] = 0
      "0000000" when "00010001101111000", -- t[9080] = 0
      "0000000" when "00010001101111001", -- t[9081] = 0
      "0000000" when "00010001101111010", -- t[9082] = 0
      "0000000" when "00010001101111011", -- t[9083] = 0
      "0000000" when "00010001101111100", -- t[9084] = 0
      "0000000" when "00010001101111101", -- t[9085] = 0
      "0000000" when "00010001101111110", -- t[9086] = 0
      "0000000" when "00010001101111111", -- t[9087] = 0
      "0000000" when "00010001110000000", -- t[9088] = 0
      "0000000" when "00010001110000001", -- t[9089] = 0
      "0000000" when "00010001110000010", -- t[9090] = 0
      "0000000" when "00010001110000011", -- t[9091] = 0
      "0000000" when "00010001110000100", -- t[9092] = 0
      "0000000" when "00010001110000101", -- t[9093] = 0
      "0000000" when "00010001110000110", -- t[9094] = 0
      "0000000" when "00010001110000111", -- t[9095] = 0
      "0000000" when "00010001110001000", -- t[9096] = 0
      "0000000" when "00010001110001001", -- t[9097] = 0
      "0000000" when "00010001110001010", -- t[9098] = 0
      "0000000" when "00010001110001011", -- t[9099] = 0
      "0000000" when "00010001110001100", -- t[9100] = 0
      "0000000" when "00010001110001101", -- t[9101] = 0
      "0000000" when "00010001110001110", -- t[9102] = 0
      "0000000" when "00010001110001111", -- t[9103] = 0
      "0000000" when "00010001110010000", -- t[9104] = 0
      "0000000" when "00010001110010001", -- t[9105] = 0
      "0000000" when "00010001110010010", -- t[9106] = 0
      "0000000" when "00010001110010011", -- t[9107] = 0
      "0000000" when "00010001110010100", -- t[9108] = 0
      "0000000" when "00010001110010101", -- t[9109] = 0
      "0000000" when "00010001110010110", -- t[9110] = 0
      "0000000" when "00010001110010111", -- t[9111] = 0
      "0000000" when "00010001110011000", -- t[9112] = 0
      "0000000" when "00010001110011001", -- t[9113] = 0
      "0000000" when "00010001110011010", -- t[9114] = 0
      "0000000" when "00010001110011011", -- t[9115] = 0
      "0000000" when "00010001110011100", -- t[9116] = 0
      "0000000" when "00010001110011101", -- t[9117] = 0
      "0000000" when "00010001110011110", -- t[9118] = 0
      "0000000" when "00010001110011111", -- t[9119] = 0
      "0000000" when "00010001110100000", -- t[9120] = 0
      "0000000" when "00010001110100001", -- t[9121] = 0
      "0000000" when "00010001110100010", -- t[9122] = 0
      "0000000" when "00010001110100011", -- t[9123] = 0
      "0000000" when "00010001110100100", -- t[9124] = 0
      "0000000" when "00010001110100101", -- t[9125] = 0
      "0000000" when "00010001110100110", -- t[9126] = 0
      "0000000" when "00010001110100111", -- t[9127] = 0
      "0000000" when "00010001110101000", -- t[9128] = 0
      "0000000" when "00010001110101001", -- t[9129] = 0
      "0000000" when "00010001110101010", -- t[9130] = 0
      "0000000" when "00010001110101011", -- t[9131] = 0
      "0000000" when "00010001110101100", -- t[9132] = 0
      "0000000" when "00010001110101101", -- t[9133] = 0
      "0000000" when "00010001110101110", -- t[9134] = 0
      "0000000" when "00010001110101111", -- t[9135] = 0
      "0000000" when "00010001110110000", -- t[9136] = 0
      "0000000" when "00010001110110001", -- t[9137] = 0
      "0000000" when "00010001110110010", -- t[9138] = 0
      "0000000" when "00010001110110011", -- t[9139] = 0
      "0000000" when "00010001110110100", -- t[9140] = 0
      "0000000" when "00010001110110101", -- t[9141] = 0
      "0000000" when "00010001110110110", -- t[9142] = 0
      "0000000" when "00010001110110111", -- t[9143] = 0
      "0000000" when "00010001110111000", -- t[9144] = 0
      "0000000" when "00010001110111001", -- t[9145] = 0
      "0000000" when "00010001110111010", -- t[9146] = 0
      "0000000" when "00010001110111011", -- t[9147] = 0
      "0000000" when "00010001110111100", -- t[9148] = 0
      "0000000" when "00010001110111101", -- t[9149] = 0
      "0000000" when "00010001110111110", -- t[9150] = 0
      "0000000" when "00010001110111111", -- t[9151] = 0
      "0000000" when "00010001111000000", -- t[9152] = 0
      "0000000" when "00010001111000001", -- t[9153] = 0
      "0000000" when "00010001111000010", -- t[9154] = 0
      "0000000" when "00010001111000011", -- t[9155] = 0
      "0000000" when "00010001111000100", -- t[9156] = 0
      "0000000" when "00010001111000101", -- t[9157] = 0
      "0000000" when "00010001111000110", -- t[9158] = 0
      "0000000" when "00010001111000111", -- t[9159] = 0
      "0000000" when "00010001111001000", -- t[9160] = 0
      "0000000" when "00010001111001001", -- t[9161] = 0
      "0000000" when "00010001111001010", -- t[9162] = 0
      "0000000" when "00010001111001011", -- t[9163] = 0
      "0000000" when "00010001111001100", -- t[9164] = 0
      "0000000" when "00010001111001101", -- t[9165] = 0
      "0000000" when "00010001111001110", -- t[9166] = 0
      "0000000" when "00010001111001111", -- t[9167] = 0
      "0000000" when "00010001111010000", -- t[9168] = 0
      "0000000" when "00010001111010001", -- t[9169] = 0
      "0000000" when "00010001111010010", -- t[9170] = 0
      "0000000" when "00010001111010011", -- t[9171] = 0
      "0000000" when "00010001111010100", -- t[9172] = 0
      "0000000" when "00010001111010101", -- t[9173] = 0
      "0000000" when "00010001111010110", -- t[9174] = 0
      "0000000" when "00010001111010111", -- t[9175] = 0
      "0000000" when "00010001111011000", -- t[9176] = 0
      "0000000" when "00010001111011001", -- t[9177] = 0
      "0000000" when "00010001111011010", -- t[9178] = 0
      "0000000" when "00010001111011011", -- t[9179] = 0
      "0000000" when "00010001111011100", -- t[9180] = 0
      "0000000" when "00010001111011101", -- t[9181] = 0
      "0000000" when "00010001111011110", -- t[9182] = 0
      "0000000" when "00010001111011111", -- t[9183] = 0
      "0000000" when "00010001111100000", -- t[9184] = 0
      "0000000" when "00010001111100001", -- t[9185] = 0
      "0000000" when "00010001111100010", -- t[9186] = 0
      "0000000" when "00010001111100011", -- t[9187] = 0
      "0000000" when "00010001111100100", -- t[9188] = 0
      "0000000" when "00010001111100101", -- t[9189] = 0
      "0000000" when "00010001111100110", -- t[9190] = 0
      "0000000" when "00010001111100111", -- t[9191] = 0
      "0000000" when "00010001111101000", -- t[9192] = 0
      "0000000" when "00010001111101001", -- t[9193] = 0
      "0000000" when "00010001111101010", -- t[9194] = 0
      "0000000" when "00010001111101011", -- t[9195] = 0
      "0000000" when "00010001111101100", -- t[9196] = 0
      "0000000" when "00010001111101101", -- t[9197] = 0
      "0000000" when "00010001111101110", -- t[9198] = 0
      "0000000" when "00010001111101111", -- t[9199] = 0
      "0000000" when "00010001111110000", -- t[9200] = 0
      "0000000" when "00010001111110001", -- t[9201] = 0
      "0000000" when "00010001111110010", -- t[9202] = 0
      "0000000" when "00010001111110011", -- t[9203] = 0
      "0000000" when "00010001111110100", -- t[9204] = 0
      "0000000" when "00010001111110101", -- t[9205] = 0
      "0000000" when "00010001111110110", -- t[9206] = 0
      "0000000" when "00010001111110111", -- t[9207] = 0
      "0000000" when "00010001111111000", -- t[9208] = 0
      "0000000" when "00010001111111001", -- t[9209] = 0
      "0000000" when "00010001111111010", -- t[9210] = 0
      "0000000" when "00010001111111011", -- t[9211] = 0
      "0000000" when "00010001111111100", -- t[9212] = 0
      "0000000" when "00010001111111101", -- t[9213] = 0
      "0000000" when "00010001111111110", -- t[9214] = 0
      "0000000" when "00010001111111111", -- t[9215] = 0
      "0000000" when "00010010000000000", -- t[9216] = 0
      "0000000" when "00010010000000001", -- t[9217] = 0
      "0000000" when "00010010000000010", -- t[9218] = 0
      "0000000" when "00010010000000011", -- t[9219] = 0
      "0000000" when "00010010000000100", -- t[9220] = 0
      "0000000" when "00010010000000101", -- t[9221] = 0
      "0000000" when "00010010000000110", -- t[9222] = 0
      "0000000" when "00010010000000111", -- t[9223] = 0
      "0000000" when "00010010000001000", -- t[9224] = 0
      "0000000" when "00010010000001001", -- t[9225] = 0
      "0000000" when "00010010000001010", -- t[9226] = 0
      "0000000" when "00010010000001011", -- t[9227] = 0
      "0000000" when "00010010000001100", -- t[9228] = 0
      "0000000" when "00010010000001101", -- t[9229] = 0
      "0000000" when "00010010000001110", -- t[9230] = 0
      "0000000" when "00010010000001111", -- t[9231] = 0
      "0000000" when "00010010000010000", -- t[9232] = 0
      "0000000" when "00010010000010001", -- t[9233] = 0
      "0000000" when "00010010000010010", -- t[9234] = 0
      "0000000" when "00010010000010011", -- t[9235] = 0
      "0000000" when "00010010000010100", -- t[9236] = 0
      "0000000" when "00010010000010101", -- t[9237] = 0
      "0000000" when "00010010000010110", -- t[9238] = 0
      "0000000" when "00010010000010111", -- t[9239] = 0
      "0000000" when "00010010000011000", -- t[9240] = 0
      "0000000" when "00010010000011001", -- t[9241] = 0
      "0000000" when "00010010000011010", -- t[9242] = 0
      "0000000" when "00010010000011011", -- t[9243] = 0
      "0000000" when "00010010000011100", -- t[9244] = 0
      "0000000" when "00010010000011101", -- t[9245] = 0
      "0000000" when "00010010000011110", -- t[9246] = 0
      "0000000" when "00010010000011111", -- t[9247] = 0
      "0000000" when "00010010000100000", -- t[9248] = 0
      "0000000" when "00010010000100001", -- t[9249] = 0
      "0000000" when "00010010000100010", -- t[9250] = 0
      "0000000" when "00010010000100011", -- t[9251] = 0
      "0000000" when "00010010000100100", -- t[9252] = 0
      "0000000" when "00010010000100101", -- t[9253] = 0
      "0000000" when "00010010000100110", -- t[9254] = 0
      "0000000" when "00010010000100111", -- t[9255] = 0
      "0000000" when "00010010000101000", -- t[9256] = 0
      "0000000" when "00010010000101001", -- t[9257] = 0
      "0000000" when "00010010000101010", -- t[9258] = 0
      "0000000" when "00010010000101011", -- t[9259] = 0
      "0000000" when "00010010000101100", -- t[9260] = 0
      "0000000" when "00010010000101101", -- t[9261] = 0
      "0000000" when "00010010000101110", -- t[9262] = 0
      "0000000" when "00010010000101111", -- t[9263] = 0
      "0000000" when "00010010000110000", -- t[9264] = 0
      "0000000" when "00010010000110001", -- t[9265] = 0
      "0000000" when "00010010000110010", -- t[9266] = 0
      "0000000" when "00010010000110011", -- t[9267] = 0
      "0000000" when "00010010000110100", -- t[9268] = 0
      "0000000" when "00010010000110101", -- t[9269] = 0
      "0000000" when "00010010000110110", -- t[9270] = 0
      "0000000" when "00010010000110111", -- t[9271] = 0
      "0000000" when "00010010000111000", -- t[9272] = 0
      "0000000" when "00010010000111001", -- t[9273] = 0
      "0000000" when "00010010000111010", -- t[9274] = 0
      "0000000" when "00010010000111011", -- t[9275] = 0
      "0000000" when "00010010000111100", -- t[9276] = 0
      "0000000" when "00010010000111101", -- t[9277] = 0
      "0000000" when "00010010000111110", -- t[9278] = 0
      "0000000" when "00010010000111111", -- t[9279] = 0
      "0000000" when "00010010001000000", -- t[9280] = 0
      "0000000" when "00010010001000001", -- t[9281] = 0
      "0000000" when "00010010001000010", -- t[9282] = 0
      "0000000" when "00010010001000011", -- t[9283] = 0
      "0000000" when "00010010001000100", -- t[9284] = 0
      "0000000" when "00010010001000101", -- t[9285] = 0
      "0000000" when "00010010001000110", -- t[9286] = 0
      "0000000" when "00010010001000111", -- t[9287] = 0
      "0000000" when "00010010001001000", -- t[9288] = 0
      "0000000" when "00010010001001001", -- t[9289] = 0
      "0000000" when "00010010001001010", -- t[9290] = 0
      "0000000" when "00010010001001011", -- t[9291] = 0
      "0000000" when "00010010001001100", -- t[9292] = 0
      "0000000" when "00010010001001101", -- t[9293] = 0
      "0000000" when "00010010001001110", -- t[9294] = 0
      "0000000" when "00010010001001111", -- t[9295] = 0
      "0000000" when "00010010001010000", -- t[9296] = 0
      "0000000" when "00010010001010001", -- t[9297] = 0
      "0000000" when "00010010001010010", -- t[9298] = 0
      "0000000" when "00010010001010011", -- t[9299] = 0
      "0000000" when "00010010001010100", -- t[9300] = 0
      "0000000" when "00010010001010101", -- t[9301] = 0
      "0000000" when "00010010001010110", -- t[9302] = 0
      "0000000" when "00010010001010111", -- t[9303] = 0
      "0000000" when "00010010001011000", -- t[9304] = 0
      "0000000" when "00010010001011001", -- t[9305] = 0
      "0000000" when "00010010001011010", -- t[9306] = 0
      "0000000" when "00010010001011011", -- t[9307] = 0
      "0000000" when "00010010001011100", -- t[9308] = 0
      "0000000" when "00010010001011101", -- t[9309] = 0
      "0000000" when "00010010001011110", -- t[9310] = 0
      "0000000" when "00010010001011111", -- t[9311] = 0
      "0000000" when "00010010001100000", -- t[9312] = 0
      "0000000" when "00010010001100001", -- t[9313] = 0
      "0000000" when "00010010001100010", -- t[9314] = 0
      "0000000" when "00010010001100011", -- t[9315] = 0
      "0000000" when "00010010001100100", -- t[9316] = 0
      "0000000" when "00010010001100101", -- t[9317] = 0
      "0000000" when "00010010001100110", -- t[9318] = 0
      "0000000" when "00010010001100111", -- t[9319] = 0
      "0000000" when "00010010001101000", -- t[9320] = 0
      "0000000" when "00010010001101001", -- t[9321] = 0
      "0000000" when "00010010001101010", -- t[9322] = 0
      "0000000" when "00010010001101011", -- t[9323] = 0
      "0000000" when "00010010001101100", -- t[9324] = 0
      "0000000" when "00010010001101101", -- t[9325] = 0
      "0000000" when "00010010001101110", -- t[9326] = 0
      "0000000" when "00010010001101111", -- t[9327] = 0
      "0000000" when "00010010001110000", -- t[9328] = 0
      "0000000" when "00010010001110001", -- t[9329] = 0
      "0000000" when "00010010001110010", -- t[9330] = 0
      "0000000" when "00010010001110011", -- t[9331] = 0
      "0000000" when "00010010001110100", -- t[9332] = 0
      "0000000" when "00010010001110101", -- t[9333] = 0
      "0000000" when "00010010001110110", -- t[9334] = 0
      "0000000" when "00010010001110111", -- t[9335] = 0
      "0000000" when "00010010001111000", -- t[9336] = 0
      "0000000" when "00010010001111001", -- t[9337] = 0
      "0000000" when "00010010001111010", -- t[9338] = 0
      "0000000" when "00010010001111011", -- t[9339] = 0
      "0000000" when "00010010001111100", -- t[9340] = 0
      "0000000" when "00010010001111101", -- t[9341] = 0
      "0000000" when "00010010001111110", -- t[9342] = 0
      "0000000" when "00010010001111111", -- t[9343] = 0
      "0000000" when "00010010010000000", -- t[9344] = 0
      "0000000" when "00010010010000001", -- t[9345] = 0
      "0000000" when "00010010010000010", -- t[9346] = 0
      "0000000" when "00010010010000011", -- t[9347] = 0
      "0000000" when "00010010010000100", -- t[9348] = 0
      "0000000" when "00010010010000101", -- t[9349] = 0
      "0000000" when "00010010010000110", -- t[9350] = 0
      "0000000" when "00010010010000111", -- t[9351] = 0
      "0000000" when "00010010010001000", -- t[9352] = 0
      "0000000" when "00010010010001001", -- t[9353] = 0
      "0000000" when "00010010010001010", -- t[9354] = 0
      "0000000" when "00010010010001011", -- t[9355] = 0
      "0000000" when "00010010010001100", -- t[9356] = 0
      "0000000" when "00010010010001101", -- t[9357] = 0
      "0000000" when "00010010010001110", -- t[9358] = 0
      "0000000" when "00010010010001111", -- t[9359] = 0
      "0000000" when "00010010010010000", -- t[9360] = 0
      "0000000" when "00010010010010001", -- t[9361] = 0
      "0000000" when "00010010010010010", -- t[9362] = 0
      "0000000" when "00010010010010011", -- t[9363] = 0
      "0000000" when "00010010010010100", -- t[9364] = 0
      "0000000" when "00010010010010101", -- t[9365] = 0
      "0000000" when "00010010010010110", -- t[9366] = 0
      "0000000" when "00010010010010111", -- t[9367] = 0
      "0000000" when "00010010010011000", -- t[9368] = 0
      "0000000" when "00010010010011001", -- t[9369] = 0
      "0000000" when "00010010010011010", -- t[9370] = 0
      "0000000" when "00010010010011011", -- t[9371] = 0
      "0000000" when "00010010010011100", -- t[9372] = 0
      "0000000" when "00010010010011101", -- t[9373] = 0
      "0000000" when "00010010010011110", -- t[9374] = 0
      "0000000" when "00010010010011111", -- t[9375] = 0
      "0000000" when "00010010010100000", -- t[9376] = 0
      "0000000" when "00010010010100001", -- t[9377] = 0
      "0000000" when "00010010010100010", -- t[9378] = 0
      "0000000" when "00010010010100011", -- t[9379] = 0
      "0000000" when "00010010010100100", -- t[9380] = 0
      "0000000" when "00010010010100101", -- t[9381] = 0
      "0000000" when "00010010010100110", -- t[9382] = 0
      "0000000" when "00010010010100111", -- t[9383] = 0
      "0000000" when "00010010010101000", -- t[9384] = 0
      "0000000" when "00010010010101001", -- t[9385] = 0
      "0000000" when "00010010010101010", -- t[9386] = 0
      "0000000" when "00010010010101011", -- t[9387] = 0
      "0000000" when "00010010010101100", -- t[9388] = 0
      "0000000" when "00010010010101101", -- t[9389] = 0
      "0000000" when "00010010010101110", -- t[9390] = 0
      "0000000" when "00010010010101111", -- t[9391] = 0
      "0000000" when "00010010010110000", -- t[9392] = 0
      "0000000" when "00010010010110001", -- t[9393] = 0
      "0000000" when "00010010010110010", -- t[9394] = 0
      "0000000" when "00010010010110011", -- t[9395] = 0
      "0000000" when "00010010010110100", -- t[9396] = 0
      "0000000" when "00010010010110101", -- t[9397] = 0
      "0000000" when "00010010010110110", -- t[9398] = 0
      "0000000" when "00010010010110111", -- t[9399] = 0
      "0000000" when "00010010010111000", -- t[9400] = 0
      "0000000" when "00010010010111001", -- t[9401] = 0
      "0000000" when "00010010010111010", -- t[9402] = 0
      "0000000" when "00010010010111011", -- t[9403] = 0
      "0000000" when "00010010010111100", -- t[9404] = 0
      "0000000" when "00010010010111101", -- t[9405] = 0
      "0000000" when "00010010010111110", -- t[9406] = 0
      "0000000" when "00010010010111111", -- t[9407] = 0
      "0000000" when "00010010011000000", -- t[9408] = 0
      "0000000" when "00010010011000001", -- t[9409] = 0
      "0000000" when "00010010011000010", -- t[9410] = 0
      "0000000" when "00010010011000011", -- t[9411] = 0
      "0000000" when "00010010011000100", -- t[9412] = 0
      "0000000" when "00010010011000101", -- t[9413] = 0
      "0000000" when "00010010011000110", -- t[9414] = 0
      "0000000" when "00010010011000111", -- t[9415] = 0
      "0000000" when "00010010011001000", -- t[9416] = 0
      "0000000" when "00010010011001001", -- t[9417] = 0
      "0000000" when "00010010011001010", -- t[9418] = 0
      "0000000" when "00010010011001011", -- t[9419] = 0
      "0000000" when "00010010011001100", -- t[9420] = 0
      "0000000" when "00010010011001101", -- t[9421] = 0
      "0000000" when "00010010011001110", -- t[9422] = 0
      "0000000" when "00010010011001111", -- t[9423] = 0
      "0000000" when "00010010011010000", -- t[9424] = 0
      "0000000" when "00010010011010001", -- t[9425] = 0
      "0000000" when "00010010011010010", -- t[9426] = 0
      "0000000" when "00010010011010011", -- t[9427] = 0
      "0000000" when "00010010011010100", -- t[9428] = 0
      "0000000" when "00010010011010101", -- t[9429] = 0
      "0000000" when "00010010011010110", -- t[9430] = 0
      "0000000" when "00010010011010111", -- t[9431] = 0
      "0000000" when "00010010011011000", -- t[9432] = 0
      "0000000" when "00010010011011001", -- t[9433] = 0
      "0000000" when "00010010011011010", -- t[9434] = 0
      "0000000" when "00010010011011011", -- t[9435] = 0
      "0000000" when "00010010011011100", -- t[9436] = 0
      "0000000" when "00010010011011101", -- t[9437] = 0
      "0000000" when "00010010011011110", -- t[9438] = 0
      "0000000" when "00010010011011111", -- t[9439] = 0
      "0000000" when "00010010011100000", -- t[9440] = 0
      "0000000" when "00010010011100001", -- t[9441] = 0
      "0000000" when "00010010011100010", -- t[9442] = 0
      "0000000" when "00010010011100011", -- t[9443] = 0
      "0000000" when "00010010011100100", -- t[9444] = 0
      "0000000" when "00010010011100101", -- t[9445] = 0
      "0000000" when "00010010011100110", -- t[9446] = 0
      "0000000" when "00010010011100111", -- t[9447] = 0
      "0000000" when "00010010011101000", -- t[9448] = 0
      "0000000" when "00010010011101001", -- t[9449] = 0
      "0000000" when "00010010011101010", -- t[9450] = 0
      "0000000" when "00010010011101011", -- t[9451] = 0
      "0000000" when "00010010011101100", -- t[9452] = 0
      "0000000" when "00010010011101101", -- t[9453] = 0
      "0000000" when "00010010011101110", -- t[9454] = 0
      "0000000" when "00010010011101111", -- t[9455] = 0
      "0000000" when "00010010011110000", -- t[9456] = 0
      "0000000" when "00010010011110001", -- t[9457] = 0
      "0000000" when "00010010011110010", -- t[9458] = 0
      "0000000" when "00010010011110011", -- t[9459] = 0
      "0000000" when "00010010011110100", -- t[9460] = 0
      "0000000" when "00010010011110101", -- t[9461] = 0
      "0000000" when "00010010011110110", -- t[9462] = 0
      "0000000" when "00010010011110111", -- t[9463] = 0
      "0000000" when "00010010011111000", -- t[9464] = 0
      "0000000" when "00010010011111001", -- t[9465] = 0
      "0000000" when "00010010011111010", -- t[9466] = 0
      "0000000" when "00010010011111011", -- t[9467] = 0
      "0000000" when "00010010011111100", -- t[9468] = 0
      "0000000" when "00010010011111101", -- t[9469] = 0
      "0000000" when "00010010011111110", -- t[9470] = 0
      "0000000" when "00010010011111111", -- t[9471] = 0
      "0000000" when "00010010100000000", -- t[9472] = 0
      "0000000" when "00010010100000001", -- t[9473] = 0
      "0000000" when "00010010100000010", -- t[9474] = 0
      "0000000" when "00010010100000011", -- t[9475] = 0
      "0000000" when "00010010100000100", -- t[9476] = 0
      "0000000" when "00010010100000101", -- t[9477] = 0
      "0000000" when "00010010100000110", -- t[9478] = 0
      "0000000" when "00010010100000111", -- t[9479] = 0
      "0000000" when "00010010100001000", -- t[9480] = 0
      "0000000" when "00010010100001001", -- t[9481] = 0
      "0000000" when "00010010100001010", -- t[9482] = 0
      "0000000" when "00010010100001011", -- t[9483] = 0
      "0000000" when "00010010100001100", -- t[9484] = 0
      "0000000" when "00010010100001101", -- t[9485] = 0
      "0000000" when "00010010100001110", -- t[9486] = 0
      "0000000" when "00010010100001111", -- t[9487] = 0
      "0000000" when "00010010100010000", -- t[9488] = 0
      "0000000" when "00010010100010001", -- t[9489] = 0
      "0000000" when "00010010100010010", -- t[9490] = 0
      "0000000" when "00010010100010011", -- t[9491] = 0
      "0000000" when "00010010100010100", -- t[9492] = 0
      "0000000" when "00010010100010101", -- t[9493] = 0
      "0000000" when "00010010100010110", -- t[9494] = 0
      "0000000" when "00010010100010111", -- t[9495] = 0
      "0000000" when "00010010100011000", -- t[9496] = 0
      "0000000" when "00010010100011001", -- t[9497] = 0
      "0000000" when "00010010100011010", -- t[9498] = 0
      "0000000" when "00010010100011011", -- t[9499] = 0
      "0000000" when "00010010100011100", -- t[9500] = 0
      "0000000" when "00010010100011101", -- t[9501] = 0
      "0000000" when "00010010100011110", -- t[9502] = 0
      "0000000" when "00010010100011111", -- t[9503] = 0
      "0000000" when "00010010100100000", -- t[9504] = 0
      "0000000" when "00010010100100001", -- t[9505] = 0
      "0000000" when "00010010100100010", -- t[9506] = 0
      "0000000" when "00010010100100011", -- t[9507] = 0
      "0000000" when "00010010100100100", -- t[9508] = 0
      "0000000" when "00010010100100101", -- t[9509] = 0
      "0000000" when "00010010100100110", -- t[9510] = 0
      "0000000" when "00010010100100111", -- t[9511] = 0
      "0000000" when "00010010100101000", -- t[9512] = 0
      "0000000" when "00010010100101001", -- t[9513] = 0
      "0000000" when "00010010100101010", -- t[9514] = 0
      "0000000" when "00010010100101011", -- t[9515] = 0
      "0000000" when "00010010100101100", -- t[9516] = 0
      "0000000" when "00010010100101101", -- t[9517] = 0
      "0000000" when "00010010100101110", -- t[9518] = 0
      "0000000" when "00010010100101111", -- t[9519] = 0
      "0000000" when "00010010100110000", -- t[9520] = 0
      "0000000" when "00010010100110001", -- t[9521] = 0
      "0000000" when "00010010100110010", -- t[9522] = 0
      "0000000" when "00010010100110011", -- t[9523] = 0
      "0000000" when "00010010100110100", -- t[9524] = 0
      "0000000" when "00010010100110101", -- t[9525] = 0
      "0000000" when "00010010100110110", -- t[9526] = 0
      "0000000" when "00010010100110111", -- t[9527] = 0
      "0000000" when "00010010100111000", -- t[9528] = 0
      "0000000" when "00010010100111001", -- t[9529] = 0
      "0000000" when "00010010100111010", -- t[9530] = 0
      "0000000" when "00010010100111011", -- t[9531] = 0
      "0000000" when "00010010100111100", -- t[9532] = 0
      "0000000" when "00010010100111101", -- t[9533] = 0
      "0000000" when "00010010100111110", -- t[9534] = 0
      "0000000" when "00010010100111111", -- t[9535] = 0
      "0000000" when "00010010101000000", -- t[9536] = 0
      "0000000" when "00010010101000001", -- t[9537] = 0
      "0000000" when "00010010101000010", -- t[9538] = 0
      "0000000" when "00010010101000011", -- t[9539] = 0
      "0000000" when "00010010101000100", -- t[9540] = 0
      "0000000" when "00010010101000101", -- t[9541] = 0
      "0000000" when "00010010101000110", -- t[9542] = 0
      "0000000" when "00010010101000111", -- t[9543] = 0
      "0000000" when "00010010101001000", -- t[9544] = 0
      "0000000" when "00010010101001001", -- t[9545] = 0
      "0000000" when "00010010101001010", -- t[9546] = 0
      "0000000" when "00010010101001011", -- t[9547] = 0
      "0000000" when "00010010101001100", -- t[9548] = 0
      "0000000" when "00010010101001101", -- t[9549] = 0
      "0000000" when "00010010101001110", -- t[9550] = 0
      "0000000" when "00010010101001111", -- t[9551] = 0
      "0000000" when "00010010101010000", -- t[9552] = 0
      "0000000" when "00010010101010001", -- t[9553] = 0
      "0000000" when "00010010101010010", -- t[9554] = 0
      "0000000" when "00010010101010011", -- t[9555] = 0
      "0000000" when "00010010101010100", -- t[9556] = 0
      "0000000" when "00010010101010101", -- t[9557] = 0
      "0000000" when "00010010101010110", -- t[9558] = 0
      "0000000" when "00010010101010111", -- t[9559] = 0
      "0000000" when "00010010101011000", -- t[9560] = 0
      "0000000" when "00010010101011001", -- t[9561] = 0
      "0000000" when "00010010101011010", -- t[9562] = 0
      "0000000" when "00010010101011011", -- t[9563] = 0
      "0000000" when "00010010101011100", -- t[9564] = 0
      "0000000" when "00010010101011101", -- t[9565] = 0
      "0000000" when "00010010101011110", -- t[9566] = 0
      "0000000" when "00010010101011111", -- t[9567] = 0
      "0000000" when "00010010101100000", -- t[9568] = 0
      "0000000" when "00010010101100001", -- t[9569] = 0
      "0000000" when "00010010101100010", -- t[9570] = 0
      "0000000" when "00010010101100011", -- t[9571] = 0
      "0000000" when "00010010101100100", -- t[9572] = 0
      "0000000" when "00010010101100101", -- t[9573] = 0
      "0000000" when "00010010101100110", -- t[9574] = 0
      "0000000" when "00010010101100111", -- t[9575] = 0
      "0000000" when "00010010101101000", -- t[9576] = 0
      "0000000" when "00010010101101001", -- t[9577] = 0
      "0000000" when "00010010101101010", -- t[9578] = 0
      "0000000" when "00010010101101011", -- t[9579] = 0
      "0000000" when "00010010101101100", -- t[9580] = 0
      "0000000" when "00010010101101101", -- t[9581] = 0
      "0000000" when "00010010101101110", -- t[9582] = 0
      "0000000" when "00010010101101111", -- t[9583] = 0
      "0000000" when "00010010101110000", -- t[9584] = 0
      "0000000" when "00010010101110001", -- t[9585] = 0
      "0000000" when "00010010101110010", -- t[9586] = 0
      "0000000" when "00010010101110011", -- t[9587] = 0
      "0000000" when "00010010101110100", -- t[9588] = 0
      "0000000" when "00010010101110101", -- t[9589] = 0
      "0000000" when "00010010101110110", -- t[9590] = 0
      "0000000" when "00010010101110111", -- t[9591] = 0
      "0000000" when "00010010101111000", -- t[9592] = 0
      "0000000" when "00010010101111001", -- t[9593] = 0
      "0000000" when "00010010101111010", -- t[9594] = 0
      "0000000" when "00010010101111011", -- t[9595] = 0
      "0000000" when "00010010101111100", -- t[9596] = 0
      "0000000" when "00010010101111101", -- t[9597] = 0
      "0000000" when "00010010101111110", -- t[9598] = 0
      "0000000" when "00010010101111111", -- t[9599] = 0
      "0000000" when "00010010110000000", -- t[9600] = 0
      "0000000" when "00010010110000001", -- t[9601] = 0
      "0000000" when "00010010110000010", -- t[9602] = 0
      "0000000" when "00010010110000011", -- t[9603] = 0
      "0000000" when "00010010110000100", -- t[9604] = 0
      "0000000" when "00010010110000101", -- t[9605] = 0
      "0000000" when "00010010110000110", -- t[9606] = 0
      "0000000" when "00010010110000111", -- t[9607] = 0
      "0000000" when "00010010110001000", -- t[9608] = 0
      "0000000" when "00010010110001001", -- t[9609] = 0
      "0000000" when "00010010110001010", -- t[9610] = 0
      "0000000" when "00010010110001011", -- t[9611] = 0
      "0000000" when "00010010110001100", -- t[9612] = 0
      "0000000" when "00010010110001101", -- t[9613] = 0
      "0000000" when "00010010110001110", -- t[9614] = 0
      "0000000" when "00010010110001111", -- t[9615] = 0
      "0000000" when "00010010110010000", -- t[9616] = 0
      "0000000" when "00010010110010001", -- t[9617] = 0
      "0000000" when "00010010110010010", -- t[9618] = 0
      "0000000" when "00010010110010011", -- t[9619] = 0
      "0000000" when "00010010110010100", -- t[9620] = 0
      "0000000" when "00010010110010101", -- t[9621] = 0
      "0000000" when "00010010110010110", -- t[9622] = 0
      "0000000" when "00010010110010111", -- t[9623] = 0
      "0000000" when "00010010110011000", -- t[9624] = 0
      "0000000" when "00010010110011001", -- t[9625] = 0
      "0000000" when "00010010110011010", -- t[9626] = 0
      "0000000" when "00010010110011011", -- t[9627] = 0
      "0000000" when "00010010110011100", -- t[9628] = 0
      "0000000" when "00010010110011101", -- t[9629] = 0
      "0000000" when "00010010110011110", -- t[9630] = 0
      "0000000" when "00010010110011111", -- t[9631] = 0
      "0000000" when "00010010110100000", -- t[9632] = 0
      "0000000" when "00010010110100001", -- t[9633] = 0
      "0000000" when "00010010110100010", -- t[9634] = 0
      "0000000" when "00010010110100011", -- t[9635] = 0
      "0000000" when "00010010110100100", -- t[9636] = 0
      "0000000" when "00010010110100101", -- t[9637] = 0
      "0000000" when "00010010110100110", -- t[9638] = 0
      "0000000" when "00010010110100111", -- t[9639] = 0
      "0000000" when "00010010110101000", -- t[9640] = 0
      "0000000" when "00010010110101001", -- t[9641] = 0
      "0000000" when "00010010110101010", -- t[9642] = 0
      "0000000" when "00010010110101011", -- t[9643] = 0
      "0000000" when "00010010110101100", -- t[9644] = 0
      "0000000" when "00010010110101101", -- t[9645] = 0
      "0000000" when "00010010110101110", -- t[9646] = 0
      "0000000" when "00010010110101111", -- t[9647] = 0
      "0000000" when "00010010110110000", -- t[9648] = 0
      "0000000" when "00010010110110001", -- t[9649] = 0
      "0000000" when "00010010110110010", -- t[9650] = 0
      "0000000" when "00010010110110011", -- t[9651] = 0
      "0000000" when "00010010110110100", -- t[9652] = 0
      "0000000" when "00010010110110101", -- t[9653] = 0
      "0000000" when "00010010110110110", -- t[9654] = 0
      "0000000" when "00010010110110111", -- t[9655] = 0
      "0000000" when "00010010110111000", -- t[9656] = 0
      "0000000" when "00010010110111001", -- t[9657] = 0
      "0000000" when "00010010110111010", -- t[9658] = 0
      "0000000" when "00010010110111011", -- t[9659] = 0
      "0000000" when "00010010110111100", -- t[9660] = 0
      "0000000" when "00010010110111101", -- t[9661] = 0
      "0000000" when "00010010110111110", -- t[9662] = 0
      "0000000" when "00010010110111111", -- t[9663] = 0
      "0000000" when "00010010111000000", -- t[9664] = 0
      "0000000" when "00010010111000001", -- t[9665] = 0
      "0000000" when "00010010111000010", -- t[9666] = 0
      "0000000" when "00010010111000011", -- t[9667] = 0
      "0000000" when "00010010111000100", -- t[9668] = 0
      "0000000" when "00010010111000101", -- t[9669] = 0
      "0000000" when "00010010111000110", -- t[9670] = 0
      "0000000" when "00010010111000111", -- t[9671] = 0
      "0000000" when "00010010111001000", -- t[9672] = 0
      "0000000" when "00010010111001001", -- t[9673] = 0
      "0000000" when "00010010111001010", -- t[9674] = 0
      "0000000" when "00010010111001011", -- t[9675] = 0
      "0000000" when "00010010111001100", -- t[9676] = 0
      "0000000" when "00010010111001101", -- t[9677] = 0
      "0000000" when "00010010111001110", -- t[9678] = 0
      "0000000" when "00010010111001111", -- t[9679] = 0
      "0000000" when "00010010111010000", -- t[9680] = 0
      "0000000" when "00010010111010001", -- t[9681] = 0
      "0000000" when "00010010111010010", -- t[9682] = 0
      "0000000" when "00010010111010011", -- t[9683] = 0
      "0000000" when "00010010111010100", -- t[9684] = 0
      "0000000" when "00010010111010101", -- t[9685] = 0
      "0000000" when "00010010111010110", -- t[9686] = 0
      "0000000" when "00010010111010111", -- t[9687] = 0
      "0000000" when "00010010111011000", -- t[9688] = 0
      "0000000" when "00010010111011001", -- t[9689] = 0
      "0000000" when "00010010111011010", -- t[9690] = 0
      "0000000" when "00010010111011011", -- t[9691] = 0
      "0000000" when "00010010111011100", -- t[9692] = 0
      "0000000" when "00010010111011101", -- t[9693] = 0
      "0000000" when "00010010111011110", -- t[9694] = 0
      "0000000" when "00010010111011111", -- t[9695] = 0
      "0000000" when "00010010111100000", -- t[9696] = 0
      "0000000" when "00010010111100001", -- t[9697] = 0
      "0000000" when "00010010111100010", -- t[9698] = 0
      "0000000" when "00010010111100011", -- t[9699] = 0
      "0000000" when "00010010111100100", -- t[9700] = 0
      "0000000" when "00010010111100101", -- t[9701] = 0
      "0000000" when "00010010111100110", -- t[9702] = 0
      "0000000" when "00010010111100111", -- t[9703] = 0
      "0000000" when "00010010111101000", -- t[9704] = 0
      "0000000" when "00010010111101001", -- t[9705] = 0
      "0000000" when "00010010111101010", -- t[9706] = 0
      "0000000" when "00010010111101011", -- t[9707] = 0
      "0000000" when "00010010111101100", -- t[9708] = 0
      "0000000" when "00010010111101101", -- t[9709] = 0
      "0000000" when "00010010111101110", -- t[9710] = 0
      "0000000" when "00010010111101111", -- t[9711] = 0
      "0000000" when "00010010111110000", -- t[9712] = 0
      "0000000" when "00010010111110001", -- t[9713] = 0
      "0000000" when "00010010111110010", -- t[9714] = 0
      "0000000" when "00010010111110011", -- t[9715] = 0
      "0000000" when "00010010111110100", -- t[9716] = 0
      "0000000" when "00010010111110101", -- t[9717] = 0
      "0000000" when "00010010111110110", -- t[9718] = 0
      "0000000" when "00010010111110111", -- t[9719] = 0
      "0000000" when "00010010111111000", -- t[9720] = 0
      "0000000" when "00010010111111001", -- t[9721] = 0
      "0000000" when "00010010111111010", -- t[9722] = 0
      "0000000" when "00010010111111011", -- t[9723] = 0
      "0000000" when "00010010111111100", -- t[9724] = 0
      "0000000" when "00010010111111101", -- t[9725] = 0
      "0000000" when "00010010111111110", -- t[9726] = 0
      "0000000" when "00010010111111111", -- t[9727] = 0
      "0000000" when "00010011000000000", -- t[9728] = 0
      "0000000" when "00010011000000001", -- t[9729] = 0
      "0000000" when "00010011000000010", -- t[9730] = 0
      "0000000" when "00010011000000011", -- t[9731] = 0
      "0000000" when "00010011000000100", -- t[9732] = 0
      "0000000" when "00010011000000101", -- t[9733] = 0
      "0000000" when "00010011000000110", -- t[9734] = 0
      "0000000" when "00010011000000111", -- t[9735] = 0
      "0000000" when "00010011000001000", -- t[9736] = 0
      "0000000" when "00010011000001001", -- t[9737] = 0
      "0000000" when "00010011000001010", -- t[9738] = 0
      "0000000" when "00010011000001011", -- t[9739] = 0
      "0000000" when "00010011000001100", -- t[9740] = 0
      "0000000" when "00010011000001101", -- t[9741] = 0
      "0000000" when "00010011000001110", -- t[9742] = 0
      "0000000" when "00010011000001111", -- t[9743] = 0
      "0000000" when "00010011000010000", -- t[9744] = 0
      "0000000" when "00010011000010001", -- t[9745] = 0
      "0000000" when "00010011000010010", -- t[9746] = 0
      "0000000" when "00010011000010011", -- t[9747] = 0
      "0000000" when "00010011000010100", -- t[9748] = 0
      "0000000" when "00010011000010101", -- t[9749] = 0
      "0000000" when "00010011000010110", -- t[9750] = 0
      "0000000" when "00010011000010111", -- t[9751] = 0
      "0000000" when "00010011000011000", -- t[9752] = 0
      "0000000" when "00010011000011001", -- t[9753] = 0
      "0000000" when "00010011000011010", -- t[9754] = 0
      "0000000" when "00010011000011011", -- t[9755] = 0
      "0000000" when "00010011000011100", -- t[9756] = 0
      "0000000" when "00010011000011101", -- t[9757] = 0
      "0000000" when "00010011000011110", -- t[9758] = 0
      "0000000" when "00010011000011111", -- t[9759] = 0
      "0000000" when "00010011000100000", -- t[9760] = 0
      "0000000" when "00010011000100001", -- t[9761] = 0
      "0000000" when "00010011000100010", -- t[9762] = 0
      "0000000" when "00010011000100011", -- t[9763] = 0
      "0000000" when "00010011000100100", -- t[9764] = 0
      "0000000" when "00010011000100101", -- t[9765] = 0
      "0000000" when "00010011000100110", -- t[9766] = 0
      "0000000" when "00010011000100111", -- t[9767] = 0
      "0000000" when "00010011000101000", -- t[9768] = 0
      "0000000" when "00010011000101001", -- t[9769] = 0
      "0000000" when "00010011000101010", -- t[9770] = 0
      "0000000" when "00010011000101011", -- t[9771] = 0
      "0000000" when "00010011000101100", -- t[9772] = 0
      "0000000" when "00010011000101101", -- t[9773] = 0
      "0000000" when "00010011000101110", -- t[9774] = 0
      "0000000" when "00010011000101111", -- t[9775] = 0
      "0000000" when "00010011000110000", -- t[9776] = 0
      "0000000" when "00010011000110001", -- t[9777] = 0
      "0000000" when "00010011000110010", -- t[9778] = 0
      "0000000" when "00010011000110011", -- t[9779] = 0
      "0000000" when "00010011000110100", -- t[9780] = 0
      "0000000" when "00010011000110101", -- t[9781] = 0
      "0000000" when "00010011000110110", -- t[9782] = 0
      "0000000" when "00010011000110111", -- t[9783] = 0
      "0000000" when "00010011000111000", -- t[9784] = 0
      "0000000" when "00010011000111001", -- t[9785] = 0
      "0000000" when "00010011000111010", -- t[9786] = 0
      "0000000" when "00010011000111011", -- t[9787] = 0
      "0000000" when "00010011000111100", -- t[9788] = 0
      "0000000" when "00010011000111101", -- t[9789] = 0
      "0000000" when "00010011000111110", -- t[9790] = 0
      "0000000" when "00010011000111111", -- t[9791] = 0
      "0000000" when "00010011001000000", -- t[9792] = 0
      "0000000" when "00010011001000001", -- t[9793] = 0
      "0000000" when "00010011001000010", -- t[9794] = 0
      "0000000" when "00010011001000011", -- t[9795] = 0
      "0000000" when "00010011001000100", -- t[9796] = 0
      "0000000" when "00010011001000101", -- t[9797] = 0
      "0000000" when "00010011001000110", -- t[9798] = 0
      "0000000" when "00010011001000111", -- t[9799] = 0
      "0000000" when "00010011001001000", -- t[9800] = 0
      "0000000" when "00010011001001001", -- t[9801] = 0
      "0000000" when "00010011001001010", -- t[9802] = 0
      "0000000" when "00010011001001011", -- t[9803] = 0
      "0000000" when "00010011001001100", -- t[9804] = 0
      "0000000" when "00010011001001101", -- t[9805] = 0
      "0000000" when "00010011001001110", -- t[9806] = 0
      "0000000" when "00010011001001111", -- t[9807] = 0
      "0000000" when "00010011001010000", -- t[9808] = 0
      "0000000" when "00010011001010001", -- t[9809] = 0
      "0000000" when "00010011001010010", -- t[9810] = 0
      "0000000" when "00010011001010011", -- t[9811] = 0
      "0000000" when "00010011001010100", -- t[9812] = 0
      "0000000" when "00010011001010101", -- t[9813] = 0
      "0000000" when "00010011001010110", -- t[9814] = 0
      "0000000" when "00010011001010111", -- t[9815] = 0
      "0000000" when "00010011001011000", -- t[9816] = 0
      "0000000" when "00010011001011001", -- t[9817] = 0
      "0000000" when "00010011001011010", -- t[9818] = 0
      "0000000" when "00010011001011011", -- t[9819] = 0
      "0000000" when "00010011001011100", -- t[9820] = 0
      "0000000" when "00010011001011101", -- t[9821] = 0
      "0000000" when "00010011001011110", -- t[9822] = 0
      "0000000" when "00010011001011111", -- t[9823] = 0
      "0000000" when "00010011001100000", -- t[9824] = 0
      "0000000" when "00010011001100001", -- t[9825] = 0
      "0000000" when "00010011001100010", -- t[9826] = 0
      "0000000" when "00010011001100011", -- t[9827] = 0
      "0000000" when "00010011001100100", -- t[9828] = 0
      "0000000" when "00010011001100101", -- t[9829] = 0
      "0000000" when "00010011001100110", -- t[9830] = 0
      "0000000" when "00010011001100111", -- t[9831] = 0
      "0000000" when "00010011001101000", -- t[9832] = 0
      "0000000" when "00010011001101001", -- t[9833] = 0
      "0000000" when "00010011001101010", -- t[9834] = 0
      "0000000" when "00010011001101011", -- t[9835] = 0
      "0000000" when "00010011001101100", -- t[9836] = 0
      "0000000" when "00010011001101101", -- t[9837] = 0
      "0000000" when "00010011001101110", -- t[9838] = 0
      "0000000" when "00010011001101111", -- t[9839] = 0
      "0000000" when "00010011001110000", -- t[9840] = 0
      "0000000" when "00010011001110001", -- t[9841] = 0
      "0000000" when "00010011001110010", -- t[9842] = 0
      "0000000" when "00010011001110011", -- t[9843] = 0
      "0000000" when "00010011001110100", -- t[9844] = 0
      "0000000" when "00010011001110101", -- t[9845] = 0
      "0000000" when "00010011001110110", -- t[9846] = 0
      "0000000" when "00010011001110111", -- t[9847] = 0
      "0000000" when "00010011001111000", -- t[9848] = 0
      "0000000" when "00010011001111001", -- t[9849] = 0
      "0000000" when "00010011001111010", -- t[9850] = 0
      "0000000" when "00010011001111011", -- t[9851] = 0
      "0000000" when "00010011001111100", -- t[9852] = 0
      "0000000" when "00010011001111101", -- t[9853] = 0
      "0000000" when "00010011001111110", -- t[9854] = 0
      "0000000" when "00010011001111111", -- t[9855] = 0
      "0000000" when "00010011010000000", -- t[9856] = 0
      "0000000" when "00010011010000001", -- t[9857] = 0
      "0000000" when "00010011010000010", -- t[9858] = 0
      "0000000" when "00010011010000011", -- t[9859] = 0
      "0000000" when "00010011010000100", -- t[9860] = 0
      "0000000" when "00010011010000101", -- t[9861] = 0
      "0000000" when "00010011010000110", -- t[9862] = 0
      "0000000" when "00010011010000111", -- t[9863] = 0
      "0000000" when "00010011010001000", -- t[9864] = 0
      "0000000" when "00010011010001001", -- t[9865] = 0
      "0000000" when "00010011010001010", -- t[9866] = 0
      "0000000" when "00010011010001011", -- t[9867] = 0
      "0000000" when "00010011010001100", -- t[9868] = 0
      "0000000" when "00010011010001101", -- t[9869] = 0
      "0000000" when "00010011010001110", -- t[9870] = 0
      "0000000" when "00010011010001111", -- t[9871] = 0
      "0000000" when "00010011010010000", -- t[9872] = 0
      "0000000" when "00010011010010001", -- t[9873] = 0
      "0000000" when "00010011010010010", -- t[9874] = 0
      "0000000" when "00010011010010011", -- t[9875] = 0
      "0000000" when "00010011010010100", -- t[9876] = 0
      "0000000" when "00010011010010101", -- t[9877] = 0
      "0000000" when "00010011010010110", -- t[9878] = 0
      "0000000" when "00010011010010111", -- t[9879] = 0
      "0000000" when "00010011010011000", -- t[9880] = 0
      "0000000" when "00010011010011001", -- t[9881] = 0
      "0000000" when "00010011010011010", -- t[9882] = 0
      "0000000" when "00010011010011011", -- t[9883] = 0
      "0000000" when "00010011010011100", -- t[9884] = 0
      "0000000" when "00010011010011101", -- t[9885] = 0
      "0000000" when "00010011010011110", -- t[9886] = 0
      "0000000" when "00010011010011111", -- t[9887] = 0
      "0000000" when "00010011010100000", -- t[9888] = 0
      "0000000" when "00010011010100001", -- t[9889] = 0
      "0000000" when "00010011010100010", -- t[9890] = 0
      "0000000" when "00010011010100011", -- t[9891] = 0
      "0000000" when "00010011010100100", -- t[9892] = 0
      "0000000" when "00010011010100101", -- t[9893] = 0
      "0000000" when "00010011010100110", -- t[9894] = 0
      "0000000" when "00010011010100111", -- t[9895] = 0
      "0000000" when "00010011010101000", -- t[9896] = 0
      "0000000" when "00010011010101001", -- t[9897] = 0
      "0000000" when "00010011010101010", -- t[9898] = 0
      "0000000" when "00010011010101011", -- t[9899] = 0
      "0000000" when "00010011010101100", -- t[9900] = 0
      "0000000" when "00010011010101101", -- t[9901] = 0
      "0000000" when "00010011010101110", -- t[9902] = 0
      "0000000" when "00010011010101111", -- t[9903] = 0
      "0000000" when "00010011010110000", -- t[9904] = 0
      "0000000" when "00010011010110001", -- t[9905] = 0
      "0000000" when "00010011010110010", -- t[9906] = 0
      "0000000" when "00010011010110011", -- t[9907] = 0
      "0000000" when "00010011010110100", -- t[9908] = 0
      "0000000" when "00010011010110101", -- t[9909] = 0
      "0000000" when "00010011010110110", -- t[9910] = 0
      "0000000" when "00010011010110111", -- t[9911] = 0
      "0000000" when "00010011010111000", -- t[9912] = 0
      "0000000" when "00010011010111001", -- t[9913] = 0
      "0000000" when "00010011010111010", -- t[9914] = 0
      "0000000" when "00010011010111011", -- t[9915] = 0
      "0000000" when "00010011010111100", -- t[9916] = 0
      "0000000" when "00010011010111101", -- t[9917] = 0
      "0000000" when "00010011010111110", -- t[9918] = 0
      "0000000" when "00010011010111111", -- t[9919] = 0
      "0000000" when "00010011011000000", -- t[9920] = 0
      "0000000" when "00010011011000001", -- t[9921] = 0
      "0000000" when "00010011011000010", -- t[9922] = 0
      "0000000" when "00010011011000011", -- t[9923] = 0
      "0000000" when "00010011011000100", -- t[9924] = 0
      "0000000" when "00010011011000101", -- t[9925] = 0
      "0000000" when "00010011011000110", -- t[9926] = 0
      "0000000" when "00010011011000111", -- t[9927] = 0
      "0000000" when "00010011011001000", -- t[9928] = 0
      "0000000" when "00010011011001001", -- t[9929] = 0
      "0000000" when "00010011011001010", -- t[9930] = 0
      "0000000" when "00010011011001011", -- t[9931] = 0
      "0000000" when "00010011011001100", -- t[9932] = 0
      "0000000" when "00010011011001101", -- t[9933] = 0
      "0000000" when "00010011011001110", -- t[9934] = 0
      "0000000" when "00010011011001111", -- t[9935] = 0
      "0000000" when "00010011011010000", -- t[9936] = 0
      "0000000" when "00010011011010001", -- t[9937] = 0
      "0000000" when "00010011011010010", -- t[9938] = 0
      "0000000" when "00010011011010011", -- t[9939] = 0
      "0000000" when "00010011011010100", -- t[9940] = 0
      "0000000" when "00010011011010101", -- t[9941] = 0
      "0000000" when "00010011011010110", -- t[9942] = 0
      "0000000" when "00010011011010111", -- t[9943] = 0
      "0000000" when "00010011011011000", -- t[9944] = 0
      "0000000" when "00010011011011001", -- t[9945] = 0
      "0000000" when "00010011011011010", -- t[9946] = 0
      "0000000" when "00010011011011011", -- t[9947] = 0
      "0000000" when "00010011011011100", -- t[9948] = 0
      "0000000" when "00010011011011101", -- t[9949] = 0
      "0000000" when "00010011011011110", -- t[9950] = 0
      "0000000" when "00010011011011111", -- t[9951] = 0
      "0000000" when "00010011011100000", -- t[9952] = 0
      "0000000" when "00010011011100001", -- t[9953] = 0
      "0000000" when "00010011011100010", -- t[9954] = 0
      "0000000" when "00010011011100011", -- t[9955] = 0
      "0000000" when "00010011011100100", -- t[9956] = 0
      "0000000" when "00010011011100101", -- t[9957] = 0
      "0000000" when "00010011011100110", -- t[9958] = 0
      "0000000" when "00010011011100111", -- t[9959] = 0
      "0000000" when "00010011011101000", -- t[9960] = 0
      "0000000" when "00010011011101001", -- t[9961] = 0
      "0000000" when "00010011011101010", -- t[9962] = 0
      "0000000" when "00010011011101011", -- t[9963] = 0
      "0000000" when "00010011011101100", -- t[9964] = 0
      "0000000" when "00010011011101101", -- t[9965] = 0
      "0000000" when "00010011011101110", -- t[9966] = 0
      "0000000" when "00010011011101111", -- t[9967] = 0
      "0000000" when "00010011011110000", -- t[9968] = 0
      "0000000" when "00010011011110001", -- t[9969] = 0
      "0000000" when "00010011011110010", -- t[9970] = 0
      "0000000" when "00010011011110011", -- t[9971] = 0
      "0000000" when "00010011011110100", -- t[9972] = 0
      "0000000" when "00010011011110101", -- t[9973] = 0
      "0000000" when "00010011011110110", -- t[9974] = 0
      "0000000" when "00010011011110111", -- t[9975] = 0
      "0000000" when "00010011011111000", -- t[9976] = 0
      "0000000" when "00010011011111001", -- t[9977] = 0
      "0000000" when "00010011011111010", -- t[9978] = 0
      "0000000" when "00010011011111011", -- t[9979] = 0
      "0000000" when "00010011011111100", -- t[9980] = 0
      "0000000" when "00010011011111101", -- t[9981] = 0
      "0000000" when "00010011011111110", -- t[9982] = 0
      "0000000" when "00010011011111111", -- t[9983] = 0
      "0000000" when "00010011100000000", -- t[9984] = 0
      "0000000" when "00010011100000001", -- t[9985] = 0
      "0000000" when "00010011100000010", -- t[9986] = 0
      "0000000" when "00010011100000011", -- t[9987] = 0
      "0000000" when "00010011100000100", -- t[9988] = 0
      "0000000" when "00010011100000101", -- t[9989] = 0
      "0000000" when "00010011100000110", -- t[9990] = 0
      "0000000" when "00010011100000111", -- t[9991] = 0
      "0000000" when "00010011100001000", -- t[9992] = 0
      "0000000" when "00010011100001001", -- t[9993] = 0
      "0000000" when "00010011100001010", -- t[9994] = 0
      "0000000" when "00010011100001011", -- t[9995] = 0
      "0000000" when "00010011100001100", -- t[9996] = 0
      "0000000" when "00010011100001101", -- t[9997] = 0
      "0000000" when "00010011100001110", -- t[9998] = 0
      "0000000" when "00010011100001111", -- t[9999] = 0
      "0000000" when "00010011100010000", -- t[10000] = 0
      "0000000" when "00010011100010001", -- t[10001] = 0
      "0000000" when "00010011100010010", -- t[10002] = 0
      "0000000" when "00010011100010011", -- t[10003] = 0
      "0000000" when "00010011100010100", -- t[10004] = 0
      "0000000" when "00010011100010101", -- t[10005] = 0
      "0000000" when "00010011100010110", -- t[10006] = 0
      "0000000" when "00010011100010111", -- t[10007] = 0
      "0000000" when "00010011100011000", -- t[10008] = 0
      "0000000" when "00010011100011001", -- t[10009] = 0
      "0000000" when "00010011100011010", -- t[10010] = 0
      "0000000" when "00010011100011011", -- t[10011] = 0
      "0000000" when "00010011100011100", -- t[10012] = 0
      "0000000" when "00010011100011101", -- t[10013] = 0
      "0000000" when "00010011100011110", -- t[10014] = 0
      "0000000" when "00010011100011111", -- t[10015] = 0
      "0000000" when "00010011100100000", -- t[10016] = 0
      "0000000" when "00010011100100001", -- t[10017] = 0
      "0000000" when "00010011100100010", -- t[10018] = 0
      "0000000" when "00010011100100011", -- t[10019] = 0
      "0000000" when "00010011100100100", -- t[10020] = 0
      "0000000" when "00010011100100101", -- t[10021] = 0
      "0000000" when "00010011100100110", -- t[10022] = 0
      "0000000" when "00010011100100111", -- t[10023] = 0
      "0000000" when "00010011100101000", -- t[10024] = 0
      "0000000" when "00010011100101001", -- t[10025] = 0
      "0000000" when "00010011100101010", -- t[10026] = 0
      "0000000" when "00010011100101011", -- t[10027] = 0
      "0000000" when "00010011100101100", -- t[10028] = 0
      "0000000" when "00010011100101101", -- t[10029] = 0
      "0000000" when "00010011100101110", -- t[10030] = 0
      "0000000" when "00010011100101111", -- t[10031] = 0
      "0000000" when "00010011100110000", -- t[10032] = 0
      "0000000" when "00010011100110001", -- t[10033] = 0
      "0000000" when "00010011100110010", -- t[10034] = 0
      "0000000" when "00010011100110011", -- t[10035] = 0
      "0000000" when "00010011100110100", -- t[10036] = 0
      "0000000" when "00010011100110101", -- t[10037] = 0
      "0000000" when "00010011100110110", -- t[10038] = 0
      "0000000" when "00010011100110111", -- t[10039] = 0
      "0000000" when "00010011100111000", -- t[10040] = 0
      "0000000" when "00010011100111001", -- t[10041] = 0
      "0000000" when "00010011100111010", -- t[10042] = 0
      "0000000" when "00010011100111011", -- t[10043] = 0
      "0000000" when "00010011100111100", -- t[10044] = 0
      "0000000" when "00010011100111101", -- t[10045] = 0
      "0000000" when "00010011100111110", -- t[10046] = 0
      "0000000" when "00010011100111111", -- t[10047] = 0
      "0000000" when "00010011101000000", -- t[10048] = 0
      "0000000" when "00010011101000001", -- t[10049] = 0
      "0000000" when "00010011101000010", -- t[10050] = 0
      "0000000" when "00010011101000011", -- t[10051] = 0
      "0000000" when "00010011101000100", -- t[10052] = 0
      "0000000" when "00010011101000101", -- t[10053] = 0
      "0000000" when "00010011101000110", -- t[10054] = 0
      "0000000" when "00010011101000111", -- t[10055] = 0
      "0000000" when "00010011101001000", -- t[10056] = 0
      "0000000" when "00010011101001001", -- t[10057] = 0
      "0000000" when "00010011101001010", -- t[10058] = 0
      "0000000" when "00010011101001011", -- t[10059] = 0
      "0000000" when "00010011101001100", -- t[10060] = 0
      "0000000" when "00010011101001101", -- t[10061] = 0
      "0000000" when "00010011101001110", -- t[10062] = 0
      "0000000" when "00010011101001111", -- t[10063] = 0
      "0000000" when "00010011101010000", -- t[10064] = 0
      "0000000" when "00010011101010001", -- t[10065] = 0
      "0000000" when "00010011101010010", -- t[10066] = 0
      "0000000" when "00010011101010011", -- t[10067] = 0
      "0000000" when "00010011101010100", -- t[10068] = 0
      "0000000" when "00010011101010101", -- t[10069] = 0
      "0000000" when "00010011101010110", -- t[10070] = 0
      "0000000" when "00010011101010111", -- t[10071] = 0
      "0000000" when "00010011101011000", -- t[10072] = 0
      "0000000" when "00010011101011001", -- t[10073] = 0
      "0000000" when "00010011101011010", -- t[10074] = 0
      "0000000" when "00010011101011011", -- t[10075] = 0
      "0000000" when "00010011101011100", -- t[10076] = 0
      "0000000" when "00010011101011101", -- t[10077] = 0
      "0000000" when "00010011101011110", -- t[10078] = 0
      "0000000" when "00010011101011111", -- t[10079] = 0
      "0000000" when "00010011101100000", -- t[10080] = 0
      "0000000" when "00010011101100001", -- t[10081] = 0
      "0000000" when "00010011101100010", -- t[10082] = 0
      "0000000" when "00010011101100011", -- t[10083] = 0
      "0000000" when "00010011101100100", -- t[10084] = 0
      "0000000" when "00010011101100101", -- t[10085] = 0
      "0000000" when "00010011101100110", -- t[10086] = 0
      "0000000" when "00010011101100111", -- t[10087] = 0
      "0000000" when "00010011101101000", -- t[10088] = 0
      "0000000" when "00010011101101001", -- t[10089] = 0
      "0000000" when "00010011101101010", -- t[10090] = 0
      "0000000" when "00010011101101011", -- t[10091] = 0
      "0000000" when "00010011101101100", -- t[10092] = 0
      "0000000" when "00010011101101101", -- t[10093] = 0
      "0000000" when "00010011101101110", -- t[10094] = 0
      "0000000" when "00010011101101111", -- t[10095] = 0
      "0000000" when "00010011101110000", -- t[10096] = 0
      "0000000" when "00010011101110001", -- t[10097] = 0
      "0000000" when "00010011101110010", -- t[10098] = 0
      "0000000" when "00010011101110011", -- t[10099] = 0
      "0000000" when "00010011101110100", -- t[10100] = 0
      "0000000" when "00010011101110101", -- t[10101] = 0
      "0000000" when "00010011101110110", -- t[10102] = 0
      "0000000" when "00010011101110111", -- t[10103] = 0
      "0000000" when "00010011101111000", -- t[10104] = 0
      "0000000" when "00010011101111001", -- t[10105] = 0
      "0000000" when "00010011101111010", -- t[10106] = 0
      "0000000" when "00010011101111011", -- t[10107] = 0
      "0000000" when "00010011101111100", -- t[10108] = 0
      "0000000" when "00010011101111101", -- t[10109] = 0
      "0000000" when "00010011101111110", -- t[10110] = 0
      "0000000" when "00010011101111111", -- t[10111] = 0
      "0000000" when "00010011110000000", -- t[10112] = 0
      "0000000" when "00010011110000001", -- t[10113] = 0
      "0000000" when "00010011110000010", -- t[10114] = 0
      "0000000" when "00010011110000011", -- t[10115] = 0
      "0000000" when "00010011110000100", -- t[10116] = 0
      "0000000" when "00010011110000101", -- t[10117] = 0
      "0000000" when "00010011110000110", -- t[10118] = 0
      "0000000" when "00010011110000111", -- t[10119] = 0
      "0000000" when "00010011110001000", -- t[10120] = 0
      "0000000" when "00010011110001001", -- t[10121] = 0
      "0000000" when "00010011110001010", -- t[10122] = 0
      "0000000" when "00010011110001011", -- t[10123] = 0
      "0000000" when "00010011110001100", -- t[10124] = 0
      "0000000" when "00010011110001101", -- t[10125] = 0
      "0000000" when "00010011110001110", -- t[10126] = 0
      "0000000" when "00010011110001111", -- t[10127] = 0
      "0000000" when "00010011110010000", -- t[10128] = 0
      "0000000" when "00010011110010001", -- t[10129] = 0
      "0000000" when "00010011110010010", -- t[10130] = 0
      "0000000" when "00010011110010011", -- t[10131] = 0
      "0000000" when "00010011110010100", -- t[10132] = 0
      "0000000" when "00010011110010101", -- t[10133] = 0
      "0000000" when "00010011110010110", -- t[10134] = 0
      "0000000" when "00010011110010111", -- t[10135] = 0
      "0000000" when "00010011110011000", -- t[10136] = 0
      "0000000" when "00010011110011001", -- t[10137] = 0
      "0000000" when "00010011110011010", -- t[10138] = 0
      "0000000" when "00010011110011011", -- t[10139] = 0
      "0000000" when "00010011110011100", -- t[10140] = 0
      "0000000" when "00010011110011101", -- t[10141] = 0
      "0000000" when "00010011110011110", -- t[10142] = 0
      "0000000" when "00010011110011111", -- t[10143] = 0
      "0000000" when "00010011110100000", -- t[10144] = 0
      "0000000" when "00010011110100001", -- t[10145] = 0
      "0000000" when "00010011110100010", -- t[10146] = 0
      "0000000" when "00010011110100011", -- t[10147] = 0
      "0000000" when "00010011110100100", -- t[10148] = 0
      "0000000" when "00010011110100101", -- t[10149] = 0
      "0000000" when "00010011110100110", -- t[10150] = 0
      "0000000" when "00010011110100111", -- t[10151] = 0
      "0000000" when "00010011110101000", -- t[10152] = 0
      "0000000" when "00010011110101001", -- t[10153] = 0
      "0000000" when "00010011110101010", -- t[10154] = 0
      "0000000" when "00010011110101011", -- t[10155] = 0
      "0000000" when "00010011110101100", -- t[10156] = 0
      "0000000" when "00010011110101101", -- t[10157] = 0
      "0000000" when "00010011110101110", -- t[10158] = 0
      "0000000" when "00010011110101111", -- t[10159] = 0
      "0000000" when "00010011110110000", -- t[10160] = 0
      "0000000" when "00010011110110001", -- t[10161] = 0
      "0000000" when "00010011110110010", -- t[10162] = 0
      "0000000" when "00010011110110011", -- t[10163] = 0
      "0000000" when "00010011110110100", -- t[10164] = 0
      "0000000" when "00010011110110101", -- t[10165] = 0
      "0000000" when "00010011110110110", -- t[10166] = 0
      "0000000" when "00010011110110111", -- t[10167] = 0
      "0000000" when "00010011110111000", -- t[10168] = 0
      "0000000" when "00010011110111001", -- t[10169] = 0
      "0000000" when "00010011110111010", -- t[10170] = 0
      "0000000" when "00010011110111011", -- t[10171] = 0
      "0000000" when "00010011110111100", -- t[10172] = 0
      "0000000" when "00010011110111101", -- t[10173] = 0
      "0000000" when "00010011110111110", -- t[10174] = 0
      "0000000" when "00010011110111111", -- t[10175] = 0
      "0000000" when "00010011111000000", -- t[10176] = 0
      "0000000" when "00010011111000001", -- t[10177] = 0
      "0000000" when "00010011111000010", -- t[10178] = 0
      "0000000" when "00010011111000011", -- t[10179] = 0
      "0000000" when "00010011111000100", -- t[10180] = 0
      "0000000" when "00010011111000101", -- t[10181] = 0
      "0000000" when "00010011111000110", -- t[10182] = 0
      "0000000" when "00010011111000111", -- t[10183] = 0
      "0000000" when "00010011111001000", -- t[10184] = 0
      "0000000" when "00010011111001001", -- t[10185] = 0
      "0000000" when "00010011111001010", -- t[10186] = 0
      "0000000" when "00010011111001011", -- t[10187] = 0
      "0000000" when "00010011111001100", -- t[10188] = 0
      "0000000" when "00010011111001101", -- t[10189] = 0
      "0000000" when "00010011111001110", -- t[10190] = 0
      "0000000" when "00010011111001111", -- t[10191] = 0
      "0000000" when "00010011111010000", -- t[10192] = 0
      "0000000" when "00010011111010001", -- t[10193] = 0
      "0000000" when "00010011111010010", -- t[10194] = 0
      "0000000" when "00010011111010011", -- t[10195] = 0
      "0000000" when "00010011111010100", -- t[10196] = 0
      "0000000" when "00010011111010101", -- t[10197] = 0
      "0000000" when "00010011111010110", -- t[10198] = 0
      "0000000" when "00010011111010111", -- t[10199] = 0
      "0000000" when "00010011111011000", -- t[10200] = 0
      "0000000" when "00010011111011001", -- t[10201] = 0
      "0000000" when "00010011111011010", -- t[10202] = 0
      "0000000" when "00010011111011011", -- t[10203] = 0
      "0000000" when "00010011111011100", -- t[10204] = 0
      "0000000" when "00010011111011101", -- t[10205] = 0
      "0000000" when "00010011111011110", -- t[10206] = 0
      "0000000" when "00010011111011111", -- t[10207] = 0
      "0000000" when "00010011111100000", -- t[10208] = 0
      "0000000" when "00010011111100001", -- t[10209] = 0
      "0000000" when "00010011111100010", -- t[10210] = 0
      "0000000" when "00010011111100011", -- t[10211] = 0
      "0000000" when "00010011111100100", -- t[10212] = 0
      "0000000" when "00010011111100101", -- t[10213] = 0
      "0000000" when "00010011111100110", -- t[10214] = 0
      "0000000" when "00010011111100111", -- t[10215] = 0
      "0000000" when "00010011111101000", -- t[10216] = 0
      "0000000" when "00010011111101001", -- t[10217] = 0
      "0000000" when "00010011111101010", -- t[10218] = 0
      "0000000" when "00010011111101011", -- t[10219] = 0
      "0000000" when "00010011111101100", -- t[10220] = 0
      "0000000" when "00010011111101101", -- t[10221] = 0
      "0000000" when "00010011111101110", -- t[10222] = 0
      "0000000" when "00010011111101111", -- t[10223] = 0
      "0000000" when "00010011111110000", -- t[10224] = 0
      "0000000" when "00010011111110001", -- t[10225] = 0
      "0000000" when "00010011111110010", -- t[10226] = 0
      "0000000" when "00010011111110011", -- t[10227] = 0
      "0000000" when "00010011111110100", -- t[10228] = 0
      "0000000" when "00010011111110101", -- t[10229] = 0
      "0000000" when "00010011111110110", -- t[10230] = 0
      "0000000" when "00010011111110111", -- t[10231] = 0
      "0000000" when "00010011111111000", -- t[10232] = 0
      "0000000" when "00010011111111001", -- t[10233] = 0
      "0000000" when "00010011111111010", -- t[10234] = 0
      "0000000" when "00010011111111011", -- t[10235] = 0
      "0000000" when "00010011111111100", -- t[10236] = 0
      "0000000" when "00010011111111101", -- t[10237] = 0
      "0000000" when "00010011111111110", -- t[10238] = 0
      "0000000" when "00010011111111111", -- t[10239] = 0
      "0000000" when "00010100000000000", -- t[10240] = 0
      "0000000" when "00010100000000001", -- t[10241] = 0
      "0000000" when "00010100000000010", -- t[10242] = 0
      "0000000" when "00010100000000011", -- t[10243] = 0
      "0000000" when "00010100000000100", -- t[10244] = 0
      "0000000" when "00010100000000101", -- t[10245] = 0
      "0000000" when "00010100000000110", -- t[10246] = 0
      "0000000" when "00010100000000111", -- t[10247] = 0
      "0000000" when "00010100000001000", -- t[10248] = 0
      "0000000" when "00010100000001001", -- t[10249] = 0
      "0000000" when "00010100000001010", -- t[10250] = 0
      "0000000" when "00010100000001011", -- t[10251] = 0
      "0000000" when "00010100000001100", -- t[10252] = 0
      "0000000" when "00010100000001101", -- t[10253] = 0
      "0000000" when "00010100000001110", -- t[10254] = 0
      "0000000" when "00010100000001111", -- t[10255] = 0
      "0000000" when "00010100000010000", -- t[10256] = 0
      "0000000" when "00010100000010001", -- t[10257] = 0
      "0000000" when "00010100000010010", -- t[10258] = 0
      "0000000" when "00010100000010011", -- t[10259] = 0
      "0000000" when "00010100000010100", -- t[10260] = 0
      "0000000" when "00010100000010101", -- t[10261] = 0
      "0000000" when "00010100000010110", -- t[10262] = 0
      "0000000" when "00010100000010111", -- t[10263] = 0
      "0000000" when "00010100000011000", -- t[10264] = 0
      "0000000" when "00010100000011001", -- t[10265] = 0
      "0000000" when "00010100000011010", -- t[10266] = 0
      "0000000" when "00010100000011011", -- t[10267] = 0
      "0000000" when "00010100000011100", -- t[10268] = 0
      "0000000" when "00010100000011101", -- t[10269] = 0
      "0000000" when "00010100000011110", -- t[10270] = 0
      "0000000" when "00010100000011111", -- t[10271] = 0
      "0000000" when "00010100000100000", -- t[10272] = 0
      "0000000" when "00010100000100001", -- t[10273] = 0
      "0000000" when "00010100000100010", -- t[10274] = 0
      "0000000" when "00010100000100011", -- t[10275] = 0
      "0000000" when "00010100000100100", -- t[10276] = 0
      "0000000" when "00010100000100101", -- t[10277] = 0
      "0000000" when "00010100000100110", -- t[10278] = 0
      "0000000" when "00010100000100111", -- t[10279] = 0
      "0000000" when "00010100000101000", -- t[10280] = 0
      "0000000" when "00010100000101001", -- t[10281] = 0
      "0000000" when "00010100000101010", -- t[10282] = 0
      "0000000" when "00010100000101011", -- t[10283] = 0
      "0000000" when "00010100000101100", -- t[10284] = 0
      "0000000" when "00010100000101101", -- t[10285] = 0
      "0000000" when "00010100000101110", -- t[10286] = 0
      "0000000" when "00010100000101111", -- t[10287] = 0
      "0000000" when "00010100000110000", -- t[10288] = 0
      "0000000" when "00010100000110001", -- t[10289] = 0
      "0000000" when "00010100000110010", -- t[10290] = 0
      "0000000" when "00010100000110011", -- t[10291] = 0
      "0000000" when "00010100000110100", -- t[10292] = 0
      "0000000" when "00010100000110101", -- t[10293] = 0
      "0000000" when "00010100000110110", -- t[10294] = 0
      "0000000" when "00010100000110111", -- t[10295] = 0
      "0000000" when "00010100000111000", -- t[10296] = 0
      "0000000" when "00010100000111001", -- t[10297] = 0
      "0000000" when "00010100000111010", -- t[10298] = 0
      "0000000" when "00010100000111011", -- t[10299] = 0
      "0000000" when "00010100000111100", -- t[10300] = 0
      "0000000" when "00010100000111101", -- t[10301] = 0
      "0000000" when "00010100000111110", -- t[10302] = 0
      "0000000" when "00010100000111111", -- t[10303] = 0
      "0000000" when "00010100001000000", -- t[10304] = 0
      "0000000" when "00010100001000001", -- t[10305] = 0
      "0000000" when "00010100001000010", -- t[10306] = 0
      "0000000" when "00010100001000011", -- t[10307] = 0
      "0000000" when "00010100001000100", -- t[10308] = 0
      "0000000" when "00010100001000101", -- t[10309] = 0
      "0000000" when "00010100001000110", -- t[10310] = 0
      "0000000" when "00010100001000111", -- t[10311] = 0
      "0000000" when "00010100001001000", -- t[10312] = 0
      "0000000" when "00010100001001001", -- t[10313] = 0
      "0000000" when "00010100001001010", -- t[10314] = 0
      "0000000" when "00010100001001011", -- t[10315] = 0
      "0000000" when "00010100001001100", -- t[10316] = 0
      "0000000" when "00010100001001101", -- t[10317] = 0
      "0000000" when "00010100001001110", -- t[10318] = 0
      "0000000" when "00010100001001111", -- t[10319] = 0
      "0000000" when "00010100001010000", -- t[10320] = 0
      "0000000" when "00010100001010001", -- t[10321] = 0
      "0000000" when "00010100001010010", -- t[10322] = 0
      "0000000" when "00010100001010011", -- t[10323] = 0
      "0000000" when "00010100001010100", -- t[10324] = 0
      "0000000" when "00010100001010101", -- t[10325] = 0
      "0000000" when "00010100001010110", -- t[10326] = 0
      "0000000" when "00010100001010111", -- t[10327] = 0
      "0000000" when "00010100001011000", -- t[10328] = 0
      "0000000" when "00010100001011001", -- t[10329] = 0
      "0000000" when "00010100001011010", -- t[10330] = 0
      "0000000" when "00010100001011011", -- t[10331] = 0
      "0000000" when "00010100001011100", -- t[10332] = 0
      "0000000" when "00010100001011101", -- t[10333] = 0
      "0000000" when "00010100001011110", -- t[10334] = 0
      "0000000" when "00010100001011111", -- t[10335] = 0
      "0000000" when "00010100001100000", -- t[10336] = 0
      "0000000" when "00010100001100001", -- t[10337] = 0
      "0000000" when "00010100001100010", -- t[10338] = 0
      "0000000" when "00010100001100011", -- t[10339] = 0
      "0000000" when "00010100001100100", -- t[10340] = 0
      "0000000" when "00010100001100101", -- t[10341] = 0
      "0000000" when "00010100001100110", -- t[10342] = 0
      "0000000" when "00010100001100111", -- t[10343] = 0
      "0000000" when "00010100001101000", -- t[10344] = 0
      "0000000" when "00010100001101001", -- t[10345] = 0
      "0000000" when "00010100001101010", -- t[10346] = 0
      "0000000" when "00010100001101011", -- t[10347] = 0
      "0000000" when "00010100001101100", -- t[10348] = 0
      "0000000" when "00010100001101101", -- t[10349] = 0
      "0000000" when "00010100001101110", -- t[10350] = 0
      "0000000" when "00010100001101111", -- t[10351] = 0
      "0000000" when "00010100001110000", -- t[10352] = 0
      "0000000" when "00010100001110001", -- t[10353] = 0
      "0000000" when "00010100001110010", -- t[10354] = 0
      "0000000" when "00010100001110011", -- t[10355] = 0
      "0000000" when "00010100001110100", -- t[10356] = 0
      "0000000" when "00010100001110101", -- t[10357] = 0
      "0000000" when "00010100001110110", -- t[10358] = 0
      "0000000" when "00010100001110111", -- t[10359] = 0
      "0000000" when "00010100001111000", -- t[10360] = 0
      "0000000" when "00010100001111001", -- t[10361] = 0
      "0000000" when "00010100001111010", -- t[10362] = 0
      "0000000" when "00010100001111011", -- t[10363] = 0
      "0000000" when "00010100001111100", -- t[10364] = 0
      "0000000" when "00010100001111101", -- t[10365] = 0
      "0000000" when "00010100001111110", -- t[10366] = 0
      "0000000" when "00010100001111111", -- t[10367] = 0
      "0000000" when "00010100010000000", -- t[10368] = 0
      "0000000" when "00010100010000001", -- t[10369] = 0
      "0000000" when "00010100010000010", -- t[10370] = 0
      "0000000" when "00010100010000011", -- t[10371] = 0
      "0000000" when "00010100010000100", -- t[10372] = 0
      "0000000" when "00010100010000101", -- t[10373] = 0
      "0000000" when "00010100010000110", -- t[10374] = 0
      "0000000" when "00010100010000111", -- t[10375] = 0
      "0000000" when "00010100010001000", -- t[10376] = 0
      "0000000" when "00010100010001001", -- t[10377] = 0
      "0000000" when "00010100010001010", -- t[10378] = 0
      "0000000" when "00010100010001011", -- t[10379] = 0
      "0000000" when "00010100010001100", -- t[10380] = 0
      "0000000" when "00010100010001101", -- t[10381] = 0
      "0000000" when "00010100010001110", -- t[10382] = 0
      "0000000" when "00010100010001111", -- t[10383] = 0
      "0000000" when "00010100010010000", -- t[10384] = 0
      "0000000" when "00010100010010001", -- t[10385] = 0
      "0000000" when "00010100010010010", -- t[10386] = 0
      "0000000" when "00010100010010011", -- t[10387] = 0
      "0000000" when "00010100010010100", -- t[10388] = 0
      "0000000" when "00010100010010101", -- t[10389] = 0
      "0000000" when "00010100010010110", -- t[10390] = 0
      "0000000" when "00010100010010111", -- t[10391] = 0
      "0000000" when "00010100010011000", -- t[10392] = 0
      "0000000" when "00010100010011001", -- t[10393] = 0
      "0000000" when "00010100010011010", -- t[10394] = 0
      "0000000" when "00010100010011011", -- t[10395] = 0
      "0000000" when "00010100010011100", -- t[10396] = 0
      "0000000" when "00010100010011101", -- t[10397] = 0
      "0000000" when "00010100010011110", -- t[10398] = 0
      "0000000" when "00010100010011111", -- t[10399] = 0
      "0000000" when "00010100010100000", -- t[10400] = 0
      "0000000" when "00010100010100001", -- t[10401] = 0
      "0000000" when "00010100010100010", -- t[10402] = 0
      "0000000" when "00010100010100011", -- t[10403] = 0
      "0000000" when "00010100010100100", -- t[10404] = 0
      "0000000" when "00010100010100101", -- t[10405] = 0
      "0000000" when "00010100010100110", -- t[10406] = 0
      "0000000" when "00010100010100111", -- t[10407] = 0
      "0000000" when "00010100010101000", -- t[10408] = 0
      "0000000" when "00010100010101001", -- t[10409] = 0
      "0000000" when "00010100010101010", -- t[10410] = 0
      "0000000" when "00010100010101011", -- t[10411] = 0
      "0000000" when "00010100010101100", -- t[10412] = 0
      "0000000" when "00010100010101101", -- t[10413] = 0
      "0000000" when "00010100010101110", -- t[10414] = 0
      "0000000" when "00010100010101111", -- t[10415] = 0
      "0000000" when "00010100010110000", -- t[10416] = 0
      "0000000" when "00010100010110001", -- t[10417] = 0
      "0000000" when "00010100010110010", -- t[10418] = 0
      "0000000" when "00010100010110011", -- t[10419] = 0
      "0000000" when "00010100010110100", -- t[10420] = 0
      "0000000" when "00010100010110101", -- t[10421] = 0
      "0000000" when "00010100010110110", -- t[10422] = 0
      "0000000" when "00010100010110111", -- t[10423] = 0
      "0000000" when "00010100010111000", -- t[10424] = 0
      "0000000" when "00010100010111001", -- t[10425] = 0
      "0000000" when "00010100010111010", -- t[10426] = 0
      "0000000" when "00010100010111011", -- t[10427] = 0
      "0000000" when "00010100010111100", -- t[10428] = 0
      "0000000" when "00010100010111101", -- t[10429] = 0
      "0000000" when "00010100010111110", -- t[10430] = 0
      "0000000" when "00010100010111111", -- t[10431] = 0
      "0000000" when "00010100011000000", -- t[10432] = 0
      "0000000" when "00010100011000001", -- t[10433] = 0
      "0000000" when "00010100011000010", -- t[10434] = 0
      "0000000" when "00010100011000011", -- t[10435] = 0
      "0000000" when "00010100011000100", -- t[10436] = 0
      "0000000" when "00010100011000101", -- t[10437] = 0
      "0000000" when "00010100011000110", -- t[10438] = 0
      "0000000" when "00010100011000111", -- t[10439] = 0
      "0000000" when "00010100011001000", -- t[10440] = 0
      "0000000" when "00010100011001001", -- t[10441] = 0
      "0000000" when "00010100011001010", -- t[10442] = 0
      "0000000" when "00010100011001011", -- t[10443] = 0
      "0000000" when "00010100011001100", -- t[10444] = 0
      "0000000" when "00010100011001101", -- t[10445] = 0
      "0000000" when "00010100011001110", -- t[10446] = 0
      "0000000" when "00010100011001111", -- t[10447] = 0
      "0000000" when "00010100011010000", -- t[10448] = 0
      "0000000" when "00010100011010001", -- t[10449] = 0
      "0000000" when "00010100011010010", -- t[10450] = 0
      "0000000" when "00010100011010011", -- t[10451] = 0
      "0000000" when "00010100011010100", -- t[10452] = 0
      "0000000" when "00010100011010101", -- t[10453] = 0
      "0000000" when "00010100011010110", -- t[10454] = 0
      "0000000" when "00010100011010111", -- t[10455] = 0
      "0000000" when "00010100011011000", -- t[10456] = 0
      "0000000" when "00010100011011001", -- t[10457] = 0
      "0000000" when "00010100011011010", -- t[10458] = 0
      "0000000" when "00010100011011011", -- t[10459] = 0
      "0000000" when "00010100011011100", -- t[10460] = 0
      "0000000" when "00010100011011101", -- t[10461] = 0
      "0000000" when "00010100011011110", -- t[10462] = 0
      "0000000" when "00010100011011111", -- t[10463] = 0
      "0000000" when "00010100011100000", -- t[10464] = 0
      "0000000" when "00010100011100001", -- t[10465] = 0
      "0000000" when "00010100011100010", -- t[10466] = 0
      "0000000" when "00010100011100011", -- t[10467] = 0
      "0000000" when "00010100011100100", -- t[10468] = 0
      "0000000" when "00010100011100101", -- t[10469] = 0
      "0000000" when "00010100011100110", -- t[10470] = 0
      "0000000" when "00010100011100111", -- t[10471] = 0
      "0000000" when "00010100011101000", -- t[10472] = 0
      "0000000" when "00010100011101001", -- t[10473] = 0
      "0000000" when "00010100011101010", -- t[10474] = 0
      "0000000" when "00010100011101011", -- t[10475] = 0
      "0000000" when "00010100011101100", -- t[10476] = 0
      "0000000" when "00010100011101101", -- t[10477] = 0
      "0000000" when "00010100011101110", -- t[10478] = 0
      "0000000" when "00010100011101111", -- t[10479] = 0
      "0000000" when "00010100011110000", -- t[10480] = 0
      "0000000" when "00010100011110001", -- t[10481] = 0
      "0000000" when "00010100011110010", -- t[10482] = 0
      "0000000" when "00010100011110011", -- t[10483] = 0
      "0000000" when "00010100011110100", -- t[10484] = 0
      "0000000" when "00010100011110101", -- t[10485] = 0
      "0000000" when "00010100011110110", -- t[10486] = 0
      "0000000" when "00010100011110111", -- t[10487] = 0
      "0000000" when "00010100011111000", -- t[10488] = 0
      "0000000" when "00010100011111001", -- t[10489] = 0
      "0000000" when "00010100011111010", -- t[10490] = 0
      "0000000" when "00010100011111011", -- t[10491] = 0
      "0000000" when "00010100011111100", -- t[10492] = 0
      "0000000" when "00010100011111101", -- t[10493] = 0
      "0000000" when "00010100011111110", -- t[10494] = 0
      "0000000" when "00010100011111111", -- t[10495] = 0
      "0000000" when "00010100100000000", -- t[10496] = 0
      "0000000" when "00010100100000001", -- t[10497] = 0
      "0000000" when "00010100100000010", -- t[10498] = 0
      "0000000" when "00010100100000011", -- t[10499] = 0
      "0000000" when "00010100100000100", -- t[10500] = 0
      "0000000" when "00010100100000101", -- t[10501] = 0
      "0000000" when "00010100100000110", -- t[10502] = 0
      "0000000" when "00010100100000111", -- t[10503] = 0
      "0000000" when "00010100100001000", -- t[10504] = 0
      "0000000" when "00010100100001001", -- t[10505] = 0
      "0000000" when "00010100100001010", -- t[10506] = 0
      "0000000" when "00010100100001011", -- t[10507] = 0
      "0000000" when "00010100100001100", -- t[10508] = 0
      "0000000" when "00010100100001101", -- t[10509] = 0
      "0000000" when "00010100100001110", -- t[10510] = 0
      "0000000" when "00010100100001111", -- t[10511] = 0
      "0000000" when "00010100100010000", -- t[10512] = 0
      "0000000" when "00010100100010001", -- t[10513] = 0
      "0000000" when "00010100100010010", -- t[10514] = 0
      "0000000" when "00010100100010011", -- t[10515] = 0
      "0000000" when "00010100100010100", -- t[10516] = 0
      "0000000" when "00010100100010101", -- t[10517] = 0
      "0000000" when "00010100100010110", -- t[10518] = 0
      "0000000" when "00010100100010111", -- t[10519] = 0
      "0000000" when "00010100100011000", -- t[10520] = 0
      "0000000" when "00010100100011001", -- t[10521] = 0
      "0000000" when "00010100100011010", -- t[10522] = 0
      "0000000" when "00010100100011011", -- t[10523] = 0
      "0000000" when "00010100100011100", -- t[10524] = 0
      "0000000" when "00010100100011101", -- t[10525] = 0
      "0000000" when "00010100100011110", -- t[10526] = 0
      "0000000" when "00010100100011111", -- t[10527] = 0
      "0000000" when "00010100100100000", -- t[10528] = 0
      "0000000" when "00010100100100001", -- t[10529] = 0
      "0000000" when "00010100100100010", -- t[10530] = 0
      "0000000" when "00010100100100011", -- t[10531] = 0
      "0000000" when "00010100100100100", -- t[10532] = 0
      "0000000" when "00010100100100101", -- t[10533] = 0
      "0000000" when "00010100100100110", -- t[10534] = 0
      "0000000" when "00010100100100111", -- t[10535] = 0
      "0000000" when "00010100100101000", -- t[10536] = 0
      "0000000" when "00010100100101001", -- t[10537] = 0
      "0000000" when "00010100100101010", -- t[10538] = 0
      "0000000" when "00010100100101011", -- t[10539] = 0
      "0000000" when "00010100100101100", -- t[10540] = 0
      "0000000" when "00010100100101101", -- t[10541] = 0
      "0000000" when "00010100100101110", -- t[10542] = 0
      "0000000" when "00010100100101111", -- t[10543] = 0
      "0000000" when "00010100100110000", -- t[10544] = 0
      "0000000" when "00010100100110001", -- t[10545] = 0
      "0000000" when "00010100100110010", -- t[10546] = 0
      "0000000" when "00010100100110011", -- t[10547] = 0
      "0000000" when "00010100100110100", -- t[10548] = 0
      "0000000" when "00010100100110101", -- t[10549] = 0
      "0000000" when "00010100100110110", -- t[10550] = 0
      "0000000" when "00010100100110111", -- t[10551] = 0
      "0000000" when "00010100100111000", -- t[10552] = 0
      "0000000" when "00010100100111001", -- t[10553] = 0
      "0000000" when "00010100100111010", -- t[10554] = 0
      "0000000" when "00010100100111011", -- t[10555] = 0
      "0000000" when "00010100100111100", -- t[10556] = 0
      "0000000" when "00010100100111101", -- t[10557] = 0
      "0000000" when "00010100100111110", -- t[10558] = 0
      "0000000" when "00010100100111111", -- t[10559] = 0
      "0000000" when "00010100101000000", -- t[10560] = 0
      "0000000" when "00010100101000001", -- t[10561] = 0
      "0000000" when "00010100101000010", -- t[10562] = 0
      "0000000" when "00010100101000011", -- t[10563] = 0
      "0000000" when "00010100101000100", -- t[10564] = 0
      "0000000" when "00010100101000101", -- t[10565] = 0
      "0000000" when "00010100101000110", -- t[10566] = 0
      "0000000" when "00010100101000111", -- t[10567] = 0
      "0000000" when "00010100101001000", -- t[10568] = 0
      "0000000" when "00010100101001001", -- t[10569] = 0
      "0000000" when "00010100101001010", -- t[10570] = 0
      "0000000" when "00010100101001011", -- t[10571] = 0
      "0000000" when "00010100101001100", -- t[10572] = 0
      "0000000" when "00010100101001101", -- t[10573] = 0
      "0000000" when "00010100101001110", -- t[10574] = 0
      "0000000" when "00010100101001111", -- t[10575] = 0
      "0000000" when "00010100101010000", -- t[10576] = 0
      "0000000" when "00010100101010001", -- t[10577] = 0
      "0000000" when "00010100101010010", -- t[10578] = 0
      "0000000" when "00010100101010011", -- t[10579] = 0
      "0000000" when "00010100101010100", -- t[10580] = 0
      "0000000" when "00010100101010101", -- t[10581] = 0
      "0000000" when "00010100101010110", -- t[10582] = 0
      "0000000" when "00010100101010111", -- t[10583] = 0
      "0000000" when "00010100101011000", -- t[10584] = 0
      "0000000" when "00010100101011001", -- t[10585] = 0
      "0000000" when "00010100101011010", -- t[10586] = 0
      "0000000" when "00010100101011011", -- t[10587] = 0
      "0000000" when "00010100101011100", -- t[10588] = 0
      "0000000" when "00010100101011101", -- t[10589] = 0
      "0000000" when "00010100101011110", -- t[10590] = 0
      "0000000" when "00010100101011111", -- t[10591] = 0
      "0000000" when "00010100101100000", -- t[10592] = 0
      "0000000" when "00010100101100001", -- t[10593] = 0
      "0000000" when "00010100101100010", -- t[10594] = 0
      "0000000" when "00010100101100011", -- t[10595] = 0
      "0000000" when "00010100101100100", -- t[10596] = 0
      "0000000" when "00010100101100101", -- t[10597] = 0
      "0000000" when "00010100101100110", -- t[10598] = 0
      "0000000" when "00010100101100111", -- t[10599] = 0
      "0000000" when "00010100101101000", -- t[10600] = 0
      "0000000" when "00010100101101001", -- t[10601] = 0
      "0000000" when "00010100101101010", -- t[10602] = 0
      "0000000" when "00010100101101011", -- t[10603] = 0
      "0000000" when "00010100101101100", -- t[10604] = 0
      "0000000" when "00010100101101101", -- t[10605] = 0
      "0000000" when "00010100101101110", -- t[10606] = 0
      "0000000" when "00010100101101111", -- t[10607] = 0
      "0000000" when "00010100101110000", -- t[10608] = 0
      "0000000" when "00010100101110001", -- t[10609] = 0
      "0000000" when "00010100101110010", -- t[10610] = 0
      "0000000" when "00010100101110011", -- t[10611] = 0
      "0000000" when "00010100101110100", -- t[10612] = 0
      "0000000" when "00010100101110101", -- t[10613] = 0
      "0000000" when "00010100101110110", -- t[10614] = 0
      "0000000" when "00010100101110111", -- t[10615] = 0
      "0000000" when "00010100101111000", -- t[10616] = 0
      "0000000" when "00010100101111001", -- t[10617] = 0
      "0000000" when "00010100101111010", -- t[10618] = 0
      "0000000" when "00010100101111011", -- t[10619] = 0
      "0000000" when "00010100101111100", -- t[10620] = 0
      "0000000" when "00010100101111101", -- t[10621] = 0
      "0000000" when "00010100101111110", -- t[10622] = 0
      "0000000" when "00010100101111111", -- t[10623] = 0
      "0000000" when "00010100110000000", -- t[10624] = 0
      "0000000" when "00010100110000001", -- t[10625] = 0
      "0000000" when "00010100110000010", -- t[10626] = 0
      "0000000" when "00010100110000011", -- t[10627] = 0
      "0000000" when "00010100110000100", -- t[10628] = 0
      "0000000" when "00010100110000101", -- t[10629] = 0
      "0000000" when "00010100110000110", -- t[10630] = 0
      "0000000" when "00010100110000111", -- t[10631] = 0
      "0000000" when "00010100110001000", -- t[10632] = 0
      "0000000" when "00010100110001001", -- t[10633] = 0
      "0000000" when "00010100110001010", -- t[10634] = 0
      "0000000" when "00010100110001011", -- t[10635] = 0
      "0000000" when "00010100110001100", -- t[10636] = 0
      "0000000" when "00010100110001101", -- t[10637] = 0
      "0000000" when "00010100110001110", -- t[10638] = 0
      "0000000" when "00010100110001111", -- t[10639] = 0
      "0000000" when "00010100110010000", -- t[10640] = 0
      "0000000" when "00010100110010001", -- t[10641] = 0
      "0000000" when "00010100110010010", -- t[10642] = 0
      "0000000" when "00010100110010011", -- t[10643] = 0
      "0000000" when "00010100110010100", -- t[10644] = 0
      "0000000" when "00010100110010101", -- t[10645] = 0
      "0000000" when "00010100110010110", -- t[10646] = 0
      "0000000" when "00010100110010111", -- t[10647] = 0
      "0000000" when "00010100110011000", -- t[10648] = 0
      "0000000" when "00010100110011001", -- t[10649] = 0
      "0000000" when "00010100110011010", -- t[10650] = 0
      "0000000" when "00010100110011011", -- t[10651] = 0
      "0000000" when "00010100110011100", -- t[10652] = 0
      "0000000" when "00010100110011101", -- t[10653] = 0
      "0000000" when "00010100110011110", -- t[10654] = 0
      "0000000" when "00010100110011111", -- t[10655] = 0
      "0000000" when "00010100110100000", -- t[10656] = 0
      "0000000" when "00010100110100001", -- t[10657] = 0
      "0000000" when "00010100110100010", -- t[10658] = 0
      "0000000" when "00010100110100011", -- t[10659] = 0
      "0000000" when "00010100110100100", -- t[10660] = 0
      "0000000" when "00010100110100101", -- t[10661] = 0
      "0000000" when "00010100110100110", -- t[10662] = 0
      "0000000" when "00010100110100111", -- t[10663] = 0
      "0000000" when "00010100110101000", -- t[10664] = 0
      "0000000" when "00010100110101001", -- t[10665] = 0
      "0000000" when "00010100110101010", -- t[10666] = 0
      "0000000" when "00010100110101011", -- t[10667] = 0
      "0000000" when "00010100110101100", -- t[10668] = 0
      "0000000" when "00010100110101101", -- t[10669] = 0
      "0000000" when "00010100110101110", -- t[10670] = 0
      "0000000" when "00010100110101111", -- t[10671] = 0
      "0000000" when "00010100110110000", -- t[10672] = 0
      "0000000" when "00010100110110001", -- t[10673] = 0
      "0000000" when "00010100110110010", -- t[10674] = 0
      "0000000" when "00010100110110011", -- t[10675] = 0
      "0000000" when "00010100110110100", -- t[10676] = 0
      "0000000" when "00010100110110101", -- t[10677] = 0
      "0000000" when "00010100110110110", -- t[10678] = 0
      "0000000" when "00010100110110111", -- t[10679] = 0
      "0000000" when "00010100110111000", -- t[10680] = 0
      "0000000" when "00010100110111001", -- t[10681] = 0
      "0000000" when "00010100110111010", -- t[10682] = 0
      "0000000" when "00010100110111011", -- t[10683] = 0
      "0000000" when "00010100110111100", -- t[10684] = 0
      "0000000" when "00010100110111101", -- t[10685] = 0
      "0000000" when "00010100110111110", -- t[10686] = 0
      "0000000" when "00010100110111111", -- t[10687] = 0
      "0000000" when "00010100111000000", -- t[10688] = 0
      "0000000" when "00010100111000001", -- t[10689] = 0
      "0000000" when "00010100111000010", -- t[10690] = 0
      "0000000" when "00010100111000011", -- t[10691] = 0
      "0000000" when "00010100111000100", -- t[10692] = 0
      "0000000" when "00010100111000101", -- t[10693] = 0
      "0000000" when "00010100111000110", -- t[10694] = 0
      "0000000" when "00010100111000111", -- t[10695] = 0
      "0000000" when "00010100111001000", -- t[10696] = 0
      "0000000" when "00010100111001001", -- t[10697] = 0
      "0000000" when "00010100111001010", -- t[10698] = 0
      "0000000" when "00010100111001011", -- t[10699] = 0
      "0000000" when "00010100111001100", -- t[10700] = 0
      "0000000" when "00010100111001101", -- t[10701] = 0
      "0000000" when "00010100111001110", -- t[10702] = 0
      "0000000" when "00010100111001111", -- t[10703] = 0
      "0000000" when "00010100111010000", -- t[10704] = 0
      "0000000" when "00010100111010001", -- t[10705] = 0
      "0000000" when "00010100111010010", -- t[10706] = 0
      "0000000" when "00010100111010011", -- t[10707] = 0
      "0000000" when "00010100111010100", -- t[10708] = 0
      "0000000" when "00010100111010101", -- t[10709] = 0
      "0000000" when "00010100111010110", -- t[10710] = 0
      "0000000" when "00010100111010111", -- t[10711] = 0
      "0000000" when "00010100111011000", -- t[10712] = 0
      "0000000" when "00010100111011001", -- t[10713] = 0
      "0000000" when "00010100111011010", -- t[10714] = 0
      "0000000" when "00010100111011011", -- t[10715] = 0
      "0000000" when "00010100111011100", -- t[10716] = 0
      "0000000" when "00010100111011101", -- t[10717] = 0
      "0000000" when "00010100111011110", -- t[10718] = 0
      "0000000" when "00010100111011111", -- t[10719] = 0
      "0000000" when "00010100111100000", -- t[10720] = 0
      "0000000" when "00010100111100001", -- t[10721] = 0
      "0000000" when "00010100111100010", -- t[10722] = 0
      "0000000" when "00010100111100011", -- t[10723] = 0
      "0000000" when "00010100111100100", -- t[10724] = 0
      "0000000" when "00010100111100101", -- t[10725] = 0
      "0000000" when "00010100111100110", -- t[10726] = 0
      "0000000" when "00010100111100111", -- t[10727] = 0
      "0000000" when "00010100111101000", -- t[10728] = 0
      "0000000" when "00010100111101001", -- t[10729] = 0
      "0000000" when "00010100111101010", -- t[10730] = 0
      "0000000" when "00010100111101011", -- t[10731] = 0
      "0000000" when "00010100111101100", -- t[10732] = 0
      "0000000" when "00010100111101101", -- t[10733] = 0
      "0000000" when "00010100111101110", -- t[10734] = 0
      "0000000" when "00010100111101111", -- t[10735] = 0
      "0000000" when "00010100111110000", -- t[10736] = 0
      "0000000" when "00010100111110001", -- t[10737] = 0
      "0000000" when "00010100111110010", -- t[10738] = 0
      "0000000" when "00010100111110011", -- t[10739] = 0
      "0000000" when "00010100111110100", -- t[10740] = 0
      "0000000" when "00010100111110101", -- t[10741] = 0
      "0000000" when "00010100111110110", -- t[10742] = 0
      "0000000" when "00010100111110111", -- t[10743] = 0
      "0000000" when "00010100111111000", -- t[10744] = 0
      "0000000" when "00010100111111001", -- t[10745] = 0
      "0000000" when "00010100111111010", -- t[10746] = 0
      "0000000" when "00010100111111011", -- t[10747] = 0
      "0000000" when "00010100111111100", -- t[10748] = 0
      "0000000" when "00010100111111101", -- t[10749] = 0
      "0000000" when "00010100111111110", -- t[10750] = 0
      "0000000" when "00010100111111111", -- t[10751] = 0
      "0000000" when "00010101000000000", -- t[10752] = 0
      "0000000" when "00010101000000001", -- t[10753] = 0
      "0000000" when "00010101000000010", -- t[10754] = 0
      "0000000" when "00010101000000011", -- t[10755] = 0
      "0000000" when "00010101000000100", -- t[10756] = 0
      "0000000" when "00010101000000101", -- t[10757] = 0
      "0000000" when "00010101000000110", -- t[10758] = 0
      "0000000" when "00010101000000111", -- t[10759] = 0
      "0000000" when "00010101000001000", -- t[10760] = 0
      "0000000" when "00010101000001001", -- t[10761] = 0
      "0000000" when "00010101000001010", -- t[10762] = 0
      "0000000" when "00010101000001011", -- t[10763] = 0
      "0000000" when "00010101000001100", -- t[10764] = 0
      "0000000" when "00010101000001101", -- t[10765] = 0
      "0000000" when "00010101000001110", -- t[10766] = 0
      "0000000" when "00010101000001111", -- t[10767] = 0
      "0000000" when "00010101000010000", -- t[10768] = 0
      "0000000" when "00010101000010001", -- t[10769] = 0
      "0000000" when "00010101000010010", -- t[10770] = 0
      "0000000" when "00010101000010011", -- t[10771] = 0
      "0000000" when "00010101000010100", -- t[10772] = 0
      "0000000" when "00010101000010101", -- t[10773] = 0
      "0000000" when "00010101000010110", -- t[10774] = 0
      "0000000" when "00010101000010111", -- t[10775] = 0
      "0000000" when "00010101000011000", -- t[10776] = 0
      "0000000" when "00010101000011001", -- t[10777] = 0
      "0000000" when "00010101000011010", -- t[10778] = 0
      "0000000" when "00010101000011011", -- t[10779] = 0
      "0000000" when "00010101000011100", -- t[10780] = 0
      "0000000" when "00010101000011101", -- t[10781] = 0
      "0000000" when "00010101000011110", -- t[10782] = 0
      "0000000" when "00010101000011111", -- t[10783] = 0
      "0000000" when "00010101000100000", -- t[10784] = 0
      "0000000" when "00010101000100001", -- t[10785] = 0
      "0000000" when "00010101000100010", -- t[10786] = 0
      "0000000" when "00010101000100011", -- t[10787] = 0
      "0000000" when "00010101000100100", -- t[10788] = 0
      "0000000" when "00010101000100101", -- t[10789] = 0
      "0000000" when "00010101000100110", -- t[10790] = 0
      "0000000" when "00010101000100111", -- t[10791] = 0
      "0000000" when "00010101000101000", -- t[10792] = 0
      "0000000" when "00010101000101001", -- t[10793] = 0
      "0000000" when "00010101000101010", -- t[10794] = 0
      "0000000" when "00010101000101011", -- t[10795] = 0
      "0000000" when "00010101000101100", -- t[10796] = 0
      "0000000" when "00010101000101101", -- t[10797] = 0
      "0000000" when "00010101000101110", -- t[10798] = 0
      "0000000" when "00010101000101111", -- t[10799] = 0
      "0000000" when "00010101000110000", -- t[10800] = 0
      "0000000" when "00010101000110001", -- t[10801] = 0
      "0000000" when "00010101000110010", -- t[10802] = 0
      "0000000" when "00010101000110011", -- t[10803] = 0
      "0000000" when "00010101000110100", -- t[10804] = 0
      "0000000" when "00010101000110101", -- t[10805] = 0
      "0000000" when "00010101000110110", -- t[10806] = 0
      "0000000" when "00010101000110111", -- t[10807] = 0
      "0000000" when "00010101000111000", -- t[10808] = 0
      "0000000" when "00010101000111001", -- t[10809] = 0
      "0000000" when "00010101000111010", -- t[10810] = 0
      "0000000" when "00010101000111011", -- t[10811] = 0
      "0000000" when "00010101000111100", -- t[10812] = 0
      "0000000" when "00010101000111101", -- t[10813] = 0
      "0000000" when "00010101000111110", -- t[10814] = 0
      "0000000" when "00010101000111111", -- t[10815] = 0
      "0000000" when "00010101001000000", -- t[10816] = 0
      "0000000" when "00010101001000001", -- t[10817] = 0
      "0000000" when "00010101001000010", -- t[10818] = 0
      "0000000" when "00010101001000011", -- t[10819] = 0
      "0000000" when "00010101001000100", -- t[10820] = 0
      "0000000" when "00010101001000101", -- t[10821] = 0
      "0000000" when "00010101001000110", -- t[10822] = 0
      "0000000" when "00010101001000111", -- t[10823] = 0
      "0000000" when "00010101001001000", -- t[10824] = 0
      "0000000" when "00010101001001001", -- t[10825] = 0
      "0000000" when "00010101001001010", -- t[10826] = 0
      "0000000" when "00010101001001011", -- t[10827] = 0
      "0000000" when "00010101001001100", -- t[10828] = 0
      "0000000" when "00010101001001101", -- t[10829] = 0
      "0000000" when "00010101001001110", -- t[10830] = 0
      "0000000" when "00010101001001111", -- t[10831] = 0
      "0000000" when "00010101001010000", -- t[10832] = 0
      "0000000" when "00010101001010001", -- t[10833] = 0
      "0000000" when "00010101001010010", -- t[10834] = 0
      "0000000" when "00010101001010011", -- t[10835] = 0
      "0000000" when "00010101001010100", -- t[10836] = 0
      "0000000" when "00010101001010101", -- t[10837] = 0
      "0000000" when "00010101001010110", -- t[10838] = 0
      "0000000" when "00010101001010111", -- t[10839] = 0
      "0000000" when "00010101001011000", -- t[10840] = 0
      "0000000" when "00010101001011001", -- t[10841] = 0
      "0000000" when "00010101001011010", -- t[10842] = 0
      "0000000" when "00010101001011011", -- t[10843] = 0
      "0000000" when "00010101001011100", -- t[10844] = 0
      "0000000" when "00010101001011101", -- t[10845] = 0
      "0000000" when "00010101001011110", -- t[10846] = 0
      "0000000" when "00010101001011111", -- t[10847] = 0
      "0000000" when "00010101001100000", -- t[10848] = 0
      "0000000" when "00010101001100001", -- t[10849] = 0
      "0000000" when "00010101001100010", -- t[10850] = 0
      "0000000" when "00010101001100011", -- t[10851] = 0
      "0000000" when "00010101001100100", -- t[10852] = 0
      "0000000" when "00010101001100101", -- t[10853] = 0
      "0000000" when "00010101001100110", -- t[10854] = 0
      "0000000" when "00010101001100111", -- t[10855] = 0
      "0000000" when "00010101001101000", -- t[10856] = 0
      "0000000" when "00010101001101001", -- t[10857] = 0
      "0000000" when "00010101001101010", -- t[10858] = 0
      "0000000" when "00010101001101011", -- t[10859] = 0
      "0000000" when "00010101001101100", -- t[10860] = 0
      "0000000" when "00010101001101101", -- t[10861] = 0
      "0000000" when "00010101001101110", -- t[10862] = 0
      "0000000" when "00010101001101111", -- t[10863] = 0
      "0000000" when "00010101001110000", -- t[10864] = 0
      "0000000" when "00010101001110001", -- t[10865] = 0
      "0000000" when "00010101001110010", -- t[10866] = 0
      "0000000" when "00010101001110011", -- t[10867] = 0
      "0000000" when "00010101001110100", -- t[10868] = 0
      "0000000" when "00010101001110101", -- t[10869] = 0
      "0000000" when "00010101001110110", -- t[10870] = 0
      "0000000" when "00010101001110111", -- t[10871] = 0
      "0000000" when "00010101001111000", -- t[10872] = 0
      "0000000" when "00010101001111001", -- t[10873] = 0
      "0000000" when "00010101001111010", -- t[10874] = 0
      "0000000" when "00010101001111011", -- t[10875] = 0
      "0000000" when "00010101001111100", -- t[10876] = 0
      "0000000" when "00010101001111101", -- t[10877] = 0
      "0000000" when "00010101001111110", -- t[10878] = 0
      "0000000" when "00010101001111111", -- t[10879] = 0
      "0000000" when "00010101010000000", -- t[10880] = 0
      "0000000" when "00010101010000001", -- t[10881] = 0
      "0000000" when "00010101010000010", -- t[10882] = 0
      "0000000" when "00010101010000011", -- t[10883] = 0
      "0000000" when "00010101010000100", -- t[10884] = 0
      "0000000" when "00010101010000101", -- t[10885] = 0
      "0000000" when "00010101010000110", -- t[10886] = 0
      "0000000" when "00010101010000111", -- t[10887] = 0
      "0000000" when "00010101010001000", -- t[10888] = 0
      "0000000" when "00010101010001001", -- t[10889] = 0
      "0000000" when "00010101010001010", -- t[10890] = 0
      "0000000" when "00010101010001011", -- t[10891] = 0
      "0000000" when "00010101010001100", -- t[10892] = 0
      "0000000" when "00010101010001101", -- t[10893] = 0
      "0000000" when "00010101010001110", -- t[10894] = 0
      "0000000" when "00010101010001111", -- t[10895] = 0
      "0000000" when "00010101010010000", -- t[10896] = 0
      "0000000" when "00010101010010001", -- t[10897] = 0
      "0000000" when "00010101010010010", -- t[10898] = 0
      "0000000" when "00010101010010011", -- t[10899] = 0
      "0000000" when "00010101010010100", -- t[10900] = 0
      "0000000" when "00010101010010101", -- t[10901] = 0
      "0000000" when "00010101010010110", -- t[10902] = 0
      "0000000" when "00010101010010111", -- t[10903] = 0
      "0000000" when "00010101010011000", -- t[10904] = 0
      "0000000" when "00010101010011001", -- t[10905] = 0
      "0000000" when "00010101010011010", -- t[10906] = 0
      "0000000" when "00010101010011011", -- t[10907] = 0
      "0000000" when "00010101010011100", -- t[10908] = 0
      "0000000" when "00010101010011101", -- t[10909] = 0
      "0000000" when "00010101010011110", -- t[10910] = 0
      "0000000" when "00010101010011111", -- t[10911] = 0
      "0000000" when "00010101010100000", -- t[10912] = 0
      "0000000" when "00010101010100001", -- t[10913] = 0
      "0000000" when "00010101010100010", -- t[10914] = 0
      "0000000" when "00010101010100011", -- t[10915] = 0
      "0000000" when "00010101010100100", -- t[10916] = 0
      "0000000" when "00010101010100101", -- t[10917] = 0
      "0000000" when "00010101010100110", -- t[10918] = 0
      "0000000" when "00010101010100111", -- t[10919] = 0
      "0000000" when "00010101010101000", -- t[10920] = 0
      "0000000" when "00010101010101001", -- t[10921] = 0
      "0000000" when "00010101010101010", -- t[10922] = 0
      "0000000" when "00010101010101011", -- t[10923] = 0
      "0000000" when "00010101010101100", -- t[10924] = 0
      "0000000" when "00010101010101101", -- t[10925] = 0
      "0000000" when "00010101010101110", -- t[10926] = 0
      "0000000" when "00010101010101111", -- t[10927] = 0
      "0000000" when "00010101010110000", -- t[10928] = 0
      "0000000" when "00010101010110001", -- t[10929] = 0
      "0000000" when "00010101010110010", -- t[10930] = 0
      "0000000" when "00010101010110011", -- t[10931] = 0
      "0000000" when "00010101010110100", -- t[10932] = 0
      "0000000" when "00010101010110101", -- t[10933] = 0
      "0000000" when "00010101010110110", -- t[10934] = 0
      "0000000" when "00010101010110111", -- t[10935] = 0
      "0000000" when "00010101010111000", -- t[10936] = 0
      "0000000" when "00010101010111001", -- t[10937] = 0
      "0000000" when "00010101010111010", -- t[10938] = 0
      "0000000" when "00010101010111011", -- t[10939] = 0
      "0000000" when "00010101010111100", -- t[10940] = 0
      "0000000" when "00010101010111101", -- t[10941] = 0
      "0000000" when "00010101010111110", -- t[10942] = 0
      "0000000" when "00010101010111111", -- t[10943] = 0
      "0000000" when "00010101011000000", -- t[10944] = 0
      "0000000" when "00010101011000001", -- t[10945] = 0
      "0000000" when "00010101011000010", -- t[10946] = 0
      "0000000" when "00010101011000011", -- t[10947] = 0
      "0000000" when "00010101011000100", -- t[10948] = 0
      "0000000" when "00010101011000101", -- t[10949] = 0
      "0000000" when "00010101011000110", -- t[10950] = 0
      "0000000" when "00010101011000111", -- t[10951] = 0
      "0000000" when "00010101011001000", -- t[10952] = 0
      "0000000" when "00010101011001001", -- t[10953] = 0
      "0000000" when "00010101011001010", -- t[10954] = 0
      "0000000" when "00010101011001011", -- t[10955] = 0
      "0000000" when "00010101011001100", -- t[10956] = 0
      "0000000" when "00010101011001101", -- t[10957] = 0
      "0000000" when "00010101011001110", -- t[10958] = 0
      "0000000" when "00010101011001111", -- t[10959] = 0
      "0000000" when "00010101011010000", -- t[10960] = 0
      "0000000" when "00010101011010001", -- t[10961] = 0
      "0000000" when "00010101011010010", -- t[10962] = 0
      "0000000" when "00010101011010011", -- t[10963] = 0
      "0000000" when "00010101011010100", -- t[10964] = 0
      "0000000" when "00010101011010101", -- t[10965] = 0
      "0000000" when "00010101011010110", -- t[10966] = 0
      "0000000" when "00010101011010111", -- t[10967] = 0
      "0000000" when "00010101011011000", -- t[10968] = 0
      "0000000" when "00010101011011001", -- t[10969] = 0
      "0000000" when "00010101011011010", -- t[10970] = 0
      "0000000" when "00010101011011011", -- t[10971] = 0
      "0000000" when "00010101011011100", -- t[10972] = 0
      "0000000" when "00010101011011101", -- t[10973] = 0
      "0000000" when "00010101011011110", -- t[10974] = 0
      "0000000" when "00010101011011111", -- t[10975] = 0
      "0000000" when "00010101011100000", -- t[10976] = 0
      "0000000" when "00010101011100001", -- t[10977] = 0
      "0000000" when "00010101011100010", -- t[10978] = 0
      "0000000" when "00010101011100011", -- t[10979] = 0
      "0000000" when "00010101011100100", -- t[10980] = 0
      "0000000" when "00010101011100101", -- t[10981] = 0
      "0000000" when "00010101011100110", -- t[10982] = 0
      "0000000" when "00010101011100111", -- t[10983] = 0
      "0000000" when "00010101011101000", -- t[10984] = 0
      "0000000" when "00010101011101001", -- t[10985] = 0
      "0000000" when "00010101011101010", -- t[10986] = 0
      "0000000" when "00010101011101011", -- t[10987] = 0
      "0000000" when "00010101011101100", -- t[10988] = 0
      "0000000" when "00010101011101101", -- t[10989] = 0
      "0000000" when "00010101011101110", -- t[10990] = 0
      "0000000" when "00010101011101111", -- t[10991] = 0
      "0000000" when "00010101011110000", -- t[10992] = 0
      "0000000" when "00010101011110001", -- t[10993] = 0
      "0000000" when "00010101011110010", -- t[10994] = 0
      "0000000" when "00010101011110011", -- t[10995] = 0
      "0000000" when "00010101011110100", -- t[10996] = 0
      "0000000" when "00010101011110101", -- t[10997] = 0
      "0000000" when "00010101011110110", -- t[10998] = 0
      "0000000" when "00010101011110111", -- t[10999] = 0
      "0000000" when "00010101011111000", -- t[11000] = 0
      "0000000" when "00010101011111001", -- t[11001] = 0
      "0000000" when "00010101011111010", -- t[11002] = 0
      "0000000" when "00010101011111011", -- t[11003] = 0
      "0000000" when "00010101011111100", -- t[11004] = 0
      "0000000" when "00010101011111101", -- t[11005] = 0
      "0000000" when "00010101011111110", -- t[11006] = 0
      "0000000" when "00010101011111111", -- t[11007] = 0
      "0000000" when "00010101100000000", -- t[11008] = 0
      "0000000" when "00010101100000001", -- t[11009] = 0
      "0000000" when "00010101100000010", -- t[11010] = 0
      "0000000" when "00010101100000011", -- t[11011] = 0
      "0000000" when "00010101100000100", -- t[11012] = 0
      "0000000" when "00010101100000101", -- t[11013] = 0
      "0000000" when "00010101100000110", -- t[11014] = 0
      "0000000" when "00010101100000111", -- t[11015] = 0
      "0000000" when "00010101100001000", -- t[11016] = 0
      "0000000" when "00010101100001001", -- t[11017] = 0
      "0000000" when "00010101100001010", -- t[11018] = 0
      "0000000" when "00010101100001011", -- t[11019] = 0
      "0000000" when "00010101100001100", -- t[11020] = 0
      "0000000" when "00010101100001101", -- t[11021] = 0
      "0000000" when "00010101100001110", -- t[11022] = 0
      "0000000" when "00010101100001111", -- t[11023] = 0
      "0000000" when "00010101100010000", -- t[11024] = 0
      "0000000" when "00010101100010001", -- t[11025] = 0
      "0000000" when "00010101100010010", -- t[11026] = 0
      "0000000" when "00010101100010011", -- t[11027] = 0
      "0000000" when "00010101100010100", -- t[11028] = 0
      "0000000" when "00010101100010101", -- t[11029] = 0
      "0000000" when "00010101100010110", -- t[11030] = 0
      "0000000" when "00010101100010111", -- t[11031] = 0
      "0000000" when "00010101100011000", -- t[11032] = 0
      "0000000" when "00010101100011001", -- t[11033] = 0
      "0000000" when "00010101100011010", -- t[11034] = 0
      "0000000" when "00010101100011011", -- t[11035] = 0
      "0000000" when "00010101100011100", -- t[11036] = 0
      "0000000" when "00010101100011101", -- t[11037] = 0
      "0000000" when "00010101100011110", -- t[11038] = 0
      "0000000" when "00010101100011111", -- t[11039] = 0
      "0000000" when "00010101100100000", -- t[11040] = 0
      "0000000" when "00010101100100001", -- t[11041] = 0
      "0000000" when "00010101100100010", -- t[11042] = 0
      "0000000" when "00010101100100011", -- t[11043] = 0
      "0000000" when "00010101100100100", -- t[11044] = 0
      "0000000" when "00010101100100101", -- t[11045] = 0
      "0000000" when "00010101100100110", -- t[11046] = 0
      "0000000" when "00010101100100111", -- t[11047] = 0
      "0000000" when "00010101100101000", -- t[11048] = 0
      "0000000" when "00010101100101001", -- t[11049] = 0
      "0000000" when "00010101100101010", -- t[11050] = 0
      "0000000" when "00010101100101011", -- t[11051] = 0
      "0000000" when "00010101100101100", -- t[11052] = 0
      "0000000" when "00010101100101101", -- t[11053] = 0
      "0000000" when "00010101100101110", -- t[11054] = 0
      "0000000" when "00010101100101111", -- t[11055] = 0
      "0000000" when "00010101100110000", -- t[11056] = 0
      "0000000" when "00010101100110001", -- t[11057] = 0
      "0000000" when "00010101100110010", -- t[11058] = 0
      "0000000" when "00010101100110011", -- t[11059] = 0
      "0000000" when "00010101100110100", -- t[11060] = 0
      "0000000" when "00010101100110101", -- t[11061] = 0
      "0000000" when "00010101100110110", -- t[11062] = 0
      "0000000" when "00010101100110111", -- t[11063] = 0
      "0000000" when "00010101100111000", -- t[11064] = 0
      "0000000" when "00010101100111001", -- t[11065] = 0
      "0000000" when "00010101100111010", -- t[11066] = 0
      "0000000" when "00010101100111011", -- t[11067] = 0
      "0000000" when "00010101100111100", -- t[11068] = 0
      "0000000" when "00010101100111101", -- t[11069] = 0
      "0000000" when "00010101100111110", -- t[11070] = 0
      "0000000" when "00010101100111111", -- t[11071] = 0
      "0000000" when "00010101101000000", -- t[11072] = 0
      "0000000" when "00010101101000001", -- t[11073] = 0
      "0000000" when "00010101101000010", -- t[11074] = 0
      "0000000" when "00010101101000011", -- t[11075] = 0
      "0000000" when "00010101101000100", -- t[11076] = 0
      "0000000" when "00010101101000101", -- t[11077] = 0
      "0000000" when "00010101101000110", -- t[11078] = 0
      "0000000" when "00010101101000111", -- t[11079] = 0
      "0000000" when "00010101101001000", -- t[11080] = 0
      "0000000" when "00010101101001001", -- t[11081] = 0
      "0000000" when "00010101101001010", -- t[11082] = 0
      "0000000" when "00010101101001011", -- t[11083] = 0
      "0000000" when "00010101101001100", -- t[11084] = 0
      "0000000" when "00010101101001101", -- t[11085] = 0
      "0000000" when "00010101101001110", -- t[11086] = 0
      "0000000" when "00010101101001111", -- t[11087] = 0
      "0000000" when "00010101101010000", -- t[11088] = 0
      "0000000" when "00010101101010001", -- t[11089] = 0
      "0000000" when "00010101101010010", -- t[11090] = 0
      "0000000" when "00010101101010011", -- t[11091] = 0
      "0000000" when "00010101101010100", -- t[11092] = 0
      "0000000" when "00010101101010101", -- t[11093] = 0
      "0000000" when "00010101101010110", -- t[11094] = 0
      "0000000" when "00010101101010111", -- t[11095] = 0
      "0000000" when "00010101101011000", -- t[11096] = 0
      "0000000" when "00010101101011001", -- t[11097] = 0
      "0000000" when "00010101101011010", -- t[11098] = 0
      "0000000" when "00010101101011011", -- t[11099] = 0
      "0000000" when "00010101101011100", -- t[11100] = 0
      "0000000" when "00010101101011101", -- t[11101] = 0
      "0000000" when "00010101101011110", -- t[11102] = 0
      "0000000" when "00010101101011111", -- t[11103] = 0
      "0000000" when "00010101101100000", -- t[11104] = 0
      "0000000" when "00010101101100001", -- t[11105] = 0
      "0000000" when "00010101101100010", -- t[11106] = 0
      "0000000" when "00010101101100011", -- t[11107] = 0
      "0000000" when "00010101101100100", -- t[11108] = 0
      "0000000" when "00010101101100101", -- t[11109] = 0
      "0000000" when "00010101101100110", -- t[11110] = 0
      "0000000" when "00010101101100111", -- t[11111] = 0
      "0000000" when "00010101101101000", -- t[11112] = 0
      "0000000" when "00010101101101001", -- t[11113] = 0
      "0000000" when "00010101101101010", -- t[11114] = 0
      "0000000" when "00010101101101011", -- t[11115] = 0
      "0000000" when "00010101101101100", -- t[11116] = 0
      "0000000" when "00010101101101101", -- t[11117] = 0
      "0000000" when "00010101101101110", -- t[11118] = 0
      "0000000" when "00010101101101111", -- t[11119] = 0
      "0000000" when "00010101101110000", -- t[11120] = 0
      "0000000" when "00010101101110001", -- t[11121] = 0
      "0000000" when "00010101101110010", -- t[11122] = 0
      "0000000" when "00010101101110011", -- t[11123] = 0
      "0000000" when "00010101101110100", -- t[11124] = 0
      "0000000" when "00010101101110101", -- t[11125] = 0
      "0000000" when "00010101101110110", -- t[11126] = 0
      "0000000" when "00010101101110111", -- t[11127] = 0
      "0000000" when "00010101101111000", -- t[11128] = 0
      "0000000" when "00010101101111001", -- t[11129] = 0
      "0000000" when "00010101101111010", -- t[11130] = 0
      "0000000" when "00010101101111011", -- t[11131] = 0
      "0000000" when "00010101101111100", -- t[11132] = 0
      "0000000" when "00010101101111101", -- t[11133] = 0
      "0000000" when "00010101101111110", -- t[11134] = 0
      "0000000" when "00010101101111111", -- t[11135] = 0
      "0000000" when "00010101110000000", -- t[11136] = 0
      "0000000" when "00010101110000001", -- t[11137] = 0
      "0000000" when "00010101110000010", -- t[11138] = 0
      "0000000" when "00010101110000011", -- t[11139] = 0
      "0000000" when "00010101110000100", -- t[11140] = 0
      "0000000" when "00010101110000101", -- t[11141] = 0
      "0000000" when "00010101110000110", -- t[11142] = 0
      "0000000" when "00010101110000111", -- t[11143] = 0
      "0000000" when "00010101110001000", -- t[11144] = 0
      "0000000" when "00010101110001001", -- t[11145] = 0
      "0000000" when "00010101110001010", -- t[11146] = 0
      "0000000" when "00010101110001011", -- t[11147] = 0
      "0000000" when "00010101110001100", -- t[11148] = 0
      "0000000" when "00010101110001101", -- t[11149] = 0
      "0000000" when "00010101110001110", -- t[11150] = 0
      "0000000" when "00010101110001111", -- t[11151] = 0
      "0000000" when "00010101110010000", -- t[11152] = 0
      "0000000" when "00010101110010001", -- t[11153] = 0
      "0000000" when "00010101110010010", -- t[11154] = 0
      "0000000" when "00010101110010011", -- t[11155] = 0
      "0000000" when "00010101110010100", -- t[11156] = 0
      "0000000" when "00010101110010101", -- t[11157] = 0
      "0000000" when "00010101110010110", -- t[11158] = 0
      "0000000" when "00010101110010111", -- t[11159] = 0
      "0000000" when "00010101110011000", -- t[11160] = 0
      "0000000" when "00010101110011001", -- t[11161] = 0
      "0000000" when "00010101110011010", -- t[11162] = 0
      "0000000" when "00010101110011011", -- t[11163] = 0
      "0000000" when "00010101110011100", -- t[11164] = 0
      "0000000" when "00010101110011101", -- t[11165] = 0
      "0000000" when "00010101110011110", -- t[11166] = 0
      "0000000" when "00010101110011111", -- t[11167] = 0
      "0000000" when "00010101110100000", -- t[11168] = 0
      "0000000" when "00010101110100001", -- t[11169] = 0
      "0000000" when "00010101110100010", -- t[11170] = 0
      "0000000" when "00010101110100011", -- t[11171] = 0
      "0000000" when "00010101110100100", -- t[11172] = 0
      "0000000" when "00010101110100101", -- t[11173] = 0
      "0000000" when "00010101110100110", -- t[11174] = 0
      "0000000" when "00010101110100111", -- t[11175] = 0
      "0000000" when "00010101110101000", -- t[11176] = 0
      "0000000" when "00010101110101001", -- t[11177] = 0
      "0000000" when "00010101110101010", -- t[11178] = 0
      "0000000" when "00010101110101011", -- t[11179] = 0
      "0000000" when "00010101110101100", -- t[11180] = 0
      "0000000" when "00010101110101101", -- t[11181] = 0
      "0000000" when "00010101110101110", -- t[11182] = 0
      "0000000" when "00010101110101111", -- t[11183] = 0
      "0000000" when "00010101110110000", -- t[11184] = 0
      "0000000" when "00010101110110001", -- t[11185] = 0
      "0000000" when "00010101110110010", -- t[11186] = 0
      "0000000" when "00010101110110011", -- t[11187] = 0
      "0000000" when "00010101110110100", -- t[11188] = 0
      "0000000" when "00010101110110101", -- t[11189] = 0
      "0000000" when "00010101110110110", -- t[11190] = 0
      "0000000" when "00010101110110111", -- t[11191] = 0
      "0000000" when "00010101110111000", -- t[11192] = 0
      "0000000" when "00010101110111001", -- t[11193] = 0
      "0000000" when "00010101110111010", -- t[11194] = 0
      "0000000" when "00010101110111011", -- t[11195] = 0
      "0000000" when "00010101110111100", -- t[11196] = 0
      "0000000" when "00010101110111101", -- t[11197] = 0
      "0000000" when "00010101110111110", -- t[11198] = 0
      "0000000" when "00010101110111111", -- t[11199] = 0
      "0000000" when "00010101111000000", -- t[11200] = 0
      "0000000" when "00010101111000001", -- t[11201] = 0
      "0000000" when "00010101111000010", -- t[11202] = 0
      "0000000" when "00010101111000011", -- t[11203] = 0
      "0000000" when "00010101111000100", -- t[11204] = 0
      "0000000" when "00010101111000101", -- t[11205] = 0
      "0000000" when "00010101111000110", -- t[11206] = 0
      "0000000" when "00010101111000111", -- t[11207] = 0
      "0000000" when "00010101111001000", -- t[11208] = 0
      "0000000" when "00010101111001001", -- t[11209] = 0
      "0000000" when "00010101111001010", -- t[11210] = 0
      "0000000" when "00010101111001011", -- t[11211] = 0
      "0000000" when "00010101111001100", -- t[11212] = 0
      "0000000" when "00010101111001101", -- t[11213] = 0
      "0000000" when "00010101111001110", -- t[11214] = 0
      "0000000" when "00010101111001111", -- t[11215] = 0
      "0000000" when "00010101111010000", -- t[11216] = 0
      "0000000" when "00010101111010001", -- t[11217] = 0
      "0000000" when "00010101111010010", -- t[11218] = 0
      "0000000" when "00010101111010011", -- t[11219] = 0
      "0000000" when "00010101111010100", -- t[11220] = 0
      "0000000" when "00010101111010101", -- t[11221] = 0
      "0000000" when "00010101111010110", -- t[11222] = 0
      "0000000" when "00010101111010111", -- t[11223] = 0
      "0000000" when "00010101111011000", -- t[11224] = 0
      "0000000" when "00010101111011001", -- t[11225] = 0
      "0000000" when "00010101111011010", -- t[11226] = 0
      "0000000" when "00010101111011011", -- t[11227] = 0
      "0000000" when "00010101111011100", -- t[11228] = 0
      "0000000" when "00010101111011101", -- t[11229] = 0
      "0000000" when "00010101111011110", -- t[11230] = 0
      "0000000" when "00010101111011111", -- t[11231] = 0
      "0000000" when "00010101111100000", -- t[11232] = 0
      "0000000" when "00010101111100001", -- t[11233] = 0
      "0000000" when "00010101111100010", -- t[11234] = 0
      "0000000" when "00010101111100011", -- t[11235] = 0
      "0000000" when "00010101111100100", -- t[11236] = 0
      "0000000" when "00010101111100101", -- t[11237] = 0
      "0000000" when "00010101111100110", -- t[11238] = 0
      "0000000" when "00010101111100111", -- t[11239] = 0
      "0000000" when "00010101111101000", -- t[11240] = 0
      "0000000" when "00010101111101001", -- t[11241] = 0
      "0000000" when "00010101111101010", -- t[11242] = 0
      "0000000" when "00010101111101011", -- t[11243] = 0
      "0000000" when "00010101111101100", -- t[11244] = 0
      "0000000" when "00010101111101101", -- t[11245] = 0
      "0000000" when "00010101111101110", -- t[11246] = 0
      "0000000" when "00010101111101111", -- t[11247] = 0
      "0000000" when "00010101111110000", -- t[11248] = 0
      "0000000" when "00010101111110001", -- t[11249] = 0
      "0000000" when "00010101111110010", -- t[11250] = 0
      "0000000" when "00010101111110011", -- t[11251] = 0
      "0000000" when "00010101111110100", -- t[11252] = 0
      "0000000" when "00010101111110101", -- t[11253] = 0
      "0000000" when "00010101111110110", -- t[11254] = 0
      "0000000" when "00010101111110111", -- t[11255] = 0
      "0000000" when "00010101111111000", -- t[11256] = 0
      "0000000" when "00010101111111001", -- t[11257] = 0
      "0000000" when "00010101111111010", -- t[11258] = 0
      "0000000" when "00010101111111011", -- t[11259] = 0
      "0000000" when "00010101111111100", -- t[11260] = 0
      "0000000" when "00010101111111101", -- t[11261] = 0
      "0000000" when "00010101111111110", -- t[11262] = 0
      "0000000" when "00010101111111111", -- t[11263] = 0
      "0000000" when "00010110000000000", -- t[11264] = 0
      "0000000" when "00010110000000001", -- t[11265] = 0
      "0000000" when "00010110000000010", -- t[11266] = 0
      "0000000" when "00010110000000011", -- t[11267] = 0
      "0000000" when "00010110000000100", -- t[11268] = 0
      "0000000" when "00010110000000101", -- t[11269] = 0
      "0000000" when "00010110000000110", -- t[11270] = 0
      "0000000" when "00010110000000111", -- t[11271] = 0
      "0000000" when "00010110000001000", -- t[11272] = 0
      "0000000" when "00010110000001001", -- t[11273] = 0
      "0000000" when "00010110000001010", -- t[11274] = 0
      "0000000" when "00010110000001011", -- t[11275] = 0
      "0000000" when "00010110000001100", -- t[11276] = 0
      "0000000" when "00010110000001101", -- t[11277] = 0
      "0000000" when "00010110000001110", -- t[11278] = 0
      "0000000" when "00010110000001111", -- t[11279] = 0
      "0000000" when "00010110000010000", -- t[11280] = 0
      "0000000" when "00010110000010001", -- t[11281] = 0
      "0000000" when "00010110000010010", -- t[11282] = 0
      "0000000" when "00010110000010011", -- t[11283] = 0
      "0000000" when "00010110000010100", -- t[11284] = 0
      "0000000" when "00010110000010101", -- t[11285] = 0
      "0000000" when "00010110000010110", -- t[11286] = 0
      "0000000" when "00010110000010111", -- t[11287] = 0
      "0000000" when "00010110000011000", -- t[11288] = 0
      "0000000" when "00010110000011001", -- t[11289] = 0
      "0000000" when "00010110000011010", -- t[11290] = 0
      "0000000" when "00010110000011011", -- t[11291] = 0
      "0000000" when "00010110000011100", -- t[11292] = 0
      "0000000" when "00010110000011101", -- t[11293] = 0
      "0000000" when "00010110000011110", -- t[11294] = 0
      "0000000" when "00010110000011111", -- t[11295] = 0
      "0000000" when "00010110000100000", -- t[11296] = 0
      "0000000" when "00010110000100001", -- t[11297] = 0
      "0000000" when "00010110000100010", -- t[11298] = 0
      "0000000" when "00010110000100011", -- t[11299] = 0
      "0000000" when "00010110000100100", -- t[11300] = 0
      "0000000" when "00010110000100101", -- t[11301] = 0
      "0000000" when "00010110000100110", -- t[11302] = 0
      "0000000" when "00010110000100111", -- t[11303] = 0
      "0000000" when "00010110000101000", -- t[11304] = 0
      "0000000" when "00010110000101001", -- t[11305] = 0
      "0000000" when "00010110000101010", -- t[11306] = 0
      "0000000" when "00010110000101011", -- t[11307] = 0
      "0000000" when "00010110000101100", -- t[11308] = 0
      "0000000" when "00010110000101101", -- t[11309] = 0
      "0000000" when "00010110000101110", -- t[11310] = 0
      "0000000" when "00010110000101111", -- t[11311] = 0
      "0000000" when "00010110000110000", -- t[11312] = 0
      "0000000" when "00010110000110001", -- t[11313] = 0
      "0000000" when "00010110000110010", -- t[11314] = 0
      "0000000" when "00010110000110011", -- t[11315] = 0
      "0000000" when "00010110000110100", -- t[11316] = 0
      "0000000" when "00010110000110101", -- t[11317] = 0
      "0000000" when "00010110000110110", -- t[11318] = 0
      "0000000" when "00010110000110111", -- t[11319] = 0
      "0000000" when "00010110000111000", -- t[11320] = 0
      "0000000" when "00010110000111001", -- t[11321] = 0
      "0000000" when "00010110000111010", -- t[11322] = 0
      "0000000" when "00010110000111011", -- t[11323] = 0
      "0000000" when "00010110000111100", -- t[11324] = 0
      "0000000" when "00010110000111101", -- t[11325] = 0
      "0000000" when "00010110000111110", -- t[11326] = 0
      "0000000" when "00010110000111111", -- t[11327] = 0
      "0000000" when "00010110001000000", -- t[11328] = 0
      "0000000" when "00010110001000001", -- t[11329] = 0
      "0000000" when "00010110001000010", -- t[11330] = 0
      "0000000" when "00010110001000011", -- t[11331] = 0
      "0000000" when "00010110001000100", -- t[11332] = 0
      "0000000" when "00010110001000101", -- t[11333] = 0
      "0000000" when "00010110001000110", -- t[11334] = 0
      "0000000" when "00010110001000111", -- t[11335] = 0
      "0000000" when "00010110001001000", -- t[11336] = 0
      "0000000" when "00010110001001001", -- t[11337] = 0
      "0000000" when "00010110001001010", -- t[11338] = 0
      "0000000" when "00010110001001011", -- t[11339] = 0
      "0000000" when "00010110001001100", -- t[11340] = 0
      "0000000" when "00010110001001101", -- t[11341] = 0
      "0000000" when "00010110001001110", -- t[11342] = 0
      "0000000" when "00010110001001111", -- t[11343] = 0
      "0000000" when "00010110001010000", -- t[11344] = 0
      "0000000" when "00010110001010001", -- t[11345] = 0
      "0000000" when "00010110001010010", -- t[11346] = 0
      "0000000" when "00010110001010011", -- t[11347] = 0
      "0000000" when "00010110001010100", -- t[11348] = 0
      "0000000" when "00010110001010101", -- t[11349] = 0
      "0000000" when "00010110001010110", -- t[11350] = 0
      "0000000" when "00010110001010111", -- t[11351] = 0
      "0000000" when "00010110001011000", -- t[11352] = 0
      "0000000" when "00010110001011001", -- t[11353] = 0
      "0000000" when "00010110001011010", -- t[11354] = 0
      "0000000" when "00010110001011011", -- t[11355] = 0
      "0000000" when "00010110001011100", -- t[11356] = 0
      "0000000" when "00010110001011101", -- t[11357] = 0
      "0000000" when "00010110001011110", -- t[11358] = 0
      "0000000" when "00010110001011111", -- t[11359] = 0
      "0000000" when "00010110001100000", -- t[11360] = 0
      "0000000" when "00010110001100001", -- t[11361] = 0
      "0000000" when "00010110001100010", -- t[11362] = 0
      "0000000" when "00010110001100011", -- t[11363] = 0
      "0000000" when "00010110001100100", -- t[11364] = 0
      "0000000" when "00010110001100101", -- t[11365] = 0
      "0000000" when "00010110001100110", -- t[11366] = 0
      "0000000" when "00010110001100111", -- t[11367] = 0
      "0000000" when "00010110001101000", -- t[11368] = 0
      "0000000" when "00010110001101001", -- t[11369] = 0
      "0000000" when "00010110001101010", -- t[11370] = 0
      "0000000" when "00010110001101011", -- t[11371] = 0
      "0000000" when "00010110001101100", -- t[11372] = 0
      "0000000" when "00010110001101101", -- t[11373] = 0
      "0000000" when "00010110001101110", -- t[11374] = 0
      "0000000" when "00010110001101111", -- t[11375] = 0
      "0000000" when "00010110001110000", -- t[11376] = 0
      "0000000" when "00010110001110001", -- t[11377] = 0
      "0000000" when "00010110001110010", -- t[11378] = 0
      "0000000" when "00010110001110011", -- t[11379] = 0
      "0000000" when "00010110001110100", -- t[11380] = 0
      "0000000" when "00010110001110101", -- t[11381] = 0
      "0000000" when "00010110001110110", -- t[11382] = 0
      "0000000" when "00010110001110111", -- t[11383] = 0
      "0000000" when "00010110001111000", -- t[11384] = 0
      "0000000" when "00010110001111001", -- t[11385] = 0
      "0000000" when "00010110001111010", -- t[11386] = 0
      "0000000" when "00010110001111011", -- t[11387] = 0
      "0000000" when "00010110001111100", -- t[11388] = 0
      "0000000" when "00010110001111101", -- t[11389] = 0
      "0000000" when "00010110001111110", -- t[11390] = 0
      "0000000" when "00010110001111111", -- t[11391] = 0
      "0000000" when "00010110010000000", -- t[11392] = 0
      "0000000" when "00010110010000001", -- t[11393] = 0
      "0000000" when "00010110010000010", -- t[11394] = 0
      "0000000" when "00010110010000011", -- t[11395] = 0
      "0000000" when "00010110010000100", -- t[11396] = 0
      "0000000" when "00010110010000101", -- t[11397] = 0
      "0000000" when "00010110010000110", -- t[11398] = 0
      "0000000" when "00010110010000111", -- t[11399] = 0
      "0000000" when "00010110010001000", -- t[11400] = 0
      "0000000" when "00010110010001001", -- t[11401] = 0
      "0000000" when "00010110010001010", -- t[11402] = 0
      "0000000" when "00010110010001011", -- t[11403] = 0
      "0000000" when "00010110010001100", -- t[11404] = 0
      "0000000" when "00010110010001101", -- t[11405] = 0
      "0000000" when "00010110010001110", -- t[11406] = 0
      "0000000" when "00010110010001111", -- t[11407] = 0
      "0000000" when "00010110010010000", -- t[11408] = 0
      "0000000" when "00010110010010001", -- t[11409] = 0
      "0000000" when "00010110010010010", -- t[11410] = 0
      "0000000" when "00010110010010011", -- t[11411] = 0
      "0000000" when "00010110010010100", -- t[11412] = 0
      "0000000" when "00010110010010101", -- t[11413] = 0
      "0000000" when "00010110010010110", -- t[11414] = 0
      "0000000" when "00010110010010111", -- t[11415] = 0
      "0000000" when "00010110010011000", -- t[11416] = 0
      "0000000" when "00010110010011001", -- t[11417] = 0
      "0000000" when "00010110010011010", -- t[11418] = 0
      "0000000" when "00010110010011011", -- t[11419] = 0
      "0000000" when "00010110010011100", -- t[11420] = 0
      "0000000" when "00010110010011101", -- t[11421] = 0
      "0000000" when "00010110010011110", -- t[11422] = 0
      "0000000" when "00010110010011111", -- t[11423] = 0
      "0000000" when "00010110010100000", -- t[11424] = 0
      "0000000" when "00010110010100001", -- t[11425] = 0
      "0000000" when "00010110010100010", -- t[11426] = 0
      "0000000" when "00010110010100011", -- t[11427] = 0
      "0000000" when "00010110010100100", -- t[11428] = 0
      "0000000" when "00010110010100101", -- t[11429] = 0
      "0000000" when "00010110010100110", -- t[11430] = 0
      "0000000" when "00010110010100111", -- t[11431] = 0
      "0000000" when "00010110010101000", -- t[11432] = 0
      "0000000" when "00010110010101001", -- t[11433] = 0
      "0000000" when "00010110010101010", -- t[11434] = 0
      "0000000" when "00010110010101011", -- t[11435] = 0
      "0000000" when "00010110010101100", -- t[11436] = 0
      "0000000" when "00010110010101101", -- t[11437] = 0
      "0000000" when "00010110010101110", -- t[11438] = 0
      "0000000" when "00010110010101111", -- t[11439] = 0
      "0000000" when "00010110010110000", -- t[11440] = 0
      "0000000" when "00010110010110001", -- t[11441] = 0
      "0000000" when "00010110010110010", -- t[11442] = 0
      "0000000" when "00010110010110011", -- t[11443] = 0
      "0000000" when "00010110010110100", -- t[11444] = 0
      "0000000" when "00010110010110101", -- t[11445] = 0
      "0000000" when "00010110010110110", -- t[11446] = 0
      "0000000" when "00010110010110111", -- t[11447] = 0
      "0000000" when "00010110010111000", -- t[11448] = 0
      "0000000" when "00010110010111001", -- t[11449] = 0
      "0000000" when "00010110010111010", -- t[11450] = 0
      "0000000" when "00010110010111011", -- t[11451] = 0
      "0000000" when "00010110010111100", -- t[11452] = 0
      "0000000" when "00010110010111101", -- t[11453] = 0
      "0000000" when "00010110010111110", -- t[11454] = 0
      "0000000" when "00010110010111111", -- t[11455] = 0
      "0000000" when "00010110011000000", -- t[11456] = 0
      "0000000" when "00010110011000001", -- t[11457] = 0
      "0000000" when "00010110011000010", -- t[11458] = 0
      "0000000" when "00010110011000011", -- t[11459] = 0
      "0000000" when "00010110011000100", -- t[11460] = 0
      "0000000" when "00010110011000101", -- t[11461] = 0
      "0000000" when "00010110011000110", -- t[11462] = 0
      "0000000" when "00010110011000111", -- t[11463] = 0
      "0000000" when "00010110011001000", -- t[11464] = 0
      "0000000" when "00010110011001001", -- t[11465] = 0
      "0000000" when "00010110011001010", -- t[11466] = 0
      "0000000" when "00010110011001011", -- t[11467] = 0
      "0000000" when "00010110011001100", -- t[11468] = 0
      "0000000" when "00010110011001101", -- t[11469] = 0
      "0000000" when "00010110011001110", -- t[11470] = 0
      "0000000" when "00010110011001111", -- t[11471] = 0
      "0000000" when "00010110011010000", -- t[11472] = 0
      "0000000" when "00010110011010001", -- t[11473] = 0
      "0000000" when "00010110011010010", -- t[11474] = 0
      "0000000" when "00010110011010011", -- t[11475] = 0
      "0000000" when "00010110011010100", -- t[11476] = 0
      "0000000" when "00010110011010101", -- t[11477] = 0
      "0000000" when "00010110011010110", -- t[11478] = 0
      "0000000" when "00010110011010111", -- t[11479] = 0
      "0000000" when "00010110011011000", -- t[11480] = 0
      "0000000" when "00010110011011001", -- t[11481] = 0
      "0000000" when "00010110011011010", -- t[11482] = 0
      "0000000" when "00010110011011011", -- t[11483] = 0
      "0000000" when "00010110011011100", -- t[11484] = 0
      "0000000" when "00010110011011101", -- t[11485] = 0
      "0000000" when "00010110011011110", -- t[11486] = 0
      "0000000" when "00010110011011111", -- t[11487] = 0
      "0000000" when "00010110011100000", -- t[11488] = 0
      "0000000" when "00010110011100001", -- t[11489] = 0
      "0000000" when "00010110011100010", -- t[11490] = 0
      "0000000" when "00010110011100011", -- t[11491] = 0
      "0000000" when "00010110011100100", -- t[11492] = 0
      "0000000" when "00010110011100101", -- t[11493] = 0
      "0000000" when "00010110011100110", -- t[11494] = 0
      "0000000" when "00010110011100111", -- t[11495] = 0
      "0000000" when "00010110011101000", -- t[11496] = 0
      "0000000" when "00010110011101001", -- t[11497] = 0
      "0000000" when "00010110011101010", -- t[11498] = 0
      "0000000" when "00010110011101011", -- t[11499] = 0
      "0000000" when "00010110011101100", -- t[11500] = 0
      "0000000" when "00010110011101101", -- t[11501] = 0
      "0000000" when "00010110011101110", -- t[11502] = 0
      "0000000" when "00010110011101111", -- t[11503] = 0
      "0000000" when "00010110011110000", -- t[11504] = 0
      "0000000" when "00010110011110001", -- t[11505] = 0
      "0000000" when "00010110011110010", -- t[11506] = 0
      "0000000" when "00010110011110011", -- t[11507] = 0
      "0000000" when "00010110011110100", -- t[11508] = 0
      "0000000" when "00010110011110101", -- t[11509] = 0
      "0000000" when "00010110011110110", -- t[11510] = 0
      "0000000" when "00010110011110111", -- t[11511] = 0
      "0000000" when "00010110011111000", -- t[11512] = 0
      "0000000" when "00010110011111001", -- t[11513] = 0
      "0000000" when "00010110011111010", -- t[11514] = 0
      "0000000" when "00010110011111011", -- t[11515] = 0
      "0000000" when "00010110011111100", -- t[11516] = 0
      "0000000" when "00010110011111101", -- t[11517] = 0
      "0000000" when "00010110011111110", -- t[11518] = 0
      "0000000" when "00010110011111111", -- t[11519] = 0
      "0000000" when "00010110100000000", -- t[11520] = 0
      "0000000" when "00010110100000001", -- t[11521] = 0
      "0000000" when "00010110100000010", -- t[11522] = 0
      "0000000" when "00010110100000011", -- t[11523] = 0
      "0000000" when "00010110100000100", -- t[11524] = 0
      "0000000" when "00010110100000101", -- t[11525] = 0
      "0000000" when "00010110100000110", -- t[11526] = 0
      "0000000" when "00010110100000111", -- t[11527] = 0
      "0000000" when "00010110100001000", -- t[11528] = 0
      "0000000" when "00010110100001001", -- t[11529] = 0
      "0000000" when "00010110100001010", -- t[11530] = 0
      "0000000" when "00010110100001011", -- t[11531] = 0
      "0000000" when "00010110100001100", -- t[11532] = 0
      "0000000" when "00010110100001101", -- t[11533] = 0
      "0000000" when "00010110100001110", -- t[11534] = 0
      "0000000" when "00010110100001111", -- t[11535] = 0
      "0000000" when "00010110100010000", -- t[11536] = 0
      "0000000" when "00010110100010001", -- t[11537] = 0
      "0000000" when "00010110100010010", -- t[11538] = 0
      "0000000" when "00010110100010011", -- t[11539] = 0
      "0000000" when "00010110100010100", -- t[11540] = 0
      "0000000" when "00010110100010101", -- t[11541] = 0
      "0000000" when "00010110100010110", -- t[11542] = 0
      "0000000" when "00010110100010111", -- t[11543] = 0
      "0000000" when "00010110100011000", -- t[11544] = 0
      "0000000" when "00010110100011001", -- t[11545] = 0
      "0000000" when "00010110100011010", -- t[11546] = 0
      "0000000" when "00010110100011011", -- t[11547] = 0
      "0000000" when "00010110100011100", -- t[11548] = 0
      "0000000" when "00010110100011101", -- t[11549] = 0
      "0000000" when "00010110100011110", -- t[11550] = 0
      "0000000" when "00010110100011111", -- t[11551] = 0
      "0000000" when "00010110100100000", -- t[11552] = 0
      "0000000" when "00010110100100001", -- t[11553] = 0
      "0000000" when "00010110100100010", -- t[11554] = 0
      "0000000" when "00010110100100011", -- t[11555] = 0
      "0000000" when "00010110100100100", -- t[11556] = 0
      "0000000" when "00010110100100101", -- t[11557] = 0
      "0000000" when "00010110100100110", -- t[11558] = 0
      "0000000" when "00010110100100111", -- t[11559] = 0
      "0000000" when "00010110100101000", -- t[11560] = 0
      "0000000" when "00010110100101001", -- t[11561] = 0
      "0000000" when "00010110100101010", -- t[11562] = 0
      "0000000" when "00010110100101011", -- t[11563] = 0
      "0000000" when "00010110100101100", -- t[11564] = 0
      "0000000" when "00010110100101101", -- t[11565] = 0
      "0000000" when "00010110100101110", -- t[11566] = 0
      "0000000" when "00010110100101111", -- t[11567] = 0
      "0000000" when "00010110100110000", -- t[11568] = 0
      "0000000" when "00010110100110001", -- t[11569] = 0
      "0000000" when "00010110100110010", -- t[11570] = 0
      "0000000" when "00010110100110011", -- t[11571] = 0
      "0000000" when "00010110100110100", -- t[11572] = 0
      "0000000" when "00010110100110101", -- t[11573] = 0
      "0000000" when "00010110100110110", -- t[11574] = 0
      "0000000" when "00010110100110111", -- t[11575] = 0
      "0000000" when "00010110100111000", -- t[11576] = 0
      "0000000" when "00010110100111001", -- t[11577] = 0
      "0000000" when "00010110100111010", -- t[11578] = 0
      "0000000" when "00010110100111011", -- t[11579] = 0
      "0000000" when "00010110100111100", -- t[11580] = 0
      "0000000" when "00010110100111101", -- t[11581] = 0
      "0000000" when "00010110100111110", -- t[11582] = 0
      "0000000" when "00010110100111111", -- t[11583] = 0
      "0000000" when "00010110101000000", -- t[11584] = 0
      "0000000" when "00010110101000001", -- t[11585] = 0
      "0000000" when "00010110101000010", -- t[11586] = 0
      "0000000" when "00010110101000011", -- t[11587] = 0
      "0000000" when "00010110101000100", -- t[11588] = 0
      "0000000" when "00010110101000101", -- t[11589] = 0
      "0000000" when "00010110101000110", -- t[11590] = 0
      "0000000" when "00010110101000111", -- t[11591] = 0
      "0000000" when "00010110101001000", -- t[11592] = 0
      "0000000" when "00010110101001001", -- t[11593] = 0
      "0000000" when "00010110101001010", -- t[11594] = 0
      "0000000" when "00010110101001011", -- t[11595] = 0
      "0000000" when "00010110101001100", -- t[11596] = 0
      "0000000" when "00010110101001101", -- t[11597] = 0
      "0000000" when "00010110101001110", -- t[11598] = 0
      "0000000" when "00010110101001111", -- t[11599] = 0
      "0000000" when "00010110101010000", -- t[11600] = 0
      "0000000" when "00010110101010001", -- t[11601] = 0
      "0000000" when "00010110101010010", -- t[11602] = 0
      "0000000" when "00010110101010011", -- t[11603] = 0
      "0000000" when "00010110101010100", -- t[11604] = 0
      "0000000" when "00010110101010101", -- t[11605] = 0
      "0000000" when "00010110101010110", -- t[11606] = 0
      "0000000" when "00010110101010111", -- t[11607] = 0
      "0000000" when "00010110101011000", -- t[11608] = 0
      "0000000" when "00010110101011001", -- t[11609] = 0
      "0000000" when "00010110101011010", -- t[11610] = 0
      "0000000" when "00010110101011011", -- t[11611] = 0
      "0000000" when "00010110101011100", -- t[11612] = 0
      "0000000" when "00010110101011101", -- t[11613] = 0
      "0000000" when "00010110101011110", -- t[11614] = 0
      "0000000" when "00010110101011111", -- t[11615] = 0
      "0000000" when "00010110101100000", -- t[11616] = 0
      "0000000" when "00010110101100001", -- t[11617] = 0
      "0000000" when "00010110101100010", -- t[11618] = 0
      "0000000" when "00010110101100011", -- t[11619] = 0
      "0000000" when "00010110101100100", -- t[11620] = 0
      "0000000" when "00010110101100101", -- t[11621] = 0
      "0000000" when "00010110101100110", -- t[11622] = 0
      "0000000" when "00010110101100111", -- t[11623] = 0
      "0000000" when "00010110101101000", -- t[11624] = 0
      "0000000" when "00010110101101001", -- t[11625] = 0
      "0000000" when "00010110101101010", -- t[11626] = 0
      "0000000" when "00010110101101011", -- t[11627] = 0
      "0000000" when "00010110101101100", -- t[11628] = 0
      "0000000" when "00010110101101101", -- t[11629] = 0
      "0000000" when "00010110101101110", -- t[11630] = 0
      "0000000" when "00010110101101111", -- t[11631] = 0
      "0000000" when "00010110101110000", -- t[11632] = 0
      "0000000" when "00010110101110001", -- t[11633] = 0
      "0000000" when "00010110101110010", -- t[11634] = 0
      "0000000" when "00010110101110011", -- t[11635] = 0
      "0000000" when "00010110101110100", -- t[11636] = 0
      "0000000" when "00010110101110101", -- t[11637] = 0
      "0000000" when "00010110101110110", -- t[11638] = 0
      "0000000" when "00010110101110111", -- t[11639] = 0
      "0000000" when "00010110101111000", -- t[11640] = 0
      "0000000" when "00010110101111001", -- t[11641] = 0
      "0000000" when "00010110101111010", -- t[11642] = 0
      "0000000" when "00010110101111011", -- t[11643] = 0
      "0000000" when "00010110101111100", -- t[11644] = 0
      "0000000" when "00010110101111101", -- t[11645] = 0
      "0000000" when "00010110101111110", -- t[11646] = 0
      "0000000" when "00010110101111111", -- t[11647] = 0
      "0000000" when "00010110110000000", -- t[11648] = 0
      "0000000" when "00010110110000001", -- t[11649] = 0
      "0000000" when "00010110110000010", -- t[11650] = 0
      "0000000" when "00010110110000011", -- t[11651] = 0
      "0000000" when "00010110110000100", -- t[11652] = 0
      "0000000" when "00010110110000101", -- t[11653] = 0
      "0000000" when "00010110110000110", -- t[11654] = 0
      "0000000" when "00010110110000111", -- t[11655] = 0
      "0000000" when "00010110110001000", -- t[11656] = 0
      "0000000" when "00010110110001001", -- t[11657] = 0
      "0000000" when "00010110110001010", -- t[11658] = 0
      "0000000" when "00010110110001011", -- t[11659] = 0
      "0000000" when "00010110110001100", -- t[11660] = 0
      "0000000" when "00010110110001101", -- t[11661] = 0
      "0000000" when "00010110110001110", -- t[11662] = 0
      "0000000" when "00010110110001111", -- t[11663] = 0
      "0000000" when "00010110110010000", -- t[11664] = 0
      "0000000" when "00010110110010001", -- t[11665] = 0
      "0000000" when "00010110110010010", -- t[11666] = 0
      "0000000" when "00010110110010011", -- t[11667] = 0
      "0000000" when "00010110110010100", -- t[11668] = 0
      "0000000" when "00010110110010101", -- t[11669] = 0
      "0000000" when "00010110110010110", -- t[11670] = 0
      "0000000" when "00010110110010111", -- t[11671] = 0
      "0000000" when "00010110110011000", -- t[11672] = 0
      "0000000" when "00010110110011001", -- t[11673] = 0
      "0000000" when "00010110110011010", -- t[11674] = 0
      "0000000" when "00010110110011011", -- t[11675] = 0
      "0000000" when "00010110110011100", -- t[11676] = 0
      "0000000" when "00010110110011101", -- t[11677] = 0
      "0000000" when "00010110110011110", -- t[11678] = 0
      "0000000" when "00010110110011111", -- t[11679] = 0
      "0000000" when "00010110110100000", -- t[11680] = 0
      "0000000" when "00010110110100001", -- t[11681] = 0
      "0000000" when "00010110110100010", -- t[11682] = 0
      "0000000" when "00010110110100011", -- t[11683] = 0
      "0000000" when "00010110110100100", -- t[11684] = 0
      "0000000" when "00010110110100101", -- t[11685] = 0
      "0000000" when "00010110110100110", -- t[11686] = 0
      "0000000" when "00010110110100111", -- t[11687] = 0
      "0000000" when "00010110110101000", -- t[11688] = 0
      "0000000" when "00010110110101001", -- t[11689] = 0
      "0000000" when "00010110110101010", -- t[11690] = 0
      "0000000" when "00010110110101011", -- t[11691] = 0
      "0000000" when "00010110110101100", -- t[11692] = 0
      "0000000" when "00010110110101101", -- t[11693] = 0
      "0000000" when "00010110110101110", -- t[11694] = 0
      "0000000" when "00010110110101111", -- t[11695] = 0
      "0000000" when "00010110110110000", -- t[11696] = 0
      "0000000" when "00010110110110001", -- t[11697] = 0
      "0000000" when "00010110110110010", -- t[11698] = 0
      "0000000" when "00010110110110011", -- t[11699] = 0
      "0000000" when "00010110110110100", -- t[11700] = 0
      "0000000" when "00010110110110101", -- t[11701] = 0
      "0000000" when "00010110110110110", -- t[11702] = 0
      "0000000" when "00010110110110111", -- t[11703] = 0
      "0000000" when "00010110110111000", -- t[11704] = 0
      "0000000" when "00010110110111001", -- t[11705] = 0
      "0000000" when "00010110110111010", -- t[11706] = 0
      "0000000" when "00010110110111011", -- t[11707] = 0
      "0000000" when "00010110110111100", -- t[11708] = 0
      "0000000" when "00010110110111101", -- t[11709] = 0
      "0000000" when "00010110110111110", -- t[11710] = 0
      "0000000" when "00010110110111111", -- t[11711] = 0
      "0000000" when "00010110111000000", -- t[11712] = 0
      "0000000" when "00010110111000001", -- t[11713] = 0
      "0000000" when "00010110111000010", -- t[11714] = 0
      "0000000" when "00010110111000011", -- t[11715] = 0
      "0000000" when "00010110111000100", -- t[11716] = 0
      "0000000" when "00010110111000101", -- t[11717] = 0
      "0000000" when "00010110111000110", -- t[11718] = 0
      "0000000" when "00010110111000111", -- t[11719] = 0
      "0000000" when "00010110111001000", -- t[11720] = 0
      "0000000" when "00010110111001001", -- t[11721] = 0
      "0000000" when "00010110111001010", -- t[11722] = 0
      "0000000" when "00010110111001011", -- t[11723] = 0
      "0000000" when "00010110111001100", -- t[11724] = 0
      "0000000" when "00010110111001101", -- t[11725] = 0
      "0000000" when "00010110111001110", -- t[11726] = 0
      "0000000" when "00010110111001111", -- t[11727] = 0
      "0000000" when "00010110111010000", -- t[11728] = 0
      "0000000" when "00010110111010001", -- t[11729] = 0
      "0000000" when "00010110111010010", -- t[11730] = 0
      "0000000" when "00010110111010011", -- t[11731] = 0
      "0000000" when "00010110111010100", -- t[11732] = 0
      "0000000" when "00010110111010101", -- t[11733] = 0
      "0000000" when "00010110111010110", -- t[11734] = 0
      "0000000" when "00010110111010111", -- t[11735] = 0
      "0000000" when "00010110111011000", -- t[11736] = 0
      "0000000" when "00010110111011001", -- t[11737] = 0
      "0000000" when "00010110111011010", -- t[11738] = 0
      "0000000" when "00010110111011011", -- t[11739] = 0
      "0000000" when "00010110111011100", -- t[11740] = 0
      "0000000" when "00010110111011101", -- t[11741] = 0
      "0000000" when "00010110111011110", -- t[11742] = 0
      "0000000" when "00010110111011111", -- t[11743] = 0
      "0000000" when "00010110111100000", -- t[11744] = 0
      "0000000" when "00010110111100001", -- t[11745] = 0
      "0000000" when "00010110111100010", -- t[11746] = 0
      "0000000" when "00010110111100011", -- t[11747] = 0
      "0000000" when "00010110111100100", -- t[11748] = 0
      "0000000" when "00010110111100101", -- t[11749] = 0
      "0000000" when "00010110111100110", -- t[11750] = 0
      "0000000" when "00010110111100111", -- t[11751] = 0
      "0000000" when "00010110111101000", -- t[11752] = 0
      "0000000" when "00010110111101001", -- t[11753] = 0
      "0000000" when "00010110111101010", -- t[11754] = 0
      "0000000" when "00010110111101011", -- t[11755] = 0
      "0000000" when "00010110111101100", -- t[11756] = 0
      "0000000" when "00010110111101101", -- t[11757] = 0
      "0000000" when "00010110111101110", -- t[11758] = 0
      "0000000" when "00010110111101111", -- t[11759] = 0
      "0000000" when "00010110111110000", -- t[11760] = 0
      "0000000" when "00010110111110001", -- t[11761] = 0
      "0000000" when "00010110111110010", -- t[11762] = 0
      "0000000" when "00010110111110011", -- t[11763] = 0
      "0000000" when "00010110111110100", -- t[11764] = 0
      "0000000" when "00010110111110101", -- t[11765] = 0
      "0000000" when "00010110111110110", -- t[11766] = 0
      "0000000" when "00010110111110111", -- t[11767] = 0
      "0000000" when "00010110111111000", -- t[11768] = 0
      "0000000" when "00010110111111001", -- t[11769] = 0
      "0000000" when "00010110111111010", -- t[11770] = 0
      "0000000" when "00010110111111011", -- t[11771] = 0
      "0000000" when "00010110111111100", -- t[11772] = 0
      "0000000" when "00010110111111101", -- t[11773] = 0
      "0000000" when "00010110111111110", -- t[11774] = 0
      "0000000" when "00010110111111111", -- t[11775] = 0
      "0000000" when "00010111000000000", -- t[11776] = 0
      "0000000" when "00010111000000001", -- t[11777] = 0
      "0000000" when "00010111000000010", -- t[11778] = 0
      "0000000" when "00010111000000011", -- t[11779] = 0
      "0000000" when "00010111000000100", -- t[11780] = 0
      "0000000" when "00010111000000101", -- t[11781] = 0
      "0000000" when "00010111000000110", -- t[11782] = 0
      "0000000" when "00010111000000111", -- t[11783] = 0
      "0000000" when "00010111000001000", -- t[11784] = 0
      "0000000" when "00010111000001001", -- t[11785] = 0
      "0000000" when "00010111000001010", -- t[11786] = 0
      "0000000" when "00010111000001011", -- t[11787] = 0
      "0000000" when "00010111000001100", -- t[11788] = 0
      "0000000" when "00010111000001101", -- t[11789] = 0
      "0000000" when "00010111000001110", -- t[11790] = 0
      "0000000" when "00010111000001111", -- t[11791] = 0
      "0000000" when "00010111000010000", -- t[11792] = 0
      "0000000" when "00010111000010001", -- t[11793] = 0
      "0000000" when "00010111000010010", -- t[11794] = 0
      "0000000" when "00010111000010011", -- t[11795] = 0
      "0000000" when "00010111000010100", -- t[11796] = 0
      "0000000" when "00010111000010101", -- t[11797] = 0
      "0000000" when "00010111000010110", -- t[11798] = 0
      "0000000" when "00010111000010111", -- t[11799] = 0
      "0000000" when "00010111000011000", -- t[11800] = 0
      "0000000" when "00010111000011001", -- t[11801] = 0
      "0000000" when "00010111000011010", -- t[11802] = 0
      "0000000" when "00010111000011011", -- t[11803] = 0
      "0000000" when "00010111000011100", -- t[11804] = 0
      "0000000" when "00010111000011101", -- t[11805] = 0
      "0000000" when "00010111000011110", -- t[11806] = 0
      "0000000" when "00010111000011111", -- t[11807] = 0
      "0000000" when "00010111000100000", -- t[11808] = 0
      "0000000" when "00010111000100001", -- t[11809] = 0
      "0000000" when "00010111000100010", -- t[11810] = 0
      "0000000" when "00010111000100011", -- t[11811] = 0
      "0000000" when "00010111000100100", -- t[11812] = 0
      "0000000" when "00010111000100101", -- t[11813] = 0
      "0000000" when "00010111000100110", -- t[11814] = 0
      "0000000" when "00010111000100111", -- t[11815] = 0
      "0000000" when "00010111000101000", -- t[11816] = 0
      "0000000" when "00010111000101001", -- t[11817] = 0
      "0000000" when "00010111000101010", -- t[11818] = 0
      "0000000" when "00010111000101011", -- t[11819] = 0
      "0000000" when "00010111000101100", -- t[11820] = 0
      "0000000" when "00010111000101101", -- t[11821] = 0
      "0000000" when "00010111000101110", -- t[11822] = 0
      "0000000" when "00010111000101111", -- t[11823] = 0
      "0000000" when "00010111000110000", -- t[11824] = 0
      "0000000" when "00010111000110001", -- t[11825] = 0
      "0000000" when "00010111000110010", -- t[11826] = 0
      "0000000" when "00010111000110011", -- t[11827] = 0
      "0000000" when "00010111000110100", -- t[11828] = 0
      "0000000" when "00010111000110101", -- t[11829] = 0
      "0000000" when "00010111000110110", -- t[11830] = 0
      "0000000" when "00010111000110111", -- t[11831] = 0
      "0000000" when "00010111000111000", -- t[11832] = 0
      "0000000" when "00010111000111001", -- t[11833] = 0
      "0000000" when "00010111000111010", -- t[11834] = 0
      "0000000" when "00010111000111011", -- t[11835] = 0
      "0000000" when "00010111000111100", -- t[11836] = 0
      "0000000" when "00010111000111101", -- t[11837] = 0
      "0000000" when "00010111000111110", -- t[11838] = 0
      "0000000" when "00010111000111111", -- t[11839] = 0
      "0000000" when "00010111001000000", -- t[11840] = 0
      "0000000" when "00010111001000001", -- t[11841] = 0
      "0000000" when "00010111001000010", -- t[11842] = 0
      "0000000" when "00010111001000011", -- t[11843] = 0
      "0000000" when "00010111001000100", -- t[11844] = 0
      "0000000" when "00010111001000101", -- t[11845] = 0
      "0000000" when "00010111001000110", -- t[11846] = 0
      "0000000" when "00010111001000111", -- t[11847] = 0
      "0000000" when "00010111001001000", -- t[11848] = 0
      "0000000" when "00010111001001001", -- t[11849] = 0
      "0000000" when "00010111001001010", -- t[11850] = 0
      "0000000" when "00010111001001011", -- t[11851] = 0
      "0000000" when "00010111001001100", -- t[11852] = 0
      "0000000" when "00010111001001101", -- t[11853] = 0
      "0000000" when "00010111001001110", -- t[11854] = 0
      "0000000" when "00010111001001111", -- t[11855] = 0
      "0000000" when "00010111001010000", -- t[11856] = 0
      "0000000" when "00010111001010001", -- t[11857] = 0
      "0000000" when "00010111001010010", -- t[11858] = 0
      "0000000" when "00010111001010011", -- t[11859] = 0
      "0000000" when "00010111001010100", -- t[11860] = 0
      "0000000" when "00010111001010101", -- t[11861] = 0
      "0000000" when "00010111001010110", -- t[11862] = 0
      "0000000" when "00010111001010111", -- t[11863] = 0
      "0000000" when "00010111001011000", -- t[11864] = 0
      "0000000" when "00010111001011001", -- t[11865] = 0
      "0000000" when "00010111001011010", -- t[11866] = 0
      "0000000" when "00010111001011011", -- t[11867] = 0
      "0000000" when "00010111001011100", -- t[11868] = 0
      "0000000" when "00010111001011101", -- t[11869] = 0
      "0000000" when "00010111001011110", -- t[11870] = 0
      "0000000" when "00010111001011111", -- t[11871] = 0
      "0000000" when "00010111001100000", -- t[11872] = 0
      "0000000" when "00010111001100001", -- t[11873] = 0
      "0000000" when "00010111001100010", -- t[11874] = 0
      "0000000" when "00010111001100011", -- t[11875] = 0
      "0000000" when "00010111001100100", -- t[11876] = 0
      "0000000" when "00010111001100101", -- t[11877] = 0
      "0000000" when "00010111001100110", -- t[11878] = 0
      "0000000" when "00010111001100111", -- t[11879] = 0
      "0000000" when "00010111001101000", -- t[11880] = 0
      "0000000" when "00010111001101001", -- t[11881] = 0
      "0000000" when "00010111001101010", -- t[11882] = 0
      "0000000" when "00010111001101011", -- t[11883] = 0
      "0000000" when "00010111001101100", -- t[11884] = 0
      "0000000" when "00010111001101101", -- t[11885] = 0
      "0000000" when "00010111001101110", -- t[11886] = 0
      "0000000" when "00010111001101111", -- t[11887] = 0
      "0000000" when "00010111001110000", -- t[11888] = 0
      "0000000" when "00010111001110001", -- t[11889] = 0
      "0000000" when "00010111001110010", -- t[11890] = 0
      "0000000" when "00010111001110011", -- t[11891] = 0
      "0000000" when "00010111001110100", -- t[11892] = 0
      "0000000" when "00010111001110101", -- t[11893] = 0
      "0000000" when "00010111001110110", -- t[11894] = 0
      "0000000" when "00010111001110111", -- t[11895] = 0
      "0000000" when "00010111001111000", -- t[11896] = 0
      "0000000" when "00010111001111001", -- t[11897] = 0
      "0000000" when "00010111001111010", -- t[11898] = 0
      "0000000" when "00010111001111011", -- t[11899] = 0
      "0000000" when "00010111001111100", -- t[11900] = 0
      "0000000" when "00010111001111101", -- t[11901] = 0
      "0000000" when "00010111001111110", -- t[11902] = 0
      "0000000" when "00010111001111111", -- t[11903] = 0
      "0000000" when "00010111010000000", -- t[11904] = 0
      "0000000" when "00010111010000001", -- t[11905] = 0
      "0000000" when "00010111010000010", -- t[11906] = 0
      "0000000" when "00010111010000011", -- t[11907] = 0
      "0000000" when "00010111010000100", -- t[11908] = 0
      "0000000" when "00010111010000101", -- t[11909] = 0
      "0000000" when "00010111010000110", -- t[11910] = 0
      "0000000" when "00010111010000111", -- t[11911] = 0
      "0000000" when "00010111010001000", -- t[11912] = 0
      "0000000" when "00010111010001001", -- t[11913] = 0
      "0000000" when "00010111010001010", -- t[11914] = 0
      "0000000" when "00010111010001011", -- t[11915] = 0
      "0000000" when "00010111010001100", -- t[11916] = 0
      "0000000" when "00010111010001101", -- t[11917] = 0
      "0000000" when "00010111010001110", -- t[11918] = 0
      "0000000" when "00010111010001111", -- t[11919] = 0
      "0000000" when "00010111010010000", -- t[11920] = 0
      "0000000" when "00010111010010001", -- t[11921] = 0
      "0000000" when "00010111010010010", -- t[11922] = 0
      "0000000" when "00010111010010011", -- t[11923] = 0
      "0000000" when "00010111010010100", -- t[11924] = 0
      "0000000" when "00010111010010101", -- t[11925] = 0
      "0000000" when "00010111010010110", -- t[11926] = 0
      "0000000" when "00010111010010111", -- t[11927] = 0
      "0000000" when "00010111010011000", -- t[11928] = 0
      "0000000" when "00010111010011001", -- t[11929] = 0
      "0000000" when "00010111010011010", -- t[11930] = 0
      "0000000" when "00010111010011011", -- t[11931] = 0
      "0000000" when "00010111010011100", -- t[11932] = 0
      "0000000" when "00010111010011101", -- t[11933] = 0
      "0000000" when "00010111010011110", -- t[11934] = 0
      "0000000" when "00010111010011111", -- t[11935] = 0
      "0000000" when "00010111010100000", -- t[11936] = 0
      "0000000" when "00010111010100001", -- t[11937] = 0
      "0000000" when "00010111010100010", -- t[11938] = 0
      "0000000" when "00010111010100011", -- t[11939] = 0
      "0000000" when "00010111010100100", -- t[11940] = 0
      "0000000" when "00010111010100101", -- t[11941] = 0
      "0000000" when "00010111010100110", -- t[11942] = 0
      "0000000" when "00010111010100111", -- t[11943] = 0
      "0000000" when "00010111010101000", -- t[11944] = 0
      "0000000" when "00010111010101001", -- t[11945] = 0
      "0000000" when "00010111010101010", -- t[11946] = 0
      "0000000" when "00010111010101011", -- t[11947] = 0
      "0000000" when "00010111010101100", -- t[11948] = 0
      "0000000" when "00010111010101101", -- t[11949] = 0
      "0000000" when "00010111010101110", -- t[11950] = 0
      "0000000" when "00010111010101111", -- t[11951] = 0
      "0000000" when "00010111010110000", -- t[11952] = 0
      "0000000" when "00010111010110001", -- t[11953] = 0
      "0000000" when "00010111010110010", -- t[11954] = 0
      "0000000" when "00010111010110011", -- t[11955] = 0
      "0000000" when "00010111010110100", -- t[11956] = 0
      "0000000" when "00010111010110101", -- t[11957] = 0
      "0000000" when "00010111010110110", -- t[11958] = 0
      "0000000" when "00010111010110111", -- t[11959] = 0
      "0000000" when "00010111010111000", -- t[11960] = 0
      "0000000" when "00010111010111001", -- t[11961] = 0
      "0000000" when "00010111010111010", -- t[11962] = 0
      "0000000" when "00010111010111011", -- t[11963] = 0
      "0000000" when "00010111010111100", -- t[11964] = 0
      "0000000" when "00010111010111101", -- t[11965] = 0
      "0000000" when "00010111010111110", -- t[11966] = 0
      "0000000" when "00010111010111111", -- t[11967] = 0
      "0000000" when "00010111011000000", -- t[11968] = 0
      "0000000" when "00010111011000001", -- t[11969] = 0
      "0000000" when "00010111011000010", -- t[11970] = 0
      "0000000" when "00010111011000011", -- t[11971] = 0
      "0000000" when "00010111011000100", -- t[11972] = 0
      "0000000" when "00010111011000101", -- t[11973] = 0
      "0000000" when "00010111011000110", -- t[11974] = 0
      "0000000" when "00010111011000111", -- t[11975] = 0
      "0000000" when "00010111011001000", -- t[11976] = 0
      "0000000" when "00010111011001001", -- t[11977] = 0
      "0000000" when "00010111011001010", -- t[11978] = 0
      "0000000" when "00010111011001011", -- t[11979] = 0
      "0000000" when "00010111011001100", -- t[11980] = 0
      "0000000" when "00010111011001101", -- t[11981] = 0
      "0000000" when "00010111011001110", -- t[11982] = 0
      "0000000" when "00010111011001111", -- t[11983] = 0
      "0000000" when "00010111011010000", -- t[11984] = 0
      "0000000" when "00010111011010001", -- t[11985] = 0
      "0000000" when "00010111011010010", -- t[11986] = 0
      "0000000" when "00010111011010011", -- t[11987] = 0
      "0000000" when "00010111011010100", -- t[11988] = 0
      "0000000" when "00010111011010101", -- t[11989] = 0
      "0000000" when "00010111011010110", -- t[11990] = 0
      "0000000" when "00010111011010111", -- t[11991] = 0
      "0000000" when "00010111011011000", -- t[11992] = 0
      "0000000" when "00010111011011001", -- t[11993] = 0
      "0000000" when "00010111011011010", -- t[11994] = 0
      "0000000" when "00010111011011011", -- t[11995] = 0
      "0000000" when "00010111011011100", -- t[11996] = 0
      "0000000" when "00010111011011101", -- t[11997] = 0
      "0000000" when "00010111011011110", -- t[11998] = 0
      "0000000" when "00010111011011111", -- t[11999] = 0
      "0000000" when "00010111011100000", -- t[12000] = 0
      "0000000" when "00010111011100001", -- t[12001] = 0
      "0000000" when "00010111011100010", -- t[12002] = 0
      "0000000" when "00010111011100011", -- t[12003] = 0
      "0000000" when "00010111011100100", -- t[12004] = 0
      "0000000" when "00010111011100101", -- t[12005] = 0
      "0000000" when "00010111011100110", -- t[12006] = 0
      "0000000" when "00010111011100111", -- t[12007] = 0
      "0000000" when "00010111011101000", -- t[12008] = 0
      "0000000" when "00010111011101001", -- t[12009] = 0
      "0000000" when "00010111011101010", -- t[12010] = 0
      "0000000" when "00010111011101011", -- t[12011] = 0
      "0000000" when "00010111011101100", -- t[12012] = 0
      "0000000" when "00010111011101101", -- t[12013] = 0
      "0000000" when "00010111011101110", -- t[12014] = 0
      "0000000" when "00010111011101111", -- t[12015] = 0
      "0000000" when "00010111011110000", -- t[12016] = 0
      "0000000" when "00010111011110001", -- t[12017] = 0
      "0000000" when "00010111011110010", -- t[12018] = 0
      "0000000" when "00010111011110011", -- t[12019] = 0
      "0000000" when "00010111011110100", -- t[12020] = 0
      "0000000" when "00010111011110101", -- t[12021] = 0
      "0000000" when "00010111011110110", -- t[12022] = 0
      "0000000" when "00010111011110111", -- t[12023] = 0
      "0000000" when "00010111011111000", -- t[12024] = 0
      "0000000" when "00010111011111001", -- t[12025] = 0
      "0000000" when "00010111011111010", -- t[12026] = 0
      "0000000" when "00010111011111011", -- t[12027] = 0
      "0000000" when "00010111011111100", -- t[12028] = 0
      "0000000" when "00010111011111101", -- t[12029] = 0
      "0000000" when "00010111011111110", -- t[12030] = 0
      "0000000" when "00010111011111111", -- t[12031] = 0
      "0000000" when "00010111100000000", -- t[12032] = 0
      "0000000" when "00010111100000001", -- t[12033] = 0
      "0000000" when "00010111100000010", -- t[12034] = 0
      "0000000" when "00010111100000011", -- t[12035] = 0
      "0000000" when "00010111100000100", -- t[12036] = 0
      "0000000" when "00010111100000101", -- t[12037] = 0
      "0000000" when "00010111100000110", -- t[12038] = 0
      "0000000" when "00010111100000111", -- t[12039] = 0
      "0000000" when "00010111100001000", -- t[12040] = 0
      "0000000" when "00010111100001001", -- t[12041] = 0
      "0000000" when "00010111100001010", -- t[12042] = 0
      "0000000" when "00010111100001011", -- t[12043] = 0
      "0000000" when "00010111100001100", -- t[12044] = 0
      "0000000" when "00010111100001101", -- t[12045] = 0
      "0000000" when "00010111100001110", -- t[12046] = 0
      "0000000" when "00010111100001111", -- t[12047] = 0
      "0000000" when "00010111100010000", -- t[12048] = 0
      "0000000" when "00010111100010001", -- t[12049] = 0
      "0000000" when "00010111100010010", -- t[12050] = 0
      "0000000" when "00010111100010011", -- t[12051] = 0
      "0000000" when "00010111100010100", -- t[12052] = 0
      "0000001" when "00010111100010101", -- t[12053] = 1
      "0000001" when "00010111100010110", -- t[12054] = 1
      "0000001" when "00010111100010111", -- t[12055] = 1
      "0000001" when "00010111100011000", -- t[12056] = 1
      "0000001" when "00010111100011001", -- t[12057] = 1
      "0000001" when "00010111100011010", -- t[12058] = 1
      "0000001" when "00010111100011011", -- t[12059] = 1
      "0000001" when "00010111100011100", -- t[12060] = 1
      "0000001" when "00010111100011101", -- t[12061] = 1
      "0000001" when "00010111100011110", -- t[12062] = 1
      "0000001" when "00010111100011111", -- t[12063] = 1
      "0000001" when "00010111100100000", -- t[12064] = 1
      "0000001" when "00010111100100001", -- t[12065] = 1
      "0000001" when "00010111100100010", -- t[12066] = 1
      "0000001" when "00010111100100011", -- t[12067] = 1
      "0000001" when "00010111100100100", -- t[12068] = 1
      "0000001" when "00010111100100101", -- t[12069] = 1
      "0000001" when "00010111100100110", -- t[12070] = 1
      "0000001" when "00010111100100111", -- t[12071] = 1
      "0000001" when "00010111100101000", -- t[12072] = 1
      "0000001" when "00010111100101001", -- t[12073] = 1
      "0000001" when "00010111100101010", -- t[12074] = 1
      "0000001" when "00010111100101011", -- t[12075] = 1
      "0000001" when "00010111100101100", -- t[12076] = 1
      "0000001" when "00010111100101101", -- t[12077] = 1
      "0000001" when "00010111100101110", -- t[12078] = 1
      "0000001" when "00010111100101111", -- t[12079] = 1
      "0000001" when "00010111100110000", -- t[12080] = 1
      "0000001" when "00010111100110001", -- t[12081] = 1
      "0000001" when "00010111100110010", -- t[12082] = 1
      "0000001" when "00010111100110011", -- t[12083] = 1
      "0000001" when "00010111100110100", -- t[12084] = 1
      "0000001" when "00010111100110101", -- t[12085] = 1
      "0000001" when "00010111100110110", -- t[12086] = 1
      "0000001" when "00010111100110111", -- t[12087] = 1
      "0000001" when "00010111100111000", -- t[12088] = 1
      "0000001" when "00010111100111001", -- t[12089] = 1
      "0000001" when "00010111100111010", -- t[12090] = 1
      "0000001" when "00010111100111011", -- t[12091] = 1
      "0000001" when "00010111100111100", -- t[12092] = 1
      "0000001" when "00010111100111101", -- t[12093] = 1
      "0000001" when "00010111100111110", -- t[12094] = 1
      "0000001" when "00010111100111111", -- t[12095] = 1
      "0000001" when "00010111101000000", -- t[12096] = 1
      "0000001" when "00010111101000001", -- t[12097] = 1
      "0000001" when "00010111101000010", -- t[12098] = 1
      "0000001" when "00010111101000011", -- t[12099] = 1
      "0000001" when "00010111101000100", -- t[12100] = 1
      "0000001" when "00010111101000101", -- t[12101] = 1
      "0000001" when "00010111101000110", -- t[12102] = 1
      "0000001" when "00010111101000111", -- t[12103] = 1
      "0000001" when "00010111101001000", -- t[12104] = 1
      "0000001" when "00010111101001001", -- t[12105] = 1
      "0000001" when "00010111101001010", -- t[12106] = 1
      "0000001" when "00010111101001011", -- t[12107] = 1
      "0000001" when "00010111101001100", -- t[12108] = 1
      "0000001" when "00010111101001101", -- t[12109] = 1
      "0000001" when "00010111101001110", -- t[12110] = 1
      "0000001" when "00010111101001111", -- t[12111] = 1
      "0000001" when "00010111101010000", -- t[12112] = 1
      "0000001" when "00010111101010001", -- t[12113] = 1
      "0000001" when "00010111101010010", -- t[12114] = 1
      "0000001" when "00010111101010011", -- t[12115] = 1
      "0000001" when "00010111101010100", -- t[12116] = 1
      "0000001" when "00010111101010101", -- t[12117] = 1
      "0000001" when "00010111101010110", -- t[12118] = 1
      "0000001" when "00010111101010111", -- t[12119] = 1
      "0000001" when "00010111101011000", -- t[12120] = 1
      "0000001" when "00010111101011001", -- t[12121] = 1
      "0000001" when "00010111101011010", -- t[12122] = 1
      "0000001" when "00010111101011011", -- t[12123] = 1
      "0000001" when "00010111101011100", -- t[12124] = 1
      "0000001" when "00010111101011101", -- t[12125] = 1
      "0000001" when "00010111101011110", -- t[12126] = 1
      "0000001" when "00010111101011111", -- t[12127] = 1
      "0000001" when "00010111101100000", -- t[12128] = 1
      "0000001" when "00010111101100001", -- t[12129] = 1
      "0000001" when "00010111101100010", -- t[12130] = 1
      "0000001" when "00010111101100011", -- t[12131] = 1
      "0000001" when "00010111101100100", -- t[12132] = 1
      "0000001" when "00010111101100101", -- t[12133] = 1
      "0000001" when "00010111101100110", -- t[12134] = 1
      "0000001" when "00010111101100111", -- t[12135] = 1
      "0000001" when "00010111101101000", -- t[12136] = 1
      "0000001" when "00010111101101001", -- t[12137] = 1
      "0000001" when "00010111101101010", -- t[12138] = 1
      "0000001" when "00010111101101011", -- t[12139] = 1
      "0000001" when "00010111101101100", -- t[12140] = 1
      "0000001" when "00010111101101101", -- t[12141] = 1
      "0000001" when "00010111101101110", -- t[12142] = 1
      "0000001" when "00010111101101111", -- t[12143] = 1
      "0000001" when "00010111101110000", -- t[12144] = 1
      "0000001" when "00010111101110001", -- t[12145] = 1
      "0000001" when "00010111101110010", -- t[12146] = 1
      "0000001" when "00010111101110011", -- t[12147] = 1
      "0000001" when "00010111101110100", -- t[12148] = 1
      "0000001" when "00010111101110101", -- t[12149] = 1
      "0000001" when "00010111101110110", -- t[12150] = 1
      "0000001" when "00010111101110111", -- t[12151] = 1
      "0000001" when "00010111101111000", -- t[12152] = 1
      "0000001" when "00010111101111001", -- t[12153] = 1
      "0000001" when "00010111101111010", -- t[12154] = 1
      "0000001" when "00010111101111011", -- t[12155] = 1
      "0000001" when "00010111101111100", -- t[12156] = 1
      "0000001" when "00010111101111101", -- t[12157] = 1
      "0000001" when "00010111101111110", -- t[12158] = 1
      "0000001" when "00010111101111111", -- t[12159] = 1
      "0000001" when "00010111110000000", -- t[12160] = 1
      "0000001" when "00010111110000001", -- t[12161] = 1
      "0000001" when "00010111110000010", -- t[12162] = 1
      "0000001" when "00010111110000011", -- t[12163] = 1
      "0000001" when "00010111110000100", -- t[12164] = 1
      "0000001" when "00010111110000101", -- t[12165] = 1
      "0000001" when "00010111110000110", -- t[12166] = 1
      "0000001" when "00010111110000111", -- t[12167] = 1
      "0000001" when "00010111110001000", -- t[12168] = 1
      "0000001" when "00010111110001001", -- t[12169] = 1
      "0000001" when "00010111110001010", -- t[12170] = 1
      "0000001" when "00010111110001011", -- t[12171] = 1
      "0000001" when "00010111110001100", -- t[12172] = 1
      "0000001" when "00010111110001101", -- t[12173] = 1
      "0000001" when "00010111110001110", -- t[12174] = 1
      "0000001" when "00010111110001111", -- t[12175] = 1
      "0000001" when "00010111110010000", -- t[12176] = 1
      "0000001" when "00010111110010001", -- t[12177] = 1
      "0000001" when "00010111110010010", -- t[12178] = 1
      "0000001" when "00010111110010011", -- t[12179] = 1
      "0000001" when "00010111110010100", -- t[12180] = 1
      "0000001" when "00010111110010101", -- t[12181] = 1
      "0000001" when "00010111110010110", -- t[12182] = 1
      "0000001" when "00010111110010111", -- t[12183] = 1
      "0000001" when "00010111110011000", -- t[12184] = 1
      "0000001" when "00010111110011001", -- t[12185] = 1
      "0000001" when "00010111110011010", -- t[12186] = 1
      "0000001" when "00010111110011011", -- t[12187] = 1
      "0000001" when "00010111110011100", -- t[12188] = 1
      "0000001" when "00010111110011101", -- t[12189] = 1
      "0000001" when "00010111110011110", -- t[12190] = 1
      "0000001" when "00010111110011111", -- t[12191] = 1
      "0000001" when "00010111110100000", -- t[12192] = 1
      "0000001" when "00010111110100001", -- t[12193] = 1
      "0000001" when "00010111110100010", -- t[12194] = 1
      "0000001" when "00010111110100011", -- t[12195] = 1
      "0000001" when "00010111110100100", -- t[12196] = 1
      "0000001" when "00010111110100101", -- t[12197] = 1
      "0000001" when "00010111110100110", -- t[12198] = 1
      "0000001" when "00010111110100111", -- t[12199] = 1
      "0000001" when "00010111110101000", -- t[12200] = 1
      "0000001" when "00010111110101001", -- t[12201] = 1
      "0000001" when "00010111110101010", -- t[12202] = 1
      "0000001" when "00010111110101011", -- t[12203] = 1
      "0000001" when "00010111110101100", -- t[12204] = 1
      "0000001" when "00010111110101101", -- t[12205] = 1
      "0000001" when "00010111110101110", -- t[12206] = 1
      "0000001" when "00010111110101111", -- t[12207] = 1
      "0000001" when "00010111110110000", -- t[12208] = 1
      "0000001" when "00010111110110001", -- t[12209] = 1
      "0000001" when "00010111110110010", -- t[12210] = 1
      "0000001" when "00010111110110011", -- t[12211] = 1
      "0000001" when "00010111110110100", -- t[12212] = 1
      "0000001" when "00010111110110101", -- t[12213] = 1
      "0000001" when "00010111110110110", -- t[12214] = 1
      "0000001" when "00010111110110111", -- t[12215] = 1
      "0000001" when "00010111110111000", -- t[12216] = 1
      "0000001" when "00010111110111001", -- t[12217] = 1
      "0000001" when "00010111110111010", -- t[12218] = 1
      "0000001" when "00010111110111011", -- t[12219] = 1
      "0000001" when "00010111110111100", -- t[12220] = 1
      "0000001" when "00010111110111101", -- t[12221] = 1
      "0000001" when "00010111110111110", -- t[12222] = 1
      "0000001" when "00010111110111111", -- t[12223] = 1
      "0000001" when "00010111111000000", -- t[12224] = 1
      "0000001" when "00010111111000001", -- t[12225] = 1
      "0000001" when "00010111111000010", -- t[12226] = 1
      "0000001" when "00010111111000011", -- t[12227] = 1
      "0000001" when "00010111111000100", -- t[12228] = 1
      "0000001" when "00010111111000101", -- t[12229] = 1
      "0000001" when "00010111111000110", -- t[12230] = 1
      "0000001" when "00010111111000111", -- t[12231] = 1
      "0000001" when "00010111111001000", -- t[12232] = 1
      "0000001" when "00010111111001001", -- t[12233] = 1
      "0000001" when "00010111111001010", -- t[12234] = 1
      "0000001" when "00010111111001011", -- t[12235] = 1
      "0000001" when "00010111111001100", -- t[12236] = 1
      "0000001" when "00010111111001101", -- t[12237] = 1
      "0000001" when "00010111111001110", -- t[12238] = 1
      "0000001" when "00010111111001111", -- t[12239] = 1
      "0000001" when "00010111111010000", -- t[12240] = 1
      "0000001" when "00010111111010001", -- t[12241] = 1
      "0000001" when "00010111111010010", -- t[12242] = 1
      "0000001" when "00010111111010011", -- t[12243] = 1
      "0000001" when "00010111111010100", -- t[12244] = 1
      "0000001" when "00010111111010101", -- t[12245] = 1
      "0000001" when "00010111111010110", -- t[12246] = 1
      "0000001" when "00010111111010111", -- t[12247] = 1
      "0000001" when "00010111111011000", -- t[12248] = 1
      "0000001" when "00010111111011001", -- t[12249] = 1
      "0000001" when "00010111111011010", -- t[12250] = 1
      "0000001" when "00010111111011011", -- t[12251] = 1
      "0000001" when "00010111111011100", -- t[12252] = 1
      "0000001" when "00010111111011101", -- t[12253] = 1
      "0000001" when "00010111111011110", -- t[12254] = 1
      "0000001" when "00010111111011111", -- t[12255] = 1
      "0000001" when "00010111111100000", -- t[12256] = 1
      "0000001" when "00010111111100001", -- t[12257] = 1
      "0000001" when "00010111111100010", -- t[12258] = 1
      "0000001" when "00010111111100011", -- t[12259] = 1
      "0000001" when "00010111111100100", -- t[12260] = 1
      "0000001" when "00010111111100101", -- t[12261] = 1
      "0000001" when "00010111111100110", -- t[12262] = 1
      "0000001" when "00010111111100111", -- t[12263] = 1
      "0000001" when "00010111111101000", -- t[12264] = 1
      "0000001" when "00010111111101001", -- t[12265] = 1
      "0000001" when "00010111111101010", -- t[12266] = 1
      "0000001" when "00010111111101011", -- t[12267] = 1
      "0000001" when "00010111111101100", -- t[12268] = 1
      "0000001" when "00010111111101101", -- t[12269] = 1
      "0000001" when "00010111111101110", -- t[12270] = 1
      "0000001" when "00010111111101111", -- t[12271] = 1
      "0000001" when "00010111111110000", -- t[12272] = 1
      "0000001" when "00010111111110001", -- t[12273] = 1
      "0000001" when "00010111111110010", -- t[12274] = 1
      "0000001" when "00010111111110011", -- t[12275] = 1
      "0000001" when "00010111111110100", -- t[12276] = 1
      "0000001" when "00010111111110101", -- t[12277] = 1
      "0000001" when "00010111111110110", -- t[12278] = 1
      "0000001" when "00010111111110111", -- t[12279] = 1
      "0000001" when "00010111111111000", -- t[12280] = 1
      "0000001" when "00010111111111001", -- t[12281] = 1
      "0000001" when "00010111111111010", -- t[12282] = 1
      "0000001" when "00010111111111011", -- t[12283] = 1
      "0000001" when "00010111111111100", -- t[12284] = 1
      "0000001" when "00010111111111101", -- t[12285] = 1
      "0000001" when "00010111111111110", -- t[12286] = 1
      "0000001" when "00010111111111111", -- t[12287] = 1
      "0000001" when "00011000000000000", -- t[12288] = 1
      "0000001" when "00011000000000001", -- t[12289] = 1
      "0000001" when "00011000000000010", -- t[12290] = 1
      "0000001" when "00011000000000011", -- t[12291] = 1
      "0000001" when "00011000000000100", -- t[12292] = 1
      "0000001" when "00011000000000101", -- t[12293] = 1
      "0000001" when "00011000000000110", -- t[12294] = 1
      "0000001" when "00011000000000111", -- t[12295] = 1
      "0000001" when "00011000000001000", -- t[12296] = 1
      "0000001" when "00011000000001001", -- t[12297] = 1
      "0000001" when "00011000000001010", -- t[12298] = 1
      "0000001" when "00011000000001011", -- t[12299] = 1
      "0000001" when "00011000000001100", -- t[12300] = 1
      "0000001" when "00011000000001101", -- t[12301] = 1
      "0000001" when "00011000000001110", -- t[12302] = 1
      "0000001" when "00011000000001111", -- t[12303] = 1
      "0000001" when "00011000000010000", -- t[12304] = 1
      "0000001" when "00011000000010001", -- t[12305] = 1
      "0000001" when "00011000000010010", -- t[12306] = 1
      "0000001" when "00011000000010011", -- t[12307] = 1
      "0000001" when "00011000000010100", -- t[12308] = 1
      "0000001" when "00011000000010101", -- t[12309] = 1
      "0000001" when "00011000000010110", -- t[12310] = 1
      "0000001" when "00011000000010111", -- t[12311] = 1
      "0000001" when "00011000000011000", -- t[12312] = 1
      "0000001" when "00011000000011001", -- t[12313] = 1
      "0000001" when "00011000000011010", -- t[12314] = 1
      "0000001" when "00011000000011011", -- t[12315] = 1
      "0000001" when "00011000000011100", -- t[12316] = 1
      "0000001" when "00011000000011101", -- t[12317] = 1
      "0000001" when "00011000000011110", -- t[12318] = 1
      "0000001" when "00011000000011111", -- t[12319] = 1
      "0000001" when "00011000000100000", -- t[12320] = 1
      "0000001" when "00011000000100001", -- t[12321] = 1
      "0000001" when "00011000000100010", -- t[12322] = 1
      "0000001" when "00011000000100011", -- t[12323] = 1
      "0000001" when "00011000000100100", -- t[12324] = 1
      "0000001" when "00011000000100101", -- t[12325] = 1
      "0000001" when "00011000000100110", -- t[12326] = 1
      "0000001" when "00011000000100111", -- t[12327] = 1
      "0000001" when "00011000000101000", -- t[12328] = 1
      "0000001" when "00011000000101001", -- t[12329] = 1
      "0000001" when "00011000000101010", -- t[12330] = 1
      "0000001" when "00011000000101011", -- t[12331] = 1
      "0000001" when "00011000000101100", -- t[12332] = 1
      "0000001" when "00011000000101101", -- t[12333] = 1
      "0000001" when "00011000000101110", -- t[12334] = 1
      "0000001" when "00011000000101111", -- t[12335] = 1
      "0000001" when "00011000000110000", -- t[12336] = 1
      "0000001" when "00011000000110001", -- t[12337] = 1
      "0000001" when "00011000000110010", -- t[12338] = 1
      "0000001" when "00011000000110011", -- t[12339] = 1
      "0000001" when "00011000000110100", -- t[12340] = 1
      "0000001" when "00011000000110101", -- t[12341] = 1
      "0000001" when "00011000000110110", -- t[12342] = 1
      "0000001" when "00011000000110111", -- t[12343] = 1
      "0000001" when "00011000000111000", -- t[12344] = 1
      "0000001" when "00011000000111001", -- t[12345] = 1
      "0000001" when "00011000000111010", -- t[12346] = 1
      "0000001" when "00011000000111011", -- t[12347] = 1
      "0000001" when "00011000000111100", -- t[12348] = 1
      "0000001" when "00011000000111101", -- t[12349] = 1
      "0000001" when "00011000000111110", -- t[12350] = 1
      "0000001" when "00011000000111111", -- t[12351] = 1
      "0000001" when "00011000001000000", -- t[12352] = 1
      "0000001" when "00011000001000001", -- t[12353] = 1
      "0000001" when "00011000001000010", -- t[12354] = 1
      "0000001" when "00011000001000011", -- t[12355] = 1
      "0000001" when "00011000001000100", -- t[12356] = 1
      "0000001" when "00011000001000101", -- t[12357] = 1
      "0000001" when "00011000001000110", -- t[12358] = 1
      "0000001" when "00011000001000111", -- t[12359] = 1
      "0000001" when "00011000001001000", -- t[12360] = 1
      "0000001" when "00011000001001001", -- t[12361] = 1
      "0000001" when "00011000001001010", -- t[12362] = 1
      "0000001" when "00011000001001011", -- t[12363] = 1
      "0000001" when "00011000001001100", -- t[12364] = 1
      "0000001" when "00011000001001101", -- t[12365] = 1
      "0000001" when "00011000001001110", -- t[12366] = 1
      "0000001" when "00011000001001111", -- t[12367] = 1
      "0000001" when "00011000001010000", -- t[12368] = 1
      "0000001" when "00011000001010001", -- t[12369] = 1
      "0000001" when "00011000001010010", -- t[12370] = 1
      "0000001" when "00011000001010011", -- t[12371] = 1
      "0000001" when "00011000001010100", -- t[12372] = 1
      "0000001" when "00011000001010101", -- t[12373] = 1
      "0000001" when "00011000001010110", -- t[12374] = 1
      "0000001" when "00011000001010111", -- t[12375] = 1
      "0000001" when "00011000001011000", -- t[12376] = 1
      "0000001" when "00011000001011001", -- t[12377] = 1
      "0000001" when "00011000001011010", -- t[12378] = 1
      "0000001" when "00011000001011011", -- t[12379] = 1
      "0000001" when "00011000001011100", -- t[12380] = 1
      "0000001" when "00011000001011101", -- t[12381] = 1
      "0000001" when "00011000001011110", -- t[12382] = 1
      "0000001" when "00011000001011111", -- t[12383] = 1
      "0000001" when "00011000001100000", -- t[12384] = 1
      "0000001" when "00011000001100001", -- t[12385] = 1
      "0000001" when "00011000001100010", -- t[12386] = 1
      "0000001" when "00011000001100011", -- t[12387] = 1
      "0000001" when "00011000001100100", -- t[12388] = 1
      "0000001" when "00011000001100101", -- t[12389] = 1
      "0000001" when "00011000001100110", -- t[12390] = 1
      "0000001" when "00011000001100111", -- t[12391] = 1
      "0000001" when "00011000001101000", -- t[12392] = 1
      "0000001" when "00011000001101001", -- t[12393] = 1
      "0000001" when "00011000001101010", -- t[12394] = 1
      "0000001" when "00011000001101011", -- t[12395] = 1
      "0000001" when "00011000001101100", -- t[12396] = 1
      "0000001" when "00011000001101101", -- t[12397] = 1
      "0000001" when "00011000001101110", -- t[12398] = 1
      "0000001" when "00011000001101111", -- t[12399] = 1
      "0000001" when "00011000001110000", -- t[12400] = 1
      "0000001" when "00011000001110001", -- t[12401] = 1
      "0000001" when "00011000001110010", -- t[12402] = 1
      "0000001" when "00011000001110011", -- t[12403] = 1
      "0000001" when "00011000001110100", -- t[12404] = 1
      "0000001" when "00011000001110101", -- t[12405] = 1
      "0000001" when "00011000001110110", -- t[12406] = 1
      "0000001" when "00011000001110111", -- t[12407] = 1
      "0000001" when "00011000001111000", -- t[12408] = 1
      "0000001" when "00011000001111001", -- t[12409] = 1
      "0000001" when "00011000001111010", -- t[12410] = 1
      "0000001" when "00011000001111011", -- t[12411] = 1
      "0000001" when "00011000001111100", -- t[12412] = 1
      "0000001" when "00011000001111101", -- t[12413] = 1
      "0000001" when "00011000001111110", -- t[12414] = 1
      "0000001" when "00011000001111111", -- t[12415] = 1
      "0000001" when "00011000010000000", -- t[12416] = 1
      "0000001" when "00011000010000001", -- t[12417] = 1
      "0000001" when "00011000010000010", -- t[12418] = 1
      "0000001" when "00011000010000011", -- t[12419] = 1
      "0000001" when "00011000010000100", -- t[12420] = 1
      "0000001" when "00011000010000101", -- t[12421] = 1
      "0000001" when "00011000010000110", -- t[12422] = 1
      "0000001" when "00011000010000111", -- t[12423] = 1
      "0000001" when "00011000010001000", -- t[12424] = 1
      "0000001" when "00011000010001001", -- t[12425] = 1
      "0000001" when "00011000010001010", -- t[12426] = 1
      "0000001" when "00011000010001011", -- t[12427] = 1
      "0000001" when "00011000010001100", -- t[12428] = 1
      "0000001" when "00011000010001101", -- t[12429] = 1
      "0000001" when "00011000010001110", -- t[12430] = 1
      "0000001" when "00011000010001111", -- t[12431] = 1
      "0000001" when "00011000010010000", -- t[12432] = 1
      "0000001" when "00011000010010001", -- t[12433] = 1
      "0000001" when "00011000010010010", -- t[12434] = 1
      "0000001" when "00011000010010011", -- t[12435] = 1
      "0000001" when "00011000010010100", -- t[12436] = 1
      "0000001" when "00011000010010101", -- t[12437] = 1
      "0000001" when "00011000010010110", -- t[12438] = 1
      "0000001" when "00011000010010111", -- t[12439] = 1
      "0000001" when "00011000010011000", -- t[12440] = 1
      "0000001" when "00011000010011001", -- t[12441] = 1
      "0000001" when "00011000010011010", -- t[12442] = 1
      "0000001" when "00011000010011011", -- t[12443] = 1
      "0000001" when "00011000010011100", -- t[12444] = 1
      "0000001" when "00011000010011101", -- t[12445] = 1
      "0000001" when "00011000010011110", -- t[12446] = 1
      "0000001" when "00011000010011111", -- t[12447] = 1
      "0000001" when "00011000010100000", -- t[12448] = 1
      "0000001" when "00011000010100001", -- t[12449] = 1
      "0000001" when "00011000010100010", -- t[12450] = 1
      "0000001" when "00011000010100011", -- t[12451] = 1
      "0000001" when "00011000010100100", -- t[12452] = 1
      "0000001" when "00011000010100101", -- t[12453] = 1
      "0000001" when "00011000010100110", -- t[12454] = 1
      "0000001" when "00011000010100111", -- t[12455] = 1
      "0000001" when "00011000010101000", -- t[12456] = 1
      "0000001" when "00011000010101001", -- t[12457] = 1
      "0000001" when "00011000010101010", -- t[12458] = 1
      "0000001" when "00011000010101011", -- t[12459] = 1
      "0000001" when "00011000010101100", -- t[12460] = 1
      "0000001" when "00011000010101101", -- t[12461] = 1
      "0000001" when "00011000010101110", -- t[12462] = 1
      "0000001" when "00011000010101111", -- t[12463] = 1
      "0000001" when "00011000010110000", -- t[12464] = 1
      "0000001" when "00011000010110001", -- t[12465] = 1
      "0000001" when "00011000010110010", -- t[12466] = 1
      "0000001" when "00011000010110011", -- t[12467] = 1
      "0000001" when "00011000010110100", -- t[12468] = 1
      "0000001" when "00011000010110101", -- t[12469] = 1
      "0000001" when "00011000010110110", -- t[12470] = 1
      "0000001" when "00011000010110111", -- t[12471] = 1
      "0000001" when "00011000010111000", -- t[12472] = 1
      "0000001" when "00011000010111001", -- t[12473] = 1
      "0000001" when "00011000010111010", -- t[12474] = 1
      "0000001" when "00011000010111011", -- t[12475] = 1
      "0000001" when "00011000010111100", -- t[12476] = 1
      "0000001" when "00011000010111101", -- t[12477] = 1
      "0000001" when "00011000010111110", -- t[12478] = 1
      "0000001" when "00011000010111111", -- t[12479] = 1
      "0000001" when "00011000011000000", -- t[12480] = 1
      "0000001" when "00011000011000001", -- t[12481] = 1
      "0000001" when "00011000011000010", -- t[12482] = 1
      "0000001" when "00011000011000011", -- t[12483] = 1
      "0000001" when "00011000011000100", -- t[12484] = 1
      "0000001" when "00011000011000101", -- t[12485] = 1
      "0000001" when "00011000011000110", -- t[12486] = 1
      "0000001" when "00011000011000111", -- t[12487] = 1
      "0000001" when "00011000011001000", -- t[12488] = 1
      "0000001" when "00011000011001001", -- t[12489] = 1
      "0000001" when "00011000011001010", -- t[12490] = 1
      "0000001" when "00011000011001011", -- t[12491] = 1
      "0000001" when "00011000011001100", -- t[12492] = 1
      "0000001" when "00011000011001101", -- t[12493] = 1
      "0000001" when "00011000011001110", -- t[12494] = 1
      "0000001" when "00011000011001111", -- t[12495] = 1
      "0000001" when "00011000011010000", -- t[12496] = 1
      "0000001" when "00011000011010001", -- t[12497] = 1
      "0000001" when "00011000011010010", -- t[12498] = 1
      "0000001" when "00011000011010011", -- t[12499] = 1
      "0000001" when "00011000011010100", -- t[12500] = 1
      "0000001" when "00011000011010101", -- t[12501] = 1
      "0000001" when "00011000011010110", -- t[12502] = 1
      "0000001" when "00011000011010111", -- t[12503] = 1
      "0000001" when "00011000011011000", -- t[12504] = 1
      "0000001" when "00011000011011001", -- t[12505] = 1
      "0000001" when "00011000011011010", -- t[12506] = 1
      "0000001" when "00011000011011011", -- t[12507] = 1
      "0000001" when "00011000011011100", -- t[12508] = 1
      "0000001" when "00011000011011101", -- t[12509] = 1
      "0000001" when "00011000011011110", -- t[12510] = 1
      "0000001" when "00011000011011111", -- t[12511] = 1
      "0000001" when "00011000011100000", -- t[12512] = 1
      "0000001" when "00011000011100001", -- t[12513] = 1
      "0000001" when "00011000011100010", -- t[12514] = 1
      "0000001" when "00011000011100011", -- t[12515] = 1
      "0000001" when "00011000011100100", -- t[12516] = 1
      "0000001" when "00011000011100101", -- t[12517] = 1
      "0000001" when "00011000011100110", -- t[12518] = 1
      "0000001" when "00011000011100111", -- t[12519] = 1
      "0000001" when "00011000011101000", -- t[12520] = 1
      "0000001" when "00011000011101001", -- t[12521] = 1
      "0000001" when "00011000011101010", -- t[12522] = 1
      "0000001" when "00011000011101011", -- t[12523] = 1
      "0000001" when "00011000011101100", -- t[12524] = 1
      "0000001" when "00011000011101101", -- t[12525] = 1
      "0000001" when "00011000011101110", -- t[12526] = 1
      "0000001" when "00011000011101111", -- t[12527] = 1
      "0000001" when "00011000011110000", -- t[12528] = 1
      "0000001" when "00011000011110001", -- t[12529] = 1
      "0000001" when "00011000011110010", -- t[12530] = 1
      "0000001" when "00011000011110011", -- t[12531] = 1
      "0000001" when "00011000011110100", -- t[12532] = 1
      "0000001" when "00011000011110101", -- t[12533] = 1
      "0000001" when "00011000011110110", -- t[12534] = 1
      "0000001" when "00011000011110111", -- t[12535] = 1
      "0000001" when "00011000011111000", -- t[12536] = 1
      "0000001" when "00011000011111001", -- t[12537] = 1
      "0000001" when "00011000011111010", -- t[12538] = 1
      "0000001" when "00011000011111011", -- t[12539] = 1
      "0000001" when "00011000011111100", -- t[12540] = 1
      "0000001" when "00011000011111101", -- t[12541] = 1
      "0000001" when "00011000011111110", -- t[12542] = 1
      "0000001" when "00011000011111111", -- t[12543] = 1
      "0000001" when "00011000100000000", -- t[12544] = 1
      "0000001" when "00011000100000001", -- t[12545] = 1
      "0000001" when "00011000100000010", -- t[12546] = 1
      "0000001" when "00011000100000011", -- t[12547] = 1
      "0000001" when "00011000100000100", -- t[12548] = 1
      "0000001" when "00011000100000101", -- t[12549] = 1
      "0000001" when "00011000100000110", -- t[12550] = 1
      "0000001" when "00011000100000111", -- t[12551] = 1
      "0000001" when "00011000100001000", -- t[12552] = 1
      "0000001" when "00011000100001001", -- t[12553] = 1
      "0000001" when "00011000100001010", -- t[12554] = 1
      "0000001" when "00011000100001011", -- t[12555] = 1
      "0000001" when "00011000100001100", -- t[12556] = 1
      "0000001" when "00011000100001101", -- t[12557] = 1
      "0000001" when "00011000100001110", -- t[12558] = 1
      "0000001" when "00011000100001111", -- t[12559] = 1
      "0000001" when "00011000100010000", -- t[12560] = 1
      "0000001" when "00011000100010001", -- t[12561] = 1
      "0000001" when "00011000100010010", -- t[12562] = 1
      "0000001" when "00011000100010011", -- t[12563] = 1
      "0000001" when "00011000100010100", -- t[12564] = 1
      "0000001" when "00011000100010101", -- t[12565] = 1
      "0000001" when "00011000100010110", -- t[12566] = 1
      "0000001" when "00011000100010111", -- t[12567] = 1
      "0000001" when "00011000100011000", -- t[12568] = 1
      "0000001" when "00011000100011001", -- t[12569] = 1
      "0000001" when "00011000100011010", -- t[12570] = 1
      "0000001" when "00011000100011011", -- t[12571] = 1
      "0000001" when "00011000100011100", -- t[12572] = 1
      "0000001" when "00011000100011101", -- t[12573] = 1
      "0000001" when "00011000100011110", -- t[12574] = 1
      "0000001" when "00011000100011111", -- t[12575] = 1
      "0000001" when "00011000100100000", -- t[12576] = 1
      "0000001" when "00011000100100001", -- t[12577] = 1
      "0000001" when "00011000100100010", -- t[12578] = 1
      "0000001" when "00011000100100011", -- t[12579] = 1
      "0000001" when "00011000100100100", -- t[12580] = 1
      "0000001" when "00011000100100101", -- t[12581] = 1
      "0000001" when "00011000100100110", -- t[12582] = 1
      "0000001" when "00011000100100111", -- t[12583] = 1
      "0000001" when "00011000100101000", -- t[12584] = 1
      "0000001" when "00011000100101001", -- t[12585] = 1
      "0000001" when "00011000100101010", -- t[12586] = 1
      "0000001" when "00011000100101011", -- t[12587] = 1
      "0000001" when "00011000100101100", -- t[12588] = 1
      "0000001" when "00011000100101101", -- t[12589] = 1
      "0000001" when "00011000100101110", -- t[12590] = 1
      "0000001" when "00011000100101111", -- t[12591] = 1
      "0000001" when "00011000100110000", -- t[12592] = 1
      "0000001" when "00011000100110001", -- t[12593] = 1
      "0000001" when "00011000100110010", -- t[12594] = 1
      "0000001" when "00011000100110011", -- t[12595] = 1
      "0000001" when "00011000100110100", -- t[12596] = 1
      "0000001" when "00011000100110101", -- t[12597] = 1
      "0000001" when "00011000100110110", -- t[12598] = 1
      "0000001" when "00011000100110111", -- t[12599] = 1
      "0000001" when "00011000100111000", -- t[12600] = 1
      "0000001" when "00011000100111001", -- t[12601] = 1
      "0000001" when "00011000100111010", -- t[12602] = 1
      "0000001" when "00011000100111011", -- t[12603] = 1
      "0000001" when "00011000100111100", -- t[12604] = 1
      "0000001" when "00011000100111101", -- t[12605] = 1
      "0000001" when "00011000100111110", -- t[12606] = 1
      "0000001" when "00011000100111111", -- t[12607] = 1
      "0000001" when "00011000101000000", -- t[12608] = 1
      "0000001" when "00011000101000001", -- t[12609] = 1
      "0000001" when "00011000101000010", -- t[12610] = 1
      "0000001" when "00011000101000011", -- t[12611] = 1
      "0000001" when "00011000101000100", -- t[12612] = 1
      "0000001" when "00011000101000101", -- t[12613] = 1
      "0000001" when "00011000101000110", -- t[12614] = 1
      "0000001" when "00011000101000111", -- t[12615] = 1
      "0000001" when "00011000101001000", -- t[12616] = 1
      "0000001" when "00011000101001001", -- t[12617] = 1
      "0000001" when "00011000101001010", -- t[12618] = 1
      "0000001" when "00011000101001011", -- t[12619] = 1
      "0000001" when "00011000101001100", -- t[12620] = 1
      "0000001" when "00011000101001101", -- t[12621] = 1
      "0000001" when "00011000101001110", -- t[12622] = 1
      "0000001" when "00011000101001111", -- t[12623] = 1
      "0000001" when "00011000101010000", -- t[12624] = 1
      "0000001" when "00011000101010001", -- t[12625] = 1
      "0000001" when "00011000101010010", -- t[12626] = 1
      "0000001" when "00011000101010011", -- t[12627] = 1
      "0000001" when "00011000101010100", -- t[12628] = 1
      "0000001" when "00011000101010101", -- t[12629] = 1
      "0000001" when "00011000101010110", -- t[12630] = 1
      "0000001" when "00011000101010111", -- t[12631] = 1
      "0000001" when "00011000101011000", -- t[12632] = 1
      "0000001" when "00011000101011001", -- t[12633] = 1
      "0000001" when "00011000101011010", -- t[12634] = 1
      "0000001" when "00011000101011011", -- t[12635] = 1
      "0000001" when "00011000101011100", -- t[12636] = 1
      "0000001" when "00011000101011101", -- t[12637] = 1
      "0000001" when "00011000101011110", -- t[12638] = 1
      "0000001" when "00011000101011111", -- t[12639] = 1
      "0000001" when "00011000101100000", -- t[12640] = 1
      "0000001" when "00011000101100001", -- t[12641] = 1
      "0000001" when "00011000101100010", -- t[12642] = 1
      "0000001" when "00011000101100011", -- t[12643] = 1
      "0000001" when "00011000101100100", -- t[12644] = 1
      "0000001" when "00011000101100101", -- t[12645] = 1
      "0000001" when "00011000101100110", -- t[12646] = 1
      "0000001" when "00011000101100111", -- t[12647] = 1
      "0000001" when "00011000101101000", -- t[12648] = 1
      "0000001" when "00011000101101001", -- t[12649] = 1
      "0000001" when "00011000101101010", -- t[12650] = 1
      "0000001" when "00011000101101011", -- t[12651] = 1
      "0000001" when "00011000101101100", -- t[12652] = 1
      "0000001" when "00011000101101101", -- t[12653] = 1
      "0000001" when "00011000101101110", -- t[12654] = 1
      "0000001" when "00011000101101111", -- t[12655] = 1
      "0000001" when "00011000101110000", -- t[12656] = 1
      "0000001" when "00011000101110001", -- t[12657] = 1
      "0000001" when "00011000101110010", -- t[12658] = 1
      "0000001" when "00011000101110011", -- t[12659] = 1
      "0000001" when "00011000101110100", -- t[12660] = 1
      "0000001" when "00011000101110101", -- t[12661] = 1
      "0000001" when "00011000101110110", -- t[12662] = 1
      "0000001" when "00011000101110111", -- t[12663] = 1
      "0000001" when "00011000101111000", -- t[12664] = 1
      "0000001" when "00011000101111001", -- t[12665] = 1
      "0000001" when "00011000101111010", -- t[12666] = 1
      "0000001" when "00011000101111011", -- t[12667] = 1
      "0000001" when "00011000101111100", -- t[12668] = 1
      "0000001" when "00011000101111101", -- t[12669] = 1
      "0000001" when "00011000101111110", -- t[12670] = 1
      "0000001" when "00011000101111111", -- t[12671] = 1
      "0000001" when "00011000110000000", -- t[12672] = 1
      "0000001" when "00011000110000001", -- t[12673] = 1
      "0000001" when "00011000110000010", -- t[12674] = 1
      "0000001" when "00011000110000011", -- t[12675] = 1
      "0000001" when "00011000110000100", -- t[12676] = 1
      "0000001" when "00011000110000101", -- t[12677] = 1
      "0000001" when "00011000110000110", -- t[12678] = 1
      "0000001" when "00011000110000111", -- t[12679] = 1
      "0000001" when "00011000110001000", -- t[12680] = 1
      "0000001" when "00011000110001001", -- t[12681] = 1
      "0000001" when "00011000110001010", -- t[12682] = 1
      "0000001" when "00011000110001011", -- t[12683] = 1
      "0000001" when "00011000110001100", -- t[12684] = 1
      "0000001" when "00011000110001101", -- t[12685] = 1
      "0000001" when "00011000110001110", -- t[12686] = 1
      "0000001" when "00011000110001111", -- t[12687] = 1
      "0000001" when "00011000110010000", -- t[12688] = 1
      "0000001" when "00011000110010001", -- t[12689] = 1
      "0000001" when "00011000110010010", -- t[12690] = 1
      "0000001" when "00011000110010011", -- t[12691] = 1
      "0000001" when "00011000110010100", -- t[12692] = 1
      "0000001" when "00011000110010101", -- t[12693] = 1
      "0000001" when "00011000110010110", -- t[12694] = 1
      "0000001" when "00011000110010111", -- t[12695] = 1
      "0000001" when "00011000110011000", -- t[12696] = 1
      "0000001" when "00011000110011001", -- t[12697] = 1
      "0000001" when "00011000110011010", -- t[12698] = 1
      "0000001" when "00011000110011011", -- t[12699] = 1
      "0000001" when "00011000110011100", -- t[12700] = 1
      "0000001" when "00011000110011101", -- t[12701] = 1
      "0000001" when "00011000110011110", -- t[12702] = 1
      "0000001" when "00011000110011111", -- t[12703] = 1
      "0000001" when "00011000110100000", -- t[12704] = 1
      "0000001" when "00011000110100001", -- t[12705] = 1
      "0000001" when "00011000110100010", -- t[12706] = 1
      "0000001" when "00011000110100011", -- t[12707] = 1
      "0000001" when "00011000110100100", -- t[12708] = 1
      "0000001" when "00011000110100101", -- t[12709] = 1
      "0000001" when "00011000110100110", -- t[12710] = 1
      "0000001" when "00011000110100111", -- t[12711] = 1
      "0000001" when "00011000110101000", -- t[12712] = 1
      "0000001" when "00011000110101001", -- t[12713] = 1
      "0000001" when "00011000110101010", -- t[12714] = 1
      "0000001" when "00011000110101011", -- t[12715] = 1
      "0000001" when "00011000110101100", -- t[12716] = 1
      "0000001" when "00011000110101101", -- t[12717] = 1
      "0000001" when "00011000110101110", -- t[12718] = 1
      "0000001" when "00011000110101111", -- t[12719] = 1
      "0000001" when "00011000110110000", -- t[12720] = 1
      "0000001" when "00011000110110001", -- t[12721] = 1
      "0000001" when "00011000110110010", -- t[12722] = 1
      "0000001" when "00011000110110011", -- t[12723] = 1
      "0000001" when "00011000110110100", -- t[12724] = 1
      "0000001" when "00011000110110101", -- t[12725] = 1
      "0000001" when "00011000110110110", -- t[12726] = 1
      "0000001" when "00011000110110111", -- t[12727] = 1
      "0000001" when "00011000110111000", -- t[12728] = 1
      "0000001" when "00011000110111001", -- t[12729] = 1
      "0000001" when "00011000110111010", -- t[12730] = 1
      "0000001" when "00011000110111011", -- t[12731] = 1
      "0000001" when "00011000110111100", -- t[12732] = 1
      "0000001" when "00011000110111101", -- t[12733] = 1
      "0000001" when "00011000110111110", -- t[12734] = 1
      "0000001" when "00011000110111111", -- t[12735] = 1
      "0000001" when "00011000111000000", -- t[12736] = 1
      "0000001" when "00011000111000001", -- t[12737] = 1
      "0000001" when "00011000111000010", -- t[12738] = 1
      "0000001" when "00011000111000011", -- t[12739] = 1
      "0000001" when "00011000111000100", -- t[12740] = 1
      "0000001" when "00011000111000101", -- t[12741] = 1
      "0000001" when "00011000111000110", -- t[12742] = 1
      "0000001" when "00011000111000111", -- t[12743] = 1
      "0000001" when "00011000111001000", -- t[12744] = 1
      "0000001" when "00011000111001001", -- t[12745] = 1
      "0000001" when "00011000111001010", -- t[12746] = 1
      "0000001" when "00011000111001011", -- t[12747] = 1
      "0000001" when "00011000111001100", -- t[12748] = 1
      "0000001" when "00011000111001101", -- t[12749] = 1
      "0000001" when "00011000111001110", -- t[12750] = 1
      "0000001" when "00011000111001111", -- t[12751] = 1
      "0000001" when "00011000111010000", -- t[12752] = 1
      "0000001" when "00011000111010001", -- t[12753] = 1
      "0000001" when "00011000111010010", -- t[12754] = 1
      "0000001" when "00011000111010011", -- t[12755] = 1
      "0000001" when "00011000111010100", -- t[12756] = 1
      "0000001" when "00011000111010101", -- t[12757] = 1
      "0000001" when "00011000111010110", -- t[12758] = 1
      "0000001" when "00011000111010111", -- t[12759] = 1
      "0000001" when "00011000111011000", -- t[12760] = 1
      "0000001" when "00011000111011001", -- t[12761] = 1
      "0000001" when "00011000111011010", -- t[12762] = 1
      "0000001" when "00011000111011011", -- t[12763] = 1
      "0000001" when "00011000111011100", -- t[12764] = 1
      "0000001" when "00011000111011101", -- t[12765] = 1
      "0000001" when "00011000111011110", -- t[12766] = 1
      "0000001" when "00011000111011111", -- t[12767] = 1
      "0000001" when "00011000111100000", -- t[12768] = 1
      "0000001" when "00011000111100001", -- t[12769] = 1
      "0000001" when "00011000111100010", -- t[12770] = 1
      "0000001" when "00011000111100011", -- t[12771] = 1
      "0000001" when "00011000111100100", -- t[12772] = 1
      "0000001" when "00011000111100101", -- t[12773] = 1
      "0000001" when "00011000111100110", -- t[12774] = 1
      "0000001" when "00011000111100111", -- t[12775] = 1
      "0000001" when "00011000111101000", -- t[12776] = 1
      "0000001" when "00011000111101001", -- t[12777] = 1
      "0000001" when "00011000111101010", -- t[12778] = 1
      "0000001" when "00011000111101011", -- t[12779] = 1
      "0000001" when "00011000111101100", -- t[12780] = 1
      "0000001" when "00011000111101101", -- t[12781] = 1
      "0000001" when "00011000111101110", -- t[12782] = 1
      "0000001" when "00011000111101111", -- t[12783] = 1
      "0000001" when "00011000111110000", -- t[12784] = 1
      "0000001" when "00011000111110001", -- t[12785] = 1
      "0000001" when "00011000111110010", -- t[12786] = 1
      "0000001" when "00011000111110011", -- t[12787] = 1
      "0000001" when "00011000111110100", -- t[12788] = 1
      "0000001" when "00011000111110101", -- t[12789] = 1
      "0000001" when "00011000111110110", -- t[12790] = 1
      "0000001" when "00011000111110111", -- t[12791] = 1
      "0000001" when "00011000111111000", -- t[12792] = 1
      "0000001" when "00011000111111001", -- t[12793] = 1
      "0000001" when "00011000111111010", -- t[12794] = 1
      "0000001" when "00011000111111011", -- t[12795] = 1
      "0000001" when "00011000111111100", -- t[12796] = 1
      "0000001" when "00011000111111101", -- t[12797] = 1
      "0000001" when "00011000111111110", -- t[12798] = 1
      "0000001" when "00011000111111111", -- t[12799] = 1
      "0000001" when "00011001000000000", -- t[12800] = 1
      "0000001" when "00011001000000001", -- t[12801] = 1
      "0000001" when "00011001000000010", -- t[12802] = 1
      "0000001" when "00011001000000011", -- t[12803] = 1
      "0000001" when "00011001000000100", -- t[12804] = 1
      "0000001" when "00011001000000101", -- t[12805] = 1
      "0000001" when "00011001000000110", -- t[12806] = 1
      "0000001" when "00011001000000111", -- t[12807] = 1
      "0000001" when "00011001000001000", -- t[12808] = 1
      "0000001" when "00011001000001001", -- t[12809] = 1
      "0000001" when "00011001000001010", -- t[12810] = 1
      "0000001" when "00011001000001011", -- t[12811] = 1
      "0000001" when "00011001000001100", -- t[12812] = 1
      "0000001" when "00011001000001101", -- t[12813] = 1
      "0000001" when "00011001000001110", -- t[12814] = 1
      "0000001" when "00011001000001111", -- t[12815] = 1
      "0000001" when "00011001000010000", -- t[12816] = 1
      "0000001" when "00011001000010001", -- t[12817] = 1
      "0000001" when "00011001000010010", -- t[12818] = 1
      "0000001" when "00011001000010011", -- t[12819] = 1
      "0000001" when "00011001000010100", -- t[12820] = 1
      "0000001" when "00011001000010101", -- t[12821] = 1
      "0000001" when "00011001000010110", -- t[12822] = 1
      "0000001" when "00011001000010111", -- t[12823] = 1
      "0000001" when "00011001000011000", -- t[12824] = 1
      "0000001" when "00011001000011001", -- t[12825] = 1
      "0000001" when "00011001000011010", -- t[12826] = 1
      "0000001" when "00011001000011011", -- t[12827] = 1
      "0000001" when "00011001000011100", -- t[12828] = 1
      "0000001" when "00011001000011101", -- t[12829] = 1
      "0000001" when "00011001000011110", -- t[12830] = 1
      "0000001" when "00011001000011111", -- t[12831] = 1
      "0000001" when "00011001000100000", -- t[12832] = 1
      "0000001" when "00011001000100001", -- t[12833] = 1
      "0000001" when "00011001000100010", -- t[12834] = 1
      "0000001" when "00011001000100011", -- t[12835] = 1
      "0000001" when "00011001000100100", -- t[12836] = 1
      "0000001" when "00011001000100101", -- t[12837] = 1
      "0000001" when "00011001000100110", -- t[12838] = 1
      "0000001" when "00011001000100111", -- t[12839] = 1
      "0000001" when "00011001000101000", -- t[12840] = 1
      "0000001" when "00011001000101001", -- t[12841] = 1
      "0000001" when "00011001000101010", -- t[12842] = 1
      "0000001" when "00011001000101011", -- t[12843] = 1
      "0000001" when "00011001000101100", -- t[12844] = 1
      "0000001" when "00011001000101101", -- t[12845] = 1
      "0000001" when "00011001000101110", -- t[12846] = 1
      "0000001" when "00011001000101111", -- t[12847] = 1
      "0000001" when "00011001000110000", -- t[12848] = 1
      "0000001" when "00011001000110001", -- t[12849] = 1
      "0000001" when "00011001000110010", -- t[12850] = 1
      "0000001" when "00011001000110011", -- t[12851] = 1
      "0000001" when "00011001000110100", -- t[12852] = 1
      "0000001" when "00011001000110101", -- t[12853] = 1
      "0000001" when "00011001000110110", -- t[12854] = 1
      "0000001" when "00011001000110111", -- t[12855] = 1
      "0000001" when "00011001000111000", -- t[12856] = 1
      "0000001" when "00011001000111001", -- t[12857] = 1
      "0000001" when "00011001000111010", -- t[12858] = 1
      "0000001" when "00011001000111011", -- t[12859] = 1
      "0000001" when "00011001000111100", -- t[12860] = 1
      "0000001" when "00011001000111101", -- t[12861] = 1
      "0000001" when "00011001000111110", -- t[12862] = 1
      "0000001" when "00011001000111111", -- t[12863] = 1
      "0000001" when "00011001001000000", -- t[12864] = 1
      "0000001" when "00011001001000001", -- t[12865] = 1
      "0000001" when "00011001001000010", -- t[12866] = 1
      "0000001" when "00011001001000011", -- t[12867] = 1
      "0000001" when "00011001001000100", -- t[12868] = 1
      "0000001" when "00011001001000101", -- t[12869] = 1
      "0000001" when "00011001001000110", -- t[12870] = 1
      "0000001" when "00011001001000111", -- t[12871] = 1
      "0000001" when "00011001001001000", -- t[12872] = 1
      "0000001" when "00011001001001001", -- t[12873] = 1
      "0000001" when "00011001001001010", -- t[12874] = 1
      "0000001" when "00011001001001011", -- t[12875] = 1
      "0000001" when "00011001001001100", -- t[12876] = 1
      "0000001" when "00011001001001101", -- t[12877] = 1
      "0000001" when "00011001001001110", -- t[12878] = 1
      "0000001" when "00011001001001111", -- t[12879] = 1
      "0000001" when "00011001001010000", -- t[12880] = 1
      "0000001" when "00011001001010001", -- t[12881] = 1
      "0000001" when "00011001001010010", -- t[12882] = 1
      "0000001" when "00011001001010011", -- t[12883] = 1
      "0000001" when "00011001001010100", -- t[12884] = 1
      "0000001" when "00011001001010101", -- t[12885] = 1
      "0000001" when "00011001001010110", -- t[12886] = 1
      "0000001" when "00011001001010111", -- t[12887] = 1
      "0000001" when "00011001001011000", -- t[12888] = 1
      "0000001" when "00011001001011001", -- t[12889] = 1
      "0000001" when "00011001001011010", -- t[12890] = 1
      "0000001" when "00011001001011011", -- t[12891] = 1
      "0000001" when "00011001001011100", -- t[12892] = 1
      "0000001" when "00011001001011101", -- t[12893] = 1
      "0000001" when "00011001001011110", -- t[12894] = 1
      "0000001" when "00011001001011111", -- t[12895] = 1
      "0000001" when "00011001001100000", -- t[12896] = 1
      "0000001" when "00011001001100001", -- t[12897] = 1
      "0000001" when "00011001001100010", -- t[12898] = 1
      "0000001" when "00011001001100011", -- t[12899] = 1
      "0000001" when "00011001001100100", -- t[12900] = 1
      "0000001" when "00011001001100101", -- t[12901] = 1
      "0000001" when "00011001001100110", -- t[12902] = 1
      "0000001" when "00011001001100111", -- t[12903] = 1
      "0000001" when "00011001001101000", -- t[12904] = 1
      "0000001" when "00011001001101001", -- t[12905] = 1
      "0000001" when "00011001001101010", -- t[12906] = 1
      "0000001" when "00011001001101011", -- t[12907] = 1
      "0000001" when "00011001001101100", -- t[12908] = 1
      "0000001" when "00011001001101101", -- t[12909] = 1
      "0000001" when "00011001001101110", -- t[12910] = 1
      "0000001" when "00011001001101111", -- t[12911] = 1
      "0000001" when "00011001001110000", -- t[12912] = 1
      "0000001" when "00011001001110001", -- t[12913] = 1
      "0000001" when "00011001001110010", -- t[12914] = 1
      "0000001" when "00011001001110011", -- t[12915] = 1
      "0000001" when "00011001001110100", -- t[12916] = 1
      "0000001" when "00011001001110101", -- t[12917] = 1
      "0000001" when "00011001001110110", -- t[12918] = 1
      "0000001" when "00011001001110111", -- t[12919] = 1
      "0000001" when "00011001001111000", -- t[12920] = 1
      "0000001" when "00011001001111001", -- t[12921] = 1
      "0000001" when "00011001001111010", -- t[12922] = 1
      "0000001" when "00011001001111011", -- t[12923] = 1
      "0000001" when "00011001001111100", -- t[12924] = 1
      "0000001" when "00011001001111101", -- t[12925] = 1
      "0000001" when "00011001001111110", -- t[12926] = 1
      "0000001" when "00011001001111111", -- t[12927] = 1
      "0000001" when "00011001010000000", -- t[12928] = 1
      "0000001" when "00011001010000001", -- t[12929] = 1
      "0000001" when "00011001010000010", -- t[12930] = 1
      "0000001" when "00011001010000011", -- t[12931] = 1
      "0000001" when "00011001010000100", -- t[12932] = 1
      "0000001" when "00011001010000101", -- t[12933] = 1
      "0000001" when "00011001010000110", -- t[12934] = 1
      "0000001" when "00011001010000111", -- t[12935] = 1
      "0000001" when "00011001010001000", -- t[12936] = 1
      "0000001" when "00011001010001001", -- t[12937] = 1
      "0000001" when "00011001010001010", -- t[12938] = 1
      "0000001" when "00011001010001011", -- t[12939] = 1
      "0000001" when "00011001010001100", -- t[12940] = 1
      "0000001" when "00011001010001101", -- t[12941] = 1
      "0000001" when "00011001010001110", -- t[12942] = 1
      "0000001" when "00011001010001111", -- t[12943] = 1
      "0000001" when "00011001010010000", -- t[12944] = 1
      "0000001" when "00011001010010001", -- t[12945] = 1
      "0000001" when "00011001010010010", -- t[12946] = 1
      "0000001" when "00011001010010011", -- t[12947] = 1
      "0000001" when "00011001010010100", -- t[12948] = 1
      "0000001" when "00011001010010101", -- t[12949] = 1
      "0000001" when "00011001010010110", -- t[12950] = 1
      "0000001" when "00011001010010111", -- t[12951] = 1
      "0000001" when "00011001010011000", -- t[12952] = 1
      "0000001" when "00011001010011001", -- t[12953] = 1
      "0000001" when "00011001010011010", -- t[12954] = 1
      "0000001" when "00011001010011011", -- t[12955] = 1
      "0000001" when "00011001010011100", -- t[12956] = 1
      "0000001" when "00011001010011101", -- t[12957] = 1
      "0000001" when "00011001010011110", -- t[12958] = 1
      "0000001" when "00011001010011111", -- t[12959] = 1
      "0000001" when "00011001010100000", -- t[12960] = 1
      "0000001" when "00011001010100001", -- t[12961] = 1
      "0000001" when "00011001010100010", -- t[12962] = 1
      "0000001" when "00011001010100011", -- t[12963] = 1
      "0000001" when "00011001010100100", -- t[12964] = 1
      "0000001" when "00011001010100101", -- t[12965] = 1
      "0000001" when "00011001010100110", -- t[12966] = 1
      "0000001" when "00011001010100111", -- t[12967] = 1
      "0000001" when "00011001010101000", -- t[12968] = 1
      "0000001" when "00011001010101001", -- t[12969] = 1
      "0000001" when "00011001010101010", -- t[12970] = 1
      "0000001" when "00011001010101011", -- t[12971] = 1
      "0000001" when "00011001010101100", -- t[12972] = 1
      "0000001" when "00011001010101101", -- t[12973] = 1
      "0000001" when "00011001010101110", -- t[12974] = 1
      "0000001" when "00011001010101111", -- t[12975] = 1
      "0000001" when "00011001010110000", -- t[12976] = 1
      "0000001" when "00011001010110001", -- t[12977] = 1
      "0000001" when "00011001010110010", -- t[12978] = 1
      "0000001" when "00011001010110011", -- t[12979] = 1
      "0000001" when "00011001010110100", -- t[12980] = 1
      "0000001" when "00011001010110101", -- t[12981] = 1
      "0000001" when "00011001010110110", -- t[12982] = 1
      "0000001" when "00011001010110111", -- t[12983] = 1
      "0000001" when "00011001010111000", -- t[12984] = 1
      "0000001" when "00011001010111001", -- t[12985] = 1
      "0000001" when "00011001010111010", -- t[12986] = 1
      "0000001" when "00011001010111011", -- t[12987] = 1
      "0000001" when "00011001010111100", -- t[12988] = 1
      "0000001" when "00011001010111101", -- t[12989] = 1
      "0000001" when "00011001010111110", -- t[12990] = 1
      "0000001" when "00011001010111111", -- t[12991] = 1
      "0000001" when "00011001011000000", -- t[12992] = 1
      "0000001" when "00011001011000001", -- t[12993] = 1
      "0000001" when "00011001011000010", -- t[12994] = 1
      "0000001" when "00011001011000011", -- t[12995] = 1
      "0000001" when "00011001011000100", -- t[12996] = 1
      "0000001" when "00011001011000101", -- t[12997] = 1
      "0000001" when "00011001011000110", -- t[12998] = 1
      "0000001" when "00011001011000111", -- t[12999] = 1
      "0000001" when "00011001011001000", -- t[13000] = 1
      "0000001" when "00011001011001001", -- t[13001] = 1
      "0000001" when "00011001011001010", -- t[13002] = 1
      "0000001" when "00011001011001011", -- t[13003] = 1
      "0000001" when "00011001011001100", -- t[13004] = 1
      "0000001" when "00011001011001101", -- t[13005] = 1
      "0000001" when "00011001011001110", -- t[13006] = 1
      "0000001" when "00011001011001111", -- t[13007] = 1
      "0000001" when "00011001011010000", -- t[13008] = 1
      "0000001" when "00011001011010001", -- t[13009] = 1
      "0000001" when "00011001011010010", -- t[13010] = 1
      "0000001" when "00011001011010011", -- t[13011] = 1
      "0000001" when "00011001011010100", -- t[13012] = 1
      "0000001" when "00011001011010101", -- t[13013] = 1
      "0000001" when "00011001011010110", -- t[13014] = 1
      "0000001" when "00011001011010111", -- t[13015] = 1
      "0000001" when "00011001011011000", -- t[13016] = 1
      "0000001" when "00011001011011001", -- t[13017] = 1
      "0000001" when "00011001011011010", -- t[13018] = 1
      "0000001" when "00011001011011011", -- t[13019] = 1
      "0000001" when "00011001011011100", -- t[13020] = 1
      "0000001" when "00011001011011101", -- t[13021] = 1
      "0000001" when "00011001011011110", -- t[13022] = 1
      "0000001" when "00011001011011111", -- t[13023] = 1
      "0000001" when "00011001011100000", -- t[13024] = 1
      "0000001" when "00011001011100001", -- t[13025] = 1
      "0000001" when "00011001011100010", -- t[13026] = 1
      "0000001" when "00011001011100011", -- t[13027] = 1
      "0000001" when "00011001011100100", -- t[13028] = 1
      "0000001" when "00011001011100101", -- t[13029] = 1
      "0000001" when "00011001011100110", -- t[13030] = 1
      "0000001" when "00011001011100111", -- t[13031] = 1
      "0000001" when "00011001011101000", -- t[13032] = 1
      "0000001" when "00011001011101001", -- t[13033] = 1
      "0000001" when "00011001011101010", -- t[13034] = 1
      "0000001" when "00011001011101011", -- t[13035] = 1
      "0000001" when "00011001011101100", -- t[13036] = 1
      "0000001" when "00011001011101101", -- t[13037] = 1
      "0000001" when "00011001011101110", -- t[13038] = 1
      "0000001" when "00011001011101111", -- t[13039] = 1
      "0000001" when "00011001011110000", -- t[13040] = 1
      "0000001" when "00011001011110001", -- t[13041] = 1
      "0000001" when "00011001011110010", -- t[13042] = 1
      "0000001" when "00011001011110011", -- t[13043] = 1
      "0000001" when "00011001011110100", -- t[13044] = 1
      "0000001" when "00011001011110101", -- t[13045] = 1
      "0000001" when "00011001011110110", -- t[13046] = 1
      "0000001" when "00011001011110111", -- t[13047] = 1
      "0000001" when "00011001011111000", -- t[13048] = 1
      "0000001" when "00011001011111001", -- t[13049] = 1
      "0000001" when "00011001011111010", -- t[13050] = 1
      "0000001" when "00011001011111011", -- t[13051] = 1
      "0000001" when "00011001011111100", -- t[13052] = 1
      "0000001" when "00011001011111101", -- t[13053] = 1
      "0000001" when "00011001011111110", -- t[13054] = 1
      "0000001" when "00011001011111111", -- t[13055] = 1
      "0000001" when "00011001100000000", -- t[13056] = 1
      "0000001" when "00011001100000001", -- t[13057] = 1
      "0000001" when "00011001100000010", -- t[13058] = 1
      "0000001" when "00011001100000011", -- t[13059] = 1
      "0000001" when "00011001100000100", -- t[13060] = 1
      "0000001" when "00011001100000101", -- t[13061] = 1
      "0000001" when "00011001100000110", -- t[13062] = 1
      "0000001" when "00011001100000111", -- t[13063] = 1
      "0000001" when "00011001100001000", -- t[13064] = 1
      "0000001" when "00011001100001001", -- t[13065] = 1
      "0000001" when "00011001100001010", -- t[13066] = 1
      "0000001" when "00011001100001011", -- t[13067] = 1
      "0000001" when "00011001100001100", -- t[13068] = 1
      "0000001" when "00011001100001101", -- t[13069] = 1
      "0000001" when "00011001100001110", -- t[13070] = 1
      "0000001" when "00011001100001111", -- t[13071] = 1
      "0000001" when "00011001100010000", -- t[13072] = 1
      "0000001" when "00011001100010001", -- t[13073] = 1
      "0000001" when "00011001100010010", -- t[13074] = 1
      "0000001" when "00011001100010011", -- t[13075] = 1
      "0000001" when "00011001100010100", -- t[13076] = 1
      "0000001" when "00011001100010101", -- t[13077] = 1
      "0000001" when "00011001100010110", -- t[13078] = 1
      "0000001" when "00011001100010111", -- t[13079] = 1
      "0000001" when "00011001100011000", -- t[13080] = 1
      "0000001" when "00011001100011001", -- t[13081] = 1
      "0000001" when "00011001100011010", -- t[13082] = 1
      "0000001" when "00011001100011011", -- t[13083] = 1
      "0000001" when "00011001100011100", -- t[13084] = 1
      "0000001" when "00011001100011101", -- t[13085] = 1
      "0000001" when "00011001100011110", -- t[13086] = 1
      "0000001" when "00011001100011111", -- t[13087] = 1
      "0000001" when "00011001100100000", -- t[13088] = 1
      "0000001" when "00011001100100001", -- t[13089] = 1
      "0000001" when "00011001100100010", -- t[13090] = 1
      "0000001" when "00011001100100011", -- t[13091] = 1
      "0000001" when "00011001100100100", -- t[13092] = 1
      "0000001" when "00011001100100101", -- t[13093] = 1
      "0000001" when "00011001100100110", -- t[13094] = 1
      "0000001" when "00011001100100111", -- t[13095] = 1
      "0000001" when "00011001100101000", -- t[13096] = 1
      "0000001" when "00011001100101001", -- t[13097] = 1
      "0000001" when "00011001100101010", -- t[13098] = 1
      "0000001" when "00011001100101011", -- t[13099] = 1
      "0000001" when "00011001100101100", -- t[13100] = 1
      "0000001" when "00011001100101101", -- t[13101] = 1
      "0000001" when "00011001100101110", -- t[13102] = 1
      "0000001" when "00011001100101111", -- t[13103] = 1
      "0000001" when "00011001100110000", -- t[13104] = 1
      "0000001" when "00011001100110001", -- t[13105] = 1
      "0000001" when "00011001100110010", -- t[13106] = 1
      "0000001" when "00011001100110011", -- t[13107] = 1
      "0000001" when "00011001100110100", -- t[13108] = 1
      "0000001" when "00011001100110101", -- t[13109] = 1
      "0000001" when "00011001100110110", -- t[13110] = 1
      "0000001" when "00011001100110111", -- t[13111] = 1
      "0000001" when "00011001100111000", -- t[13112] = 1
      "0000001" when "00011001100111001", -- t[13113] = 1
      "0000001" when "00011001100111010", -- t[13114] = 1
      "0000001" when "00011001100111011", -- t[13115] = 1
      "0000001" when "00011001100111100", -- t[13116] = 1
      "0000001" when "00011001100111101", -- t[13117] = 1
      "0000001" when "00011001100111110", -- t[13118] = 1
      "0000001" when "00011001100111111", -- t[13119] = 1
      "0000001" when "00011001101000000", -- t[13120] = 1
      "0000001" when "00011001101000001", -- t[13121] = 1
      "0000001" when "00011001101000010", -- t[13122] = 1
      "0000001" when "00011001101000011", -- t[13123] = 1
      "0000001" when "00011001101000100", -- t[13124] = 1
      "0000001" when "00011001101000101", -- t[13125] = 1
      "0000001" when "00011001101000110", -- t[13126] = 1
      "0000001" when "00011001101000111", -- t[13127] = 1
      "0000001" when "00011001101001000", -- t[13128] = 1
      "0000001" when "00011001101001001", -- t[13129] = 1
      "0000001" when "00011001101001010", -- t[13130] = 1
      "0000001" when "00011001101001011", -- t[13131] = 1
      "0000001" when "00011001101001100", -- t[13132] = 1
      "0000001" when "00011001101001101", -- t[13133] = 1
      "0000001" when "00011001101001110", -- t[13134] = 1
      "0000001" when "00011001101001111", -- t[13135] = 1
      "0000001" when "00011001101010000", -- t[13136] = 1
      "0000001" when "00011001101010001", -- t[13137] = 1
      "0000001" when "00011001101010010", -- t[13138] = 1
      "0000001" when "00011001101010011", -- t[13139] = 1
      "0000001" when "00011001101010100", -- t[13140] = 1
      "0000001" when "00011001101010101", -- t[13141] = 1
      "0000001" when "00011001101010110", -- t[13142] = 1
      "0000001" when "00011001101010111", -- t[13143] = 1
      "0000001" when "00011001101011000", -- t[13144] = 1
      "0000001" when "00011001101011001", -- t[13145] = 1
      "0000001" when "00011001101011010", -- t[13146] = 1
      "0000001" when "00011001101011011", -- t[13147] = 1
      "0000001" when "00011001101011100", -- t[13148] = 1
      "0000001" when "00011001101011101", -- t[13149] = 1
      "0000001" when "00011001101011110", -- t[13150] = 1
      "0000001" when "00011001101011111", -- t[13151] = 1
      "0000001" when "00011001101100000", -- t[13152] = 1
      "0000001" when "00011001101100001", -- t[13153] = 1
      "0000001" when "00011001101100010", -- t[13154] = 1
      "0000001" when "00011001101100011", -- t[13155] = 1
      "0000001" when "00011001101100100", -- t[13156] = 1
      "0000001" when "00011001101100101", -- t[13157] = 1
      "0000001" when "00011001101100110", -- t[13158] = 1
      "0000001" when "00011001101100111", -- t[13159] = 1
      "0000001" when "00011001101101000", -- t[13160] = 1
      "0000001" when "00011001101101001", -- t[13161] = 1
      "0000001" when "00011001101101010", -- t[13162] = 1
      "0000001" when "00011001101101011", -- t[13163] = 1
      "0000001" when "00011001101101100", -- t[13164] = 1
      "0000001" when "00011001101101101", -- t[13165] = 1
      "0000001" when "00011001101101110", -- t[13166] = 1
      "0000001" when "00011001101101111", -- t[13167] = 1
      "0000001" when "00011001101110000", -- t[13168] = 1
      "0000001" when "00011001101110001", -- t[13169] = 1
      "0000001" when "00011001101110010", -- t[13170] = 1
      "0000001" when "00011001101110011", -- t[13171] = 1
      "0000001" when "00011001101110100", -- t[13172] = 1
      "0000001" when "00011001101110101", -- t[13173] = 1
      "0000001" when "00011001101110110", -- t[13174] = 1
      "0000001" when "00011001101110111", -- t[13175] = 1
      "0000001" when "00011001101111000", -- t[13176] = 1
      "0000001" when "00011001101111001", -- t[13177] = 1
      "0000001" when "00011001101111010", -- t[13178] = 1
      "0000001" when "00011001101111011", -- t[13179] = 1
      "0000001" when "00011001101111100", -- t[13180] = 1
      "0000001" when "00011001101111101", -- t[13181] = 1
      "0000001" when "00011001101111110", -- t[13182] = 1
      "0000001" when "00011001101111111", -- t[13183] = 1
      "0000001" when "00011001110000000", -- t[13184] = 1
      "0000001" when "00011001110000001", -- t[13185] = 1
      "0000001" when "00011001110000010", -- t[13186] = 1
      "0000001" when "00011001110000011", -- t[13187] = 1
      "0000001" when "00011001110000100", -- t[13188] = 1
      "0000001" when "00011001110000101", -- t[13189] = 1
      "0000001" when "00011001110000110", -- t[13190] = 1
      "0000001" when "00011001110000111", -- t[13191] = 1
      "0000001" when "00011001110001000", -- t[13192] = 1
      "0000001" when "00011001110001001", -- t[13193] = 1
      "0000001" when "00011001110001010", -- t[13194] = 1
      "0000001" when "00011001110001011", -- t[13195] = 1
      "0000001" when "00011001110001100", -- t[13196] = 1
      "0000001" when "00011001110001101", -- t[13197] = 1
      "0000001" when "00011001110001110", -- t[13198] = 1
      "0000001" when "00011001110001111", -- t[13199] = 1
      "0000001" when "00011001110010000", -- t[13200] = 1
      "0000001" when "00011001110010001", -- t[13201] = 1
      "0000001" when "00011001110010010", -- t[13202] = 1
      "0000001" when "00011001110010011", -- t[13203] = 1
      "0000001" when "00011001110010100", -- t[13204] = 1
      "0000001" when "00011001110010101", -- t[13205] = 1
      "0000001" when "00011001110010110", -- t[13206] = 1
      "0000001" when "00011001110010111", -- t[13207] = 1
      "0000001" when "00011001110011000", -- t[13208] = 1
      "0000001" when "00011001110011001", -- t[13209] = 1
      "0000001" when "00011001110011010", -- t[13210] = 1
      "0000001" when "00011001110011011", -- t[13211] = 1
      "0000001" when "00011001110011100", -- t[13212] = 1
      "0000001" when "00011001110011101", -- t[13213] = 1
      "0000001" when "00011001110011110", -- t[13214] = 1
      "0000001" when "00011001110011111", -- t[13215] = 1
      "0000001" when "00011001110100000", -- t[13216] = 1
      "0000001" when "00011001110100001", -- t[13217] = 1
      "0000001" when "00011001110100010", -- t[13218] = 1
      "0000001" when "00011001110100011", -- t[13219] = 1
      "0000001" when "00011001110100100", -- t[13220] = 1
      "0000001" when "00011001110100101", -- t[13221] = 1
      "0000001" when "00011001110100110", -- t[13222] = 1
      "0000001" when "00011001110100111", -- t[13223] = 1
      "0000001" when "00011001110101000", -- t[13224] = 1
      "0000001" when "00011001110101001", -- t[13225] = 1
      "0000001" when "00011001110101010", -- t[13226] = 1
      "0000001" when "00011001110101011", -- t[13227] = 1
      "0000001" when "00011001110101100", -- t[13228] = 1
      "0000001" when "00011001110101101", -- t[13229] = 1
      "0000001" when "00011001110101110", -- t[13230] = 1
      "0000001" when "00011001110101111", -- t[13231] = 1
      "0000001" when "00011001110110000", -- t[13232] = 1
      "0000001" when "00011001110110001", -- t[13233] = 1
      "0000001" when "00011001110110010", -- t[13234] = 1
      "0000001" when "00011001110110011", -- t[13235] = 1
      "0000001" when "00011001110110100", -- t[13236] = 1
      "0000001" when "00011001110110101", -- t[13237] = 1
      "0000001" when "00011001110110110", -- t[13238] = 1
      "0000001" when "00011001110110111", -- t[13239] = 1
      "0000001" when "00011001110111000", -- t[13240] = 1
      "0000001" when "00011001110111001", -- t[13241] = 1
      "0000001" when "00011001110111010", -- t[13242] = 1
      "0000001" when "00011001110111011", -- t[13243] = 1
      "0000001" when "00011001110111100", -- t[13244] = 1
      "0000001" when "00011001110111101", -- t[13245] = 1
      "0000001" when "00011001110111110", -- t[13246] = 1
      "0000001" when "00011001110111111", -- t[13247] = 1
      "0000001" when "00011001111000000", -- t[13248] = 1
      "0000001" when "00011001111000001", -- t[13249] = 1
      "0000001" when "00011001111000010", -- t[13250] = 1
      "0000001" when "00011001111000011", -- t[13251] = 1
      "0000001" when "00011001111000100", -- t[13252] = 1
      "0000001" when "00011001111000101", -- t[13253] = 1
      "0000001" when "00011001111000110", -- t[13254] = 1
      "0000001" when "00011001111000111", -- t[13255] = 1
      "0000001" when "00011001111001000", -- t[13256] = 1
      "0000001" when "00011001111001001", -- t[13257] = 1
      "0000001" when "00011001111001010", -- t[13258] = 1
      "0000001" when "00011001111001011", -- t[13259] = 1
      "0000001" when "00011001111001100", -- t[13260] = 1
      "0000001" when "00011001111001101", -- t[13261] = 1
      "0000001" when "00011001111001110", -- t[13262] = 1
      "0000001" when "00011001111001111", -- t[13263] = 1
      "0000001" when "00011001111010000", -- t[13264] = 1
      "0000001" when "00011001111010001", -- t[13265] = 1
      "0000001" when "00011001111010010", -- t[13266] = 1
      "0000001" when "00011001111010011", -- t[13267] = 1
      "0000001" when "00011001111010100", -- t[13268] = 1
      "0000001" when "00011001111010101", -- t[13269] = 1
      "0000001" when "00011001111010110", -- t[13270] = 1
      "0000001" when "00011001111010111", -- t[13271] = 1
      "0000001" when "00011001111011000", -- t[13272] = 1
      "0000001" when "00011001111011001", -- t[13273] = 1
      "0000001" when "00011001111011010", -- t[13274] = 1
      "0000001" when "00011001111011011", -- t[13275] = 1
      "0000001" when "00011001111011100", -- t[13276] = 1
      "0000001" when "00011001111011101", -- t[13277] = 1
      "0000001" when "00011001111011110", -- t[13278] = 1
      "0000001" when "00011001111011111", -- t[13279] = 1
      "0000001" when "00011001111100000", -- t[13280] = 1
      "0000001" when "00011001111100001", -- t[13281] = 1
      "0000001" when "00011001111100010", -- t[13282] = 1
      "0000001" when "00011001111100011", -- t[13283] = 1
      "0000001" when "00011001111100100", -- t[13284] = 1
      "0000001" when "00011001111100101", -- t[13285] = 1
      "0000001" when "00011001111100110", -- t[13286] = 1
      "0000001" when "00011001111100111", -- t[13287] = 1
      "0000001" when "00011001111101000", -- t[13288] = 1
      "0000001" when "00011001111101001", -- t[13289] = 1
      "0000001" when "00011001111101010", -- t[13290] = 1
      "0000001" when "00011001111101011", -- t[13291] = 1
      "0000001" when "00011001111101100", -- t[13292] = 1
      "0000001" when "00011001111101101", -- t[13293] = 1
      "0000001" when "00011001111101110", -- t[13294] = 1
      "0000001" when "00011001111101111", -- t[13295] = 1
      "0000001" when "00011001111110000", -- t[13296] = 1
      "0000001" when "00011001111110001", -- t[13297] = 1
      "0000001" when "00011001111110010", -- t[13298] = 1
      "0000001" when "00011001111110011", -- t[13299] = 1
      "0000001" when "00011001111110100", -- t[13300] = 1
      "0000001" when "00011001111110101", -- t[13301] = 1
      "0000001" when "00011001111110110", -- t[13302] = 1
      "0000001" when "00011001111110111", -- t[13303] = 1
      "0000001" when "00011001111111000", -- t[13304] = 1
      "0000001" when "00011001111111001", -- t[13305] = 1
      "0000001" when "00011001111111010", -- t[13306] = 1
      "0000001" when "00011001111111011", -- t[13307] = 1
      "0000001" when "00011001111111100", -- t[13308] = 1
      "0000001" when "00011001111111101", -- t[13309] = 1
      "0000001" when "00011001111111110", -- t[13310] = 1
      "0000001" when "00011001111111111", -- t[13311] = 1
      "0000001" when "00011010000000000", -- t[13312] = 1
      "0000001" when "00011010000000001", -- t[13313] = 1
      "0000001" when "00011010000000010", -- t[13314] = 1
      "0000001" when "00011010000000011", -- t[13315] = 1
      "0000001" when "00011010000000100", -- t[13316] = 1
      "0000001" when "00011010000000101", -- t[13317] = 1
      "0000001" when "00011010000000110", -- t[13318] = 1
      "0000001" when "00011010000000111", -- t[13319] = 1
      "0000001" when "00011010000001000", -- t[13320] = 1
      "0000001" when "00011010000001001", -- t[13321] = 1
      "0000001" when "00011010000001010", -- t[13322] = 1
      "0000001" when "00011010000001011", -- t[13323] = 1
      "0000001" when "00011010000001100", -- t[13324] = 1
      "0000001" when "00011010000001101", -- t[13325] = 1
      "0000001" when "00011010000001110", -- t[13326] = 1
      "0000001" when "00011010000001111", -- t[13327] = 1
      "0000001" when "00011010000010000", -- t[13328] = 1
      "0000001" when "00011010000010001", -- t[13329] = 1
      "0000001" when "00011010000010010", -- t[13330] = 1
      "0000001" when "00011010000010011", -- t[13331] = 1
      "0000001" when "00011010000010100", -- t[13332] = 1
      "0000001" when "00011010000010101", -- t[13333] = 1
      "0000001" when "00011010000010110", -- t[13334] = 1
      "0000001" when "00011010000010111", -- t[13335] = 1
      "0000001" when "00011010000011000", -- t[13336] = 1
      "0000001" when "00011010000011001", -- t[13337] = 1
      "0000001" when "00011010000011010", -- t[13338] = 1
      "0000001" when "00011010000011011", -- t[13339] = 1
      "0000001" when "00011010000011100", -- t[13340] = 1
      "0000001" when "00011010000011101", -- t[13341] = 1
      "0000001" when "00011010000011110", -- t[13342] = 1
      "0000001" when "00011010000011111", -- t[13343] = 1
      "0000001" when "00011010000100000", -- t[13344] = 1
      "0000001" when "00011010000100001", -- t[13345] = 1
      "0000001" when "00011010000100010", -- t[13346] = 1
      "0000001" when "00011010000100011", -- t[13347] = 1
      "0000001" when "00011010000100100", -- t[13348] = 1
      "0000001" when "00011010000100101", -- t[13349] = 1
      "0000001" when "00011010000100110", -- t[13350] = 1
      "0000001" when "00011010000100111", -- t[13351] = 1
      "0000001" when "00011010000101000", -- t[13352] = 1
      "0000001" when "00011010000101001", -- t[13353] = 1
      "0000001" when "00011010000101010", -- t[13354] = 1
      "0000001" when "00011010000101011", -- t[13355] = 1
      "0000001" when "00011010000101100", -- t[13356] = 1
      "0000001" when "00011010000101101", -- t[13357] = 1
      "0000001" when "00011010000101110", -- t[13358] = 1
      "0000001" when "00011010000101111", -- t[13359] = 1
      "0000001" when "00011010000110000", -- t[13360] = 1
      "0000001" when "00011010000110001", -- t[13361] = 1
      "0000001" when "00011010000110010", -- t[13362] = 1
      "0000001" when "00011010000110011", -- t[13363] = 1
      "0000001" when "00011010000110100", -- t[13364] = 1
      "0000001" when "00011010000110101", -- t[13365] = 1
      "0000001" when "00011010000110110", -- t[13366] = 1
      "0000001" when "00011010000110111", -- t[13367] = 1
      "0000001" when "00011010000111000", -- t[13368] = 1
      "0000001" when "00011010000111001", -- t[13369] = 1
      "0000001" when "00011010000111010", -- t[13370] = 1
      "0000001" when "00011010000111011", -- t[13371] = 1
      "0000001" when "00011010000111100", -- t[13372] = 1
      "0000001" when "00011010000111101", -- t[13373] = 1
      "0000001" when "00011010000111110", -- t[13374] = 1
      "0000001" when "00011010000111111", -- t[13375] = 1
      "0000001" when "00011010001000000", -- t[13376] = 1
      "0000001" when "00011010001000001", -- t[13377] = 1
      "0000001" when "00011010001000010", -- t[13378] = 1
      "0000001" when "00011010001000011", -- t[13379] = 1
      "0000001" when "00011010001000100", -- t[13380] = 1
      "0000001" when "00011010001000101", -- t[13381] = 1
      "0000001" when "00011010001000110", -- t[13382] = 1
      "0000001" when "00011010001000111", -- t[13383] = 1
      "0000001" when "00011010001001000", -- t[13384] = 1
      "0000001" when "00011010001001001", -- t[13385] = 1
      "0000001" when "00011010001001010", -- t[13386] = 1
      "0000001" when "00011010001001011", -- t[13387] = 1
      "0000001" when "00011010001001100", -- t[13388] = 1
      "0000001" when "00011010001001101", -- t[13389] = 1
      "0000001" when "00011010001001110", -- t[13390] = 1
      "0000001" when "00011010001001111", -- t[13391] = 1
      "0000001" when "00011010001010000", -- t[13392] = 1
      "0000001" when "00011010001010001", -- t[13393] = 1
      "0000001" when "00011010001010010", -- t[13394] = 1
      "0000001" when "00011010001010011", -- t[13395] = 1
      "0000001" when "00011010001010100", -- t[13396] = 1
      "0000001" when "00011010001010101", -- t[13397] = 1
      "0000001" when "00011010001010110", -- t[13398] = 1
      "0000001" when "00011010001010111", -- t[13399] = 1
      "0000001" when "00011010001011000", -- t[13400] = 1
      "0000001" when "00011010001011001", -- t[13401] = 1
      "0000001" when "00011010001011010", -- t[13402] = 1
      "0000001" when "00011010001011011", -- t[13403] = 1
      "0000001" when "00011010001011100", -- t[13404] = 1
      "0000001" when "00011010001011101", -- t[13405] = 1
      "0000001" when "00011010001011110", -- t[13406] = 1
      "0000001" when "00011010001011111", -- t[13407] = 1
      "0000001" when "00011010001100000", -- t[13408] = 1
      "0000001" when "00011010001100001", -- t[13409] = 1
      "0000001" when "00011010001100010", -- t[13410] = 1
      "0000001" when "00011010001100011", -- t[13411] = 1
      "0000001" when "00011010001100100", -- t[13412] = 1
      "0000001" when "00011010001100101", -- t[13413] = 1
      "0000001" when "00011010001100110", -- t[13414] = 1
      "0000001" when "00011010001100111", -- t[13415] = 1
      "0000001" when "00011010001101000", -- t[13416] = 1
      "0000001" when "00011010001101001", -- t[13417] = 1
      "0000001" when "00011010001101010", -- t[13418] = 1
      "0000001" when "00011010001101011", -- t[13419] = 1
      "0000001" when "00011010001101100", -- t[13420] = 1
      "0000001" when "00011010001101101", -- t[13421] = 1
      "0000001" when "00011010001101110", -- t[13422] = 1
      "0000001" when "00011010001101111", -- t[13423] = 1
      "0000001" when "00011010001110000", -- t[13424] = 1
      "0000001" when "00011010001110001", -- t[13425] = 1
      "0000001" when "00011010001110010", -- t[13426] = 1
      "0000001" when "00011010001110011", -- t[13427] = 1
      "0000001" when "00011010001110100", -- t[13428] = 1
      "0000001" when "00011010001110101", -- t[13429] = 1
      "0000001" when "00011010001110110", -- t[13430] = 1
      "0000001" when "00011010001110111", -- t[13431] = 1
      "0000001" when "00011010001111000", -- t[13432] = 1
      "0000001" when "00011010001111001", -- t[13433] = 1
      "0000001" when "00011010001111010", -- t[13434] = 1
      "0000001" when "00011010001111011", -- t[13435] = 1
      "0000001" when "00011010001111100", -- t[13436] = 1
      "0000001" when "00011010001111101", -- t[13437] = 1
      "0000001" when "00011010001111110", -- t[13438] = 1
      "0000001" when "00011010001111111", -- t[13439] = 1
      "0000001" when "00011010010000000", -- t[13440] = 1
      "0000001" when "00011010010000001", -- t[13441] = 1
      "0000001" when "00011010010000010", -- t[13442] = 1
      "0000001" when "00011010010000011", -- t[13443] = 1
      "0000001" when "00011010010000100", -- t[13444] = 1
      "0000001" when "00011010010000101", -- t[13445] = 1
      "0000001" when "00011010010000110", -- t[13446] = 1
      "0000001" when "00011010010000111", -- t[13447] = 1
      "0000001" when "00011010010001000", -- t[13448] = 1
      "0000001" when "00011010010001001", -- t[13449] = 1
      "0000001" when "00011010010001010", -- t[13450] = 1
      "0000001" when "00011010010001011", -- t[13451] = 1
      "0000001" when "00011010010001100", -- t[13452] = 1
      "0000001" when "00011010010001101", -- t[13453] = 1
      "0000001" when "00011010010001110", -- t[13454] = 1
      "0000001" when "00011010010001111", -- t[13455] = 1
      "0000001" when "00011010010010000", -- t[13456] = 1
      "0000001" when "00011010010010001", -- t[13457] = 1
      "0000001" when "00011010010010010", -- t[13458] = 1
      "0000001" when "00011010010010011", -- t[13459] = 1
      "0000001" when "00011010010010100", -- t[13460] = 1
      "0000001" when "00011010010010101", -- t[13461] = 1
      "0000001" when "00011010010010110", -- t[13462] = 1
      "0000001" when "00011010010010111", -- t[13463] = 1
      "0000001" when "00011010010011000", -- t[13464] = 1
      "0000001" when "00011010010011001", -- t[13465] = 1
      "0000001" when "00011010010011010", -- t[13466] = 1
      "0000001" when "00011010010011011", -- t[13467] = 1
      "0000001" when "00011010010011100", -- t[13468] = 1
      "0000001" when "00011010010011101", -- t[13469] = 1
      "0000001" when "00011010010011110", -- t[13470] = 1
      "0000001" when "00011010010011111", -- t[13471] = 1
      "0000001" when "00011010010100000", -- t[13472] = 1
      "0000001" when "00011010010100001", -- t[13473] = 1
      "0000001" when "00011010010100010", -- t[13474] = 1
      "0000001" when "00011010010100011", -- t[13475] = 1
      "0000001" when "00011010010100100", -- t[13476] = 1
      "0000001" when "00011010010100101", -- t[13477] = 1
      "0000001" when "00011010010100110", -- t[13478] = 1
      "0000001" when "00011010010100111", -- t[13479] = 1
      "0000001" when "00011010010101000", -- t[13480] = 1
      "0000001" when "00011010010101001", -- t[13481] = 1
      "0000001" when "00011010010101010", -- t[13482] = 1
      "0000001" when "00011010010101011", -- t[13483] = 1
      "0000001" when "00011010010101100", -- t[13484] = 1
      "0000001" when "00011010010101101", -- t[13485] = 1
      "0000001" when "00011010010101110", -- t[13486] = 1
      "0000001" when "00011010010101111", -- t[13487] = 1
      "0000001" when "00011010010110000", -- t[13488] = 1
      "0000001" when "00011010010110001", -- t[13489] = 1
      "0000001" when "00011010010110010", -- t[13490] = 1
      "0000001" when "00011010010110011", -- t[13491] = 1
      "0000001" when "00011010010110100", -- t[13492] = 1
      "0000001" when "00011010010110101", -- t[13493] = 1
      "0000001" when "00011010010110110", -- t[13494] = 1
      "0000001" when "00011010010110111", -- t[13495] = 1
      "0000001" when "00011010010111000", -- t[13496] = 1
      "0000001" when "00011010010111001", -- t[13497] = 1
      "0000001" when "00011010010111010", -- t[13498] = 1
      "0000001" when "00011010010111011", -- t[13499] = 1
      "0000001" when "00011010010111100", -- t[13500] = 1
      "0000001" when "00011010010111101", -- t[13501] = 1
      "0000001" when "00011010010111110", -- t[13502] = 1
      "0000001" when "00011010010111111", -- t[13503] = 1
      "0000001" when "00011010011000000", -- t[13504] = 1
      "0000001" when "00011010011000001", -- t[13505] = 1
      "0000001" when "00011010011000010", -- t[13506] = 1
      "0000001" when "00011010011000011", -- t[13507] = 1
      "0000001" when "00011010011000100", -- t[13508] = 1
      "0000001" when "00011010011000101", -- t[13509] = 1
      "0000001" when "00011010011000110", -- t[13510] = 1
      "0000001" when "00011010011000111", -- t[13511] = 1
      "0000001" when "00011010011001000", -- t[13512] = 1
      "0000001" when "00011010011001001", -- t[13513] = 1
      "0000001" when "00011010011001010", -- t[13514] = 1
      "0000001" when "00011010011001011", -- t[13515] = 1
      "0000001" when "00011010011001100", -- t[13516] = 1
      "0000001" when "00011010011001101", -- t[13517] = 1
      "0000001" when "00011010011001110", -- t[13518] = 1
      "0000001" when "00011010011001111", -- t[13519] = 1
      "0000001" when "00011010011010000", -- t[13520] = 1
      "0000001" when "00011010011010001", -- t[13521] = 1
      "0000001" when "00011010011010010", -- t[13522] = 1
      "0000001" when "00011010011010011", -- t[13523] = 1
      "0000001" when "00011010011010100", -- t[13524] = 1
      "0000001" when "00011010011010101", -- t[13525] = 1
      "0000001" when "00011010011010110", -- t[13526] = 1
      "0000001" when "00011010011010111", -- t[13527] = 1
      "0000001" when "00011010011011000", -- t[13528] = 1
      "0000001" when "00011010011011001", -- t[13529] = 1
      "0000001" when "00011010011011010", -- t[13530] = 1
      "0000001" when "00011010011011011", -- t[13531] = 1
      "0000001" when "00011010011011100", -- t[13532] = 1
      "0000001" when "00011010011011101", -- t[13533] = 1
      "0000001" when "00011010011011110", -- t[13534] = 1
      "0000001" when "00011010011011111", -- t[13535] = 1
      "0000001" when "00011010011100000", -- t[13536] = 1
      "0000001" when "00011010011100001", -- t[13537] = 1
      "0000001" when "00011010011100010", -- t[13538] = 1
      "0000001" when "00011010011100011", -- t[13539] = 1
      "0000001" when "00011010011100100", -- t[13540] = 1
      "0000001" when "00011010011100101", -- t[13541] = 1
      "0000001" when "00011010011100110", -- t[13542] = 1
      "0000001" when "00011010011100111", -- t[13543] = 1
      "0000001" when "00011010011101000", -- t[13544] = 1
      "0000001" when "00011010011101001", -- t[13545] = 1
      "0000001" when "00011010011101010", -- t[13546] = 1
      "0000001" when "00011010011101011", -- t[13547] = 1
      "0000001" when "00011010011101100", -- t[13548] = 1
      "0000001" when "00011010011101101", -- t[13549] = 1
      "0000001" when "00011010011101110", -- t[13550] = 1
      "0000001" when "00011010011101111", -- t[13551] = 1
      "0000001" when "00011010011110000", -- t[13552] = 1
      "0000001" when "00011010011110001", -- t[13553] = 1
      "0000001" when "00011010011110010", -- t[13554] = 1
      "0000001" when "00011010011110011", -- t[13555] = 1
      "0000001" when "00011010011110100", -- t[13556] = 1
      "0000001" when "00011010011110101", -- t[13557] = 1
      "0000001" when "00011010011110110", -- t[13558] = 1
      "0000001" when "00011010011110111", -- t[13559] = 1
      "0000001" when "00011010011111000", -- t[13560] = 1
      "0000001" when "00011010011111001", -- t[13561] = 1
      "0000001" when "00011010011111010", -- t[13562] = 1
      "0000001" when "00011010011111011", -- t[13563] = 1
      "0000001" when "00011010011111100", -- t[13564] = 1
      "0000001" when "00011010011111101", -- t[13565] = 1
      "0000001" when "00011010011111110", -- t[13566] = 1
      "0000001" when "00011010011111111", -- t[13567] = 1
      "0000001" when "00011010100000000", -- t[13568] = 1
      "0000001" when "00011010100000001", -- t[13569] = 1
      "0000001" when "00011010100000010", -- t[13570] = 1
      "0000001" when "00011010100000011", -- t[13571] = 1
      "0000001" when "00011010100000100", -- t[13572] = 1
      "0000001" when "00011010100000101", -- t[13573] = 1
      "0000001" when "00011010100000110", -- t[13574] = 1
      "0000001" when "00011010100000111", -- t[13575] = 1
      "0000001" when "00011010100001000", -- t[13576] = 1
      "0000001" when "00011010100001001", -- t[13577] = 1
      "0000001" when "00011010100001010", -- t[13578] = 1
      "0000001" when "00011010100001011", -- t[13579] = 1
      "0000001" when "00011010100001100", -- t[13580] = 1
      "0000001" when "00011010100001101", -- t[13581] = 1
      "0000001" when "00011010100001110", -- t[13582] = 1
      "0000001" when "00011010100001111", -- t[13583] = 1
      "0000001" when "00011010100010000", -- t[13584] = 1
      "0000001" when "00011010100010001", -- t[13585] = 1
      "0000001" when "00011010100010010", -- t[13586] = 1
      "0000001" when "00011010100010011", -- t[13587] = 1
      "0000001" when "00011010100010100", -- t[13588] = 1
      "0000001" when "00011010100010101", -- t[13589] = 1
      "0000001" when "00011010100010110", -- t[13590] = 1
      "0000001" when "00011010100010111", -- t[13591] = 1
      "0000001" when "00011010100011000", -- t[13592] = 1
      "0000001" when "00011010100011001", -- t[13593] = 1
      "0000001" when "00011010100011010", -- t[13594] = 1
      "0000001" when "00011010100011011", -- t[13595] = 1
      "0000001" when "00011010100011100", -- t[13596] = 1
      "0000001" when "00011010100011101", -- t[13597] = 1
      "0000001" when "00011010100011110", -- t[13598] = 1
      "0000001" when "00011010100011111", -- t[13599] = 1
      "0000001" when "00011010100100000", -- t[13600] = 1
      "0000001" when "00011010100100001", -- t[13601] = 1
      "0000001" when "00011010100100010", -- t[13602] = 1
      "0000001" when "00011010100100011", -- t[13603] = 1
      "0000001" when "00011010100100100", -- t[13604] = 1
      "0000001" when "00011010100100101", -- t[13605] = 1
      "0000001" when "00011010100100110", -- t[13606] = 1
      "0000001" when "00011010100100111", -- t[13607] = 1
      "0000001" when "00011010100101000", -- t[13608] = 1
      "0000001" when "00011010100101001", -- t[13609] = 1
      "0000001" when "00011010100101010", -- t[13610] = 1
      "0000001" when "00011010100101011", -- t[13611] = 1
      "0000001" when "00011010100101100", -- t[13612] = 1
      "0000001" when "00011010100101101", -- t[13613] = 1
      "0000001" when "00011010100101110", -- t[13614] = 1
      "0000001" when "00011010100101111", -- t[13615] = 1
      "0000001" when "00011010100110000", -- t[13616] = 1
      "0000001" when "00011010100110001", -- t[13617] = 1
      "0000001" when "00011010100110010", -- t[13618] = 1
      "0000001" when "00011010100110011", -- t[13619] = 1
      "0000001" when "00011010100110100", -- t[13620] = 1
      "0000001" when "00011010100110101", -- t[13621] = 1
      "0000001" when "00011010100110110", -- t[13622] = 1
      "0000001" when "00011010100110111", -- t[13623] = 1
      "0000001" when "00011010100111000", -- t[13624] = 1
      "0000001" when "00011010100111001", -- t[13625] = 1
      "0000001" when "00011010100111010", -- t[13626] = 1
      "0000001" when "00011010100111011", -- t[13627] = 1
      "0000001" when "00011010100111100", -- t[13628] = 1
      "0000001" when "00011010100111101", -- t[13629] = 1
      "0000001" when "00011010100111110", -- t[13630] = 1
      "0000001" when "00011010100111111", -- t[13631] = 1
      "0000001" when "00011010101000000", -- t[13632] = 1
      "0000001" when "00011010101000001", -- t[13633] = 1
      "0000001" when "00011010101000010", -- t[13634] = 1
      "0000001" when "00011010101000011", -- t[13635] = 1
      "0000001" when "00011010101000100", -- t[13636] = 1
      "0000001" when "00011010101000101", -- t[13637] = 1
      "0000001" when "00011010101000110", -- t[13638] = 1
      "0000001" when "00011010101000111", -- t[13639] = 1
      "0000001" when "00011010101001000", -- t[13640] = 1
      "0000001" when "00011010101001001", -- t[13641] = 1
      "0000001" when "00011010101001010", -- t[13642] = 1
      "0000001" when "00011010101001011", -- t[13643] = 1
      "0000001" when "00011010101001100", -- t[13644] = 1
      "0000001" when "00011010101001101", -- t[13645] = 1
      "0000001" when "00011010101001110", -- t[13646] = 1
      "0000001" when "00011010101001111", -- t[13647] = 1
      "0000001" when "00011010101010000", -- t[13648] = 1
      "0000001" when "00011010101010001", -- t[13649] = 1
      "0000001" when "00011010101010010", -- t[13650] = 1
      "0000001" when "00011010101010011", -- t[13651] = 1
      "0000001" when "00011010101010100", -- t[13652] = 1
      "0000001" when "00011010101010101", -- t[13653] = 1
      "0000001" when "00011010101010110", -- t[13654] = 1
      "0000001" when "00011010101010111", -- t[13655] = 1
      "0000001" when "00011010101011000", -- t[13656] = 1
      "0000001" when "00011010101011001", -- t[13657] = 1
      "0000001" when "00011010101011010", -- t[13658] = 1
      "0000001" when "00011010101011011", -- t[13659] = 1
      "0000001" when "00011010101011100", -- t[13660] = 1
      "0000001" when "00011010101011101", -- t[13661] = 1
      "0000001" when "00011010101011110", -- t[13662] = 1
      "0000001" when "00011010101011111", -- t[13663] = 1
      "0000001" when "00011010101100000", -- t[13664] = 1
      "0000001" when "00011010101100001", -- t[13665] = 1
      "0000001" when "00011010101100010", -- t[13666] = 1
      "0000001" when "00011010101100011", -- t[13667] = 1
      "0000001" when "00011010101100100", -- t[13668] = 1
      "0000001" when "00011010101100101", -- t[13669] = 1
      "0000001" when "00011010101100110", -- t[13670] = 1
      "0000001" when "00011010101100111", -- t[13671] = 1
      "0000001" when "00011010101101000", -- t[13672] = 1
      "0000001" when "00011010101101001", -- t[13673] = 1
      "0000001" when "00011010101101010", -- t[13674] = 1
      "0000001" when "00011010101101011", -- t[13675] = 1
      "0000001" when "00011010101101100", -- t[13676] = 1
      "0000001" when "00011010101101101", -- t[13677] = 1
      "0000001" when "00011010101101110", -- t[13678] = 1
      "0000001" when "00011010101101111", -- t[13679] = 1
      "0000001" when "00011010101110000", -- t[13680] = 1
      "0000001" when "00011010101110001", -- t[13681] = 1
      "0000001" when "00011010101110010", -- t[13682] = 1
      "0000001" when "00011010101110011", -- t[13683] = 1
      "0000001" when "00011010101110100", -- t[13684] = 1
      "0000001" when "00011010101110101", -- t[13685] = 1
      "0000001" when "00011010101110110", -- t[13686] = 1
      "0000001" when "00011010101110111", -- t[13687] = 1
      "0000001" when "00011010101111000", -- t[13688] = 1
      "0000001" when "00011010101111001", -- t[13689] = 1
      "0000001" when "00011010101111010", -- t[13690] = 1
      "0000001" when "00011010101111011", -- t[13691] = 1
      "0000001" when "00011010101111100", -- t[13692] = 1
      "0000001" when "00011010101111101", -- t[13693] = 1
      "0000001" when "00011010101111110", -- t[13694] = 1
      "0000001" when "00011010101111111", -- t[13695] = 1
      "0000001" when "00011010110000000", -- t[13696] = 1
      "0000001" when "00011010110000001", -- t[13697] = 1
      "0000001" when "00011010110000010", -- t[13698] = 1
      "0000001" when "00011010110000011", -- t[13699] = 1
      "0000001" when "00011010110000100", -- t[13700] = 1
      "0000001" when "00011010110000101", -- t[13701] = 1
      "0000001" when "00011010110000110", -- t[13702] = 1
      "0000001" when "00011010110000111", -- t[13703] = 1
      "0000001" when "00011010110001000", -- t[13704] = 1
      "0000001" when "00011010110001001", -- t[13705] = 1
      "0000001" when "00011010110001010", -- t[13706] = 1
      "0000001" when "00011010110001011", -- t[13707] = 1
      "0000001" when "00011010110001100", -- t[13708] = 1
      "0000001" when "00011010110001101", -- t[13709] = 1
      "0000001" when "00011010110001110", -- t[13710] = 1
      "0000001" when "00011010110001111", -- t[13711] = 1
      "0000001" when "00011010110010000", -- t[13712] = 1
      "0000001" when "00011010110010001", -- t[13713] = 1
      "0000001" when "00011010110010010", -- t[13714] = 1
      "0000001" when "00011010110010011", -- t[13715] = 1
      "0000001" when "00011010110010100", -- t[13716] = 1
      "0000001" when "00011010110010101", -- t[13717] = 1
      "0000001" when "00011010110010110", -- t[13718] = 1
      "0000001" when "00011010110010111", -- t[13719] = 1
      "0000001" when "00011010110011000", -- t[13720] = 1
      "0000001" when "00011010110011001", -- t[13721] = 1
      "0000001" when "00011010110011010", -- t[13722] = 1
      "0000001" when "00011010110011011", -- t[13723] = 1
      "0000001" when "00011010110011100", -- t[13724] = 1
      "0000001" when "00011010110011101", -- t[13725] = 1
      "0000001" when "00011010110011110", -- t[13726] = 1
      "0000001" when "00011010110011111", -- t[13727] = 1
      "0000001" when "00011010110100000", -- t[13728] = 1
      "0000001" when "00011010110100001", -- t[13729] = 1
      "0000001" when "00011010110100010", -- t[13730] = 1
      "0000001" when "00011010110100011", -- t[13731] = 1
      "0000001" when "00011010110100100", -- t[13732] = 1
      "0000001" when "00011010110100101", -- t[13733] = 1
      "0000001" when "00011010110100110", -- t[13734] = 1
      "0000001" when "00011010110100111", -- t[13735] = 1
      "0000001" when "00011010110101000", -- t[13736] = 1
      "0000001" when "00011010110101001", -- t[13737] = 1
      "0000001" when "00011010110101010", -- t[13738] = 1
      "0000001" when "00011010110101011", -- t[13739] = 1
      "0000001" when "00011010110101100", -- t[13740] = 1
      "0000001" when "00011010110101101", -- t[13741] = 1
      "0000001" when "00011010110101110", -- t[13742] = 1
      "0000001" when "00011010110101111", -- t[13743] = 1
      "0000001" when "00011010110110000", -- t[13744] = 1
      "0000001" when "00011010110110001", -- t[13745] = 1
      "0000001" when "00011010110110010", -- t[13746] = 1
      "0000001" when "00011010110110011", -- t[13747] = 1
      "0000001" when "00011010110110100", -- t[13748] = 1
      "0000001" when "00011010110110101", -- t[13749] = 1
      "0000001" when "00011010110110110", -- t[13750] = 1
      "0000001" when "00011010110110111", -- t[13751] = 1
      "0000001" when "00011010110111000", -- t[13752] = 1
      "0000001" when "00011010110111001", -- t[13753] = 1
      "0000001" when "00011010110111010", -- t[13754] = 1
      "0000001" when "00011010110111011", -- t[13755] = 1
      "0000001" when "00011010110111100", -- t[13756] = 1
      "0000001" when "00011010110111101", -- t[13757] = 1
      "0000001" when "00011010110111110", -- t[13758] = 1
      "0000001" when "00011010110111111", -- t[13759] = 1
      "0000001" when "00011010111000000", -- t[13760] = 1
      "0000001" when "00011010111000001", -- t[13761] = 1
      "0000001" when "00011010111000010", -- t[13762] = 1
      "0000001" when "00011010111000011", -- t[13763] = 1
      "0000001" when "00011010111000100", -- t[13764] = 1
      "0000001" when "00011010111000101", -- t[13765] = 1
      "0000001" when "00011010111000110", -- t[13766] = 1
      "0000001" when "00011010111000111", -- t[13767] = 1
      "0000001" when "00011010111001000", -- t[13768] = 1
      "0000001" when "00011010111001001", -- t[13769] = 1
      "0000001" when "00011010111001010", -- t[13770] = 1
      "0000001" when "00011010111001011", -- t[13771] = 1
      "0000001" when "00011010111001100", -- t[13772] = 1
      "0000001" when "00011010111001101", -- t[13773] = 1
      "0000001" when "00011010111001110", -- t[13774] = 1
      "0000001" when "00011010111001111", -- t[13775] = 1
      "0000001" when "00011010111010000", -- t[13776] = 1
      "0000001" when "00011010111010001", -- t[13777] = 1
      "0000001" when "00011010111010010", -- t[13778] = 1
      "0000001" when "00011010111010011", -- t[13779] = 1
      "0000001" when "00011010111010100", -- t[13780] = 1
      "0000001" when "00011010111010101", -- t[13781] = 1
      "0000001" when "00011010111010110", -- t[13782] = 1
      "0000001" when "00011010111010111", -- t[13783] = 1
      "0000001" when "00011010111011000", -- t[13784] = 1
      "0000001" when "00011010111011001", -- t[13785] = 1
      "0000001" when "00011010111011010", -- t[13786] = 1
      "0000001" when "00011010111011011", -- t[13787] = 1
      "0000001" when "00011010111011100", -- t[13788] = 1
      "0000001" when "00011010111011101", -- t[13789] = 1
      "0000001" when "00011010111011110", -- t[13790] = 1
      "0000001" when "00011010111011111", -- t[13791] = 1
      "0000001" when "00011010111100000", -- t[13792] = 1
      "0000001" when "00011010111100001", -- t[13793] = 1
      "0000001" when "00011010111100010", -- t[13794] = 1
      "0000001" when "00011010111100011", -- t[13795] = 1
      "0000001" when "00011010111100100", -- t[13796] = 1
      "0000001" when "00011010111100101", -- t[13797] = 1
      "0000001" when "00011010111100110", -- t[13798] = 1
      "0000001" when "00011010111100111", -- t[13799] = 1
      "0000001" when "00011010111101000", -- t[13800] = 1
      "0000001" when "00011010111101001", -- t[13801] = 1
      "0000001" when "00011010111101010", -- t[13802] = 1
      "0000001" when "00011010111101011", -- t[13803] = 1
      "0000001" when "00011010111101100", -- t[13804] = 1
      "0000001" when "00011010111101101", -- t[13805] = 1
      "0000001" when "00011010111101110", -- t[13806] = 1
      "0000001" when "00011010111101111", -- t[13807] = 1
      "0000001" when "00011010111110000", -- t[13808] = 1
      "0000001" when "00011010111110001", -- t[13809] = 1
      "0000001" when "00011010111110010", -- t[13810] = 1
      "0000001" when "00011010111110011", -- t[13811] = 1
      "0000001" when "00011010111110100", -- t[13812] = 1
      "0000001" when "00011010111110101", -- t[13813] = 1
      "0000001" when "00011010111110110", -- t[13814] = 1
      "0000001" when "00011010111110111", -- t[13815] = 1
      "0000001" when "00011010111111000", -- t[13816] = 1
      "0000001" when "00011010111111001", -- t[13817] = 1
      "0000001" when "00011010111111010", -- t[13818] = 1
      "0000001" when "00011010111111011", -- t[13819] = 1
      "0000001" when "00011010111111100", -- t[13820] = 1
      "0000001" when "00011010111111101", -- t[13821] = 1
      "0000001" when "00011010111111110", -- t[13822] = 1
      "0000001" when "00011010111111111", -- t[13823] = 1
      "0000001" when "00011011000000000", -- t[13824] = 1
      "0000001" when "00011011000000001", -- t[13825] = 1
      "0000001" when "00011011000000010", -- t[13826] = 1
      "0000001" when "00011011000000011", -- t[13827] = 1
      "0000001" when "00011011000000100", -- t[13828] = 1
      "0000001" when "00011011000000101", -- t[13829] = 1
      "0000001" when "00011011000000110", -- t[13830] = 1
      "0000001" when "00011011000000111", -- t[13831] = 1
      "0000001" when "00011011000001000", -- t[13832] = 1
      "0000001" when "00011011000001001", -- t[13833] = 1
      "0000001" when "00011011000001010", -- t[13834] = 1
      "0000001" when "00011011000001011", -- t[13835] = 1
      "0000001" when "00011011000001100", -- t[13836] = 1
      "0000001" when "00011011000001101", -- t[13837] = 1
      "0000001" when "00011011000001110", -- t[13838] = 1
      "0000001" when "00011011000001111", -- t[13839] = 1
      "0000001" when "00011011000010000", -- t[13840] = 1
      "0000001" when "00011011000010001", -- t[13841] = 1
      "0000001" when "00011011000010010", -- t[13842] = 1
      "0000001" when "00011011000010011", -- t[13843] = 1
      "0000001" when "00011011000010100", -- t[13844] = 1
      "0000001" when "00011011000010101", -- t[13845] = 1
      "0000001" when "00011011000010110", -- t[13846] = 1
      "0000001" when "00011011000010111", -- t[13847] = 1
      "0000001" when "00011011000011000", -- t[13848] = 1
      "0000001" when "00011011000011001", -- t[13849] = 1
      "0000001" when "00011011000011010", -- t[13850] = 1
      "0000001" when "00011011000011011", -- t[13851] = 1
      "0000001" when "00011011000011100", -- t[13852] = 1
      "0000001" when "00011011000011101", -- t[13853] = 1
      "0000001" when "00011011000011110", -- t[13854] = 1
      "0000001" when "00011011000011111", -- t[13855] = 1
      "0000001" when "00011011000100000", -- t[13856] = 1
      "0000001" when "00011011000100001", -- t[13857] = 1
      "0000001" when "00011011000100010", -- t[13858] = 1
      "0000001" when "00011011000100011", -- t[13859] = 1
      "0000001" when "00011011000100100", -- t[13860] = 1
      "0000001" when "00011011000100101", -- t[13861] = 1
      "0000001" when "00011011000100110", -- t[13862] = 1
      "0000001" when "00011011000100111", -- t[13863] = 1
      "0000001" when "00011011000101000", -- t[13864] = 1
      "0000001" when "00011011000101001", -- t[13865] = 1
      "0000001" when "00011011000101010", -- t[13866] = 1
      "0000001" when "00011011000101011", -- t[13867] = 1
      "0000001" when "00011011000101100", -- t[13868] = 1
      "0000001" when "00011011000101101", -- t[13869] = 1
      "0000001" when "00011011000101110", -- t[13870] = 1
      "0000001" when "00011011000101111", -- t[13871] = 1
      "0000001" when "00011011000110000", -- t[13872] = 1
      "0000001" when "00011011000110001", -- t[13873] = 1
      "0000001" when "00011011000110010", -- t[13874] = 1
      "0000001" when "00011011000110011", -- t[13875] = 1
      "0000001" when "00011011000110100", -- t[13876] = 1
      "0000001" when "00011011000110101", -- t[13877] = 1
      "0000001" when "00011011000110110", -- t[13878] = 1
      "0000001" when "00011011000110111", -- t[13879] = 1
      "0000001" when "00011011000111000", -- t[13880] = 1
      "0000001" when "00011011000111001", -- t[13881] = 1
      "0000001" when "00011011000111010", -- t[13882] = 1
      "0000001" when "00011011000111011", -- t[13883] = 1
      "0000001" when "00011011000111100", -- t[13884] = 1
      "0000001" when "00011011000111101", -- t[13885] = 1
      "0000001" when "00011011000111110", -- t[13886] = 1
      "0000001" when "00011011000111111", -- t[13887] = 1
      "0000001" when "00011011001000000", -- t[13888] = 1
      "0000001" when "00011011001000001", -- t[13889] = 1
      "0000001" when "00011011001000010", -- t[13890] = 1
      "0000001" when "00011011001000011", -- t[13891] = 1
      "0000001" when "00011011001000100", -- t[13892] = 1
      "0000001" when "00011011001000101", -- t[13893] = 1
      "0000001" when "00011011001000110", -- t[13894] = 1
      "0000001" when "00011011001000111", -- t[13895] = 1
      "0000001" when "00011011001001000", -- t[13896] = 1
      "0000001" when "00011011001001001", -- t[13897] = 1
      "0000001" when "00011011001001010", -- t[13898] = 1
      "0000001" when "00011011001001011", -- t[13899] = 1
      "0000001" when "00011011001001100", -- t[13900] = 1
      "0000001" when "00011011001001101", -- t[13901] = 1
      "0000001" when "00011011001001110", -- t[13902] = 1
      "0000001" when "00011011001001111", -- t[13903] = 1
      "0000001" when "00011011001010000", -- t[13904] = 1
      "0000001" when "00011011001010001", -- t[13905] = 1
      "0000001" when "00011011001010010", -- t[13906] = 1
      "0000001" when "00011011001010011", -- t[13907] = 1
      "0000001" when "00011011001010100", -- t[13908] = 1
      "0000001" when "00011011001010101", -- t[13909] = 1
      "0000001" when "00011011001010110", -- t[13910] = 1
      "0000001" when "00011011001010111", -- t[13911] = 1
      "0000001" when "00011011001011000", -- t[13912] = 1
      "0000001" when "00011011001011001", -- t[13913] = 1
      "0000001" when "00011011001011010", -- t[13914] = 1
      "0000001" when "00011011001011011", -- t[13915] = 1
      "0000001" when "00011011001011100", -- t[13916] = 1
      "0000001" when "00011011001011101", -- t[13917] = 1
      "0000001" when "00011011001011110", -- t[13918] = 1
      "0000001" when "00011011001011111", -- t[13919] = 1
      "0000001" when "00011011001100000", -- t[13920] = 1
      "0000001" when "00011011001100001", -- t[13921] = 1
      "0000001" when "00011011001100010", -- t[13922] = 1
      "0000001" when "00011011001100011", -- t[13923] = 1
      "0000001" when "00011011001100100", -- t[13924] = 1
      "0000001" when "00011011001100101", -- t[13925] = 1
      "0000001" when "00011011001100110", -- t[13926] = 1
      "0000001" when "00011011001100111", -- t[13927] = 1
      "0000001" when "00011011001101000", -- t[13928] = 1
      "0000001" when "00011011001101001", -- t[13929] = 1
      "0000001" when "00011011001101010", -- t[13930] = 1
      "0000001" when "00011011001101011", -- t[13931] = 1
      "0000001" when "00011011001101100", -- t[13932] = 1
      "0000001" when "00011011001101101", -- t[13933] = 1
      "0000001" when "00011011001101110", -- t[13934] = 1
      "0000001" when "00011011001101111", -- t[13935] = 1
      "0000001" when "00011011001110000", -- t[13936] = 1
      "0000001" when "00011011001110001", -- t[13937] = 1
      "0000001" when "00011011001110010", -- t[13938] = 1
      "0000001" when "00011011001110011", -- t[13939] = 1
      "0000001" when "00011011001110100", -- t[13940] = 1
      "0000001" when "00011011001110101", -- t[13941] = 1
      "0000001" when "00011011001110110", -- t[13942] = 1
      "0000001" when "00011011001110111", -- t[13943] = 1
      "0000001" when "00011011001111000", -- t[13944] = 1
      "0000001" when "00011011001111001", -- t[13945] = 1
      "0000001" when "00011011001111010", -- t[13946] = 1
      "0000001" when "00011011001111011", -- t[13947] = 1
      "0000001" when "00011011001111100", -- t[13948] = 1
      "0000001" when "00011011001111101", -- t[13949] = 1
      "0000001" when "00011011001111110", -- t[13950] = 1
      "0000001" when "00011011001111111", -- t[13951] = 1
      "0000001" when "00011011010000000", -- t[13952] = 1
      "0000001" when "00011011010000001", -- t[13953] = 1
      "0000001" when "00011011010000010", -- t[13954] = 1
      "0000001" when "00011011010000011", -- t[13955] = 1
      "0000001" when "00011011010000100", -- t[13956] = 1
      "0000001" when "00011011010000101", -- t[13957] = 1
      "0000001" when "00011011010000110", -- t[13958] = 1
      "0000001" when "00011011010000111", -- t[13959] = 1
      "0000001" when "00011011010001000", -- t[13960] = 1
      "0000001" when "00011011010001001", -- t[13961] = 1
      "0000001" when "00011011010001010", -- t[13962] = 1
      "0000001" when "00011011010001011", -- t[13963] = 1
      "0000001" when "00011011010001100", -- t[13964] = 1
      "0000001" when "00011011010001101", -- t[13965] = 1
      "0000001" when "00011011010001110", -- t[13966] = 1
      "0000001" when "00011011010001111", -- t[13967] = 1
      "0000001" when "00011011010010000", -- t[13968] = 1
      "0000001" when "00011011010010001", -- t[13969] = 1
      "0000001" when "00011011010010010", -- t[13970] = 1
      "0000001" when "00011011010010011", -- t[13971] = 1
      "0000001" when "00011011010010100", -- t[13972] = 1
      "0000001" when "00011011010010101", -- t[13973] = 1
      "0000001" when "00011011010010110", -- t[13974] = 1
      "0000001" when "00011011010010111", -- t[13975] = 1
      "0000001" when "00011011010011000", -- t[13976] = 1
      "0000001" when "00011011010011001", -- t[13977] = 1
      "0000001" when "00011011010011010", -- t[13978] = 1
      "0000001" when "00011011010011011", -- t[13979] = 1
      "0000001" when "00011011010011100", -- t[13980] = 1
      "0000001" when "00011011010011101", -- t[13981] = 1
      "0000001" when "00011011010011110", -- t[13982] = 1
      "0000001" when "00011011010011111", -- t[13983] = 1
      "0000001" when "00011011010100000", -- t[13984] = 1
      "0000001" when "00011011010100001", -- t[13985] = 1
      "0000001" when "00011011010100010", -- t[13986] = 1
      "0000001" when "00011011010100011", -- t[13987] = 1
      "0000001" when "00011011010100100", -- t[13988] = 1
      "0000001" when "00011011010100101", -- t[13989] = 1
      "0000001" when "00011011010100110", -- t[13990] = 1
      "0000001" when "00011011010100111", -- t[13991] = 1
      "0000001" when "00011011010101000", -- t[13992] = 1
      "0000001" when "00011011010101001", -- t[13993] = 1
      "0000001" when "00011011010101010", -- t[13994] = 1
      "0000001" when "00011011010101011", -- t[13995] = 1
      "0000001" when "00011011010101100", -- t[13996] = 1
      "0000001" when "00011011010101101", -- t[13997] = 1
      "0000001" when "00011011010101110", -- t[13998] = 1
      "0000001" when "00011011010101111", -- t[13999] = 1
      "0000001" when "00011011010110000", -- t[14000] = 1
      "0000001" when "00011011010110001", -- t[14001] = 1
      "0000001" when "00011011010110010", -- t[14002] = 1
      "0000001" when "00011011010110011", -- t[14003] = 1
      "0000001" when "00011011010110100", -- t[14004] = 1
      "0000001" when "00011011010110101", -- t[14005] = 1
      "0000001" when "00011011010110110", -- t[14006] = 1
      "0000001" when "00011011010110111", -- t[14007] = 1
      "0000001" when "00011011010111000", -- t[14008] = 1
      "0000001" when "00011011010111001", -- t[14009] = 1
      "0000001" when "00011011010111010", -- t[14010] = 1
      "0000001" when "00011011010111011", -- t[14011] = 1
      "0000001" when "00011011010111100", -- t[14012] = 1
      "0000001" when "00011011010111101", -- t[14013] = 1
      "0000001" when "00011011010111110", -- t[14014] = 1
      "0000001" when "00011011010111111", -- t[14015] = 1
      "0000001" when "00011011011000000", -- t[14016] = 1
      "0000001" when "00011011011000001", -- t[14017] = 1
      "0000001" when "00011011011000010", -- t[14018] = 1
      "0000001" when "00011011011000011", -- t[14019] = 1
      "0000001" when "00011011011000100", -- t[14020] = 1
      "0000001" when "00011011011000101", -- t[14021] = 1
      "0000001" when "00011011011000110", -- t[14022] = 1
      "0000001" when "00011011011000111", -- t[14023] = 1
      "0000001" when "00011011011001000", -- t[14024] = 1
      "0000001" when "00011011011001001", -- t[14025] = 1
      "0000001" when "00011011011001010", -- t[14026] = 1
      "0000001" when "00011011011001011", -- t[14027] = 1
      "0000001" when "00011011011001100", -- t[14028] = 1
      "0000001" when "00011011011001101", -- t[14029] = 1
      "0000001" when "00011011011001110", -- t[14030] = 1
      "0000001" when "00011011011001111", -- t[14031] = 1
      "0000001" when "00011011011010000", -- t[14032] = 1
      "0000001" when "00011011011010001", -- t[14033] = 1
      "0000001" when "00011011011010010", -- t[14034] = 1
      "0000001" when "00011011011010011", -- t[14035] = 1
      "0000001" when "00011011011010100", -- t[14036] = 1
      "0000001" when "00011011011010101", -- t[14037] = 1
      "0000001" when "00011011011010110", -- t[14038] = 1
      "0000001" when "00011011011010111", -- t[14039] = 1
      "0000001" when "00011011011011000", -- t[14040] = 1
      "0000001" when "00011011011011001", -- t[14041] = 1
      "0000001" when "00011011011011010", -- t[14042] = 1
      "0000001" when "00011011011011011", -- t[14043] = 1
      "0000001" when "00011011011011100", -- t[14044] = 1
      "0000001" when "00011011011011101", -- t[14045] = 1
      "0000001" when "00011011011011110", -- t[14046] = 1
      "0000001" when "00011011011011111", -- t[14047] = 1
      "0000001" when "00011011011100000", -- t[14048] = 1
      "0000001" when "00011011011100001", -- t[14049] = 1
      "0000001" when "00011011011100010", -- t[14050] = 1
      "0000001" when "00011011011100011", -- t[14051] = 1
      "0000001" when "00011011011100100", -- t[14052] = 1
      "0000001" when "00011011011100101", -- t[14053] = 1
      "0000001" when "00011011011100110", -- t[14054] = 1
      "0000001" when "00011011011100111", -- t[14055] = 1
      "0000001" when "00011011011101000", -- t[14056] = 1
      "0000001" when "00011011011101001", -- t[14057] = 1
      "0000001" when "00011011011101010", -- t[14058] = 1
      "0000001" when "00011011011101011", -- t[14059] = 1
      "0000001" when "00011011011101100", -- t[14060] = 1
      "0000001" when "00011011011101101", -- t[14061] = 1
      "0000001" when "00011011011101110", -- t[14062] = 1
      "0000001" when "00011011011101111", -- t[14063] = 1
      "0000001" when "00011011011110000", -- t[14064] = 1
      "0000001" when "00011011011110001", -- t[14065] = 1
      "0000001" when "00011011011110010", -- t[14066] = 1
      "0000001" when "00011011011110011", -- t[14067] = 1
      "0000001" when "00011011011110100", -- t[14068] = 1
      "0000001" when "00011011011110101", -- t[14069] = 1
      "0000001" when "00011011011110110", -- t[14070] = 1
      "0000001" when "00011011011110111", -- t[14071] = 1
      "0000001" when "00011011011111000", -- t[14072] = 1
      "0000001" when "00011011011111001", -- t[14073] = 1
      "0000001" when "00011011011111010", -- t[14074] = 1
      "0000001" when "00011011011111011", -- t[14075] = 1
      "0000001" when "00011011011111100", -- t[14076] = 1
      "0000001" when "00011011011111101", -- t[14077] = 1
      "0000001" when "00011011011111110", -- t[14078] = 1
      "0000001" when "00011011011111111", -- t[14079] = 1
      "0000001" when "00011011100000000", -- t[14080] = 1
      "0000001" when "00011011100000001", -- t[14081] = 1
      "0000001" when "00011011100000010", -- t[14082] = 1
      "0000001" when "00011011100000011", -- t[14083] = 1
      "0000001" when "00011011100000100", -- t[14084] = 1
      "0000001" when "00011011100000101", -- t[14085] = 1
      "0000001" when "00011011100000110", -- t[14086] = 1
      "0000001" when "00011011100000111", -- t[14087] = 1
      "0000001" when "00011011100001000", -- t[14088] = 1
      "0000001" when "00011011100001001", -- t[14089] = 1
      "0000001" when "00011011100001010", -- t[14090] = 1
      "0000001" when "00011011100001011", -- t[14091] = 1
      "0000001" when "00011011100001100", -- t[14092] = 1
      "0000001" when "00011011100001101", -- t[14093] = 1
      "0000001" when "00011011100001110", -- t[14094] = 1
      "0000001" when "00011011100001111", -- t[14095] = 1
      "0000001" when "00011011100010000", -- t[14096] = 1
      "0000001" when "00011011100010001", -- t[14097] = 1
      "0000001" when "00011011100010010", -- t[14098] = 1
      "0000001" when "00011011100010011", -- t[14099] = 1
      "0000001" when "00011011100010100", -- t[14100] = 1
      "0000001" when "00011011100010101", -- t[14101] = 1
      "0000001" when "00011011100010110", -- t[14102] = 1
      "0000001" when "00011011100010111", -- t[14103] = 1
      "0000001" when "00011011100011000", -- t[14104] = 1
      "0000001" when "00011011100011001", -- t[14105] = 1
      "0000001" when "00011011100011010", -- t[14106] = 1
      "0000001" when "00011011100011011", -- t[14107] = 1
      "0000001" when "00011011100011100", -- t[14108] = 1
      "0000001" when "00011011100011101", -- t[14109] = 1
      "0000001" when "00011011100011110", -- t[14110] = 1
      "0000001" when "00011011100011111", -- t[14111] = 1
      "0000001" when "00011011100100000", -- t[14112] = 1
      "0000001" when "00011011100100001", -- t[14113] = 1
      "0000001" when "00011011100100010", -- t[14114] = 1
      "0000001" when "00011011100100011", -- t[14115] = 1
      "0000001" when "00011011100100100", -- t[14116] = 1
      "0000001" when "00011011100100101", -- t[14117] = 1
      "0000001" when "00011011100100110", -- t[14118] = 1
      "0000001" when "00011011100100111", -- t[14119] = 1
      "0000001" when "00011011100101000", -- t[14120] = 1
      "0000001" when "00011011100101001", -- t[14121] = 1
      "0000001" when "00011011100101010", -- t[14122] = 1
      "0000001" when "00011011100101011", -- t[14123] = 1
      "0000001" when "00011011100101100", -- t[14124] = 1
      "0000001" when "00011011100101101", -- t[14125] = 1
      "0000001" when "00011011100101110", -- t[14126] = 1
      "0000001" when "00011011100101111", -- t[14127] = 1
      "0000001" when "00011011100110000", -- t[14128] = 1
      "0000001" when "00011011100110001", -- t[14129] = 1
      "0000001" when "00011011100110010", -- t[14130] = 1
      "0000001" when "00011011100110011", -- t[14131] = 1
      "0000001" when "00011011100110100", -- t[14132] = 1
      "0000001" when "00011011100110101", -- t[14133] = 1
      "0000001" when "00011011100110110", -- t[14134] = 1
      "0000001" when "00011011100110111", -- t[14135] = 1
      "0000001" when "00011011100111000", -- t[14136] = 1
      "0000001" when "00011011100111001", -- t[14137] = 1
      "0000001" when "00011011100111010", -- t[14138] = 1
      "0000001" when "00011011100111011", -- t[14139] = 1
      "0000001" when "00011011100111100", -- t[14140] = 1
      "0000001" when "00011011100111101", -- t[14141] = 1
      "0000001" when "00011011100111110", -- t[14142] = 1
      "0000001" when "00011011100111111", -- t[14143] = 1
      "0000001" when "00011011101000000", -- t[14144] = 1
      "0000001" when "00011011101000001", -- t[14145] = 1
      "0000001" when "00011011101000010", -- t[14146] = 1
      "0000001" when "00011011101000011", -- t[14147] = 1
      "0000001" when "00011011101000100", -- t[14148] = 1
      "0000001" when "00011011101000101", -- t[14149] = 1
      "0000001" when "00011011101000110", -- t[14150] = 1
      "0000001" when "00011011101000111", -- t[14151] = 1
      "0000001" when "00011011101001000", -- t[14152] = 1
      "0000001" when "00011011101001001", -- t[14153] = 1
      "0000001" when "00011011101001010", -- t[14154] = 1
      "0000001" when "00011011101001011", -- t[14155] = 1
      "0000001" when "00011011101001100", -- t[14156] = 1
      "0000001" when "00011011101001101", -- t[14157] = 1
      "0000001" when "00011011101001110", -- t[14158] = 1
      "0000001" when "00011011101001111", -- t[14159] = 1
      "0000001" when "00011011101010000", -- t[14160] = 1
      "0000001" when "00011011101010001", -- t[14161] = 1
      "0000001" when "00011011101010010", -- t[14162] = 1
      "0000001" when "00011011101010011", -- t[14163] = 1
      "0000001" when "00011011101010100", -- t[14164] = 1
      "0000001" when "00011011101010101", -- t[14165] = 1
      "0000001" when "00011011101010110", -- t[14166] = 1
      "0000001" when "00011011101010111", -- t[14167] = 1
      "0000001" when "00011011101011000", -- t[14168] = 1
      "0000001" when "00011011101011001", -- t[14169] = 1
      "0000001" when "00011011101011010", -- t[14170] = 1
      "0000001" when "00011011101011011", -- t[14171] = 1
      "0000001" when "00011011101011100", -- t[14172] = 1
      "0000001" when "00011011101011101", -- t[14173] = 1
      "0000001" when "00011011101011110", -- t[14174] = 1
      "0000001" when "00011011101011111", -- t[14175] = 1
      "0000001" when "00011011101100000", -- t[14176] = 1
      "0000001" when "00011011101100001", -- t[14177] = 1
      "0000001" when "00011011101100010", -- t[14178] = 1
      "0000001" when "00011011101100011", -- t[14179] = 1
      "0000001" when "00011011101100100", -- t[14180] = 1
      "0000001" when "00011011101100101", -- t[14181] = 1
      "0000001" when "00011011101100110", -- t[14182] = 1
      "0000001" when "00011011101100111", -- t[14183] = 1
      "0000001" when "00011011101101000", -- t[14184] = 1
      "0000001" when "00011011101101001", -- t[14185] = 1
      "0000001" when "00011011101101010", -- t[14186] = 1
      "0000001" when "00011011101101011", -- t[14187] = 1
      "0000001" when "00011011101101100", -- t[14188] = 1
      "0000001" when "00011011101101101", -- t[14189] = 1
      "0000001" when "00011011101101110", -- t[14190] = 1
      "0000001" when "00011011101101111", -- t[14191] = 1
      "0000001" when "00011011101110000", -- t[14192] = 1
      "0000001" when "00011011101110001", -- t[14193] = 1
      "0000001" when "00011011101110010", -- t[14194] = 1
      "0000001" when "00011011101110011", -- t[14195] = 1
      "0000001" when "00011011101110100", -- t[14196] = 1
      "0000001" when "00011011101110101", -- t[14197] = 1
      "0000001" when "00011011101110110", -- t[14198] = 1
      "0000001" when "00011011101110111", -- t[14199] = 1
      "0000001" when "00011011101111000", -- t[14200] = 1
      "0000001" when "00011011101111001", -- t[14201] = 1
      "0000001" when "00011011101111010", -- t[14202] = 1
      "0000001" when "00011011101111011", -- t[14203] = 1
      "0000001" when "00011011101111100", -- t[14204] = 1
      "0000001" when "00011011101111101", -- t[14205] = 1
      "0000001" when "00011011101111110", -- t[14206] = 1
      "0000001" when "00011011101111111", -- t[14207] = 1
      "0000001" when "00011011110000000", -- t[14208] = 1
      "0000001" when "00011011110000001", -- t[14209] = 1
      "0000001" when "00011011110000010", -- t[14210] = 1
      "0000001" when "00011011110000011", -- t[14211] = 1
      "0000001" when "00011011110000100", -- t[14212] = 1
      "0000001" when "00011011110000101", -- t[14213] = 1
      "0000001" when "00011011110000110", -- t[14214] = 1
      "0000001" when "00011011110000111", -- t[14215] = 1
      "0000001" when "00011011110001000", -- t[14216] = 1
      "0000001" when "00011011110001001", -- t[14217] = 1
      "0000001" when "00011011110001010", -- t[14218] = 1
      "0000001" when "00011011110001011", -- t[14219] = 1
      "0000001" when "00011011110001100", -- t[14220] = 1
      "0000001" when "00011011110001101", -- t[14221] = 1
      "0000001" when "00011011110001110", -- t[14222] = 1
      "0000001" when "00011011110001111", -- t[14223] = 1
      "0000001" when "00011011110010000", -- t[14224] = 1
      "0000001" when "00011011110010001", -- t[14225] = 1
      "0000001" when "00011011110010010", -- t[14226] = 1
      "0000001" when "00011011110010011", -- t[14227] = 1
      "0000001" when "00011011110010100", -- t[14228] = 1
      "0000001" when "00011011110010101", -- t[14229] = 1
      "0000001" when "00011011110010110", -- t[14230] = 1
      "0000001" when "00011011110010111", -- t[14231] = 1
      "0000001" when "00011011110011000", -- t[14232] = 1
      "0000001" when "00011011110011001", -- t[14233] = 1
      "0000001" when "00011011110011010", -- t[14234] = 1
      "0000001" when "00011011110011011", -- t[14235] = 1
      "0000001" when "00011011110011100", -- t[14236] = 1
      "0000001" when "00011011110011101", -- t[14237] = 1
      "0000001" when "00011011110011110", -- t[14238] = 1
      "0000001" when "00011011110011111", -- t[14239] = 1
      "0000001" when "00011011110100000", -- t[14240] = 1
      "0000001" when "00011011110100001", -- t[14241] = 1
      "0000001" when "00011011110100010", -- t[14242] = 1
      "0000001" when "00011011110100011", -- t[14243] = 1
      "0000001" when "00011011110100100", -- t[14244] = 1
      "0000001" when "00011011110100101", -- t[14245] = 1
      "0000001" when "00011011110100110", -- t[14246] = 1
      "0000001" when "00011011110100111", -- t[14247] = 1
      "0000001" when "00011011110101000", -- t[14248] = 1
      "0000001" when "00011011110101001", -- t[14249] = 1
      "0000001" when "00011011110101010", -- t[14250] = 1
      "0000001" when "00011011110101011", -- t[14251] = 1
      "0000001" when "00011011110101100", -- t[14252] = 1
      "0000001" when "00011011110101101", -- t[14253] = 1
      "0000001" when "00011011110101110", -- t[14254] = 1
      "0000001" when "00011011110101111", -- t[14255] = 1
      "0000001" when "00011011110110000", -- t[14256] = 1
      "0000001" when "00011011110110001", -- t[14257] = 1
      "0000001" when "00011011110110010", -- t[14258] = 1
      "0000001" when "00011011110110011", -- t[14259] = 1
      "0000001" when "00011011110110100", -- t[14260] = 1
      "0000001" when "00011011110110101", -- t[14261] = 1
      "0000001" when "00011011110110110", -- t[14262] = 1
      "0000001" when "00011011110110111", -- t[14263] = 1
      "0000001" when "00011011110111000", -- t[14264] = 1
      "0000001" when "00011011110111001", -- t[14265] = 1
      "0000001" when "00011011110111010", -- t[14266] = 1
      "0000001" when "00011011110111011", -- t[14267] = 1
      "0000001" when "00011011110111100", -- t[14268] = 1
      "0000001" when "00011011110111101", -- t[14269] = 1
      "0000001" when "00011011110111110", -- t[14270] = 1
      "0000001" when "00011011110111111", -- t[14271] = 1
      "0000001" when "00011011111000000", -- t[14272] = 1
      "0000001" when "00011011111000001", -- t[14273] = 1
      "0000001" when "00011011111000010", -- t[14274] = 1
      "0000001" when "00011011111000011", -- t[14275] = 1
      "0000001" when "00011011111000100", -- t[14276] = 1
      "0000001" when "00011011111000101", -- t[14277] = 1
      "0000001" when "00011011111000110", -- t[14278] = 1
      "0000001" when "00011011111000111", -- t[14279] = 1
      "0000001" when "00011011111001000", -- t[14280] = 1
      "0000001" when "00011011111001001", -- t[14281] = 1
      "0000001" when "00011011111001010", -- t[14282] = 1
      "0000001" when "00011011111001011", -- t[14283] = 1
      "0000001" when "00011011111001100", -- t[14284] = 1
      "0000001" when "00011011111001101", -- t[14285] = 1
      "0000001" when "00011011111001110", -- t[14286] = 1
      "0000001" when "00011011111001111", -- t[14287] = 1
      "0000001" when "00011011111010000", -- t[14288] = 1
      "0000001" when "00011011111010001", -- t[14289] = 1
      "0000001" when "00011011111010010", -- t[14290] = 1
      "0000001" when "00011011111010011", -- t[14291] = 1
      "0000001" when "00011011111010100", -- t[14292] = 1
      "0000001" when "00011011111010101", -- t[14293] = 1
      "0000001" when "00011011111010110", -- t[14294] = 1
      "0000001" when "00011011111010111", -- t[14295] = 1
      "0000001" when "00011011111011000", -- t[14296] = 1
      "0000001" when "00011011111011001", -- t[14297] = 1
      "0000001" when "00011011111011010", -- t[14298] = 1
      "0000001" when "00011011111011011", -- t[14299] = 1
      "0000001" when "00011011111011100", -- t[14300] = 1
      "0000001" when "00011011111011101", -- t[14301] = 1
      "0000001" when "00011011111011110", -- t[14302] = 1
      "0000001" when "00011011111011111", -- t[14303] = 1
      "0000001" when "00011011111100000", -- t[14304] = 1
      "0000001" when "00011011111100001", -- t[14305] = 1
      "0000001" when "00011011111100010", -- t[14306] = 1
      "0000001" when "00011011111100011", -- t[14307] = 1
      "0000001" when "00011011111100100", -- t[14308] = 1
      "0000001" when "00011011111100101", -- t[14309] = 1
      "0000001" when "00011011111100110", -- t[14310] = 1
      "0000001" when "00011011111100111", -- t[14311] = 1
      "0000001" when "00011011111101000", -- t[14312] = 1
      "0000001" when "00011011111101001", -- t[14313] = 1
      "0000001" when "00011011111101010", -- t[14314] = 1
      "0000001" when "00011011111101011", -- t[14315] = 1
      "0000001" when "00011011111101100", -- t[14316] = 1
      "0000001" when "00011011111101101", -- t[14317] = 1
      "0000001" when "00011011111101110", -- t[14318] = 1
      "0000001" when "00011011111101111", -- t[14319] = 1
      "0000001" when "00011011111110000", -- t[14320] = 1
      "0000001" when "00011011111110001", -- t[14321] = 1
      "0000001" when "00011011111110010", -- t[14322] = 1
      "0000001" when "00011011111110011", -- t[14323] = 1
      "0000001" when "00011011111110100", -- t[14324] = 1
      "0000001" when "00011011111110101", -- t[14325] = 1
      "0000001" when "00011011111110110", -- t[14326] = 1
      "0000001" when "00011011111110111", -- t[14327] = 1
      "0000001" when "00011011111111000", -- t[14328] = 1
      "0000001" when "00011011111111001", -- t[14329] = 1
      "0000001" when "00011011111111010", -- t[14330] = 1
      "0000001" when "00011011111111011", -- t[14331] = 1
      "0000001" when "00011011111111100", -- t[14332] = 1
      "0000001" when "00011011111111101", -- t[14333] = 1
      "0000001" when "00011011111111110", -- t[14334] = 1
      "0000001" when "00011011111111111", -- t[14335] = 1
      "0000001" when "00011100000000000", -- t[14336] = 1
      "0000001" when "00011100000000001", -- t[14337] = 1
      "0000001" when "00011100000000010", -- t[14338] = 1
      "0000001" when "00011100000000011", -- t[14339] = 1
      "0000001" when "00011100000000100", -- t[14340] = 1
      "0000001" when "00011100000000101", -- t[14341] = 1
      "0000001" when "00011100000000110", -- t[14342] = 1
      "0000001" when "00011100000000111", -- t[14343] = 1
      "0000001" when "00011100000001000", -- t[14344] = 1
      "0000001" when "00011100000001001", -- t[14345] = 1
      "0000001" when "00011100000001010", -- t[14346] = 1
      "0000001" when "00011100000001011", -- t[14347] = 1
      "0000001" when "00011100000001100", -- t[14348] = 1
      "0000001" when "00011100000001101", -- t[14349] = 1
      "0000001" when "00011100000001110", -- t[14350] = 1
      "0000001" when "00011100000001111", -- t[14351] = 1
      "0000001" when "00011100000010000", -- t[14352] = 1
      "0000001" when "00011100000010001", -- t[14353] = 1
      "0000001" when "00011100000010010", -- t[14354] = 1
      "0000001" when "00011100000010011", -- t[14355] = 1
      "0000001" when "00011100000010100", -- t[14356] = 1
      "0000001" when "00011100000010101", -- t[14357] = 1
      "0000001" when "00011100000010110", -- t[14358] = 1
      "0000001" when "00011100000010111", -- t[14359] = 1
      "0000001" when "00011100000011000", -- t[14360] = 1
      "0000001" when "00011100000011001", -- t[14361] = 1
      "0000001" when "00011100000011010", -- t[14362] = 1
      "0000001" when "00011100000011011", -- t[14363] = 1
      "0000001" when "00011100000011100", -- t[14364] = 1
      "0000001" when "00011100000011101", -- t[14365] = 1
      "0000001" when "00011100000011110", -- t[14366] = 1
      "0000001" when "00011100000011111", -- t[14367] = 1
      "0000001" when "00011100000100000", -- t[14368] = 1
      "0000001" when "00011100000100001", -- t[14369] = 1
      "0000001" when "00011100000100010", -- t[14370] = 1
      "0000001" when "00011100000100011", -- t[14371] = 1
      "0000001" when "00011100000100100", -- t[14372] = 1
      "0000001" when "00011100000100101", -- t[14373] = 1
      "0000001" when "00011100000100110", -- t[14374] = 1
      "0000001" when "00011100000100111", -- t[14375] = 1
      "0000001" when "00011100000101000", -- t[14376] = 1
      "0000001" when "00011100000101001", -- t[14377] = 1
      "0000001" when "00011100000101010", -- t[14378] = 1
      "0000001" when "00011100000101011", -- t[14379] = 1
      "0000001" when "00011100000101100", -- t[14380] = 1
      "0000001" when "00011100000101101", -- t[14381] = 1
      "0000001" when "00011100000101110", -- t[14382] = 1
      "0000001" when "00011100000101111", -- t[14383] = 1
      "0000001" when "00011100000110000", -- t[14384] = 1
      "0000001" when "00011100000110001", -- t[14385] = 1
      "0000001" when "00011100000110010", -- t[14386] = 1
      "0000001" when "00011100000110011", -- t[14387] = 1
      "0000001" when "00011100000110100", -- t[14388] = 1
      "0000001" when "00011100000110101", -- t[14389] = 1
      "0000001" when "00011100000110110", -- t[14390] = 1
      "0000001" when "00011100000110111", -- t[14391] = 1
      "0000001" when "00011100000111000", -- t[14392] = 1
      "0000001" when "00011100000111001", -- t[14393] = 1
      "0000001" when "00011100000111010", -- t[14394] = 1
      "0000001" when "00011100000111011", -- t[14395] = 1
      "0000001" when "00011100000111100", -- t[14396] = 1
      "0000001" when "00011100000111101", -- t[14397] = 1
      "0000001" when "00011100000111110", -- t[14398] = 1
      "0000001" when "00011100000111111", -- t[14399] = 1
      "0000001" when "00011100001000000", -- t[14400] = 1
      "0000001" when "00011100001000001", -- t[14401] = 1
      "0000001" when "00011100001000010", -- t[14402] = 1
      "0000001" when "00011100001000011", -- t[14403] = 1
      "0000001" when "00011100001000100", -- t[14404] = 1
      "0000001" when "00011100001000101", -- t[14405] = 1
      "0000001" when "00011100001000110", -- t[14406] = 1
      "0000001" when "00011100001000111", -- t[14407] = 1
      "0000001" when "00011100001001000", -- t[14408] = 1
      "0000001" when "00011100001001001", -- t[14409] = 1
      "0000001" when "00011100001001010", -- t[14410] = 1
      "0000001" when "00011100001001011", -- t[14411] = 1
      "0000001" when "00011100001001100", -- t[14412] = 1
      "0000001" when "00011100001001101", -- t[14413] = 1
      "0000001" when "00011100001001110", -- t[14414] = 1
      "0000001" when "00011100001001111", -- t[14415] = 1
      "0000001" when "00011100001010000", -- t[14416] = 1
      "0000001" when "00011100001010001", -- t[14417] = 1
      "0000001" when "00011100001010010", -- t[14418] = 1
      "0000001" when "00011100001010011", -- t[14419] = 1
      "0000001" when "00011100001010100", -- t[14420] = 1
      "0000001" when "00011100001010101", -- t[14421] = 1
      "0000001" when "00011100001010110", -- t[14422] = 1
      "0000001" when "00011100001010111", -- t[14423] = 1
      "0000001" when "00011100001011000", -- t[14424] = 1
      "0000001" when "00011100001011001", -- t[14425] = 1
      "0000001" when "00011100001011010", -- t[14426] = 1
      "0000001" when "00011100001011011", -- t[14427] = 1
      "0000001" when "00011100001011100", -- t[14428] = 1
      "0000001" when "00011100001011101", -- t[14429] = 1
      "0000001" when "00011100001011110", -- t[14430] = 1
      "0000001" when "00011100001011111", -- t[14431] = 1
      "0000001" when "00011100001100000", -- t[14432] = 1
      "0000001" when "00011100001100001", -- t[14433] = 1
      "0000001" when "00011100001100010", -- t[14434] = 1
      "0000001" when "00011100001100011", -- t[14435] = 1
      "0000001" when "00011100001100100", -- t[14436] = 1
      "0000001" when "00011100001100101", -- t[14437] = 1
      "0000001" when "00011100001100110", -- t[14438] = 1
      "0000001" when "00011100001100111", -- t[14439] = 1
      "0000001" when "00011100001101000", -- t[14440] = 1
      "0000001" when "00011100001101001", -- t[14441] = 1
      "0000001" when "00011100001101010", -- t[14442] = 1
      "0000001" when "00011100001101011", -- t[14443] = 1
      "0000001" when "00011100001101100", -- t[14444] = 1
      "0000001" when "00011100001101101", -- t[14445] = 1
      "0000001" when "00011100001101110", -- t[14446] = 1
      "0000001" when "00011100001101111", -- t[14447] = 1
      "0000001" when "00011100001110000", -- t[14448] = 1
      "0000001" when "00011100001110001", -- t[14449] = 1
      "0000001" when "00011100001110010", -- t[14450] = 1
      "0000001" when "00011100001110011", -- t[14451] = 1
      "0000001" when "00011100001110100", -- t[14452] = 1
      "0000001" when "00011100001110101", -- t[14453] = 1
      "0000001" when "00011100001110110", -- t[14454] = 1
      "0000001" when "00011100001110111", -- t[14455] = 1
      "0000001" when "00011100001111000", -- t[14456] = 1
      "0000001" when "00011100001111001", -- t[14457] = 1
      "0000001" when "00011100001111010", -- t[14458] = 1
      "0000001" when "00011100001111011", -- t[14459] = 1
      "0000001" when "00011100001111100", -- t[14460] = 1
      "0000001" when "00011100001111101", -- t[14461] = 1
      "0000001" when "00011100001111110", -- t[14462] = 1
      "0000001" when "00011100001111111", -- t[14463] = 1
      "0000001" when "00011100010000000", -- t[14464] = 1
      "0000001" when "00011100010000001", -- t[14465] = 1
      "0000001" when "00011100010000010", -- t[14466] = 1
      "0000001" when "00011100010000011", -- t[14467] = 1
      "0000001" when "00011100010000100", -- t[14468] = 1
      "0000001" when "00011100010000101", -- t[14469] = 1
      "0000001" when "00011100010000110", -- t[14470] = 1
      "0000001" when "00011100010000111", -- t[14471] = 1
      "0000001" when "00011100010001000", -- t[14472] = 1
      "0000001" when "00011100010001001", -- t[14473] = 1
      "0000001" when "00011100010001010", -- t[14474] = 1
      "0000001" when "00011100010001011", -- t[14475] = 1
      "0000001" when "00011100010001100", -- t[14476] = 1
      "0000001" when "00011100010001101", -- t[14477] = 1
      "0000001" when "00011100010001110", -- t[14478] = 1
      "0000001" when "00011100010001111", -- t[14479] = 1
      "0000001" when "00011100010010000", -- t[14480] = 1
      "0000001" when "00011100010010001", -- t[14481] = 1
      "0000001" when "00011100010010010", -- t[14482] = 1
      "0000001" when "00011100010010011", -- t[14483] = 1
      "0000001" when "00011100010010100", -- t[14484] = 1
      "0000001" when "00011100010010101", -- t[14485] = 1
      "0000001" when "00011100010010110", -- t[14486] = 1
      "0000001" when "00011100010010111", -- t[14487] = 1
      "0000001" when "00011100010011000", -- t[14488] = 1
      "0000001" when "00011100010011001", -- t[14489] = 1
      "0000001" when "00011100010011010", -- t[14490] = 1
      "0000001" when "00011100010011011", -- t[14491] = 1
      "0000001" when "00011100010011100", -- t[14492] = 1
      "0000001" when "00011100010011101", -- t[14493] = 1
      "0000001" when "00011100010011110", -- t[14494] = 1
      "0000001" when "00011100010011111", -- t[14495] = 1
      "0000001" when "00011100010100000", -- t[14496] = 1
      "0000001" when "00011100010100001", -- t[14497] = 1
      "0000001" when "00011100010100010", -- t[14498] = 1
      "0000001" when "00011100010100011", -- t[14499] = 1
      "0000001" when "00011100010100100", -- t[14500] = 1
      "0000001" when "00011100010100101", -- t[14501] = 1
      "0000001" when "00011100010100110", -- t[14502] = 1
      "0000001" when "00011100010100111", -- t[14503] = 1
      "0000001" when "00011100010101000", -- t[14504] = 1
      "0000001" when "00011100010101001", -- t[14505] = 1
      "0000001" when "00011100010101010", -- t[14506] = 1
      "0000001" when "00011100010101011", -- t[14507] = 1
      "0000001" when "00011100010101100", -- t[14508] = 1
      "0000001" when "00011100010101101", -- t[14509] = 1
      "0000001" when "00011100010101110", -- t[14510] = 1
      "0000001" when "00011100010101111", -- t[14511] = 1
      "0000001" when "00011100010110000", -- t[14512] = 1
      "0000001" when "00011100010110001", -- t[14513] = 1
      "0000001" when "00011100010110010", -- t[14514] = 1
      "0000001" when "00011100010110011", -- t[14515] = 1
      "0000001" when "00011100010110100", -- t[14516] = 1
      "0000001" when "00011100010110101", -- t[14517] = 1
      "0000001" when "00011100010110110", -- t[14518] = 1
      "0000001" when "00011100010110111", -- t[14519] = 1
      "0000001" when "00011100010111000", -- t[14520] = 1
      "0000001" when "00011100010111001", -- t[14521] = 1
      "0000001" when "00011100010111010", -- t[14522] = 1
      "0000001" when "00011100010111011", -- t[14523] = 1
      "0000001" when "00011100010111100", -- t[14524] = 1
      "0000001" when "00011100010111101", -- t[14525] = 1
      "0000001" when "00011100010111110", -- t[14526] = 1
      "0000001" when "00011100010111111", -- t[14527] = 1
      "0000001" when "00011100011000000", -- t[14528] = 1
      "0000001" when "00011100011000001", -- t[14529] = 1
      "0000001" when "00011100011000010", -- t[14530] = 1
      "0000001" when "00011100011000011", -- t[14531] = 1
      "0000001" when "00011100011000100", -- t[14532] = 1
      "0000001" when "00011100011000101", -- t[14533] = 1
      "0000001" when "00011100011000110", -- t[14534] = 1
      "0000001" when "00011100011000111", -- t[14535] = 1
      "0000001" when "00011100011001000", -- t[14536] = 1
      "0000001" when "00011100011001001", -- t[14537] = 1
      "0000001" when "00011100011001010", -- t[14538] = 1
      "0000001" when "00011100011001011", -- t[14539] = 1
      "0000001" when "00011100011001100", -- t[14540] = 1
      "0000001" when "00011100011001101", -- t[14541] = 1
      "0000001" when "00011100011001110", -- t[14542] = 1
      "0000001" when "00011100011001111", -- t[14543] = 1
      "0000001" when "00011100011010000", -- t[14544] = 1
      "0000001" when "00011100011010001", -- t[14545] = 1
      "0000001" when "00011100011010010", -- t[14546] = 1
      "0000001" when "00011100011010011", -- t[14547] = 1
      "0000001" when "00011100011010100", -- t[14548] = 1
      "0000001" when "00011100011010101", -- t[14549] = 1
      "0000001" when "00011100011010110", -- t[14550] = 1
      "0000001" when "00011100011010111", -- t[14551] = 1
      "0000001" when "00011100011011000", -- t[14552] = 1
      "0000001" when "00011100011011001", -- t[14553] = 1
      "0000001" when "00011100011011010", -- t[14554] = 1
      "0000001" when "00011100011011011", -- t[14555] = 1
      "0000001" when "00011100011011100", -- t[14556] = 1
      "0000001" when "00011100011011101", -- t[14557] = 1
      "0000001" when "00011100011011110", -- t[14558] = 1
      "0000001" when "00011100011011111", -- t[14559] = 1
      "0000001" when "00011100011100000", -- t[14560] = 1
      "0000001" when "00011100011100001", -- t[14561] = 1
      "0000001" when "00011100011100010", -- t[14562] = 1
      "0000001" when "00011100011100011", -- t[14563] = 1
      "0000001" when "00011100011100100", -- t[14564] = 1
      "0000001" when "00011100011100101", -- t[14565] = 1
      "0000001" when "00011100011100110", -- t[14566] = 1
      "0000001" when "00011100011100111", -- t[14567] = 1
      "0000001" when "00011100011101000", -- t[14568] = 1
      "0000001" when "00011100011101001", -- t[14569] = 1
      "0000001" when "00011100011101010", -- t[14570] = 1
      "0000001" when "00011100011101011", -- t[14571] = 1
      "0000001" when "00011100011101100", -- t[14572] = 1
      "0000001" when "00011100011101101", -- t[14573] = 1
      "0000001" when "00011100011101110", -- t[14574] = 1
      "0000001" when "00011100011101111", -- t[14575] = 1
      "0000001" when "00011100011110000", -- t[14576] = 1
      "0000001" when "00011100011110001", -- t[14577] = 1
      "0000001" when "00011100011110010", -- t[14578] = 1
      "0000001" when "00011100011110011", -- t[14579] = 1
      "0000001" when "00011100011110100", -- t[14580] = 1
      "0000001" when "00011100011110101", -- t[14581] = 1
      "0000001" when "00011100011110110", -- t[14582] = 1
      "0000001" when "00011100011110111", -- t[14583] = 1
      "0000001" when "00011100011111000", -- t[14584] = 1
      "0000001" when "00011100011111001", -- t[14585] = 1
      "0000001" when "00011100011111010", -- t[14586] = 1
      "0000001" when "00011100011111011", -- t[14587] = 1
      "0000001" when "00011100011111100", -- t[14588] = 1
      "0000001" when "00011100011111101", -- t[14589] = 1
      "0000001" when "00011100011111110", -- t[14590] = 1
      "0000001" when "00011100011111111", -- t[14591] = 1
      "0000001" when "00011100100000000", -- t[14592] = 1
      "0000001" when "00011100100000001", -- t[14593] = 1
      "0000001" when "00011100100000010", -- t[14594] = 1
      "0000001" when "00011100100000011", -- t[14595] = 1
      "0000001" when "00011100100000100", -- t[14596] = 1
      "0000001" when "00011100100000101", -- t[14597] = 1
      "0000001" when "00011100100000110", -- t[14598] = 1
      "0000001" when "00011100100000111", -- t[14599] = 1
      "0000001" when "00011100100001000", -- t[14600] = 1
      "0000001" when "00011100100001001", -- t[14601] = 1
      "0000001" when "00011100100001010", -- t[14602] = 1
      "0000001" when "00011100100001011", -- t[14603] = 1
      "0000001" when "00011100100001100", -- t[14604] = 1
      "0000001" when "00011100100001101", -- t[14605] = 1
      "0000001" when "00011100100001110", -- t[14606] = 1
      "0000001" when "00011100100001111", -- t[14607] = 1
      "0000001" when "00011100100010000", -- t[14608] = 1
      "0000001" when "00011100100010001", -- t[14609] = 1
      "0000001" when "00011100100010010", -- t[14610] = 1
      "0000001" when "00011100100010011", -- t[14611] = 1
      "0000001" when "00011100100010100", -- t[14612] = 1
      "0000001" when "00011100100010101", -- t[14613] = 1
      "0000001" when "00011100100010110", -- t[14614] = 1
      "0000001" when "00011100100010111", -- t[14615] = 1
      "0000001" when "00011100100011000", -- t[14616] = 1
      "0000001" when "00011100100011001", -- t[14617] = 1
      "0000001" when "00011100100011010", -- t[14618] = 1
      "0000001" when "00011100100011011", -- t[14619] = 1
      "0000001" when "00011100100011100", -- t[14620] = 1
      "0000001" when "00011100100011101", -- t[14621] = 1
      "0000001" when "00011100100011110", -- t[14622] = 1
      "0000001" when "00011100100011111", -- t[14623] = 1
      "0000001" when "00011100100100000", -- t[14624] = 1
      "0000001" when "00011100100100001", -- t[14625] = 1
      "0000001" when "00011100100100010", -- t[14626] = 1
      "0000001" when "00011100100100011", -- t[14627] = 1
      "0000001" when "00011100100100100", -- t[14628] = 1
      "0000001" when "00011100100100101", -- t[14629] = 1
      "0000001" when "00011100100100110", -- t[14630] = 1
      "0000001" when "00011100100100111", -- t[14631] = 1
      "0000001" when "00011100100101000", -- t[14632] = 1
      "0000001" when "00011100100101001", -- t[14633] = 1
      "0000001" when "00011100100101010", -- t[14634] = 1
      "0000001" when "00011100100101011", -- t[14635] = 1
      "0000001" when "00011100100101100", -- t[14636] = 1
      "0000001" when "00011100100101101", -- t[14637] = 1
      "0000001" when "00011100100101110", -- t[14638] = 1
      "0000001" when "00011100100101111", -- t[14639] = 1
      "0000001" when "00011100100110000", -- t[14640] = 1
      "0000001" when "00011100100110001", -- t[14641] = 1
      "0000001" when "00011100100110010", -- t[14642] = 1
      "0000001" when "00011100100110011", -- t[14643] = 1
      "0000001" when "00011100100110100", -- t[14644] = 1
      "0000001" when "00011100100110101", -- t[14645] = 1
      "0000001" when "00011100100110110", -- t[14646] = 1
      "0000001" when "00011100100110111", -- t[14647] = 1
      "0000001" when "00011100100111000", -- t[14648] = 1
      "0000001" when "00011100100111001", -- t[14649] = 1
      "0000001" when "00011100100111010", -- t[14650] = 1
      "0000001" when "00011100100111011", -- t[14651] = 1
      "0000001" when "00011100100111100", -- t[14652] = 1
      "0000001" when "00011100100111101", -- t[14653] = 1
      "0000001" when "00011100100111110", -- t[14654] = 1
      "0000001" when "00011100100111111", -- t[14655] = 1
      "0000001" when "00011100101000000", -- t[14656] = 1
      "0000001" when "00011100101000001", -- t[14657] = 1
      "0000001" when "00011100101000010", -- t[14658] = 1
      "0000001" when "00011100101000011", -- t[14659] = 1
      "0000001" when "00011100101000100", -- t[14660] = 1
      "0000001" when "00011100101000101", -- t[14661] = 1
      "0000001" when "00011100101000110", -- t[14662] = 1
      "0000001" when "00011100101000111", -- t[14663] = 1
      "0000001" when "00011100101001000", -- t[14664] = 1
      "0000001" when "00011100101001001", -- t[14665] = 1
      "0000001" when "00011100101001010", -- t[14666] = 1
      "0000001" when "00011100101001011", -- t[14667] = 1
      "0000001" when "00011100101001100", -- t[14668] = 1
      "0000001" when "00011100101001101", -- t[14669] = 1
      "0000001" when "00011100101001110", -- t[14670] = 1
      "0000001" when "00011100101001111", -- t[14671] = 1
      "0000001" when "00011100101010000", -- t[14672] = 1
      "0000001" when "00011100101010001", -- t[14673] = 1
      "0000001" when "00011100101010010", -- t[14674] = 1
      "0000001" when "00011100101010011", -- t[14675] = 1
      "0000001" when "00011100101010100", -- t[14676] = 1
      "0000001" when "00011100101010101", -- t[14677] = 1
      "0000001" when "00011100101010110", -- t[14678] = 1
      "0000001" when "00011100101010111", -- t[14679] = 1
      "0000001" when "00011100101011000", -- t[14680] = 1
      "0000001" when "00011100101011001", -- t[14681] = 1
      "0000001" when "00011100101011010", -- t[14682] = 1
      "0000001" when "00011100101011011", -- t[14683] = 1
      "0000001" when "00011100101011100", -- t[14684] = 1
      "0000001" when "00011100101011101", -- t[14685] = 1
      "0000001" when "00011100101011110", -- t[14686] = 1
      "0000001" when "00011100101011111", -- t[14687] = 1
      "0000001" when "00011100101100000", -- t[14688] = 1
      "0000001" when "00011100101100001", -- t[14689] = 1
      "0000001" when "00011100101100010", -- t[14690] = 1
      "0000001" when "00011100101100011", -- t[14691] = 1
      "0000001" when "00011100101100100", -- t[14692] = 1
      "0000001" when "00011100101100101", -- t[14693] = 1
      "0000001" when "00011100101100110", -- t[14694] = 1
      "0000001" when "00011100101100111", -- t[14695] = 1
      "0000001" when "00011100101101000", -- t[14696] = 1
      "0000001" when "00011100101101001", -- t[14697] = 1
      "0000001" when "00011100101101010", -- t[14698] = 1
      "0000001" when "00011100101101011", -- t[14699] = 1
      "0000001" when "00011100101101100", -- t[14700] = 1
      "0000001" when "00011100101101101", -- t[14701] = 1
      "0000001" when "00011100101101110", -- t[14702] = 1
      "0000001" when "00011100101101111", -- t[14703] = 1
      "0000001" when "00011100101110000", -- t[14704] = 1
      "0000001" when "00011100101110001", -- t[14705] = 1
      "0000001" when "00011100101110010", -- t[14706] = 1
      "0000001" when "00011100101110011", -- t[14707] = 1
      "0000001" when "00011100101110100", -- t[14708] = 1
      "0000001" when "00011100101110101", -- t[14709] = 1
      "0000001" when "00011100101110110", -- t[14710] = 1
      "0000001" when "00011100101110111", -- t[14711] = 1
      "0000001" when "00011100101111000", -- t[14712] = 1
      "0000001" when "00011100101111001", -- t[14713] = 1
      "0000001" when "00011100101111010", -- t[14714] = 1
      "0000001" when "00011100101111011", -- t[14715] = 1
      "0000001" when "00011100101111100", -- t[14716] = 1
      "0000001" when "00011100101111101", -- t[14717] = 1
      "0000001" when "00011100101111110", -- t[14718] = 1
      "0000001" when "00011100101111111", -- t[14719] = 1
      "0000001" when "00011100110000000", -- t[14720] = 1
      "0000001" when "00011100110000001", -- t[14721] = 1
      "0000001" when "00011100110000010", -- t[14722] = 1
      "0000001" when "00011100110000011", -- t[14723] = 1
      "0000001" when "00011100110000100", -- t[14724] = 1
      "0000001" when "00011100110000101", -- t[14725] = 1
      "0000001" when "00011100110000110", -- t[14726] = 1
      "0000001" when "00011100110000111", -- t[14727] = 1
      "0000001" when "00011100110001000", -- t[14728] = 1
      "0000001" when "00011100110001001", -- t[14729] = 1
      "0000001" when "00011100110001010", -- t[14730] = 1
      "0000001" when "00011100110001011", -- t[14731] = 1
      "0000001" when "00011100110001100", -- t[14732] = 1
      "0000001" when "00011100110001101", -- t[14733] = 1
      "0000001" when "00011100110001110", -- t[14734] = 1
      "0000001" when "00011100110001111", -- t[14735] = 1
      "0000001" when "00011100110010000", -- t[14736] = 1
      "0000001" when "00011100110010001", -- t[14737] = 1
      "0000001" when "00011100110010010", -- t[14738] = 1
      "0000001" when "00011100110010011", -- t[14739] = 1
      "0000001" when "00011100110010100", -- t[14740] = 1
      "0000001" when "00011100110010101", -- t[14741] = 1
      "0000001" when "00011100110010110", -- t[14742] = 1
      "0000001" when "00011100110010111", -- t[14743] = 1
      "0000001" when "00011100110011000", -- t[14744] = 1
      "0000001" when "00011100110011001", -- t[14745] = 1
      "0000001" when "00011100110011010", -- t[14746] = 1
      "0000001" when "00011100110011011", -- t[14747] = 1
      "0000001" when "00011100110011100", -- t[14748] = 1
      "0000001" when "00011100110011101", -- t[14749] = 1
      "0000001" when "00011100110011110", -- t[14750] = 1
      "0000001" when "00011100110011111", -- t[14751] = 1
      "0000001" when "00011100110100000", -- t[14752] = 1
      "0000001" when "00011100110100001", -- t[14753] = 1
      "0000001" when "00011100110100010", -- t[14754] = 1
      "0000001" when "00011100110100011", -- t[14755] = 1
      "0000001" when "00011100110100100", -- t[14756] = 1
      "0000001" when "00011100110100101", -- t[14757] = 1
      "0000001" when "00011100110100110", -- t[14758] = 1
      "0000001" when "00011100110100111", -- t[14759] = 1
      "0000001" when "00011100110101000", -- t[14760] = 1
      "0000001" when "00011100110101001", -- t[14761] = 1
      "0000001" when "00011100110101010", -- t[14762] = 1
      "0000001" when "00011100110101011", -- t[14763] = 1
      "0000001" when "00011100110101100", -- t[14764] = 1
      "0000001" when "00011100110101101", -- t[14765] = 1
      "0000001" when "00011100110101110", -- t[14766] = 1
      "0000001" when "00011100110101111", -- t[14767] = 1
      "0000001" when "00011100110110000", -- t[14768] = 1
      "0000001" when "00011100110110001", -- t[14769] = 1
      "0000001" when "00011100110110010", -- t[14770] = 1
      "0000001" when "00011100110110011", -- t[14771] = 1
      "0000001" when "00011100110110100", -- t[14772] = 1
      "0000001" when "00011100110110101", -- t[14773] = 1
      "0000001" when "00011100110110110", -- t[14774] = 1
      "0000001" when "00011100110110111", -- t[14775] = 1
      "0000001" when "00011100110111000", -- t[14776] = 1
      "0000001" when "00011100110111001", -- t[14777] = 1
      "0000001" when "00011100110111010", -- t[14778] = 1
      "0000001" when "00011100110111011", -- t[14779] = 1
      "0000001" when "00011100110111100", -- t[14780] = 1
      "0000001" when "00011100110111101", -- t[14781] = 1
      "0000001" when "00011100110111110", -- t[14782] = 1
      "0000001" when "00011100110111111", -- t[14783] = 1
      "0000001" when "00011100111000000", -- t[14784] = 1
      "0000001" when "00011100111000001", -- t[14785] = 1
      "0000001" when "00011100111000010", -- t[14786] = 1
      "0000001" when "00011100111000011", -- t[14787] = 1
      "0000001" when "00011100111000100", -- t[14788] = 1
      "0000001" when "00011100111000101", -- t[14789] = 1
      "0000001" when "00011100111000110", -- t[14790] = 1
      "0000001" when "00011100111000111", -- t[14791] = 1
      "0000001" when "00011100111001000", -- t[14792] = 1
      "0000001" when "00011100111001001", -- t[14793] = 1
      "0000001" when "00011100111001010", -- t[14794] = 1
      "0000001" when "00011100111001011", -- t[14795] = 1
      "0000001" when "00011100111001100", -- t[14796] = 1
      "0000001" when "00011100111001101", -- t[14797] = 1
      "0000001" when "00011100111001110", -- t[14798] = 1
      "0000001" when "00011100111001111", -- t[14799] = 1
      "0000001" when "00011100111010000", -- t[14800] = 1
      "0000001" when "00011100111010001", -- t[14801] = 1
      "0000001" when "00011100111010010", -- t[14802] = 1
      "0000001" when "00011100111010011", -- t[14803] = 1
      "0000001" when "00011100111010100", -- t[14804] = 1
      "0000001" when "00011100111010101", -- t[14805] = 1
      "0000001" when "00011100111010110", -- t[14806] = 1
      "0000001" when "00011100111010111", -- t[14807] = 1
      "0000001" when "00011100111011000", -- t[14808] = 1
      "0000001" when "00011100111011001", -- t[14809] = 1
      "0000001" when "00011100111011010", -- t[14810] = 1
      "0000001" when "00011100111011011", -- t[14811] = 1
      "0000001" when "00011100111011100", -- t[14812] = 1
      "0000001" when "00011100111011101", -- t[14813] = 1
      "0000001" when "00011100111011110", -- t[14814] = 1
      "0000001" when "00011100111011111", -- t[14815] = 1
      "0000001" when "00011100111100000", -- t[14816] = 1
      "0000001" when "00011100111100001", -- t[14817] = 1
      "0000001" when "00011100111100010", -- t[14818] = 1
      "0000001" when "00011100111100011", -- t[14819] = 1
      "0000001" when "00011100111100100", -- t[14820] = 1
      "0000001" when "00011100111100101", -- t[14821] = 1
      "0000001" when "00011100111100110", -- t[14822] = 1
      "0000001" when "00011100111100111", -- t[14823] = 1
      "0000001" when "00011100111101000", -- t[14824] = 1
      "0000001" when "00011100111101001", -- t[14825] = 1
      "0000001" when "00011100111101010", -- t[14826] = 1
      "0000001" when "00011100111101011", -- t[14827] = 1
      "0000001" when "00011100111101100", -- t[14828] = 1
      "0000001" when "00011100111101101", -- t[14829] = 1
      "0000001" when "00011100111101110", -- t[14830] = 1
      "0000001" when "00011100111101111", -- t[14831] = 1
      "0000001" when "00011100111110000", -- t[14832] = 1
      "0000001" when "00011100111110001", -- t[14833] = 1
      "0000001" when "00011100111110010", -- t[14834] = 1
      "0000001" when "00011100111110011", -- t[14835] = 1
      "0000001" when "00011100111110100", -- t[14836] = 1
      "0000001" when "00011100111110101", -- t[14837] = 1
      "0000001" when "00011100111110110", -- t[14838] = 1
      "0000001" when "00011100111110111", -- t[14839] = 1
      "0000001" when "00011100111111000", -- t[14840] = 1
      "0000001" when "00011100111111001", -- t[14841] = 1
      "0000001" when "00011100111111010", -- t[14842] = 1
      "0000001" when "00011100111111011", -- t[14843] = 1
      "0000001" when "00011100111111100", -- t[14844] = 1
      "0000001" when "00011100111111101", -- t[14845] = 1
      "0000001" when "00011100111111110", -- t[14846] = 1
      "0000001" when "00011100111111111", -- t[14847] = 1
      "0000001" when "00011101000000000", -- t[14848] = 1
      "0000001" when "00011101000000001", -- t[14849] = 1
      "0000001" when "00011101000000010", -- t[14850] = 1
      "0000001" when "00011101000000011", -- t[14851] = 1
      "0000001" when "00011101000000100", -- t[14852] = 1
      "0000001" when "00011101000000101", -- t[14853] = 1
      "0000001" when "00011101000000110", -- t[14854] = 1
      "0000001" when "00011101000000111", -- t[14855] = 1
      "0000001" when "00011101000001000", -- t[14856] = 1
      "0000001" when "00011101000001001", -- t[14857] = 1
      "0000001" when "00011101000001010", -- t[14858] = 1
      "0000001" when "00011101000001011", -- t[14859] = 1
      "0000001" when "00011101000001100", -- t[14860] = 1
      "0000001" when "00011101000001101", -- t[14861] = 1
      "0000001" when "00011101000001110", -- t[14862] = 1
      "0000001" when "00011101000001111", -- t[14863] = 1
      "0000001" when "00011101000010000", -- t[14864] = 1
      "0000001" when "00011101000010001", -- t[14865] = 1
      "0000001" when "00011101000010010", -- t[14866] = 1
      "0000001" when "00011101000010011", -- t[14867] = 1
      "0000001" when "00011101000010100", -- t[14868] = 1
      "0000001" when "00011101000010101", -- t[14869] = 1
      "0000001" when "00011101000010110", -- t[14870] = 1
      "0000001" when "00011101000010111", -- t[14871] = 1
      "0000001" when "00011101000011000", -- t[14872] = 1
      "0000001" when "00011101000011001", -- t[14873] = 1
      "0000001" when "00011101000011010", -- t[14874] = 1
      "0000001" when "00011101000011011", -- t[14875] = 1
      "0000001" when "00011101000011100", -- t[14876] = 1
      "0000001" when "00011101000011101", -- t[14877] = 1
      "0000001" when "00011101000011110", -- t[14878] = 1
      "0000001" when "00011101000011111", -- t[14879] = 1
      "0000001" when "00011101000100000", -- t[14880] = 1
      "0000001" when "00011101000100001", -- t[14881] = 1
      "0000001" when "00011101000100010", -- t[14882] = 1
      "0000001" when "00011101000100011", -- t[14883] = 1
      "0000001" when "00011101000100100", -- t[14884] = 1
      "0000001" when "00011101000100101", -- t[14885] = 1
      "0000001" when "00011101000100110", -- t[14886] = 1
      "0000001" when "00011101000100111", -- t[14887] = 1
      "0000001" when "00011101000101000", -- t[14888] = 1
      "0000001" when "00011101000101001", -- t[14889] = 1
      "0000001" when "00011101000101010", -- t[14890] = 1
      "0000001" when "00011101000101011", -- t[14891] = 1
      "0000001" when "00011101000101100", -- t[14892] = 1
      "0000001" when "00011101000101101", -- t[14893] = 1
      "0000001" when "00011101000101110", -- t[14894] = 1
      "0000001" when "00011101000101111", -- t[14895] = 1
      "0000001" when "00011101000110000", -- t[14896] = 1
      "0000001" when "00011101000110001", -- t[14897] = 1
      "0000001" when "00011101000110010", -- t[14898] = 1
      "0000001" when "00011101000110011", -- t[14899] = 1
      "0000001" when "00011101000110100", -- t[14900] = 1
      "0000001" when "00011101000110101", -- t[14901] = 1
      "0000001" when "00011101000110110", -- t[14902] = 1
      "0000001" when "00011101000110111", -- t[14903] = 1
      "0000001" when "00011101000111000", -- t[14904] = 1
      "0000001" when "00011101000111001", -- t[14905] = 1
      "0000001" when "00011101000111010", -- t[14906] = 1
      "0000001" when "00011101000111011", -- t[14907] = 1
      "0000001" when "00011101000111100", -- t[14908] = 1
      "0000001" when "00011101000111101", -- t[14909] = 1
      "0000001" when "00011101000111110", -- t[14910] = 1
      "0000001" when "00011101000111111", -- t[14911] = 1
      "0000001" when "00011101001000000", -- t[14912] = 1
      "0000001" when "00011101001000001", -- t[14913] = 1
      "0000001" when "00011101001000010", -- t[14914] = 1
      "0000001" when "00011101001000011", -- t[14915] = 1
      "0000001" when "00011101001000100", -- t[14916] = 1
      "0000001" when "00011101001000101", -- t[14917] = 1
      "0000001" when "00011101001000110", -- t[14918] = 1
      "0000001" when "00011101001000111", -- t[14919] = 1
      "0000001" when "00011101001001000", -- t[14920] = 1
      "0000001" when "00011101001001001", -- t[14921] = 1
      "0000001" when "00011101001001010", -- t[14922] = 1
      "0000001" when "00011101001001011", -- t[14923] = 1
      "0000001" when "00011101001001100", -- t[14924] = 1
      "0000001" when "00011101001001101", -- t[14925] = 1
      "0000001" when "00011101001001110", -- t[14926] = 1
      "0000001" when "00011101001001111", -- t[14927] = 1
      "0000001" when "00011101001010000", -- t[14928] = 1
      "0000001" when "00011101001010001", -- t[14929] = 1
      "0000001" when "00011101001010010", -- t[14930] = 1
      "0000001" when "00011101001010011", -- t[14931] = 1
      "0000001" when "00011101001010100", -- t[14932] = 1
      "0000001" when "00011101001010101", -- t[14933] = 1
      "0000001" when "00011101001010110", -- t[14934] = 1
      "0000001" when "00011101001010111", -- t[14935] = 1
      "0000001" when "00011101001011000", -- t[14936] = 1
      "0000001" when "00011101001011001", -- t[14937] = 1
      "0000001" when "00011101001011010", -- t[14938] = 1
      "0000001" when "00011101001011011", -- t[14939] = 1
      "0000001" when "00011101001011100", -- t[14940] = 1
      "0000001" when "00011101001011101", -- t[14941] = 1
      "0000001" when "00011101001011110", -- t[14942] = 1
      "0000001" when "00011101001011111", -- t[14943] = 1
      "0000001" when "00011101001100000", -- t[14944] = 1
      "0000001" when "00011101001100001", -- t[14945] = 1
      "0000001" when "00011101001100010", -- t[14946] = 1
      "0000001" when "00011101001100011", -- t[14947] = 1
      "0000001" when "00011101001100100", -- t[14948] = 1
      "0000001" when "00011101001100101", -- t[14949] = 1
      "0000001" when "00011101001100110", -- t[14950] = 1
      "0000001" when "00011101001100111", -- t[14951] = 1
      "0000001" when "00011101001101000", -- t[14952] = 1
      "0000001" when "00011101001101001", -- t[14953] = 1
      "0000001" when "00011101001101010", -- t[14954] = 1
      "0000001" when "00011101001101011", -- t[14955] = 1
      "0000001" when "00011101001101100", -- t[14956] = 1
      "0000001" when "00011101001101101", -- t[14957] = 1
      "0000001" when "00011101001101110", -- t[14958] = 1
      "0000001" when "00011101001101111", -- t[14959] = 1
      "0000001" when "00011101001110000", -- t[14960] = 1
      "0000001" when "00011101001110001", -- t[14961] = 1
      "0000001" when "00011101001110010", -- t[14962] = 1
      "0000001" when "00011101001110011", -- t[14963] = 1
      "0000001" when "00011101001110100", -- t[14964] = 1
      "0000001" when "00011101001110101", -- t[14965] = 1
      "0000001" when "00011101001110110", -- t[14966] = 1
      "0000001" when "00011101001110111", -- t[14967] = 1
      "0000001" when "00011101001111000", -- t[14968] = 1
      "0000001" when "00011101001111001", -- t[14969] = 1
      "0000001" when "00011101001111010", -- t[14970] = 1
      "0000001" when "00011101001111011", -- t[14971] = 1
      "0000001" when "00011101001111100", -- t[14972] = 1
      "0000001" when "00011101001111101", -- t[14973] = 1
      "0000001" when "00011101001111110", -- t[14974] = 1
      "0000001" when "00011101001111111", -- t[14975] = 1
      "0000001" when "00011101010000000", -- t[14976] = 1
      "0000001" when "00011101010000001", -- t[14977] = 1
      "0000001" when "00011101010000010", -- t[14978] = 1
      "0000001" when "00011101010000011", -- t[14979] = 1
      "0000001" when "00011101010000100", -- t[14980] = 1
      "0000001" when "00011101010000101", -- t[14981] = 1
      "0000001" when "00011101010000110", -- t[14982] = 1
      "0000001" when "00011101010000111", -- t[14983] = 1
      "0000001" when "00011101010001000", -- t[14984] = 1
      "0000001" when "00011101010001001", -- t[14985] = 1
      "0000001" when "00011101010001010", -- t[14986] = 1
      "0000001" when "00011101010001011", -- t[14987] = 1
      "0000001" when "00011101010001100", -- t[14988] = 1
      "0000001" when "00011101010001101", -- t[14989] = 1
      "0000001" when "00011101010001110", -- t[14990] = 1
      "0000001" when "00011101010001111", -- t[14991] = 1
      "0000001" when "00011101010010000", -- t[14992] = 1
      "0000001" when "00011101010010001", -- t[14993] = 1
      "0000001" when "00011101010010010", -- t[14994] = 1
      "0000001" when "00011101010010011", -- t[14995] = 1
      "0000001" when "00011101010010100", -- t[14996] = 1
      "0000001" when "00011101010010101", -- t[14997] = 1
      "0000001" when "00011101010010110", -- t[14998] = 1
      "0000001" when "00011101010010111", -- t[14999] = 1
      "0000001" when "00011101010011000", -- t[15000] = 1
      "0000001" when "00011101010011001", -- t[15001] = 1
      "0000001" when "00011101010011010", -- t[15002] = 1
      "0000001" when "00011101010011011", -- t[15003] = 1
      "0000001" when "00011101010011100", -- t[15004] = 1
      "0000001" when "00011101010011101", -- t[15005] = 1
      "0000001" when "00011101010011110", -- t[15006] = 1
      "0000001" when "00011101010011111", -- t[15007] = 1
      "0000001" when "00011101010100000", -- t[15008] = 1
      "0000001" when "00011101010100001", -- t[15009] = 1
      "0000001" when "00011101010100010", -- t[15010] = 1
      "0000001" when "00011101010100011", -- t[15011] = 1
      "0000001" when "00011101010100100", -- t[15012] = 1
      "0000001" when "00011101010100101", -- t[15013] = 1
      "0000001" when "00011101010100110", -- t[15014] = 1
      "0000001" when "00011101010100111", -- t[15015] = 1
      "0000001" when "00011101010101000", -- t[15016] = 1
      "0000001" when "00011101010101001", -- t[15017] = 1
      "0000001" when "00011101010101010", -- t[15018] = 1
      "0000001" when "00011101010101011", -- t[15019] = 1
      "0000001" when "00011101010101100", -- t[15020] = 1
      "0000001" when "00011101010101101", -- t[15021] = 1
      "0000001" when "00011101010101110", -- t[15022] = 1
      "0000001" when "00011101010101111", -- t[15023] = 1
      "0000001" when "00011101010110000", -- t[15024] = 1
      "0000001" when "00011101010110001", -- t[15025] = 1
      "0000001" when "00011101010110010", -- t[15026] = 1
      "0000001" when "00011101010110011", -- t[15027] = 1
      "0000001" when "00011101010110100", -- t[15028] = 1
      "0000001" when "00011101010110101", -- t[15029] = 1
      "0000001" when "00011101010110110", -- t[15030] = 1
      "0000001" when "00011101010110111", -- t[15031] = 1
      "0000001" when "00011101010111000", -- t[15032] = 1
      "0000001" when "00011101010111001", -- t[15033] = 1
      "0000001" when "00011101010111010", -- t[15034] = 1
      "0000001" when "00011101010111011", -- t[15035] = 1
      "0000001" when "00011101010111100", -- t[15036] = 1
      "0000001" when "00011101010111101", -- t[15037] = 1
      "0000001" when "00011101010111110", -- t[15038] = 1
      "0000001" when "00011101010111111", -- t[15039] = 1
      "0000001" when "00011101011000000", -- t[15040] = 1
      "0000001" when "00011101011000001", -- t[15041] = 1
      "0000001" when "00011101011000010", -- t[15042] = 1
      "0000001" when "00011101011000011", -- t[15043] = 1
      "0000001" when "00011101011000100", -- t[15044] = 1
      "0000001" when "00011101011000101", -- t[15045] = 1
      "0000001" when "00011101011000110", -- t[15046] = 1
      "0000001" when "00011101011000111", -- t[15047] = 1
      "0000001" when "00011101011001000", -- t[15048] = 1
      "0000001" when "00011101011001001", -- t[15049] = 1
      "0000001" when "00011101011001010", -- t[15050] = 1
      "0000001" when "00011101011001011", -- t[15051] = 1
      "0000001" when "00011101011001100", -- t[15052] = 1
      "0000001" when "00011101011001101", -- t[15053] = 1
      "0000001" when "00011101011001110", -- t[15054] = 1
      "0000001" when "00011101011001111", -- t[15055] = 1
      "0000001" when "00011101011010000", -- t[15056] = 1
      "0000001" when "00011101011010001", -- t[15057] = 1
      "0000001" when "00011101011010010", -- t[15058] = 1
      "0000001" when "00011101011010011", -- t[15059] = 1
      "0000001" when "00011101011010100", -- t[15060] = 1
      "0000001" when "00011101011010101", -- t[15061] = 1
      "0000001" when "00011101011010110", -- t[15062] = 1
      "0000001" when "00011101011010111", -- t[15063] = 1
      "0000001" when "00011101011011000", -- t[15064] = 1
      "0000001" when "00011101011011001", -- t[15065] = 1
      "0000001" when "00011101011011010", -- t[15066] = 1
      "0000001" when "00011101011011011", -- t[15067] = 1
      "0000001" when "00011101011011100", -- t[15068] = 1
      "0000001" when "00011101011011101", -- t[15069] = 1
      "0000001" when "00011101011011110", -- t[15070] = 1
      "0000001" when "00011101011011111", -- t[15071] = 1
      "0000001" when "00011101011100000", -- t[15072] = 1
      "0000001" when "00011101011100001", -- t[15073] = 1
      "0000001" when "00011101011100010", -- t[15074] = 1
      "0000001" when "00011101011100011", -- t[15075] = 1
      "0000001" when "00011101011100100", -- t[15076] = 1
      "0000001" when "00011101011100101", -- t[15077] = 1
      "0000001" when "00011101011100110", -- t[15078] = 1
      "0000001" when "00011101011100111", -- t[15079] = 1
      "0000001" when "00011101011101000", -- t[15080] = 1
      "0000001" when "00011101011101001", -- t[15081] = 1
      "0000001" when "00011101011101010", -- t[15082] = 1
      "0000001" when "00011101011101011", -- t[15083] = 1
      "0000001" when "00011101011101100", -- t[15084] = 1
      "0000001" when "00011101011101101", -- t[15085] = 1
      "0000001" when "00011101011101110", -- t[15086] = 1
      "0000001" when "00011101011101111", -- t[15087] = 1
      "0000001" when "00011101011110000", -- t[15088] = 1
      "0000001" when "00011101011110001", -- t[15089] = 1
      "0000001" when "00011101011110010", -- t[15090] = 1
      "0000001" when "00011101011110011", -- t[15091] = 1
      "0000001" when "00011101011110100", -- t[15092] = 1
      "0000001" when "00011101011110101", -- t[15093] = 1
      "0000001" when "00011101011110110", -- t[15094] = 1
      "0000001" when "00011101011110111", -- t[15095] = 1
      "0000001" when "00011101011111000", -- t[15096] = 1
      "0000001" when "00011101011111001", -- t[15097] = 1
      "0000001" when "00011101011111010", -- t[15098] = 1
      "0000001" when "00011101011111011", -- t[15099] = 1
      "0000001" when "00011101011111100", -- t[15100] = 1
      "0000001" when "00011101011111101", -- t[15101] = 1
      "0000001" when "00011101011111110", -- t[15102] = 1
      "0000001" when "00011101011111111", -- t[15103] = 1
      "0000001" when "00011101100000000", -- t[15104] = 1
      "0000001" when "00011101100000001", -- t[15105] = 1
      "0000001" when "00011101100000010", -- t[15106] = 1
      "0000001" when "00011101100000011", -- t[15107] = 1
      "0000001" when "00011101100000100", -- t[15108] = 1
      "0000001" when "00011101100000101", -- t[15109] = 1
      "0000001" when "00011101100000110", -- t[15110] = 1
      "0000001" when "00011101100000111", -- t[15111] = 1
      "0000001" when "00011101100001000", -- t[15112] = 1
      "0000001" when "00011101100001001", -- t[15113] = 1
      "0000001" when "00011101100001010", -- t[15114] = 1
      "0000001" when "00011101100001011", -- t[15115] = 1
      "0000001" when "00011101100001100", -- t[15116] = 1
      "0000001" when "00011101100001101", -- t[15117] = 1
      "0000001" when "00011101100001110", -- t[15118] = 1
      "0000001" when "00011101100001111", -- t[15119] = 1
      "0000001" when "00011101100010000", -- t[15120] = 1
      "0000001" when "00011101100010001", -- t[15121] = 1
      "0000001" when "00011101100010010", -- t[15122] = 1
      "0000001" when "00011101100010011", -- t[15123] = 1
      "0000001" when "00011101100010100", -- t[15124] = 1
      "0000001" when "00011101100010101", -- t[15125] = 1
      "0000001" when "00011101100010110", -- t[15126] = 1
      "0000001" when "00011101100010111", -- t[15127] = 1
      "0000001" when "00011101100011000", -- t[15128] = 1
      "0000001" when "00011101100011001", -- t[15129] = 1
      "0000001" when "00011101100011010", -- t[15130] = 1
      "0000001" when "00011101100011011", -- t[15131] = 1
      "0000001" when "00011101100011100", -- t[15132] = 1
      "0000001" when "00011101100011101", -- t[15133] = 1
      "0000001" when "00011101100011110", -- t[15134] = 1
      "0000001" when "00011101100011111", -- t[15135] = 1
      "0000001" when "00011101100100000", -- t[15136] = 1
      "0000001" when "00011101100100001", -- t[15137] = 1
      "0000001" when "00011101100100010", -- t[15138] = 1
      "0000001" when "00011101100100011", -- t[15139] = 1
      "0000001" when "00011101100100100", -- t[15140] = 1
      "0000001" when "00011101100100101", -- t[15141] = 1
      "0000001" when "00011101100100110", -- t[15142] = 1
      "0000001" when "00011101100100111", -- t[15143] = 1
      "0000001" when "00011101100101000", -- t[15144] = 1
      "0000001" when "00011101100101001", -- t[15145] = 1
      "0000001" when "00011101100101010", -- t[15146] = 1
      "0000001" when "00011101100101011", -- t[15147] = 1
      "0000001" when "00011101100101100", -- t[15148] = 1
      "0000001" when "00011101100101101", -- t[15149] = 1
      "0000001" when "00011101100101110", -- t[15150] = 1
      "0000001" when "00011101100101111", -- t[15151] = 1
      "0000001" when "00011101100110000", -- t[15152] = 1
      "0000001" when "00011101100110001", -- t[15153] = 1
      "0000001" when "00011101100110010", -- t[15154] = 1
      "0000001" when "00011101100110011", -- t[15155] = 1
      "0000001" when "00011101100110100", -- t[15156] = 1
      "0000001" when "00011101100110101", -- t[15157] = 1
      "0000001" when "00011101100110110", -- t[15158] = 1
      "0000001" when "00011101100110111", -- t[15159] = 1
      "0000001" when "00011101100111000", -- t[15160] = 1
      "0000001" when "00011101100111001", -- t[15161] = 1
      "0000001" when "00011101100111010", -- t[15162] = 1
      "0000001" when "00011101100111011", -- t[15163] = 1
      "0000001" when "00011101100111100", -- t[15164] = 1
      "0000001" when "00011101100111101", -- t[15165] = 1
      "0000001" when "00011101100111110", -- t[15166] = 1
      "0000001" when "00011101100111111", -- t[15167] = 1
      "0000001" when "00011101101000000", -- t[15168] = 1
      "0000001" when "00011101101000001", -- t[15169] = 1
      "0000001" when "00011101101000010", -- t[15170] = 1
      "0000001" when "00011101101000011", -- t[15171] = 1
      "0000001" when "00011101101000100", -- t[15172] = 1
      "0000001" when "00011101101000101", -- t[15173] = 1
      "0000001" when "00011101101000110", -- t[15174] = 1
      "0000001" when "00011101101000111", -- t[15175] = 1
      "0000001" when "00011101101001000", -- t[15176] = 1
      "0000001" when "00011101101001001", -- t[15177] = 1
      "0000001" when "00011101101001010", -- t[15178] = 1
      "0000001" when "00011101101001011", -- t[15179] = 1
      "0000001" when "00011101101001100", -- t[15180] = 1
      "0000001" when "00011101101001101", -- t[15181] = 1
      "0000001" when "00011101101001110", -- t[15182] = 1
      "0000001" when "00011101101001111", -- t[15183] = 1
      "0000001" when "00011101101010000", -- t[15184] = 1
      "0000001" when "00011101101010001", -- t[15185] = 1
      "0000001" when "00011101101010010", -- t[15186] = 1
      "0000001" when "00011101101010011", -- t[15187] = 1
      "0000001" when "00011101101010100", -- t[15188] = 1
      "0000001" when "00011101101010101", -- t[15189] = 1
      "0000001" when "00011101101010110", -- t[15190] = 1
      "0000001" when "00011101101010111", -- t[15191] = 1
      "0000001" when "00011101101011000", -- t[15192] = 1
      "0000001" when "00011101101011001", -- t[15193] = 1
      "0000001" when "00011101101011010", -- t[15194] = 1
      "0000001" when "00011101101011011", -- t[15195] = 1
      "0000001" when "00011101101011100", -- t[15196] = 1
      "0000001" when "00011101101011101", -- t[15197] = 1
      "0000001" when "00011101101011110", -- t[15198] = 1
      "0000001" when "00011101101011111", -- t[15199] = 1
      "0000001" when "00011101101100000", -- t[15200] = 1
      "0000001" when "00011101101100001", -- t[15201] = 1
      "0000001" when "00011101101100010", -- t[15202] = 1
      "0000001" when "00011101101100011", -- t[15203] = 1
      "0000001" when "00011101101100100", -- t[15204] = 1
      "0000001" when "00011101101100101", -- t[15205] = 1
      "0000001" when "00011101101100110", -- t[15206] = 1
      "0000001" when "00011101101100111", -- t[15207] = 1
      "0000001" when "00011101101101000", -- t[15208] = 1
      "0000001" when "00011101101101001", -- t[15209] = 1
      "0000001" when "00011101101101010", -- t[15210] = 1
      "0000001" when "00011101101101011", -- t[15211] = 1
      "0000001" when "00011101101101100", -- t[15212] = 1
      "0000001" when "00011101101101101", -- t[15213] = 1
      "0000001" when "00011101101101110", -- t[15214] = 1
      "0000001" when "00011101101101111", -- t[15215] = 1
      "0000001" when "00011101101110000", -- t[15216] = 1
      "0000001" when "00011101101110001", -- t[15217] = 1
      "0000001" when "00011101101110010", -- t[15218] = 1
      "0000001" when "00011101101110011", -- t[15219] = 1
      "0000001" when "00011101101110100", -- t[15220] = 1
      "0000001" when "00011101101110101", -- t[15221] = 1
      "0000001" when "00011101101110110", -- t[15222] = 1
      "0000001" when "00011101101110111", -- t[15223] = 1
      "0000001" when "00011101101111000", -- t[15224] = 1
      "0000001" when "00011101101111001", -- t[15225] = 1
      "0000001" when "00011101101111010", -- t[15226] = 1
      "0000001" when "00011101101111011", -- t[15227] = 1
      "0000001" when "00011101101111100", -- t[15228] = 1
      "0000001" when "00011101101111101", -- t[15229] = 1
      "0000001" when "00011101101111110", -- t[15230] = 1
      "0000001" when "00011101101111111", -- t[15231] = 1
      "0000001" when "00011101110000000", -- t[15232] = 1
      "0000001" when "00011101110000001", -- t[15233] = 1
      "0000001" when "00011101110000010", -- t[15234] = 1
      "0000001" when "00011101110000011", -- t[15235] = 1
      "0000001" when "00011101110000100", -- t[15236] = 1
      "0000001" when "00011101110000101", -- t[15237] = 1
      "0000001" when "00011101110000110", -- t[15238] = 1
      "0000001" when "00011101110000111", -- t[15239] = 1
      "0000001" when "00011101110001000", -- t[15240] = 1
      "0000001" when "00011101110001001", -- t[15241] = 1
      "0000001" when "00011101110001010", -- t[15242] = 1
      "0000001" when "00011101110001011", -- t[15243] = 1
      "0000001" when "00011101110001100", -- t[15244] = 1
      "0000001" when "00011101110001101", -- t[15245] = 1
      "0000001" when "00011101110001110", -- t[15246] = 1
      "0000001" when "00011101110001111", -- t[15247] = 1
      "0000001" when "00011101110010000", -- t[15248] = 1
      "0000001" when "00011101110010001", -- t[15249] = 1
      "0000001" when "00011101110010010", -- t[15250] = 1
      "0000001" when "00011101110010011", -- t[15251] = 1
      "0000001" when "00011101110010100", -- t[15252] = 1
      "0000001" when "00011101110010101", -- t[15253] = 1
      "0000001" when "00011101110010110", -- t[15254] = 1
      "0000001" when "00011101110010111", -- t[15255] = 1
      "0000001" when "00011101110011000", -- t[15256] = 1
      "0000001" when "00011101110011001", -- t[15257] = 1
      "0000001" when "00011101110011010", -- t[15258] = 1
      "0000001" when "00011101110011011", -- t[15259] = 1
      "0000001" when "00011101110011100", -- t[15260] = 1
      "0000001" when "00011101110011101", -- t[15261] = 1
      "0000001" when "00011101110011110", -- t[15262] = 1
      "0000001" when "00011101110011111", -- t[15263] = 1
      "0000001" when "00011101110100000", -- t[15264] = 1
      "0000001" when "00011101110100001", -- t[15265] = 1
      "0000001" when "00011101110100010", -- t[15266] = 1
      "0000001" when "00011101110100011", -- t[15267] = 1
      "0000001" when "00011101110100100", -- t[15268] = 1
      "0000001" when "00011101110100101", -- t[15269] = 1
      "0000001" when "00011101110100110", -- t[15270] = 1
      "0000001" when "00011101110100111", -- t[15271] = 1
      "0000001" when "00011101110101000", -- t[15272] = 1
      "0000001" when "00011101110101001", -- t[15273] = 1
      "0000001" when "00011101110101010", -- t[15274] = 1
      "0000001" when "00011101110101011", -- t[15275] = 1
      "0000001" when "00011101110101100", -- t[15276] = 1
      "0000001" when "00011101110101101", -- t[15277] = 1
      "0000001" when "00011101110101110", -- t[15278] = 1
      "0000001" when "00011101110101111", -- t[15279] = 1
      "0000001" when "00011101110110000", -- t[15280] = 1
      "0000001" when "00011101110110001", -- t[15281] = 1
      "0000001" when "00011101110110010", -- t[15282] = 1
      "0000001" when "00011101110110011", -- t[15283] = 1
      "0000001" when "00011101110110100", -- t[15284] = 1
      "0000001" when "00011101110110101", -- t[15285] = 1
      "0000001" when "00011101110110110", -- t[15286] = 1
      "0000001" when "00011101110110111", -- t[15287] = 1
      "0000001" when "00011101110111000", -- t[15288] = 1
      "0000001" when "00011101110111001", -- t[15289] = 1
      "0000001" when "00011101110111010", -- t[15290] = 1
      "0000001" when "00011101110111011", -- t[15291] = 1
      "0000001" when "00011101110111100", -- t[15292] = 1
      "0000001" when "00011101110111101", -- t[15293] = 1
      "0000001" when "00011101110111110", -- t[15294] = 1
      "0000001" when "00011101110111111", -- t[15295] = 1
      "0000001" when "00011101111000000", -- t[15296] = 1
      "0000001" when "00011101111000001", -- t[15297] = 1
      "0000001" when "00011101111000010", -- t[15298] = 1
      "0000001" when "00011101111000011", -- t[15299] = 1
      "0000001" when "00011101111000100", -- t[15300] = 1
      "0000001" when "00011101111000101", -- t[15301] = 1
      "0000001" when "00011101111000110", -- t[15302] = 1
      "0000001" when "00011101111000111", -- t[15303] = 1
      "0000001" when "00011101111001000", -- t[15304] = 1
      "0000001" when "00011101111001001", -- t[15305] = 1
      "0000001" when "00011101111001010", -- t[15306] = 1
      "0000001" when "00011101111001011", -- t[15307] = 1
      "0000001" when "00011101111001100", -- t[15308] = 1
      "0000001" when "00011101111001101", -- t[15309] = 1
      "0000001" when "00011101111001110", -- t[15310] = 1
      "0000001" when "00011101111001111", -- t[15311] = 1
      "0000001" when "00011101111010000", -- t[15312] = 1
      "0000001" when "00011101111010001", -- t[15313] = 1
      "0000001" when "00011101111010010", -- t[15314] = 1
      "0000001" when "00011101111010011", -- t[15315] = 1
      "0000001" when "00011101111010100", -- t[15316] = 1
      "0000001" when "00011101111010101", -- t[15317] = 1
      "0000001" when "00011101111010110", -- t[15318] = 1
      "0000001" when "00011101111010111", -- t[15319] = 1
      "0000001" when "00011101111011000", -- t[15320] = 1
      "0000001" when "00011101111011001", -- t[15321] = 1
      "0000001" when "00011101111011010", -- t[15322] = 1
      "0000001" when "00011101111011011", -- t[15323] = 1
      "0000001" when "00011101111011100", -- t[15324] = 1
      "0000001" when "00011101111011101", -- t[15325] = 1
      "0000001" when "00011101111011110", -- t[15326] = 1
      "0000001" when "00011101111011111", -- t[15327] = 1
      "0000001" when "00011101111100000", -- t[15328] = 1
      "0000001" when "00011101111100001", -- t[15329] = 1
      "0000001" when "00011101111100010", -- t[15330] = 1
      "0000001" when "00011101111100011", -- t[15331] = 1
      "0000001" when "00011101111100100", -- t[15332] = 1
      "0000001" when "00011101111100101", -- t[15333] = 1
      "0000001" when "00011101111100110", -- t[15334] = 1
      "0000001" when "00011101111100111", -- t[15335] = 1
      "0000001" when "00011101111101000", -- t[15336] = 1
      "0000001" when "00011101111101001", -- t[15337] = 1
      "0000001" when "00011101111101010", -- t[15338] = 1
      "0000001" when "00011101111101011", -- t[15339] = 1
      "0000001" when "00011101111101100", -- t[15340] = 1
      "0000001" when "00011101111101101", -- t[15341] = 1
      "0000001" when "00011101111101110", -- t[15342] = 1
      "0000001" when "00011101111101111", -- t[15343] = 1
      "0000001" when "00011101111110000", -- t[15344] = 1
      "0000001" when "00011101111110001", -- t[15345] = 1
      "0000001" when "00011101111110010", -- t[15346] = 1
      "0000001" when "00011101111110011", -- t[15347] = 1
      "0000001" when "00011101111110100", -- t[15348] = 1
      "0000001" when "00011101111110101", -- t[15349] = 1
      "0000001" when "00011101111110110", -- t[15350] = 1
      "0000001" when "00011101111110111", -- t[15351] = 1
      "0000001" when "00011101111111000", -- t[15352] = 1
      "0000001" when "00011101111111001", -- t[15353] = 1
      "0000001" when "00011101111111010", -- t[15354] = 1
      "0000001" when "00011101111111011", -- t[15355] = 1
      "0000001" when "00011101111111100", -- t[15356] = 1
      "0000001" when "00011101111111101", -- t[15357] = 1
      "0000001" when "00011101111111110", -- t[15358] = 1
      "0000001" when "00011101111111111", -- t[15359] = 1
      "0000001" when "00011110000000000", -- t[15360] = 1
      "0000001" when "00011110000000001", -- t[15361] = 1
      "0000001" when "00011110000000010", -- t[15362] = 1
      "0000001" when "00011110000000011", -- t[15363] = 1
      "0000001" when "00011110000000100", -- t[15364] = 1
      "0000001" when "00011110000000101", -- t[15365] = 1
      "0000001" when "00011110000000110", -- t[15366] = 1
      "0000001" when "00011110000000111", -- t[15367] = 1
      "0000001" when "00011110000001000", -- t[15368] = 1
      "0000001" when "00011110000001001", -- t[15369] = 1
      "0000001" when "00011110000001010", -- t[15370] = 1
      "0000001" when "00011110000001011", -- t[15371] = 1
      "0000001" when "00011110000001100", -- t[15372] = 1
      "0000001" when "00011110000001101", -- t[15373] = 1
      "0000001" when "00011110000001110", -- t[15374] = 1
      "0000001" when "00011110000001111", -- t[15375] = 1
      "0000001" when "00011110000010000", -- t[15376] = 1
      "0000001" when "00011110000010001", -- t[15377] = 1
      "0000001" when "00011110000010010", -- t[15378] = 1
      "0000001" when "00011110000010011", -- t[15379] = 1
      "0000001" when "00011110000010100", -- t[15380] = 1
      "0000001" when "00011110000010101", -- t[15381] = 1
      "0000001" when "00011110000010110", -- t[15382] = 1
      "0000001" when "00011110000010111", -- t[15383] = 1
      "0000001" when "00011110000011000", -- t[15384] = 1
      "0000001" when "00011110000011001", -- t[15385] = 1
      "0000001" when "00011110000011010", -- t[15386] = 1
      "0000001" when "00011110000011011", -- t[15387] = 1
      "0000001" when "00011110000011100", -- t[15388] = 1
      "0000001" when "00011110000011101", -- t[15389] = 1
      "0000001" when "00011110000011110", -- t[15390] = 1
      "0000001" when "00011110000011111", -- t[15391] = 1
      "0000001" when "00011110000100000", -- t[15392] = 1
      "0000001" when "00011110000100001", -- t[15393] = 1
      "0000001" when "00011110000100010", -- t[15394] = 1
      "0000001" when "00011110000100011", -- t[15395] = 1
      "0000001" when "00011110000100100", -- t[15396] = 1
      "0000001" when "00011110000100101", -- t[15397] = 1
      "0000001" when "00011110000100110", -- t[15398] = 1
      "0000001" when "00011110000100111", -- t[15399] = 1
      "0000001" when "00011110000101000", -- t[15400] = 1
      "0000001" when "00011110000101001", -- t[15401] = 1
      "0000001" when "00011110000101010", -- t[15402] = 1
      "0000001" when "00011110000101011", -- t[15403] = 1
      "0000001" when "00011110000101100", -- t[15404] = 1
      "0000001" when "00011110000101101", -- t[15405] = 1
      "0000001" when "00011110000101110", -- t[15406] = 1
      "0000001" when "00011110000101111", -- t[15407] = 1
      "0000001" when "00011110000110000", -- t[15408] = 1
      "0000001" when "00011110000110001", -- t[15409] = 1
      "0000001" when "00011110000110010", -- t[15410] = 1
      "0000001" when "00011110000110011", -- t[15411] = 1
      "0000001" when "00011110000110100", -- t[15412] = 1
      "0000001" when "00011110000110101", -- t[15413] = 1
      "0000001" when "00011110000110110", -- t[15414] = 1
      "0000001" when "00011110000110111", -- t[15415] = 1
      "0000001" when "00011110000111000", -- t[15416] = 1
      "0000001" when "00011110000111001", -- t[15417] = 1
      "0000001" when "00011110000111010", -- t[15418] = 1
      "0000001" when "00011110000111011", -- t[15419] = 1
      "0000001" when "00011110000111100", -- t[15420] = 1
      "0000001" when "00011110000111101", -- t[15421] = 1
      "0000001" when "00011110000111110", -- t[15422] = 1
      "0000001" when "00011110000111111", -- t[15423] = 1
      "0000001" when "00011110001000000", -- t[15424] = 1
      "0000001" when "00011110001000001", -- t[15425] = 1
      "0000001" when "00011110001000010", -- t[15426] = 1
      "0000001" when "00011110001000011", -- t[15427] = 1
      "0000001" when "00011110001000100", -- t[15428] = 1
      "0000001" when "00011110001000101", -- t[15429] = 1
      "0000001" when "00011110001000110", -- t[15430] = 1
      "0000001" when "00011110001000111", -- t[15431] = 1
      "0000001" when "00011110001001000", -- t[15432] = 1
      "0000001" when "00011110001001001", -- t[15433] = 1
      "0000001" when "00011110001001010", -- t[15434] = 1
      "0000001" when "00011110001001011", -- t[15435] = 1
      "0000001" when "00011110001001100", -- t[15436] = 1
      "0000001" when "00011110001001101", -- t[15437] = 1
      "0000001" when "00011110001001110", -- t[15438] = 1
      "0000001" when "00011110001001111", -- t[15439] = 1
      "0000001" when "00011110001010000", -- t[15440] = 1
      "0000001" when "00011110001010001", -- t[15441] = 1
      "0000001" when "00011110001010010", -- t[15442] = 1
      "0000001" when "00011110001010011", -- t[15443] = 1
      "0000001" when "00011110001010100", -- t[15444] = 1
      "0000001" when "00011110001010101", -- t[15445] = 1
      "0000001" when "00011110001010110", -- t[15446] = 1
      "0000001" when "00011110001010111", -- t[15447] = 1
      "0000001" when "00011110001011000", -- t[15448] = 1
      "0000001" when "00011110001011001", -- t[15449] = 1
      "0000001" when "00011110001011010", -- t[15450] = 1
      "0000001" when "00011110001011011", -- t[15451] = 1
      "0000001" when "00011110001011100", -- t[15452] = 1
      "0000001" when "00011110001011101", -- t[15453] = 1
      "0000001" when "00011110001011110", -- t[15454] = 1
      "0000001" when "00011110001011111", -- t[15455] = 1
      "0000001" when "00011110001100000", -- t[15456] = 1
      "0000001" when "00011110001100001", -- t[15457] = 1
      "0000001" when "00011110001100010", -- t[15458] = 1
      "0000001" when "00011110001100011", -- t[15459] = 1
      "0000001" when "00011110001100100", -- t[15460] = 1
      "0000001" when "00011110001100101", -- t[15461] = 1
      "0000001" when "00011110001100110", -- t[15462] = 1
      "0000001" when "00011110001100111", -- t[15463] = 1
      "0000001" when "00011110001101000", -- t[15464] = 1
      "0000001" when "00011110001101001", -- t[15465] = 1
      "0000001" when "00011110001101010", -- t[15466] = 1
      "0000001" when "00011110001101011", -- t[15467] = 1
      "0000001" when "00011110001101100", -- t[15468] = 1
      "0000001" when "00011110001101101", -- t[15469] = 1
      "0000001" when "00011110001101110", -- t[15470] = 1
      "0000001" when "00011110001101111", -- t[15471] = 1
      "0000001" when "00011110001110000", -- t[15472] = 1
      "0000001" when "00011110001110001", -- t[15473] = 1
      "0000001" when "00011110001110010", -- t[15474] = 1
      "0000001" when "00011110001110011", -- t[15475] = 1
      "0000001" when "00011110001110100", -- t[15476] = 1
      "0000001" when "00011110001110101", -- t[15477] = 1
      "0000001" when "00011110001110110", -- t[15478] = 1
      "0000001" when "00011110001110111", -- t[15479] = 1
      "0000001" when "00011110001111000", -- t[15480] = 1
      "0000001" when "00011110001111001", -- t[15481] = 1
      "0000001" when "00011110001111010", -- t[15482] = 1
      "0000001" when "00011110001111011", -- t[15483] = 1
      "0000001" when "00011110001111100", -- t[15484] = 1
      "0000001" when "00011110001111101", -- t[15485] = 1
      "0000001" when "00011110001111110", -- t[15486] = 1
      "0000001" when "00011110001111111", -- t[15487] = 1
      "0000001" when "00011110010000000", -- t[15488] = 1
      "0000001" when "00011110010000001", -- t[15489] = 1
      "0000001" when "00011110010000010", -- t[15490] = 1
      "0000001" when "00011110010000011", -- t[15491] = 1
      "0000001" when "00011110010000100", -- t[15492] = 1
      "0000001" when "00011110010000101", -- t[15493] = 1
      "0000001" when "00011110010000110", -- t[15494] = 1
      "0000001" when "00011110010000111", -- t[15495] = 1
      "0000001" when "00011110010001000", -- t[15496] = 1
      "0000001" when "00011110010001001", -- t[15497] = 1
      "0000001" when "00011110010001010", -- t[15498] = 1
      "0000001" when "00011110010001011", -- t[15499] = 1
      "0000001" when "00011110010001100", -- t[15500] = 1
      "0000001" when "00011110010001101", -- t[15501] = 1
      "0000001" when "00011110010001110", -- t[15502] = 1
      "0000001" when "00011110010001111", -- t[15503] = 1
      "0000001" when "00011110010010000", -- t[15504] = 1
      "0000001" when "00011110010010001", -- t[15505] = 1
      "0000001" when "00011110010010010", -- t[15506] = 1
      "0000001" when "00011110010010011", -- t[15507] = 1
      "0000001" when "00011110010010100", -- t[15508] = 1
      "0000001" when "00011110010010101", -- t[15509] = 1
      "0000001" when "00011110010010110", -- t[15510] = 1
      "0000001" when "00011110010010111", -- t[15511] = 1
      "0000001" when "00011110010011000", -- t[15512] = 1
      "0000001" when "00011110010011001", -- t[15513] = 1
      "0000001" when "00011110010011010", -- t[15514] = 1
      "0000001" when "00011110010011011", -- t[15515] = 1
      "0000001" when "00011110010011100", -- t[15516] = 1
      "0000001" when "00011110010011101", -- t[15517] = 1
      "0000001" when "00011110010011110", -- t[15518] = 1
      "0000001" when "00011110010011111", -- t[15519] = 1
      "0000001" when "00011110010100000", -- t[15520] = 1
      "0000001" when "00011110010100001", -- t[15521] = 1
      "0000001" when "00011110010100010", -- t[15522] = 1
      "0000001" when "00011110010100011", -- t[15523] = 1
      "0000001" when "00011110010100100", -- t[15524] = 1
      "0000001" when "00011110010100101", -- t[15525] = 1
      "0000001" when "00011110010100110", -- t[15526] = 1
      "0000001" when "00011110010100111", -- t[15527] = 1
      "0000001" when "00011110010101000", -- t[15528] = 1
      "0000001" when "00011110010101001", -- t[15529] = 1
      "0000001" when "00011110010101010", -- t[15530] = 1
      "0000001" when "00011110010101011", -- t[15531] = 1
      "0000001" when "00011110010101100", -- t[15532] = 1
      "0000001" when "00011110010101101", -- t[15533] = 1
      "0000001" when "00011110010101110", -- t[15534] = 1
      "0000001" when "00011110010101111", -- t[15535] = 1
      "0000001" when "00011110010110000", -- t[15536] = 1
      "0000001" when "00011110010110001", -- t[15537] = 1
      "0000001" when "00011110010110010", -- t[15538] = 1
      "0000001" when "00011110010110011", -- t[15539] = 1
      "0000001" when "00011110010110100", -- t[15540] = 1
      "0000001" when "00011110010110101", -- t[15541] = 1
      "0000001" when "00011110010110110", -- t[15542] = 1
      "0000001" when "00011110010110111", -- t[15543] = 1
      "0000001" when "00011110010111000", -- t[15544] = 1
      "0000001" when "00011110010111001", -- t[15545] = 1
      "0000001" when "00011110010111010", -- t[15546] = 1
      "0000001" when "00011110010111011", -- t[15547] = 1
      "0000001" when "00011110010111100", -- t[15548] = 1
      "0000001" when "00011110010111101", -- t[15549] = 1
      "0000001" when "00011110010111110", -- t[15550] = 1
      "0000001" when "00011110010111111", -- t[15551] = 1
      "0000001" when "00011110011000000", -- t[15552] = 1
      "0000001" when "00011110011000001", -- t[15553] = 1
      "0000001" when "00011110011000010", -- t[15554] = 1
      "0000001" when "00011110011000011", -- t[15555] = 1
      "0000001" when "00011110011000100", -- t[15556] = 1
      "0000001" when "00011110011000101", -- t[15557] = 1
      "0000001" when "00011110011000110", -- t[15558] = 1
      "0000001" when "00011110011000111", -- t[15559] = 1
      "0000001" when "00011110011001000", -- t[15560] = 1
      "0000001" when "00011110011001001", -- t[15561] = 1
      "0000001" when "00011110011001010", -- t[15562] = 1
      "0000001" when "00011110011001011", -- t[15563] = 1
      "0000001" when "00011110011001100", -- t[15564] = 1
      "0000001" when "00011110011001101", -- t[15565] = 1
      "0000001" when "00011110011001110", -- t[15566] = 1
      "0000001" when "00011110011001111", -- t[15567] = 1
      "0000001" when "00011110011010000", -- t[15568] = 1
      "0000001" when "00011110011010001", -- t[15569] = 1
      "0000001" when "00011110011010010", -- t[15570] = 1
      "0000001" when "00011110011010011", -- t[15571] = 1
      "0000001" when "00011110011010100", -- t[15572] = 1
      "0000001" when "00011110011010101", -- t[15573] = 1
      "0000001" when "00011110011010110", -- t[15574] = 1
      "0000001" when "00011110011010111", -- t[15575] = 1
      "0000001" when "00011110011011000", -- t[15576] = 1
      "0000001" when "00011110011011001", -- t[15577] = 1
      "0000001" when "00011110011011010", -- t[15578] = 1
      "0000001" when "00011110011011011", -- t[15579] = 1
      "0000001" when "00011110011011100", -- t[15580] = 1
      "0000001" when "00011110011011101", -- t[15581] = 1
      "0000001" when "00011110011011110", -- t[15582] = 1
      "0000001" when "00011110011011111", -- t[15583] = 1
      "0000001" when "00011110011100000", -- t[15584] = 1
      "0000001" when "00011110011100001", -- t[15585] = 1
      "0000001" when "00011110011100010", -- t[15586] = 1
      "0000001" when "00011110011100011", -- t[15587] = 1
      "0000001" when "00011110011100100", -- t[15588] = 1
      "0000001" when "00011110011100101", -- t[15589] = 1
      "0000001" when "00011110011100110", -- t[15590] = 1
      "0000001" when "00011110011100111", -- t[15591] = 1
      "0000001" when "00011110011101000", -- t[15592] = 1
      "0000001" when "00011110011101001", -- t[15593] = 1
      "0000001" when "00011110011101010", -- t[15594] = 1
      "0000001" when "00011110011101011", -- t[15595] = 1
      "0000001" when "00011110011101100", -- t[15596] = 1
      "0000001" when "00011110011101101", -- t[15597] = 1
      "0000001" when "00011110011101110", -- t[15598] = 1
      "0000001" when "00011110011101111", -- t[15599] = 1
      "0000001" when "00011110011110000", -- t[15600] = 1
      "0000001" when "00011110011110001", -- t[15601] = 1
      "0000001" when "00011110011110010", -- t[15602] = 1
      "0000001" when "00011110011110011", -- t[15603] = 1
      "0000001" when "00011110011110100", -- t[15604] = 1
      "0000001" when "00011110011110101", -- t[15605] = 1
      "0000001" when "00011110011110110", -- t[15606] = 1
      "0000001" when "00011110011110111", -- t[15607] = 1
      "0000001" when "00011110011111000", -- t[15608] = 1
      "0000001" when "00011110011111001", -- t[15609] = 1
      "0000001" when "00011110011111010", -- t[15610] = 1
      "0000001" when "00011110011111011", -- t[15611] = 1
      "0000001" when "00011110011111100", -- t[15612] = 1
      "0000001" when "00011110011111101", -- t[15613] = 1
      "0000001" when "00011110011111110", -- t[15614] = 1
      "0000001" when "00011110011111111", -- t[15615] = 1
      "0000001" when "00011110100000000", -- t[15616] = 1
      "0000001" when "00011110100000001", -- t[15617] = 1
      "0000001" when "00011110100000010", -- t[15618] = 1
      "0000001" when "00011110100000011", -- t[15619] = 1
      "0000001" when "00011110100000100", -- t[15620] = 1
      "0000001" when "00011110100000101", -- t[15621] = 1
      "0000001" when "00011110100000110", -- t[15622] = 1
      "0000001" when "00011110100000111", -- t[15623] = 1
      "0000001" when "00011110100001000", -- t[15624] = 1
      "0000001" when "00011110100001001", -- t[15625] = 1
      "0000001" when "00011110100001010", -- t[15626] = 1
      "0000001" when "00011110100001011", -- t[15627] = 1
      "0000001" when "00011110100001100", -- t[15628] = 1
      "0000001" when "00011110100001101", -- t[15629] = 1
      "0000001" when "00011110100001110", -- t[15630] = 1
      "0000001" when "00011110100001111", -- t[15631] = 1
      "0000001" when "00011110100010000", -- t[15632] = 1
      "0000001" when "00011110100010001", -- t[15633] = 1
      "0000001" when "00011110100010010", -- t[15634] = 1
      "0000001" when "00011110100010011", -- t[15635] = 1
      "0000001" when "00011110100010100", -- t[15636] = 1
      "0000001" when "00011110100010101", -- t[15637] = 1
      "0000001" when "00011110100010110", -- t[15638] = 1
      "0000001" when "00011110100010111", -- t[15639] = 1
      "0000001" when "00011110100011000", -- t[15640] = 1
      "0000001" when "00011110100011001", -- t[15641] = 1
      "0000001" when "00011110100011010", -- t[15642] = 1
      "0000001" when "00011110100011011", -- t[15643] = 1
      "0000001" when "00011110100011100", -- t[15644] = 1
      "0000001" when "00011110100011101", -- t[15645] = 1
      "0000001" when "00011110100011110", -- t[15646] = 1
      "0000001" when "00011110100011111", -- t[15647] = 1
      "0000001" when "00011110100100000", -- t[15648] = 1
      "0000001" when "00011110100100001", -- t[15649] = 1
      "0000001" when "00011110100100010", -- t[15650] = 1
      "0000001" when "00011110100100011", -- t[15651] = 1
      "0000001" when "00011110100100100", -- t[15652] = 1
      "0000001" when "00011110100100101", -- t[15653] = 1
      "0000001" when "00011110100100110", -- t[15654] = 1
      "0000001" when "00011110100100111", -- t[15655] = 1
      "0000001" when "00011110100101000", -- t[15656] = 1
      "0000001" when "00011110100101001", -- t[15657] = 1
      "0000001" when "00011110100101010", -- t[15658] = 1
      "0000001" when "00011110100101011", -- t[15659] = 1
      "0000001" when "00011110100101100", -- t[15660] = 1
      "0000001" when "00011110100101101", -- t[15661] = 1
      "0000001" when "00011110100101110", -- t[15662] = 1
      "0000001" when "00011110100101111", -- t[15663] = 1
      "0000001" when "00011110100110000", -- t[15664] = 1
      "0000001" when "00011110100110001", -- t[15665] = 1
      "0000001" when "00011110100110010", -- t[15666] = 1
      "0000001" when "00011110100110011", -- t[15667] = 1
      "0000001" when "00011110100110100", -- t[15668] = 1
      "0000001" when "00011110100110101", -- t[15669] = 1
      "0000001" when "00011110100110110", -- t[15670] = 1
      "0000001" when "00011110100110111", -- t[15671] = 1
      "0000001" when "00011110100111000", -- t[15672] = 1
      "0000001" when "00011110100111001", -- t[15673] = 1
      "0000001" when "00011110100111010", -- t[15674] = 1
      "0000001" when "00011110100111011", -- t[15675] = 1
      "0000001" when "00011110100111100", -- t[15676] = 1
      "0000001" when "00011110100111101", -- t[15677] = 1
      "0000001" when "00011110100111110", -- t[15678] = 1
      "0000001" when "00011110100111111", -- t[15679] = 1
      "0000001" when "00011110101000000", -- t[15680] = 1
      "0000001" when "00011110101000001", -- t[15681] = 1
      "0000001" when "00011110101000010", -- t[15682] = 1
      "0000001" when "00011110101000011", -- t[15683] = 1
      "0000001" when "00011110101000100", -- t[15684] = 1
      "0000001" when "00011110101000101", -- t[15685] = 1
      "0000001" when "00011110101000110", -- t[15686] = 1
      "0000001" when "00011110101000111", -- t[15687] = 1
      "0000001" when "00011110101001000", -- t[15688] = 1
      "0000001" when "00011110101001001", -- t[15689] = 1
      "0000001" when "00011110101001010", -- t[15690] = 1
      "0000001" when "00011110101001011", -- t[15691] = 1
      "0000001" when "00011110101001100", -- t[15692] = 1
      "0000001" when "00011110101001101", -- t[15693] = 1
      "0000001" when "00011110101001110", -- t[15694] = 1
      "0000001" when "00011110101001111", -- t[15695] = 1
      "0000001" when "00011110101010000", -- t[15696] = 1
      "0000001" when "00011110101010001", -- t[15697] = 1
      "0000001" when "00011110101010010", -- t[15698] = 1
      "0000001" when "00011110101010011", -- t[15699] = 1
      "0000001" when "00011110101010100", -- t[15700] = 1
      "0000001" when "00011110101010101", -- t[15701] = 1
      "0000001" when "00011110101010110", -- t[15702] = 1
      "0000001" when "00011110101010111", -- t[15703] = 1
      "0000001" when "00011110101011000", -- t[15704] = 1
      "0000001" when "00011110101011001", -- t[15705] = 1
      "0000001" when "00011110101011010", -- t[15706] = 1
      "0000001" when "00011110101011011", -- t[15707] = 1
      "0000001" when "00011110101011100", -- t[15708] = 1
      "0000001" when "00011110101011101", -- t[15709] = 1
      "0000001" when "00011110101011110", -- t[15710] = 1
      "0000001" when "00011110101011111", -- t[15711] = 1
      "0000001" when "00011110101100000", -- t[15712] = 1
      "0000001" when "00011110101100001", -- t[15713] = 1
      "0000001" when "00011110101100010", -- t[15714] = 1
      "0000001" when "00011110101100011", -- t[15715] = 1
      "0000001" when "00011110101100100", -- t[15716] = 1
      "0000001" when "00011110101100101", -- t[15717] = 1
      "0000001" when "00011110101100110", -- t[15718] = 1
      "0000001" when "00011110101100111", -- t[15719] = 1
      "0000001" when "00011110101101000", -- t[15720] = 1
      "0000001" when "00011110101101001", -- t[15721] = 1
      "0000001" when "00011110101101010", -- t[15722] = 1
      "0000001" when "00011110101101011", -- t[15723] = 1
      "0000001" when "00011110101101100", -- t[15724] = 1
      "0000001" when "00011110101101101", -- t[15725] = 1
      "0000001" when "00011110101101110", -- t[15726] = 1
      "0000001" when "00011110101101111", -- t[15727] = 1
      "0000001" when "00011110101110000", -- t[15728] = 1
      "0000001" when "00011110101110001", -- t[15729] = 1
      "0000001" when "00011110101110010", -- t[15730] = 1
      "0000001" when "00011110101110011", -- t[15731] = 1
      "0000001" when "00011110101110100", -- t[15732] = 1
      "0000001" when "00011110101110101", -- t[15733] = 1
      "0000001" when "00011110101110110", -- t[15734] = 1
      "0000001" when "00011110101110111", -- t[15735] = 1
      "0000001" when "00011110101111000", -- t[15736] = 1
      "0000001" when "00011110101111001", -- t[15737] = 1
      "0000001" when "00011110101111010", -- t[15738] = 1
      "0000001" when "00011110101111011", -- t[15739] = 1
      "0000001" when "00011110101111100", -- t[15740] = 1
      "0000001" when "00011110101111101", -- t[15741] = 1
      "0000001" when "00011110101111110", -- t[15742] = 1
      "0000001" when "00011110101111111", -- t[15743] = 1
      "0000001" when "00011110110000000", -- t[15744] = 1
      "0000001" when "00011110110000001", -- t[15745] = 1
      "0000001" when "00011110110000010", -- t[15746] = 1
      "0000001" when "00011110110000011", -- t[15747] = 1
      "0000001" when "00011110110000100", -- t[15748] = 1
      "0000001" when "00011110110000101", -- t[15749] = 1
      "0000001" when "00011110110000110", -- t[15750] = 1
      "0000001" when "00011110110000111", -- t[15751] = 1
      "0000001" when "00011110110001000", -- t[15752] = 1
      "0000001" when "00011110110001001", -- t[15753] = 1
      "0000001" when "00011110110001010", -- t[15754] = 1
      "0000001" when "00011110110001011", -- t[15755] = 1
      "0000001" when "00011110110001100", -- t[15756] = 1
      "0000001" when "00011110110001101", -- t[15757] = 1
      "0000001" when "00011110110001110", -- t[15758] = 1
      "0000001" when "00011110110001111", -- t[15759] = 1
      "0000001" when "00011110110010000", -- t[15760] = 1
      "0000001" when "00011110110010001", -- t[15761] = 1
      "0000001" when "00011110110010010", -- t[15762] = 1
      "0000001" when "00011110110010011", -- t[15763] = 1
      "0000001" when "00011110110010100", -- t[15764] = 1
      "0000001" when "00011110110010101", -- t[15765] = 1
      "0000001" when "00011110110010110", -- t[15766] = 1
      "0000001" when "00011110110010111", -- t[15767] = 1
      "0000001" when "00011110110011000", -- t[15768] = 1
      "0000001" when "00011110110011001", -- t[15769] = 1
      "0000001" when "00011110110011010", -- t[15770] = 1
      "0000001" when "00011110110011011", -- t[15771] = 1
      "0000001" when "00011110110011100", -- t[15772] = 1
      "0000001" when "00011110110011101", -- t[15773] = 1
      "0000001" when "00011110110011110", -- t[15774] = 1
      "0000001" when "00011110110011111", -- t[15775] = 1
      "0000001" when "00011110110100000", -- t[15776] = 1
      "0000001" when "00011110110100001", -- t[15777] = 1
      "0000001" when "00011110110100010", -- t[15778] = 1
      "0000001" when "00011110110100011", -- t[15779] = 1
      "0000001" when "00011110110100100", -- t[15780] = 1
      "0000001" when "00011110110100101", -- t[15781] = 1
      "0000001" when "00011110110100110", -- t[15782] = 1
      "0000001" when "00011110110100111", -- t[15783] = 1
      "0000001" when "00011110110101000", -- t[15784] = 1
      "0000001" when "00011110110101001", -- t[15785] = 1
      "0000001" when "00011110110101010", -- t[15786] = 1
      "0000001" when "00011110110101011", -- t[15787] = 1
      "0000001" when "00011110110101100", -- t[15788] = 1
      "0000001" when "00011110110101101", -- t[15789] = 1
      "0000001" when "00011110110101110", -- t[15790] = 1
      "0000001" when "00011110110101111", -- t[15791] = 1
      "0000001" when "00011110110110000", -- t[15792] = 1
      "0000001" when "00011110110110001", -- t[15793] = 1
      "0000001" when "00011110110110010", -- t[15794] = 1
      "0000001" when "00011110110110011", -- t[15795] = 1
      "0000001" when "00011110110110100", -- t[15796] = 1
      "0000001" when "00011110110110101", -- t[15797] = 1
      "0000001" when "00011110110110110", -- t[15798] = 1
      "0000001" when "00011110110110111", -- t[15799] = 1
      "0000001" when "00011110110111000", -- t[15800] = 1
      "0000001" when "00011110110111001", -- t[15801] = 1
      "0000001" when "00011110110111010", -- t[15802] = 1
      "0000001" when "00011110110111011", -- t[15803] = 1
      "0000001" when "00011110110111100", -- t[15804] = 1
      "0000001" when "00011110110111101", -- t[15805] = 1
      "0000001" when "00011110110111110", -- t[15806] = 1
      "0000001" when "00011110110111111", -- t[15807] = 1
      "0000001" when "00011110111000000", -- t[15808] = 1
      "0000001" when "00011110111000001", -- t[15809] = 1
      "0000001" when "00011110111000010", -- t[15810] = 1
      "0000001" when "00011110111000011", -- t[15811] = 1
      "0000001" when "00011110111000100", -- t[15812] = 1
      "0000001" when "00011110111000101", -- t[15813] = 1
      "0000001" when "00011110111000110", -- t[15814] = 1
      "0000001" when "00011110111000111", -- t[15815] = 1
      "0000001" when "00011110111001000", -- t[15816] = 1
      "0000001" when "00011110111001001", -- t[15817] = 1
      "0000001" when "00011110111001010", -- t[15818] = 1
      "0000001" when "00011110111001011", -- t[15819] = 1
      "0000001" when "00011110111001100", -- t[15820] = 1
      "0000001" when "00011110111001101", -- t[15821] = 1
      "0000001" when "00011110111001110", -- t[15822] = 1
      "0000001" when "00011110111001111", -- t[15823] = 1
      "0000001" when "00011110111010000", -- t[15824] = 1
      "0000001" when "00011110111010001", -- t[15825] = 1
      "0000001" when "00011110111010010", -- t[15826] = 1
      "0000001" when "00011110111010011", -- t[15827] = 1
      "0000001" when "00011110111010100", -- t[15828] = 1
      "0000001" when "00011110111010101", -- t[15829] = 1
      "0000001" when "00011110111010110", -- t[15830] = 1
      "0000001" when "00011110111010111", -- t[15831] = 1
      "0000001" when "00011110111011000", -- t[15832] = 1
      "0000001" when "00011110111011001", -- t[15833] = 1
      "0000001" when "00011110111011010", -- t[15834] = 1
      "0000001" when "00011110111011011", -- t[15835] = 1
      "0000001" when "00011110111011100", -- t[15836] = 1
      "0000001" when "00011110111011101", -- t[15837] = 1
      "0000001" when "00011110111011110", -- t[15838] = 1
      "0000001" when "00011110111011111", -- t[15839] = 1
      "0000001" when "00011110111100000", -- t[15840] = 1
      "0000001" when "00011110111100001", -- t[15841] = 1
      "0000001" when "00011110111100010", -- t[15842] = 1
      "0000001" when "00011110111100011", -- t[15843] = 1
      "0000001" when "00011110111100100", -- t[15844] = 1
      "0000001" when "00011110111100101", -- t[15845] = 1
      "0000001" when "00011110111100110", -- t[15846] = 1
      "0000001" when "00011110111100111", -- t[15847] = 1
      "0000001" when "00011110111101000", -- t[15848] = 1
      "0000001" when "00011110111101001", -- t[15849] = 1
      "0000001" when "00011110111101010", -- t[15850] = 1
      "0000001" when "00011110111101011", -- t[15851] = 1
      "0000001" when "00011110111101100", -- t[15852] = 1
      "0000001" when "00011110111101101", -- t[15853] = 1
      "0000001" when "00011110111101110", -- t[15854] = 1
      "0000001" when "00011110111101111", -- t[15855] = 1
      "0000001" when "00011110111110000", -- t[15856] = 1
      "0000001" when "00011110111110001", -- t[15857] = 1
      "0000001" when "00011110111110010", -- t[15858] = 1
      "0000001" when "00011110111110011", -- t[15859] = 1
      "0000001" when "00011110111110100", -- t[15860] = 1
      "0000001" when "00011110111110101", -- t[15861] = 1
      "0000001" when "00011110111110110", -- t[15862] = 1
      "0000001" when "00011110111110111", -- t[15863] = 1
      "0000001" when "00011110111111000", -- t[15864] = 1
      "0000001" when "00011110111111001", -- t[15865] = 1
      "0000001" when "00011110111111010", -- t[15866] = 1
      "0000001" when "00011110111111011", -- t[15867] = 1
      "0000001" when "00011110111111100", -- t[15868] = 1
      "0000001" when "00011110111111101", -- t[15869] = 1
      "0000001" when "00011110111111110", -- t[15870] = 1
      "0000001" when "00011110111111111", -- t[15871] = 1
      "0000001" when "00011111000000000", -- t[15872] = 1
      "0000001" when "00011111000000001", -- t[15873] = 1
      "0000001" when "00011111000000010", -- t[15874] = 1
      "0000001" when "00011111000000011", -- t[15875] = 1
      "0000001" when "00011111000000100", -- t[15876] = 1
      "0000001" when "00011111000000101", -- t[15877] = 1
      "0000001" when "00011111000000110", -- t[15878] = 1
      "0000001" when "00011111000000111", -- t[15879] = 1
      "0000001" when "00011111000001000", -- t[15880] = 1
      "0000001" when "00011111000001001", -- t[15881] = 1
      "0000001" when "00011111000001010", -- t[15882] = 1
      "0000001" when "00011111000001011", -- t[15883] = 1
      "0000001" when "00011111000001100", -- t[15884] = 1
      "0000001" when "00011111000001101", -- t[15885] = 1
      "0000001" when "00011111000001110", -- t[15886] = 1
      "0000001" when "00011111000001111", -- t[15887] = 1
      "0000001" when "00011111000010000", -- t[15888] = 1
      "0000001" when "00011111000010001", -- t[15889] = 1
      "0000001" when "00011111000010010", -- t[15890] = 1
      "0000001" when "00011111000010011", -- t[15891] = 1
      "0000001" when "00011111000010100", -- t[15892] = 1
      "0000001" when "00011111000010101", -- t[15893] = 1
      "0000001" when "00011111000010110", -- t[15894] = 1
      "0000001" when "00011111000010111", -- t[15895] = 1
      "0000001" when "00011111000011000", -- t[15896] = 1
      "0000001" when "00011111000011001", -- t[15897] = 1
      "0000001" when "00011111000011010", -- t[15898] = 1
      "0000001" when "00011111000011011", -- t[15899] = 1
      "0000001" when "00011111000011100", -- t[15900] = 1
      "0000001" when "00011111000011101", -- t[15901] = 1
      "0000001" when "00011111000011110", -- t[15902] = 1
      "0000001" when "00011111000011111", -- t[15903] = 1
      "0000001" when "00011111000100000", -- t[15904] = 1
      "0000001" when "00011111000100001", -- t[15905] = 1
      "0000001" when "00011111000100010", -- t[15906] = 1
      "0000001" when "00011111000100011", -- t[15907] = 1
      "0000001" when "00011111000100100", -- t[15908] = 1
      "0000001" when "00011111000100101", -- t[15909] = 1
      "0000001" when "00011111000100110", -- t[15910] = 1
      "0000001" when "00011111000100111", -- t[15911] = 1
      "0000001" when "00011111000101000", -- t[15912] = 1
      "0000001" when "00011111000101001", -- t[15913] = 1
      "0000001" when "00011111000101010", -- t[15914] = 1
      "0000001" when "00011111000101011", -- t[15915] = 1
      "0000001" when "00011111000101100", -- t[15916] = 1
      "0000001" when "00011111000101101", -- t[15917] = 1
      "0000001" when "00011111000101110", -- t[15918] = 1
      "0000001" when "00011111000101111", -- t[15919] = 1
      "0000001" when "00011111000110000", -- t[15920] = 1
      "0000001" when "00011111000110001", -- t[15921] = 1
      "0000001" when "00011111000110010", -- t[15922] = 1
      "0000001" when "00011111000110011", -- t[15923] = 1
      "0000001" when "00011111000110100", -- t[15924] = 1
      "0000001" when "00011111000110101", -- t[15925] = 1
      "0000001" when "00011111000110110", -- t[15926] = 1
      "0000001" when "00011111000110111", -- t[15927] = 1
      "0000001" when "00011111000111000", -- t[15928] = 1
      "0000001" when "00011111000111001", -- t[15929] = 1
      "0000001" when "00011111000111010", -- t[15930] = 1
      "0000001" when "00011111000111011", -- t[15931] = 1
      "0000001" when "00011111000111100", -- t[15932] = 1
      "0000001" when "00011111000111101", -- t[15933] = 1
      "0000001" when "00011111000111110", -- t[15934] = 1
      "0000001" when "00011111000111111", -- t[15935] = 1
      "0000001" when "00011111001000000", -- t[15936] = 1
      "0000001" when "00011111001000001", -- t[15937] = 1
      "0000001" when "00011111001000010", -- t[15938] = 1
      "0000001" when "00011111001000011", -- t[15939] = 1
      "0000001" when "00011111001000100", -- t[15940] = 1
      "0000001" when "00011111001000101", -- t[15941] = 1
      "0000001" when "00011111001000110", -- t[15942] = 1
      "0000001" when "00011111001000111", -- t[15943] = 1
      "0000001" when "00011111001001000", -- t[15944] = 1
      "0000001" when "00011111001001001", -- t[15945] = 1
      "0000001" when "00011111001001010", -- t[15946] = 1
      "0000001" when "00011111001001011", -- t[15947] = 1
      "0000001" when "00011111001001100", -- t[15948] = 1
      "0000001" when "00011111001001101", -- t[15949] = 1
      "0000001" when "00011111001001110", -- t[15950] = 1
      "0000001" when "00011111001001111", -- t[15951] = 1
      "0000001" when "00011111001010000", -- t[15952] = 1
      "0000001" when "00011111001010001", -- t[15953] = 1
      "0000001" when "00011111001010010", -- t[15954] = 1
      "0000001" when "00011111001010011", -- t[15955] = 1
      "0000001" when "00011111001010100", -- t[15956] = 1
      "0000001" when "00011111001010101", -- t[15957] = 1
      "0000001" when "00011111001010110", -- t[15958] = 1
      "0000001" when "00011111001010111", -- t[15959] = 1
      "0000001" when "00011111001011000", -- t[15960] = 1
      "0000001" when "00011111001011001", -- t[15961] = 1
      "0000001" when "00011111001011010", -- t[15962] = 1
      "0000001" when "00011111001011011", -- t[15963] = 1
      "0000001" when "00011111001011100", -- t[15964] = 1
      "0000001" when "00011111001011101", -- t[15965] = 1
      "0000001" when "00011111001011110", -- t[15966] = 1
      "0000001" when "00011111001011111", -- t[15967] = 1
      "0000001" when "00011111001100000", -- t[15968] = 1
      "0000001" when "00011111001100001", -- t[15969] = 1
      "0000001" when "00011111001100010", -- t[15970] = 1
      "0000001" when "00011111001100011", -- t[15971] = 1
      "0000001" when "00011111001100100", -- t[15972] = 1
      "0000001" when "00011111001100101", -- t[15973] = 1
      "0000001" when "00011111001100110", -- t[15974] = 1
      "0000001" when "00011111001100111", -- t[15975] = 1
      "0000001" when "00011111001101000", -- t[15976] = 1
      "0000001" when "00011111001101001", -- t[15977] = 1
      "0000001" when "00011111001101010", -- t[15978] = 1
      "0000001" when "00011111001101011", -- t[15979] = 1
      "0000001" when "00011111001101100", -- t[15980] = 1
      "0000001" when "00011111001101101", -- t[15981] = 1
      "0000001" when "00011111001101110", -- t[15982] = 1
      "0000001" when "00011111001101111", -- t[15983] = 1
      "0000001" when "00011111001110000", -- t[15984] = 1
      "0000001" when "00011111001110001", -- t[15985] = 1
      "0000001" when "00011111001110010", -- t[15986] = 1
      "0000001" when "00011111001110011", -- t[15987] = 1
      "0000001" when "00011111001110100", -- t[15988] = 1
      "0000001" when "00011111001110101", -- t[15989] = 1
      "0000001" when "00011111001110110", -- t[15990] = 1
      "0000001" when "00011111001110111", -- t[15991] = 1
      "0000001" when "00011111001111000", -- t[15992] = 1
      "0000001" when "00011111001111001", -- t[15993] = 1
      "0000001" when "00011111001111010", -- t[15994] = 1
      "0000001" when "00011111001111011", -- t[15995] = 1
      "0000001" when "00011111001111100", -- t[15996] = 1
      "0000001" when "00011111001111101", -- t[15997] = 1
      "0000001" when "00011111001111110", -- t[15998] = 1
      "0000001" when "00011111001111111", -- t[15999] = 1
      "0000001" when "00011111010000000", -- t[16000] = 1
      "0000001" when "00011111010000001", -- t[16001] = 1
      "0000001" when "00011111010000010", -- t[16002] = 1
      "0000001" when "00011111010000011", -- t[16003] = 1
      "0000001" when "00011111010000100", -- t[16004] = 1
      "0000001" when "00011111010000101", -- t[16005] = 1
      "0000001" when "00011111010000110", -- t[16006] = 1
      "0000001" when "00011111010000111", -- t[16007] = 1
      "0000001" when "00011111010001000", -- t[16008] = 1
      "0000001" when "00011111010001001", -- t[16009] = 1
      "0000001" when "00011111010001010", -- t[16010] = 1
      "0000001" when "00011111010001011", -- t[16011] = 1
      "0000001" when "00011111010001100", -- t[16012] = 1
      "0000001" when "00011111010001101", -- t[16013] = 1
      "0000001" when "00011111010001110", -- t[16014] = 1
      "0000001" when "00011111010001111", -- t[16015] = 1
      "0000001" when "00011111010010000", -- t[16016] = 1
      "0000001" when "00011111010010001", -- t[16017] = 1
      "0000001" when "00011111010010010", -- t[16018] = 1
      "0000001" when "00011111010010011", -- t[16019] = 1
      "0000001" when "00011111010010100", -- t[16020] = 1
      "0000001" when "00011111010010101", -- t[16021] = 1
      "0000001" when "00011111010010110", -- t[16022] = 1
      "0000001" when "00011111010010111", -- t[16023] = 1
      "0000001" when "00011111010011000", -- t[16024] = 1
      "0000001" when "00011111010011001", -- t[16025] = 1
      "0000001" when "00011111010011010", -- t[16026] = 1
      "0000001" when "00011111010011011", -- t[16027] = 1
      "0000001" when "00011111010011100", -- t[16028] = 1
      "0000001" when "00011111010011101", -- t[16029] = 1
      "0000001" when "00011111010011110", -- t[16030] = 1
      "0000001" when "00011111010011111", -- t[16031] = 1
      "0000001" when "00011111010100000", -- t[16032] = 1
      "0000001" when "00011111010100001", -- t[16033] = 1
      "0000001" when "00011111010100010", -- t[16034] = 1
      "0000001" when "00011111010100011", -- t[16035] = 1
      "0000001" when "00011111010100100", -- t[16036] = 1
      "0000001" when "00011111010100101", -- t[16037] = 1
      "0000001" when "00011111010100110", -- t[16038] = 1
      "0000001" when "00011111010100111", -- t[16039] = 1
      "0000001" when "00011111010101000", -- t[16040] = 1
      "0000001" when "00011111010101001", -- t[16041] = 1
      "0000001" when "00011111010101010", -- t[16042] = 1
      "0000001" when "00011111010101011", -- t[16043] = 1
      "0000001" when "00011111010101100", -- t[16044] = 1
      "0000001" when "00011111010101101", -- t[16045] = 1
      "0000001" when "00011111010101110", -- t[16046] = 1
      "0000001" when "00011111010101111", -- t[16047] = 1
      "0000001" when "00011111010110000", -- t[16048] = 1
      "0000001" when "00011111010110001", -- t[16049] = 1
      "0000001" when "00011111010110010", -- t[16050] = 1
      "0000001" when "00011111010110011", -- t[16051] = 1
      "0000001" when "00011111010110100", -- t[16052] = 1
      "0000001" when "00011111010110101", -- t[16053] = 1
      "0000001" when "00011111010110110", -- t[16054] = 1
      "0000001" when "00011111010110111", -- t[16055] = 1
      "0000001" when "00011111010111000", -- t[16056] = 1
      "0000001" when "00011111010111001", -- t[16057] = 1
      "0000001" when "00011111010111010", -- t[16058] = 1
      "0000001" when "00011111010111011", -- t[16059] = 1
      "0000001" when "00011111010111100", -- t[16060] = 1
      "0000001" when "00011111010111101", -- t[16061] = 1
      "0000001" when "00011111010111110", -- t[16062] = 1
      "0000001" when "00011111010111111", -- t[16063] = 1
      "0000001" when "00011111011000000", -- t[16064] = 1
      "0000001" when "00011111011000001", -- t[16065] = 1
      "0000001" when "00011111011000010", -- t[16066] = 1
      "0000001" when "00011111011000011", -- t[16067] = 1
      "0000001" when "00011111011000100", -- t[16068] = 1
      "0000001" when "00011111011000101", -- t[16069] = 1
      "0000001" when "00011111011000110", -- t[16070] = 1
      "0000001" when "00011111011000111", -- t[16071] = 1
      "0000001" when "00011111011001000", -- t[16072] = 1
      "0000001" when "00011111011001001", -- t[16073] = 1
      "0000001" when "00011111011001010", -- t[16074] = 1
      "0000001" when "00011111011001011", -- t[16075] = 1
      "0000001" when "00011111011001100", -- t[16076] = 1
      "0000001" when "00011111011001101", -- t[16077] = 1
      "0000001" when "00011111011001110", -- t[16078] = 1
      "0000001" when "00011111011001111", -- t[16079] = 1
      "0000001" when "00011111011010000", -- t[16080] = 1
      "0000001" when "00011111011010001", -- t[16081] = 1
      "0000001" when "00011111011010010", -- t[16082] = 1
      "0000001" when "00011111011010011", -- t[16083] = 1
      "0000001" when "00011111011010100", -- t[16084] = 1
      "0000001" when "00011111011010101", -- t[16085] = 1
      "0000001" when "00011111011010110", -- t[16086] = 1
      "0000001" when "00011111011010111", -- t[16087] = 1
      "0000001" when "00011111011011000", -- t[16088] = 1
      "0000001" when "00011111011011001", -- t[16089] = 1
      "0000001" when "00011111011011010", -- t[16090] = 1
      "0000001" when "00011111011011011", -- t[16091] = 1
      "0000001" when "00011111011011100", -- t[16092] = 1
      "0000001" when "00011111011011101", -- t[16093] = 1
      "0000001" when "00011111011011110", -- t[16094] = 1
      "0000001" when "00011111011011111", -- t[16095] = 1
      "0000001" when "00011111011100000", -- t[16096] = 1
      "0000001" when "00011111011100001", -- t[16097] = 1
      "0000001" when "00011111011100010", -- t[16098] = 1
      "0000001" when "00011111011100011", -- t[16099] = 1
      "0000001" when "00011111011100100", -- t[16100] = 1
      "0000001" when "00011111011100101", -- t[16101] = 1
      "0000001" when "00011111011100110", -- t[16102] = 1
      "0000001" when "00011111011100111", -- t[16103] = 1
      "0000001" when "00011111011101000", -- t[16104] = 1
      "0000001" when "00011111011101001", -- t[16105] = 1
      "0000001" when "00011111011101010", -- t[16106] = 1
      "0000001" when "00011111011101011", -- t[16107] = 1
      "0000001" when "00011111011101100", -- t[16108] = 1
      "0000001" when "00011111011101101", -- t[16109] = 1
      "0000001" when "00011111011101110", -- t[16110] = 1
      "0000001" when "00011111011101111", -- t[16111] = 1
      "0000001" when "00011111011110000", -- t[16112] = 1
      "0000001" when "00011111011110001", -- t[16113] = 1
      "0000001" when "00011111011110010", -- t[16114] = 1
      "0000001" when "00011111011110011", -- t[16115] = 1
      "0000001" when "00011111011110100", -- t[16116] = 1
      "0000001" when "00011111011110101", -- t[16117] = 1
      "0000001" when "00011111011110110", -- t[16118] = 1
      "0000001" when "00011111011110111", -- t[16119] = 1
      "0000001" when "00011111011111000", -- t[16120] = 1
      "0000001" when "00011111011111001", -- t[16121] = 1
      "0000001" when "00011111011111010", -- t[16122] = 1
      "0000001" when "00011111011111011", -- t[16123] = 1
      "0000001" when "00011111011111100", -- t[16124] = 1
      "0000001" when "00011111011111101", -- t[16125] = 1
      "0000001" when "00011111011111110", -- t[16126] = 1
      "0000001" when "00011111011111111", -- t[16127] = 1
      "0000001" when "00011111100000000", -- t[16128] = 1
      "0000001" when "00011111100000001", -- t[16129] = 1
      "0000001" when "00011111100000010", -- t[16130] = 1
      "0000001" when "00011111100000011", -- t[16131] = 1
      "0000001" when "00011111100000100", -- t[16132] = 1
      "0000001" when "00011111100000101", -- t[16133] = 1
      "0000001" when "00011111100000110", -- t[16134] = 1
      "0000001" when "00011111100000111", -- t[16135] = 1
      "0000001" when "00011111100001000", -- t[16136] = 1
      "0000001" when "00011111100001001", -- t[16137] = 1
      "0000001" when "00011111100001010", -- t[16138] = 1
      "0000001" when "00011111100001011", -- t[16139] = 1
      "0000001" when "00011111100001100", -- t[16140] = 1
      "0000001" when "00011111100001101", -- t[16141] = 1
      "0000001" when "00011111100001110", -- t[16142] = 1
      "0000001" when "00011111100001111", -- t[16143] = 1
      "0000001" when "00011111100010000", -- t[16144] = 1
      "0000001" when "00011111100010001", -- t[16145] = 1
      "0000001" when "00011111100010010", -- t[16146] = 1
      "0000001" when "00011111100010011", -- t[16147] = 1
      "0000001" when "00011111100010100", -- t[16148] = 1
      "0000001" when "00011111100010101", -- t[16149] = 1
      "0000001" when "00011111100010110", -- t[16150] = 1
      "0000001" when "00011111100010111", -- t[16151] = 1
      "0000001" when "00011111100011000", -- t[16152] = 1
      "0000001" when "00011111100011001", -- t[16153] = 1
      "0000001" when "00011111100011010", -- t[16154] = 1
      "0000001" when "00011111100011011", -- t[16155] = 1
      "0000001" when "00011111100011100", -- t[16156] = 1
      "0000001" when "00011111100011101", -- t[16157] = 1
      "0000001" when "00011111100011110", -- t[16158] = 1
      "0000001" when "00011111100011111", -- t[16159] = 1
      "0000001" when "00011111100100000", -- t[16160] = 1
      "0000001" when "00011111100100001", -- t[16161] = 1
      "0000001" when "00011111100100010", -- t[16162] = 1
      "0000001" when "00011111100100011", -- t[16163] = 1
      "0000001" when "00011111100100100", -- t[16164] = 1
      "0000001" when "00011111100100101", -- t[16165] = 1
      "0000001" when "00011111100100110", -- t[16166] = 1
      "0000001" when "00011111100100111", -- t[16167] = 1
      "0000001" when "00011111100101000", -- t[16168] = 1
      "0000001" when "00011111100101001", -- t[16169] = 1
      "0000001" when "00011111100101010", -- t[16170] = 1
      "0000001" when "00011111100101011", -- t[16171] = 1
      "0000001" when "00011111100101100", -- t[16172] = 1
      "0000001" when "00011111100101101", -- t[16173] = 1
      "0000001" when "00011111100101110", -- t[16174] = 1
      "0000001" when "00011111100101111", -- t[16175] = 1
      "0000001" when "00011111100110000", -- t[16176] = 1
      "0000001" when "00011111100110001", -- t[16177] = 1
      "0000001" when "00011111100110010", -- t[16178] = 1
      "0000001" when "00011111100110011", -- t[16179] = 1
      "0000001" when "00011111100110100", -- t[16180] = 1
      "0000001" when "00011111100110101", -- t[16181] = 1
      "0000001" when "00011111100110110", -- t[16182] = 1
      "0000001" when "00011111100110111", -- t[16183] = 1
      "0000001" when "00011111100111000", -- t[16184] = 1
      "0000001" when "00011111100111001", -- t[16185] = 1
      "0000001" when "00011111100111010", -- t[16186] = 1
      "0000001" when "00011111100111011", -- t[16187] = 1
      "0000001" when "00011111100111100", -- t[16188] = 1
      "0000001" when "00011111100111101", -- t[16189] = 1
      "0000001" when "00011111100111110", -- t[16190] = 1
      "0000001" when "00011111100111111", -- t[16191] = 1
      "0000001" when "00011111101000000", -- t[16192] = 1
      "0000001" when "00011111101000001", -- t[16193] = 1
      "0000001" when "00011111101000010", -- t[16194] = 1
      "0000001" when "00011111101000011", -- t[16195] = 1
      "0000001" when "00011111101000100", -- t[16196] = 1
      "0000001" when "00011111101000101", -- t[16197] = 1
      "0000001" when "00011111101000110", -- t[16198] = 1
      "0000001" when "00011111101000111", -- t[16199] = 1
      "0000001" when "00011111101001000", -- t[16200] = 1
      "0000001" when "00011111101001001", -- t[16201] = 1
      "0000001" when "00011111101001010", -- t[16202] = 1
      "0000001" when "00011111101001011", -- t[16203] = 1
      "0000001" when "00011111101001100", -- t[16204] = 1
      "0000001" when "00011111101001101", -- t[16205] = 1
      "0000001" when "00011111101001110", -- t[16206] = 1
      "0000001" when "00011111101001111", -- t[16207] = 1
      "0000001" when "00011111101010000", -- t[16208] = 1
      "0000001" when "00011111101010001", -- t[16209] = 1
      "0000001" when "00011111101010010", -- t[16210] = 1
      "0000001" when "00011111101010011", -- t[16211] = 1
      "0000001" when "00011111101010100", -- t[16212] = 1
      "0000001" when "00011111101010101", -- t[16213] = 1
      "0000001" when "00011111101010110", -- t[16214] = 1
      "0000001" when "00011111101010111", -- t[16215] = 1
      "0000001" when "00011111101011000", -- t[16216] = 1
      "0000001" when "00011111101011001", -- t[16217] = 1
      "0000001" when "00011111101011010", -- t[16218] = 1
      "0000001" when "00011111101011011", -- t[16219] = 1
      "0000001" when "00011111101011100", -- t[16220] = 1
      "0000001" when "00011111101011101", -- t[16221] = 1
      "0000001" when "00011111101011110", -- t[16222] = 1
      "0000001" when "00011111101011111", -- t[16223] = 1
      "0000001" when "00011111101100000", -- t[16224] = 1
      "0000001" when "00011111101100001", -- t[16225] = 1
      "0000001" when "00011111101100010", -- t[16226] = 1
      "0000001" when "00011111101100011", -- t[16227] = 1
      "0000001" when "00011111101100100", -- t[16228] = 1
      "0000001" when "00011111101100101", -- t[16229] = 1
      "0000001" when "00011111101100110", -- t[16230] = 1
      "0000001" when "00011111101100111", -- t[16231] = 1
      "0000001" when "00011111101101000", -- t[16232] = 1
      "0000001" when "00011111101101001", -- t[16233] = 1
      "0000001" when "00011111101101010", -- t[16234] = 1
      "0000001" when "00011111101101011", -- t[16235] = 1
      "0000001" when "00011111101101100", -- t[16236] = 1
      "0000001" when "00011111101101101", -- t[16237] = 1
      "0000001" when "00011111101101110", -- t[16238] = 1
      "0000001" when "00011111101101111", -- t[16239] = 1
      "0000001" when "00011111101110000", -- t[16240] = 1
      "0000001" when "00011111101110001", -- t[16241] = 1
      "0000001" when "00011111101110010", -- t[16242] = 1
      "0000001" when "00011111101110011", -- t[16243] = 1
      "0000001" when "00011111101110100", -- t[16244] = 1
      "0000001" when "00011111101110101", -- t[16245] = 1
      "0000001" when "00011111101110110", -- t[16246] = 1
      "0000001" when "00011111101110111", -- t[16247] = 1
      "0000001" when "00011111101111000", -- t[16248] = 1
      "0000001" when "00011111101111001", -- t[16249] = 1
      "0000001" when "00011111101111010", -- t[16250] = 1
      "0000001" when "00011111101111011", -- t[16251] = 1
      "0000001" when "00011111101111100", -- t[16252] = 1
      "0000001" when "00011111101111101", -- t[16253] = 1
      "0000001" when "00011111101111110", -- t[16254] = 1
      "0000001" when "00011111101111111", -- t[16255] = 1
      "0000001" when "00011111110000000", -- t[16256] = 1
      "0000001" when "00011111110000001", -- t[16257] = 1
      "0000001" when "00011111110000010", -- t[16258] = 1
      "0000001" when "00011111110000011", -- t[16259] = 1
      "0000001" when "00011111110000100", -- t[16260] = 1
      "0000001" when "00011111110000101", -- t[16261] = 1
      "0000001" when "00011111110000110", -- t[16262] = 1
      "0000001" when "00011111110000111", -- t[16263] = 1
      "0000001" when "00011111110001000", -- t[16264] = 1
      "0000001" when "00011111110001001", -- t[16265] = 1
      "0000001" when "00011111110001010", -- t[16266] = 1
      "0000001" when "00011111110001011", -- t[16267] = 1
      "0000001" when "00011111110001100", -- t[16268] = 1
      "0000001" when "00011111110001101", -- t[16269] = 1
      "0000001" when "00011111110001110", -- t[16270] = 1
      "0000001" when "00011111110001111", -- t[16271] = 1
      "0000001" when "00011111110010000", -- t[16272] = 1
      "0000001" when "00011111110010001", -- t[16273] = 1
      "0000001" when "00011111110010010", -- t[16274] = 1
      "0000001" when "00011111110010011", -- t[16275] = 1
      "0000001" when "00011111110010100", -- t[16276] = 1
      "0000001" when "00011111110010101", -- t[16277] = 1
      "0000001" when "00011111110010110", -- t[16278] = 1
      "0000001" when "00011111110010111", -- t[16279] = 1
      "0000001" when "00011111110011000", -- t[16280] = 1
      "0000001" when "00011111110011001", -- t[16281] = 1
      "0000001" when "00011111110011010", -- t[16282] = 1
      "0000001" when "00011111110011011", -- t[16283] = 1
      "0000001" when "00011111110011100", -- t[16284] = 1
      "0000001" when "00011111110011101", -- t[16285] = 1
      "0000001" when "00011111110011110", -- t[16286] = 1
      "0000001" when "00011111110011111", -- t[16287] = 1
      "0000001" when "00011111110100000", -- t[16288] = 1
      "0000001" when "00011111110100001", -- t[16289] = 1
      "0000001" when "00011111110100010", -- t[16290] = 1
      "0000001" when "00011111110100011", -- t[16291] = 1
      "0000001" when "00011111110100100", -- t[16292] = 1
      "0000001" when "00011111110100101", -- t[16293] = 1
      "0000001" when "00011111110100110", -- t[16294] = 1
      "0000001" when "00011111110100111", -- t[16295] = 1
      "0000001" when "00011111110101000", -- t[16296] = 1
      "0000001" when "00011111110101001", -- t[16297] = 1
      "0000001" when "00011111110101010", -- t[16298] = 1
      "0000001" when "00011111110101011", -- t[16299] = 1
      "0000001" when "00011111110101100", -- t[16300] = 1
      "0000001" when "00011111110101101", -- t[16301] = 1
      "0000001" when "00011111110101110", -- t[16302] = 1
      "0000001" when "00011111110101111", -- t[16303] = 1
      "0000001" when "00011111110110000", -- t[16304] = 1
      "0000001" when "00011111110110001", -- t[16305] = 1
      "0000001" when "00011111110110010", -- t[16306] = 1
      "0000001" when "00011111110110011", -- t[16307] = 1
      "0000001" when "00011111110110100", -- t[16308] = 1
      "0000001" when "00011111110110101", -- t[16309] = 1
      "0000001" when "00011111110110110", -- t[16310] = 1
      "0000001" when "00011111110110111", -- t[16311] = 1
      "0000001" when "00011111110111000", -- t[16312] = 1
      "0000001" when "00011111110111001", -- t[16313] = 1
      "0000001" when "00011111110111010", -- t[16314] = 1
      "0000001" when "00011111110111011", -- t[16315] = 1
      "0000001" when "00011111110111100", -- t[16316] = 1
      "0000001" when "00011111110111101", -- t[16317] = 1
      "0000001" when "00011111110111110", -- t[16318] = 1
      "0000001" when "00011111110111111", -- t[16319] = 1
      "0000001" when "00011111111000000", -- t[16320] = 1
      "0000001" when "00011111111000001", -- t[16321] = 1
      "0000001" when "00011111111000010", -- t[16322] = 1
      "0000001" when "00011111111000011", -- t[16323] = 1
      "0000001" when "00011111111000100", -- t[16324] = 1
      "0000001" when "00011111111000101", -- t[16325] = 1
      "0000001" when "00011111111000110", -- t[16326] = 1
      "0000001" when "00011111111000111", -- t[16327] = 1
      "0000001" when "00011111111001000", -- t[16328] = 1
      "0000001" when "00011111111001001", -- t[16329] = 1
      "0000001" when "00011111111001010", -- t[16330] = 1
      "0000001" when "00011111111001011", -- t[16331] = 1
      "0000001" when "00011111111001100", -- t[16332] = 1
      "0000001" when "00011111111001101", -- t[16333] = 1
      "0000001" when "00011111111001110", -- t[16334] = 1
      "0000001" when "00011111111001111", -- t[16335] = 1
      "0000001" when "00011111111010000", -- t[16336] = 1
      "0000001" when "00011111111010001", -- t[16337] = 1
      "0000001" when "00011111111010010", -- t[16338] = 1
      "0000001" when "00011111111010011", -- t[16339] = 1
      "0000001" when "00011111111010100", -- t[16340] = 1
      "0000001" when "00011111111010101", -- t[16341] = 1
      "0000001" when "00011111111010110", -- t[16342] = 1
      "0000001" when "00011111111010111", -- t[16343] = 1
      "0000001" when "00011111111011000", -- t[16344] = 1
      "0000001" when "00011111111011001", -- t[16345] = 1
      "0000001" when "00011111111011010", -- t[16346] = 1
      "0000001" when "00011111111011011", -- t[16347] = 1
      "0000001" when "00011111111011100", -- t[16348] = 1
      "0000001" when "00011111111011101", -- t[16349] = 1
      "0000001" when "00011111111011110", -- t[16350] = 1
      "0000001" when "00011111111011111", -- t[16351] = 1
      "0000001" when "00011111111100000", -- t[16352] = 1
      "0000001" when "00011111111100001", -- t[16353] = 1
      "0000001" when "00011111111100010", -- t[16354] = 1
      "0000001" when "00011111111100011", -- t[16355] = 1
      "0000001" when "00011111111100100", -- t[16356] = 1
      "0000001" when "00011111111100101", -- t[16357] = 1
      "0000001" when "00011111111100110", -- t[16358] = 1
      "0000001" when "00011111111100111", -- t[16359] = 1
      "0000001" when "00011111111101000", -- t[16360] = 1
      "0000001" when "00011111111101001", -- t[16361] = 1
      "0000001" when "00011111111101010", -- t[16362] = 1
      "0000001" when "00011111111101011", -- t[16363] = 1
      "0000001" when "00011111111101100", -- t[16364] = 1
      "0000001" when "00011111111101101", -- t[16365] = 1
      "0000001" when "00011111111101110", -- t[16366] = 1
      "0000001" when "00011111111101111", -- t[16367] = 1
      "0000001" when "00011111111110000", -- t[16368] = 1
      "0000001" when "00011111111110001", -- t[16369] = 1
      "0000001" when "00011111111110010", -- t[16370] = 1
      "0000001" when "00011111111110011", -- t[16371] = 1
      "0000001" when "00011111111110100", -- t[16372] = 1
      "0000001" when "00011111111110101", -- t[16373] = 1
      "0000001" when "00011111111110110", -- t[16374] = 1
      "0000001" when "00011111111110111", -- t[16375] = 1
      "0000001" when "00011111111111000", -- t[16376] = 1
      "0000001" when "00011111111111001", -- t[16377] = 1
      "0000001" when "00011111111111010", -- t[16378] = 1
      "0000001" when "00011111111111011", -- t[16379] = 1
      "0000001" when "00011111111111100", -- t[16380] = 1
      "0000001" when "00011111111111101", -- t[16381] = 1
      "0000001" when "00011111111111110", -- t[16382] = 1
      "0000001" when "00011111111111111", -- t[16383] = 1
      "0000001" when "00100000000000000", -- t[16384] = 1
      "0000001" when "00100000000000001", -- t[16385] = 1
      "0000001" when "00100000000000010", -- t[16386] = 1
      "0000001" when "00100000000000011", -- t[16387] = 1
      "0000001" when "00100000000000100", -- t[16388] = 1
      "0000001" when "00100000000000101", -- t[16389] = 1
      "0000001" when "00100000000000110", -- t[16390] = 1
      "0000001" when "00100000000000111", -- t[16391] = 1
      "0000001" when "00100000000001000", -- t[16392] = 1
      "0000001" when "00100000000001001", -- t[16393] = 1
      "0000001" when "00100000000001010", -- t[16394] = 1
      "0000001" when "00100000000001011", -- t[16395] = 1
      "0000001" when "00100000000001100", -- t[16396] = 1
      "0000001" when "00100000000001101", -- t[16397] = 1
      "0000001" when "00100000000001110", -- t[16398] = 1
      "0000001" when "00100000000001111", -- t[16399] = 1
      "0000001" when "00100000000010000", -- t[16400] = 1
      "0000001" when "00100000000010001", -- t[16401] = 1
      "0000001" when "00100000000010010", -- t[16402] = 1
      "0000001" when "00100000000010011", -- t[16403] = 1
      "0000001" when "00100000000010100", -- t[16404] = 1
      "0000001" when "00100000000010101", -- t[16405] = 1
      "0000001" when "00100000000010110", -- t[16406] = 1
      "0000001" when "00100000000010111", -- t[16407] = 1
      "0000001" when "00100000000011000", -- t[16408] = 1
      "0000001" when "00100000000011001", -- t[16409] = 1
      "0000001" when "00100000000011010", -- t[16410] = 1
      "0000001" when "00100000000011011", -- t[16411] = 1
      "0000001" when "00100000000011100", -- t[16412] = 1
      "0000001" when "00100000000011101", -- t[16413] = 1
      "0000001" when "00100000000011110", -- t[16414] = 1
      "0000001" when "00100000000011111", -- t[16415] = 1
      "0000001" when "00100000000100000", -- t[16416] = 1
      "0000001" when "00100000000100001", -- t[16417] = 1
      "0000001" when "00100000000100010", -- t[16418] = 1
      "0000001" when "00100000000100011", -- t[16419] = 1
      "0000001" when "00100000000100100", -- t[16420] = 1
      "0000001" when "00100000000100101", -- t[16421] = 1
      "0000001" when "00100000000100110", -- t[16422] = 1
      "0000001" when "00100000000100111", -- t[16423] = 1
      "0000001" when "00100000000101000", -- t[16424] = 1
      "0000001" when "00100000000101001", -- t[16425] = 1
      "0000001" when "00100000000101010", -- t[16426] = 1
      "0000001" when "00100000000101011", -- t[16427] = 1
      "0000001" when "00100000000101100", -- t[16428] = 1
      "0000001" when "00100000000101101", -- t[16429] = 1
      "0000001" when "00100000000101110", -- t[16430] = 1
      "0000001" when "00100000000101111", -- t[16431] = 1
      "0000001" when "00100000000110000", -- t[16432] = 1
      "0000001" when "00100000000110001", -- t[16433] = 1
      "0000001" when "00100000000110010", -- t[16434] = 1
      "0000001" when "00100000000110011", -- t[16435] = 1
      "0000001" when "00100000000110100", -- t[16436] = 1
      "0000001" when "00100000000110101", -- t[16437] = 1
      "0000001" when "00100000000110110", -- t[16438] = 1
      "0000001" when "00100000000110111", -- t[16439] = 1
      "0000001" when "00100000000111000", -- t[16440] = 1
      "0000001" when "00100000000111001", -- t[16441] = 1
      "0000001" when "00100000000111010", -- t[16442] = 1
      "0000001" when "00100000000111011", -- t[16443] = 1
      "0000001" when "00100000000111100", -- t[16444] = 1
      "0000001" when "00100000000111101", -- t[16445] = 1
      "0000001" when "00100000000111110", -- t[16446] = 1
      "0000001" when "00100000000111111", -- t[16447] = 1
      "0000001" when "00100000001000000", -- t[16448] = 1
      "0000001" when "00100000001000001", -- t[16449] = 1
      "0000001" when "00100000001000010", -- t[16450] = 1
      "0000001" when "00100000001000011", -- t[16451] = 1
      "0000001" when "00100000001000100", -- t[16452] = 1
      "0000001" when "00100000001000101", -- t[16453] = 1
      "0000001" when "00100000001000110", -- t[16454] = 1
      "0000001" when "00100000001000111", -- t[16455] = 1
      "0000001" when "00100000001001000", -- t[16456] = 1
      "0000001" when "00100000001001001", -- t[16457] = 1
      "0000001" when "00100000001001010", -- t[16458] = 1
      "0000001" when "00100000001001011", -- t[16459] = 1
      "0000001" when "00100000001001100", -- t[16460] = 1
      "0000001" when "00100000001001101", -- t[16461] = 1
      "0000001" when "00100000001001110", -- t[16462] = 1
      "0000001" when "00100000001001111", -- t[16463] = 1
      "0000001" when "00100000001010000", -- t[16464] = 1
      "0000001" when "00100000001010001", -- t[16465] = 1
      "0000001" when "00100000001010010", -- t[16466] = 1
      "0000001" when "00100000001010011", -- t[16467] = 1
      "0000001" when "00100000001010100", -- t[16468] = 1
      "0000001" when "00100000001010101", -- t[16469] = 1
      "0000001" when "00100000001010110", -- t[16470] = 1
      "0000001" when "00100000001010111", -- t[16471] = 1
      "0000001" when "00100000001011000", -- t[16472] = 1
      "0000001" when "00100000001011001", -- t[16473] = 1
      "0000001" when "00100000001011010", -- t[16474] = 1
      "0000001" when "00100000001011011", -- t[16475] = 1
      "0000001" when "00100000001011100", -- t[16476] = 1
      "0000001" when "00100000001011101", -- t[16477] = 1
      "0000001" when "00100000001011110", -- t[16478] = 1
      "0000001" when "00100000001011111", -- t[16479] = 1
      "0000001" when "00100000001100000", -- t[16480] = 1
      "0000001" when "00100000001100001", -- t[16481] = 1
      "0000001" when "00100000001100010", -- t[16482] = 1
      "0000001" when "00100000001100011", -- t[16483] = 1
      "0000001" when "00100000001100100", -- t[16484] = 1
      "0000001" when "00100000001100101", -- t[16485] = 1
      "0000001" when "00100000001100110", -- t[16486] = 1
      "0000001" when "00100000001100111", -- t[16487] = 1
      "0000001" when "00100000001101000", -- t[16488] = 1
      "0000001" when "00100000001101001", -- t[16489] = 1
      "0000001" when "00100000001101010", -- t[16490] = 1
      "0000001" when "00100000001101011", -- t[16491] = 1
      "0000001" when "00100000001101100", -- t[16492] = 1
      "0000001" when "00100000001101101", -- t[16493] = 1
      "0000001" when "00100000001101110", -- t[16494] = 1
      "0000001" when "00100000001101111", -- t[16495] = 1
      "0000001" when "00100000001110000", -- t[16496] = 1
      "0000001" when "00100000001110001", -- t[16497] = 1
      "0000001" when "00100000001110010", -- t[16498] = 1
      "0000001" when "00100000001110011", -- t[16499] = 1
      "0000001" when "00100000001110100", -- t[16500] = 1
      "0000001" when "00100000001110101", -- t[16501] = 1
      "0000001" when "00100000001110110", -- t[16502] = 1
      "0000001" when "00100000001110111", -- t[16503] = 1
      "0000001" when "00100000001111000", -- t[16504] = 1
      "0000001" when "00100000001111001", -- t[16505] = 1
      "0000001" when "00100000001111010", -- t[16506] = 1
      "0000001" when "00100000001111011", -- t[16507] = 1
      "0000001" when "00100000001111100", -- t[16508] = 1
      "0000001" when "00100000001111101", -- t[16509] = 1
      "0000001" when "00100000001111110", -- t[16510] = 1
      "0000001" when "00100000001111111", -- t[16511] = 1
      "0000001" when "00100000010000000", -- t[16512] = 1
      "0000001" when "00100000010000001", -- t[16513] = 1
      "0000001" when "00100000010000010", -- t[16514] = 1
      "0000001" when "00100000010000011", -- t[16515] = 1
      "0000001" when "00100000010000100", -- t[16516] = 1
      "0000001" when "00100000010000101", -- t[16517] = 1
      "0000001" when "00100000010000110", -- t[16518] = 1
      "0000001" when "00100000010000111", -- t[16519] = 1
      "0000001" when "00100000010001000", -- t[16520] = 1
      "0000001" when "00100000010001001", -- t[16521] = 1
      "0000001" when "00100000010001010", -- t[16522] = 1
      "0000001" when "00100000010001011", -- t[16523] = 1
      "0000001" when "00100000010001100", -- t[16524] = 1
      "0000001" when "00100000010001101", -- t[16525] = 1
      "0000001" when "00100000010001110", -- t[16526] = 1
      "0000001" when "00100000010001111", -- t[16527] = 1
      "0000001" when "00100000010010000", -- t[16528] = 1
      "0000001" when "00100000010010001", -- t[16529] = 1
      "0000001" when "00100000010010010", -- t[16530] = 1
      "0000001" when "00100000010010011", -- t[16531] = 1
      "0000001" when "00100000010010100", -- t[16532] = 1
      "0000001" when "00100000010010101", -- t[16533] = 1
      "0000001" when "00100000010010110", -- t[16534] = 1
      "0000001" when "00100000010010111", -- t[16535] = 1
      "0000001" when "00100000010011000", -- t[16536] = 1
      "0000001" when "00100000010011001", -- t[16537] = 1
      "0000001" when "00100000010011010", -- t[16538] = 1
      "0000001" when "00100000010011011", -- t[16539] = 1
      "0000001" when "00100000010011100", -- t[16540] = 1
      "0000001" when "00100000010011101", -- t[16541] = 1
      "0000001" when "00100000010011110", -- t[16542] = 1
      "0000001" when "00100000010011111", -- t[16543] = 1
      "0000001" when "00100000010100000", -- t[16544] = 1
      "0000001" when "00100000010100001", -- t[16545] = 1
      "0000001" when "00100000010100010", -- t[16546] = 1
      "0000001" when "00100000010100011", -- t[16547] = 1
      "0000001" when "00100000010100100", -- t[16548] = 1
      "0000001" when "00100000010100101", -- t[16549] = 1
      "0000001" when "00100000010100110", -- t[16550] = 1
      "0000001" when "00100000010100111", -- t[16551] = 1
      "0000001" when "00100000010101000", -- t[16552] = 1
      "0000001" when "00100000010101001", -- t[16553] = 1
      "0000001" when "00100000010101010", -- t[16554] = 1
      "0000001" when "00100000010101011", -- t[16555] = 1
      "0000001" when "00100000010101100", -- t[16556] = 1
      "0000001" when "00100000010101101", -- t[16557] = 1
      "0000001" when "00100000010101110", -- t[16558] = 1
      "0000001" when "00100000010101111", -- t[16559] = 1
      "0000001" when "00100000010110000", -- t[16560] = 1
      "0000001" when "00100000010110001", -- t[16561] = 1
      "0000001" when "00100000010110010", -- t[16562] = 1
      "0000001" when "00100000010110011", -- t[16563] = 1
      "0000001" when "00100000010110100", -- t[16564] = 1
      "0000001" when "00100000010110101", -- t[16565] = 1
      "0000001" when "00100000010110110", -- t[16566] = 1
      "0000001" when "00100000010110111", -- t[16567] = 1
      "0000001" when "00100000010111000", -- t[16568] = 1
      "0000001" when "00100000010111001", -- t[16569] = 1
      "0000001" when "00100000010111010", -- t[16570] = 1
      "0000001" when "00100000010111011", -- t[16571] = 1
      "0000001" when "00100000010111100", -- t[16572] = 1
      "0000001" when "00100000010111101", -- t[16573] = 1
      "0000001" when "00100000010111110", -- t[16574] = 1
      "0000001" when "00100000010111111", -- t[16575] = 1
      "0000001" when "00100000011000000", -- t[16576] = 1
      "0000001" when "00100000011000001", -- t[16577] = 1
      "0000001" when "00100000011000010", -- t[16578] = 1
      "0000001" when "00100000011000011", -- t[16579] = 1
      "0000001" when "00100000011000100", -- t[16580] = 1
      "0000001" when "00100000011000101", -- t[16581] = 1
      "0000001" when "00100000011000110", -- t[16582] = 1
      "0000001" when "00100000011000111", -- t[16583] = 1
      "0000001" when "00100000011001000", -- t[16584] = 1
      "0000001" when "00100000011001001", -- t[16585] = 1
      "0000001" when "00100000011001010", -- t[16586] = 1
      "0000001" when "00100000011001011", -- t[16587] = 1
      "0000001" when "00100000011001100", -- t[16588] = 1
      "0000001" when "00100000011001101", -- t[16589] = 1
      "0000001" when "00100000011001110", -- t[16590] = 1
      "0000001" when "00100000011001111", -- t[16591] = 1
      "0000001" when "00100000011010000", -- t[16592] = 1
      "0000001" when "00100000011010001", -- t[16593] = 1
      "0000001" when "00100000011010010", -- t[16594] = 1
      "0000001" when "00100000011010011", -- t[16595] = 1
      "0000001" when "00100000011010100", -- t[16596] = 1
      "0000001" when "00100000011010101", -- t[16597] = 1
      "0000001" when "00100000011010110", -- t[16598] = 1
      "0000001" when "00100000011010111", -- t[16599] = 1
      "0000001" when "00100000011011000", -- t[16600] = 1
      "0000001" when "00100000011011001", -- t[16601] = 1
      "0000001" when "00100000011011010", -- t[16602] = 1
      "0000001" when "00100000011011011", -- t[16603] = 1
      "0000001" when "00100000011011100", -- t[16604] = 1
      "0000001" when "00100000011011101", -- t[16605] = 1
      "0000001" when "00100000011011110", -- t[16606] = 1
      "0000001" when "00100000011011111", -- t[16607] = 1
      "0000001" when "00100000011100000", -- t[16608] = 1
      "0000001" when "00100000011100001", -- t[16609] = 1
      "0000001" when "00100000011100010", -- t[16610] = 1
      "0000001" when "00100000011100011", -- t[16611] = 1
      "0000001" when "00100000011100100", -- t[16612] = 1
      "0000001" when "00100000011100101", -- t[16613] = 1
      "0000001" when "00100000011100110", -- t[16614] = 1
      "0000001" when "00100000011100111", -- t[16615] = 1
      "0000001" when "00100000011101000", -- t[16616] = 1
      "0000001" when "00100000011101001", -- t[16617] = 1
      "0000001" when "00100000011101010", -- t[16618] = 1
      "0000001" when "00100000011101011", -- t[16619] = 1
      "0000001" when "00100000011101100", -- t[16620] = 1
      "0000001" when "00100000011101101", -- t[16621] = 1
      "0000001" when "00100000011101110", -- t[16622] = 1
      "0000001" when "00100000011101111", -- t[16623] = 1
      "0000001" when "00100000011110000", -- t[16624] = 1
      "0000001" when "00100000011110001", -- t[16625] = 1
      "0000001" when "00100000011110010", -- t[16626] = 1
      "0000001" when "00100000011110011", -- t[16627] = 1
      "0000001" when "00100000011110100", -- t[16628] = 1
      "0000001" when "00100000011110101", -- t[16629] = 1
      "0000001" when "00100000011110110", -- t[16630] = 1
      "0000001" when "00100000011110111", -- t[16631] = 1
      "0000001" when "00100000011111000", -- t[16632] = 1
      "0000001" when "00100000011111001", -- t[16633] = 1
      "0000001" when "00100000011111010", -- t[16634] = 1
      "0000001" when "00100000011111011", -- t[16635] = 1
      "0000001" when "00100000011111100", -- t[16636] = 1
      "0000001" when "00100000011111101", -- t[16637] = 1
      "0000001" when "00100000011111110", -- t[16638] = 1
      "0000001" when "00100000011111111", -- t[16639] = 1
      "0000001" when "00100000100000000", -- t[16640] = 1
      "0000001" when "00100000100000001", -- t[16641] = 1
      "0000001" when "00100000100000010", -- t[16642] = 1
      "0000001" when "00100000100000011", -- t[16643] = 1
      "0000001" when "00100000100000100", -- t[16644] = 1
      "0000001" when "00100000100000101", -- t[16645] = 1
      "0000001" when "00100000100000110", -- t[16646] = 1
      "0000001" when "00100000100000111", -- t[16647] = 1
      "0000001" when "00100000100001000", -- t[16648] = 1
      "0000001" when "00100000100001001", -- t[16649] = 1
      "0000001" when "00100000100001010", -- t[16650] = 1
      "0000001" when "00100000100001011", -- t[16651] = 1
      "0000001" when "00100000100001100", -- t[16652] = 1
      "0000001" when "00100000100001101", -- t[16653] = 1
      "0000001" when "00100000100001110", -- t[16654] = 1
      "0000001" when "00100000100001111", -- t[16655] = 1
      "0000001" when "00100000100010000", -- t[16656] = 1
      "0000001" when "00100000100010001", -- t[16657] = 1
      "0000001" when "00100000100010010", -- t[16658] = 1
      "0000001" when "00100000100010011", -- t[16659] = 1
      "0000001" when "00100000100010100", -- t[16660] = 1
      "0000001" when "00100000100010101", -- t[16661] = 1
      "0000001" when "00100000100010110", -- t[16662] = 1
      "0000001" when "00100000100010111", -- t[16663] = 1
      "0000001" when "00100000100011000", -- t[16664] = 1
      "0000001" when "00100000100011001", -- t[16665] = 1
      "0000001" when "00100000100011010", -- t[16666] = 1
      "0000001" when "00100000100011011", -- t[16667] = 1
      "0000001" when "00100000100011100", -- t[16668] = 1
      "0000001" when "00100000100011101", -- t[16669] = 1
      "0000001" when "00100000100011110", -- t[16670] = 1
      "0000001" when "00100000100011111", -- t[16671] = 1
      "0000001" when "00100000100100000", -- t[16672] = 1
      "0000001" when "00100000100100001", -- t[16673] = 1
      "0000001" when "00100000100100010", -- t[16674] = 1
      "0000001" when "00100000100100011", -- t[16675] = 1
      "0000001" when "00100000100100100", -- t[16676] = 1
      "0000001" when "00100000100100101", -- t[16677] = 1
      "0000001" when "00100000100100110", -- t[16678] = 1
      "0000001" when "00100000100100111", -- t[16679] = 1
      "0000001" when "00100000100101000", -- t[16680] = 1
      "0000001" when "00100000100101001", -- t[16681] = 1
      "0000001" when "00100000100101010", -- t[16682] = 1
      "0000001" when "00100000100101011", -- t[16683] = 1
      "0000001" when "00100000100101100", -- t[16684] = 1
      "0000001" when "00100000100101101", -- t[16685] = 1
      "0000001" when "00100000100101110", -- t[16686] = 1
      "0000001" when "00100000100101111", -- t[16687] = 1
      "0000001" when "00100000100110000", -- t[16688] = 1
      "0000001" when "00100000100110001", -- t[16689] = 1
      "0000001" when "00100000100110010", -- t[16690] = 1
      "0000001" when "00100000100110011", -- t[16691] = 1
      "0000001" when "00100000100110100", -- t[16692] = 1
      "0000001" when "00100000100110101", -- t[16693] = 1
      "0000001" when "00100000100110110", -- t[16694] = 1
      "0000001" when "00100000100110111", -- t[16695] = 1
      "0000001" when "00100000100111000", -- t[16696] = 1
      "0000001" when "00100000100111001", -- t[16697] = 1
      "0000001" when "00100000100111010", -- t[16698] = 1
      "0000001" when "00100000100111011", -- t[16699] = 1
      "0000001" when "00100000100111100", -- t[16700] = 1
      "0000001" when "00100000100111101", -- t[16701] = 1
      "0000001" when "00100000100111110", -- t[16702] = 1
      "0000001" when "00100000100111111", -- t[16703] = 1
      "0000001" when "00100000101000000", -- t[16704] = 1
      "0000001" when "00100000101000001", -- t[16705] = 1
      "0000001" when "00100000101000010", -- t[16706] = 1
      "0000001" when "00100000101000011", -- t[16707] = 1
      "0000001" when "00100000101000100", -- t[16708] = 1
      "0000001" when "00100000101000101", -- t[16709] = 1
      "0000001" when "00100000101000110", -- t[16710] = 1
      "0000001" when "00100000101000111", -- t[16711] = 1
      "0000001" when "00100000101001000", -- t[16712] = 1
      "0000001" when "00100000101001001", -- t[16713] = 1
      "0000001" when "00100000101001010", -- t[16714] = 1
      "0000001" when "00100000101001011", -- t[16715] = 1
      "0000001" when "00100000101001100", -- t[16716] = 1
      "0000001" when "00100000101001101", -- t[16717] = 1
      "0000001" when "00100000101001110", -- t[16718] = 1
      "0000001" when "00100000101001111", -- t[16719] = 1
      "0000001" when "00100000101010000", -- t[16720] = 1
      "0000001" when "00100000101010001", -- t[16721] = 1
      "0000001" when "00100000101010010", -- t[16722] = 1
      "0000001" when "00100000101010011", -- t[16723] = 1
      "0000001" when "00100000101010100", -- t[16724] = 1
      "0000001" when "00100000101010101", -- t[16725] = 1
      "0000001" when "00100000101010110", -- t[16726] = 1
      "0000001" when "00100000101010111", -- t[16727] = 1
      "0000001" when "00100000101011000", -- t[16728] = 1
      "0000001" when "00100000101011001", -- t[16729] = 1
      "0000001" when "00100000101011010", -- t[16730] = 1
      "0000001" when "00100000101011011", -- t[16731] = 1
      "0000001" when "00100000101011100", -- t[16732] = 1
      "0000001" when "00100000101011101", -- t[16733] = 1
      "0000001" when "00100000101011110", -- t[16734] = 1
      "0000001" when "00100000101011111", -- t[16735] = 1
      "0000001" when "00100000101100000", -- t[16736] = 1
      "0000001" when "00100000101100001", -- t[16737] = 1
      "0000001" when "00100000101100010", -- t[16738] = 1
      "0000001" when "00100000101100011", -- t[16739] = 1
      "0000001" when "00100000101100100", -- t[16740] = 1
      "0000001" when "00100000101100101", -- t[16741] = 1
      "0000001" when "00100000101100110", -- t[16742] = 1
      "0000001" when "00100000101100111", -- t[16743] = 1
      "0000001" when "00100000101101000", -- t[16744] = 1
      "0000001" when "00100000101101001", -- t[16745] = 1
      "0000001" when "00100000101101010", -- t[16746] = 1
      "0000001" when "00100000101101011", -- t[16747] = 1
      "0000001" when "00100000101101100", -- t[16748] = 1
      "0000001" when "00100000101101101", -- t[16749] = 1
      "0000001" when "00100000101101110", -- t[16750] = 1
      "0000001" when "00100000101101111", -- t[16751] = 1
      "0000001" when "00100000101110000", -- t[16752] = 1
      "0000001" when "00100000101110001", -- t[16753] = 1
      "0000001" when "00100000101110010", -- t[16754] = 1
      "0000001" when "00100000101110011", -- t[16755] = 1
      "0000001" when "00100000101110100", -- t[16756] = 1
      "0000001" when "00100000101110101", -- t[16757] = 1
      "0000001" when "00100000101110110", -- t[16758] = 1
      "0000001" when "00100000101110111", -- t[16759] = 1
      "0000001" when "00100000101111000", -- t[16760] = 1
      "0000001" when "00100000101111001", -- t[16761] = 1
      "0000001" when "00100000101111010", -- t[16762] = 1
      "0000001" when "00100000101111011", -- t[16763] = 1
      "0000001" when "00100000101111100", -- t[16764] = 1
      "0000001" when "00100000101111101", -- t[16765] = 1
      "0000001" when "00100000101111110", -- t[16766] = 1
      "0000001" when "00100000101111111", -- t[16767] = 1
      "0000001" when "00100000110000000", -- t[16768] = 1
      "0000001" when "00100000110000001", -- t[16769] = 1
      "0000001" when "00100000110000010", -- t[16770] = 1
      "0000001" when "00100000110000011", -- t[16771] = 1
      "0000001" when "00100000110000100", -- t[16772] = 1
      "0000001" when "00100000110000101", -- t[16773] = 1
      "0000001" when "00100000110000110", -- t[16774] = 1
      "0000001" when "00100000110000111", -- t[16775] = 1
      "0000001" when "00100000110001000", -- t[16776] = 1
      "0000001" when "00100000110001001", -- t[16777] = 1
      "0000001" when "00100000110001010", -- t[16778] = 1
      "0000001" when "00100000110001011", -- t[16779] = 1
      "0000001" when "00100000110001100", -- t[16780] = 1
      "0000001" when "00100000110001101", -- t[16781] = 1
      "0000001" when "00100000110001110", -- t[16782] = 1
      "0000001" when "00100000110001111", -- t[16783] = 1
      "0000001" when "00100000110010000", -- t[16784] = 1
      "0000001" when "00100000110010001", -- t[16785] = 1
      "0000001" when "00100000110010010", -- t[16786] = 1
      "0000001" when "00100000110010011", -- t[16787] = 1
      "0000001" when "00100000110010100", -- t[16788] = 1
      "0000001" when "00100000110010101", -- t[16789] = 1
      "0000001" when "00100000110010110", -- t[16790] = 1
      "0000001" when "00100000110010111", -- t[16791] = 1
      "0000001" when "00100000110011000", -- t[16792] = 1
      "0000001" when "00100000110011001", -- t[16793] = 1
      "0000001" when "00100000110011010", -- t[16794] = 1
      "0000001" when "00100000110011011", -- t[16795] = 1
      "0000001" when "00100000110011100", -- t[16796] = 1
      "0000001" when "00100000110011101", -- t[16797] = 1
      "0000001" when "00100000110011110", -- t[16798] = 1
      "0000001" when "00100000110011111", -- t[16799] = 1
      "0000001" when "00100000110100000", -- t[16800] = 1
      "0000001" when "00100000110100001", -- t[16801] = 1
      "0000001" when "00100000110100010", -- t[16802] = 1
      "0000001" when "00100000110100011", -- t[16803] = 1
      "0000001" when "00100000110100100", -- t[16804] = 1
      "0000001" when "00100000110100101", -- t[16805] = 1
      "0000001" when "00100000110100110", -- t[16806] = 1
      "0000001" when "00100000110100111", -- t[16807] = 1
      "0000001" when "00100000110101000", -- t[16808] = 1
      "0000001" when "00100000110101001", -- t[16809] = 1
      "0000001" when "00100000110101010", -- t[16810] = 1
      "0000001" when "00100000110101011", -- t[16811] = 1
      "0000001" when "00100000110101100", -- t[16812] = 1
      "0000001" when "00100000110101101", -- t[16813] = 1
      "0000001" when "00100000110101110", -- t[16814] = 1
      "0000001" when "00100000110101111", -- t[16815] = 1
      "0000001" when "00100000110110000", -- t[16816] = 1
      "0000001" when "00100000110110001", -- t[16817] = 1
      "0000001" when "00100000110110010", -- t[16818] = 1
      "0000001" when "00100000110110011", -- t[16819] = 1
      "0000001" when "00100000110110100", -- t[16820] = 1
      "0000001" when "00100000110110101", -- t[16821] = 1
      "0000001" when "00100000110110110", -- t[16822] = 1
      "0000001" when "00100000110110111", -- t[16823] = 1
      "0000001" when "00100000110111000", -- t[16824] = 1
      "0000001" when "00100000110111001", -- t[16825] = 1
      "0000001" when "00100000110111010", -- t[16826] = 1
      "0000001" when "00100000110111011", -- t[16827] = 1
      "0000001" when "00100000110111100", -- t[16828] = 1
      "0000001" when "00100000110111101", -- t[16829] = 1
      "0000001" when "00100000110111110", -- t[16830] = 1
      "0000001" when "00100000110111111", -- t[16831] = 1
      "0000001" when "00100000111000000", -- t[16832] = 1
      "0000001" when "00100000111000001", -- t[16833] = 1
      "0000001" when "00100000111000010", -- t[16834] = 1
      "0000001" when "00100000111000011", -- t[16835] = 1
      "0000001" when "00100000111000100", -- t[16836] = 1
      "0000001" when "00100000111000101", -- t[16837] = 1
      "0000001" when "00100000111000110", -- t[16838] = 1
      "0000001" when "00100000111000111", -- t[16839] = 1
      "0000001" when "00100000111001000", -- t[16840] = 1
      "0000001" when "00100000111001001", -- t[16841] = 1
      "0000001" when "00100000111001010", -- t[16842] = 1
      "0000001" when "00100000111001011", -- t[16843] = 1
      "0000001" when "00100000111001100", -- t[16844] = 1
      "0000001" when "00100000111001101", -- t[16845] = 1
      "0000001" when "00100000111001110", -- t[16846] = 1
      "0000001" when "00100000111001111", -- t[16847] = 1
      "0000001" when "00100000111010000", -- t[16848] = 1
      "0000001" when "00100000111010001", -- t[16849] = 1
      "0000001" when "00100000111010010", -- t[16850] = 1
      "0000001" when "00100000111010011", -- t[16851] = 1
      "0000001" when "00100000111010100", -- t[16852] = 1
      "0000001" when "00100000111010101", -- t[16853] = 1
      "0000001" when "00100000111010110", -- t[16854] = 1
      "0000001" when "00100000111010111", -- t[16855] = 1
      "0000001" when "00100000111011000", -- t[16856] = 1
      "0000001" when "00100000111011001", -- t[16857] = 1
      "0000001" when "00100000111011010", -- t[16858] = 1
      "0000001" when "00100000111011011", -- t[16859] = 1
      "0000001" when "00100000111011100", -- t[16860] = 1
      "0000001" when "00100000111011101", -- t[16861] = 1
      "0000001" when "00100000111011110", -- t[16862] = 1
      "0000001" when "00100000111011111", -- t[16863] = 1
      "0000001" when "00100000111100000", -- t[16864] = 1
      "0000001" when "00100000111100001", -- t[16865] = 1
      "0000001" when "00100000111100010", -- t[16866] = 1
      "0000001" when "00100000111100011", -- t[16867] = 1
      "0000001" when "00100000111100100", -- t[16868] = 1
      "0000001" when "00100000111100101", -- t[16869] = 1
      "0000001" when "00100000111100110", -- t[16870] = 1
      "0000001" when "00100000111100111", -- t[16871] = 1
      "0000001" when "00100000111101000", -- t[16872] = 1
      "0000001" when "00100000111101001", -- t[16873] = 1
      "0000001" when "00100000111101010", -- t[16874] = 1
      "0000001" when "00100000111101011", -- t[16875] = 1
      "0000001" when "00100000111101100", -- t[16876] = 1
      "0000001" when "00100000111101101", -- t[16877] = 1
      "0000001" when "00100000111101110", -- t[16878] = 1
      "0000001" when "00100000111101111", -- t[16879] = 1
      "0000001" when "00100000111110000", -- t[16880] = 1
      "0000001" when "00100000111110001", -- t[16881] = 1
      "0000001" when "00100000111110010", -- t[16882] = 1
      "0000001" when "00100000111110011", -- t[16883] = 1
      "0000001" when "00100000111110100", -- t[16884] = 1
      "0000001" when "00100000111110101", -- t[16885] = 1
      "0000001" when "00100000111110110", -- t[16886] = 1
      "0000001" when "00100000111110111", -- t[16887] = 1
      "0000001" when "00100000111111000", -- t[16888] = 1
      "0000001" when "00100000111111001", -- t[16889] = 1
      "0000001" when "00100000111111010", -- t[16890] = 1
      "0000001" when "00100000111111011", -- t[16891] = 1
      "0000001" when "00100000111111100", -- t[16892] = 1
      "0000001" when "00100000111111101", -- t[16893] = 1
      "0000001" when "00100000111111110", -- t[16894] = 1
      "0000001" when "00100000111111111", -- t[16895] = 1
      "0000001" when "00100001000000000", -- t[16896] = 1
      "0000001" when "00100001000000001", -- t[16897] = 1
      "0000001" when "00100001000000010", -- t[16898] = 1
      "0000001" when "00100001000000011", -- t[16899] = 1
      "0000001" when "00100001000000100", -- t[16900] = 1
      "0000001" when "00100001000000101", -- t[16901] = 1
      "0000001" when "00100001000000110", -- t[16902] = 1
      "0000001" when "00100001000000111", -- t[16903] = 1
      "0000001" when "00100001000001000", -- t[16904] = 1
      "0000001" when "00100001000001001", -- t[16905] = 1
      "0000001" when "00100001000001010", -- t[16906] = 1
      "0000001" when "00100001000001011", -- t[16907] = 1
      "0000001" when "00100001000001100", -- t[16908] = 1
      "0000001" when "00100001000001101", -- t[16909] = 1
      "0000001" when "00100001000001110", -- t[16910] = 1
      "0000001" when "00100001000001111", -- t[16911] = 1
      "0000001" when "00100001000010000", -- t[16912] = 1
      "0000001" when "00100001000010001", -- t[16913] = 1
      "0000001" when "00100001000010010", -- t[16914] = 1
      "0000001" when "00100001000010011", -- t[16915] = 1
      "0000001" when "00100001000010100", -- t[16916] = 1
      "0000001" when "00100001000010101", -- t[16917] = 1
      "0000001" when "00100001000010110", -- t[16918] = 1
      "0000001" when "00100001000010111", -- t[16919] = 1
      "0000001" when "00100001000011000", -- t[16920] = 1
      "0000001" when "00100001000011001", -- t[16921] = 1
      "0000001" when "00100001000011010", -- t[16922] = 1
      "0000001" when "00100001000011011", -- t[16923] = 1
      "0000001" when "00100001000011100", -- t[16924] = 1
      "0000001" when "00100001000011101", -- t[16925] = 1
      "0000001" when "00100001000011110", -- t[16926] = 1
      "0000001" when "00100001000011111", -- t[16927] = 1
      "0000001" when "00100001000100000", -- t[16928] = 1
      "0000001" when "00100001000100001", -- t[16929] = 1
      "0000001" when "00100001000100010", -- t[16930] = 1
      "0000001" when "00100001000100011", -- t[16931] = 1
      "0000001" when "00100001000100100", -- t[16932] = 1
      "0000001" when "00100001000100101", -- t[16933] = 1
      "0000001" when "00100001000100110", -- t[16934] = 1
      "0000001" when "00100001000100111", -- t[16935] = 1
      "0000001" when "00100001000101000", -- t[16936] = 1
      "0000001" when "00100001000101001", -- t[16937] = 1
      "0000001" when "00100001000101010", -- t[16938] = 1
      "0000001" when "00100001000101011", -- t[16939] = 1
      "0000001" when "00100001000101100", -- t[16940] = 1
      "0000001" when "00100001000101101", -- t[16941] = 1
      "0000001" when "00100001000101110", -- t[16942] = 1
      "0000001" when "00100001000101111", -- t[16943] = 1
      "0000001" when "00100001000110000", -- t[16944] = 1
      "0000001" when "00100001000110001", -- t[16945] = 1
      "0000001" when "00100001000110010", -- t[16946] = 1
      "0000001" when "00100001000110011", -- t[16947] = 1
      "0000001" when "00100001000110100", -- t[16948] = 1
      "0000001" when "00100001000110101", -- t[16949] = 1
      "0000001" when "00100001000110110", -- t[16950] = 1
      "0000001" when "00100001000110111", -- t[16951] = 1
      "0000001" when "00100001000111000", -- t[16952] = 1
      "0000001" when "00100001000111001", -- t[16953] = 1
      "0000001" when "00100001000111010", -- t[16954] = 1
      "0000001" when "00100001000111011", -- t[16955] = 1
      "0000001" when "00100001000111100", -- t[16956] = 1
      "0000001" when "00100001000111101", -- t[16957] = 1
      "0000001" when "00100001000111110", -- t[16958] = 1
      "0000001" when "00100001000111111", -- t[16959] = 1
      "0000001" when "00100001001000000", -- t[16960] = 1
      "0000001" when "00100001001000001", -- t[16961] = 1
      "0000001" when "00100001001000010", -- t[16962] = 1
      "0000001" when "00100001001000011", -- t[16963] = 1
      "0000001" when "00100001001000100", -- t[16964] = 1
      "0000001" when "00100001001000101", -- t[16965] = 1
      "0000001" when "00100001001000110", -- t[16966] = 1
      "0000001" when "00100001001000111", -- t[16967] = 1
      "0000001" when "00100001001001000", -- t[16968] = 1
      "0000001" when "00100001001001001", -- t[16969] = 1
      "0000001" when "00100001001001010", -- t[16970] = 1
      "0000001" when "00100001001001011", -- t[16971] = 1
      "0000001" when "00100001001001100", -- t[16972] = 1
      "0000001" when "00100001001001101", -- t[16973] = 1
      "0000001" when "00100001001001110", -- t[16974] = 1
      "0000001" when "00100001001001111", -- t[16975] = 1
      "0000001" when "00100001001010000", -- t[16976] = 1
      "0000001" when "00100001001010001", -- t[16977] = 1
      "0000001" when "00100001001010010", -- t[16978] = 1
      "0000001" when "00100001001010011", -- t[16979] = 1
      "0000001" when "00100001001010100", -- t[16980] = 1
      "0000001" when "00100001001010101", -- t[16981] = 1
      "0000001" when "00100001001010110", -- t[16982] = 1
      "0000001" when "00100001001010111", -- t[16983] = 1
      "0000001" when "00100001001011000", -- t[16984] = 1
      "0000001" when "00100001001011001", -- t[16985] = 1
      "0000001" when "00100001001011010", -- t[16986] = 1
      "0000001" when "00100001001011011", -- t[16987] = 1
      "0000001" when "00100001001011100", -- t[16988] = 1
      "0000001" when "00100001001011101", -- t[16989] = 1
      "0000001" when "00100001001011110", -- t[16990] = 1
      "0000001" when "00100001001011111", -- t[16991] = 1
      "0000001" when "00100001001100000", -- t[16992] = 1
      "0000001" when "00100001001100001", -- t[16993] = 1
      "0000001" when "00100001001100010", -- t[16994] = 1
      "0000001" when "00100001001100011", -- t[16995] = 1
      "0000001" when "00100001001100100", -- t[16996] = 1
      "0000001" when "00100001001100101", -- t[16997] = 1
      "0000001" when "00100001001100110", -- t[16998] = 1
      "0000001" when "00100001001100111", -- t[16999] = 1
      "0000001" when "00100001001101000", -- t[17000] = 1
      "0000001" when "00100001001101001", -- t[17001] = 1
      "0000001" when "00100001001101010", -- t[17002] = 1
      "0000001" when "00100001001101011", -- t[17003] = 1
      "0000001" when "00100001001101100", -- t[17004] = 1
      "0000001" when "00100001001101101", -- t[17005] = 1
      "0000001" when "00100001001101110", -- t[17006] = 1
      "0000001" when "00100001001101111", -- t[17007] = 1
      "0000001" when "00100001001110000", -- t[17008] = 1
      "0000001" when "00100001001110001", -- t[17009] = 1
      "0000001" when "00100001001110010", -- t[17010] = 1
      "0000001" when "00100001001110011", -- t[17011] = 1
      "0000001" when "00100001001110100", -- t[17012] = 1
      "0000001" when "00100001001110101", -- t[17013] = 1
      "0000001" when "00100001001110110", -- t[17014] = 1
      "0000001" when "00100001001110111", -- t[17015] = 1
      "0000001" when "00100001001111000", -- t[17016] = 1
      "0000001" when "00100001001111001", -- t[17017] = 1
      "0000001" when "00100001001111010", -- t[17018] = 1
      "0000001" when "00100001001111011", -- t[17019] = 1
      "0000001" when "00100001001111100", -- t[17020] = 1
      "0000001" when "00100001001111101", -- t[17021] = 1
      "0000001" when "00100001001111110", -- t[17022] = 1
      "0000001" when "00100001001111111", -- t[17023] = 1
      "0000001" when "00100001010000000", -- t[17024] = 1
      "0000001" when "00100001010000001", -- t[17025] = 1
      "0000001" when "00100001010000010", -- t[17026] = 1
      "0000001" when "00100001010000011", -- t[17027] = 1
      "0000001" when "00100001010000100", -- t[17028] = 1
      "0000001" when "00100001010000101", -- t[17029] = 1
      "0000001" when "00100001010000110", -- t[17030] = 1
      "0000001" when "00100001010000111", -- t[17031] = 1
      "0000001" when "00100001010001000", -- t[17032] = 1
      "0000001" when "00100001010001001", -- t[17033] = 1
      "0000001" when "00100001010001010", -- t[17034] = 1
      "0000001" when "00100001010001011", -- t[17035] = 1
      "0000001" when "00100001010001100", -- t[17036] = 1
      "0000001" when "00100001010001101", -- t[17037] = 1
      "0000001" when "00100001010001110", -- t[17038] = 1
      "0000001" when "00100001010001111", -- t[17039] = 1
      "0000001" when "00100001010010000", -- t[17040] = 1
      "0000001" when "00100001010010001", -- t[17041] = 1
      "0000001" when "00100001010010010", -- t[17042] = 1
      "0000001" when "00100001010010011", -- t[17043] = 1
      "0000001" when "00100001010010100", -- t[17044] = 1
      "0000001" when "00100001010010101", -- t[17045] = 1
      "0000001" when "00100001010010110", -- t[17046] = 1
      "0000001" when "00100001010010111", -- t[17047] = 1
      "0000001" when "00100001010011000", -- t[17048] = 1
      "0000001" when "00100001010011001", -- t[17049] = 1
      "0000001" when "00100001010011010", -- t[17050] = 1
      "0000001" when "00100001010011011", -- t[17051] = 1
      "0000001" when "00100001010011100", -- t[17052] = 1
      "0000001" when "00100001010011101", -- t[17053] = 1
      "0000001" when "00100001010011110", -- t[17054] = 1
      "0000001" when "00100001010011111", -- t[17055] = 1
      "0000001" when "00100001010100000", -- t[17056] = 1
      "0000001" when "00100001010100001", -- t[17057] = 1
      "0000001" when "00100001010100010", -- t[17058] = 1
      "0000001" when "00100001010100011", -- t[17059] = 1
      "0000001" when "00100001010100100", -- t[17060] = 1
      "0000001" when "00100001010100101", -- t[17061] = 1
      "0000001" when "00100001010100110", -- t[17062] = 1
      "0000001" when "00100001010100111", -- t[17063] = 1
      "0000001" when "00100001010101000", -- t[17064] = 1
      "0000001" when "00100001010101001", -- t[17065] = 1
      "0000001" when "00100001010101010", -- t[17066] = 1
      "0000001" when "00100001010101011", -- t[17067] = 1
      "0000001" when "00100001010101100", -- t[17068] = 1
      "0000001" when "00100001010101101", -- t[17069] = 1
      "0000001" when "00100001010101110", -- t[17070] = 1
      "0000001" when "00100001010101111", -- t[17071] = 1
      "0000001" when "00100001010110000", -- t[17072] = 1
      "0000001" when "00100001010110001", -- t[17073] = 1
      "0000001" when "00100001010110010", -- t[17074] = 1
      "0000001" when "00100001010110011", -- t[17075] = 1
      "0000001" when "00100001010110100", -- t[17076] = 1
      "0000001" when "00100001010110101", -- t[17077] = 1
      "0000001" when "00100001010110110", -- t[17078] = 1
      "0000001" when "00100001010110111", -- t[17079] = 1
      "0000001" when "00100001010111000", -- t[17080] = 1
      "0000001" when "00100001010111001", -- t[17081] = 1
      "0000001" when "00100001010111010", -- t[17082] = 1
      "0000001" when "00100001010111011", -- t[17083] = 1
      "0000001" when "00100001010111100", -- t[17084] = 1
      "0000001" when "00100001010111101", -- t[17085] = 1
      "0000001" when "00100001010111110", -- t[17086] = 1
      "0000001" when "00100001010111111", -- t[17087] = 1
      "0000001" when "00100001011000000", -- t[17088] = 1
      "0000001" when "00100001011000001", -- t[17089] = 1
      "0000001" when "00100001011000010", -- t[17090] = 1
      "0000001" when "00100001011000011", -- t[17091] = 1
      "0000001" when "00100001011000100", -- t[17092] = 1
      "0000001" when "00100001011000101", -- t[17093] = 1
      "0000001" when "00100001011000110", -- t[17094] = 1
      "0000001" when "00100001011000111", -- t[17095] = 1
      "0000001" when "00100001011001000", -- t[17096] = 1
      "0000001" when "00100001011001001", -- t[17097] = 1
      "0000001" when "00100001011001010", -- t[17098] = 1
      "0000001" when "00100001011001011", -- t[17099] = 1
      "0000001" when "00100001011001100", -- t[17100] = 1
      "0000001" when "00100001011001101", -- t[17101] = 1
      "0000001" when "00100001011001110", -- t[17102] = 1
      "0000001" when "00100001011001111", -- t[17103] = 1
      "0000001" when "00100001011010000", -- t[17104] = 1
      "0000001" when "00100001011010001", -- t[17105] = 1
      "0000001" when "00100001011010010", -- t[17106] = 1
      "0000001" when "00100001011010011", -- t[17107] = 1
      "0000001" when "00100001011010100", -- t[17108] = 1
      "0000001" when "00100001011010101", -- t[17109] = 1
      "0000001" when "00100001011010110", -- t[17110] = 1
      "0000001" when "00100001011010111", -- t[17111] = 1
      "0000001" when "00100001011011000", -- t[17112] = 1
      "0000001" when "00100001011011001", -- t[17113] = 1
      "0000001" when "00100001011011010", -- t[17114] = 1
      "0000001" when "00100001011011011", -- t[17115] = 1
      "0000001" when "00100001011011100", -- t[17116] = 1
      "0000001" when "00100001011011101", -- t[17117] = 1
      "0000001" when "00100001011011110", -- t[17118] = 1
      "0000001" when "00100001011011111", -- t[17119] = 1
      "0000001" when "00100001011100000", -- t[17120] = 1
      "0000001" when "00100001011100001", -- t[17121] = 1
      "0000001" when "00100001011100010", -- t[17122] = 1
      "0000001" when "00100001011100011", -- t[17123] = 1
      "0000001" when "00100001011100100", -- t[17124] = 1
      "0000001" when "00100001011100101", -- t[17125] = 1
      "0000001" when "00100001011100110", -- t[17126] = 1
      "0000001" when "00100001011100111", -- t[17127] = 1
      "0000001" when "00100001011101000", -- t[17128] = 1
      "0000001" when "00100001011101001", -- t[17129] = 1
      "0000001" when "00100001011101010", -- t[17130] = 1
      "0000001" when "00100001011101011", -- t[17131] = 1
      "0000001" when "00100001011101100", -- t[17132] = 1
      "0000001" when "00100001011101101", -- t[17133] = 1
      "0000001" when "00100001011101110", -- t[17134] = 1
      "0000001" when "00100001011101111", -- t[17135] = 1
      "0000001" when "00100001011110000", -- t[17136] = 1
      "0000001" when "00100001011110001", -- t[17137] = 1
      "0000001" when "00100001011110010", -- t[17138] = 1
      "0000001" when "00100001011110011", -- t[17139] = 1
      "0000001" when "00100001011110100", -- t[17140] = 1
      "0000001" when "00100001011110101", -- t[17141] = 1
      "0000001" when "00100001011110110", -- t[17142] = 1
      "0000001" when "00100001011110111", -- t[17143] = 1
      "0000001" when "00100001011111000", -- t[17144] = 1
      "0000001" when "00100001011111001", -- t[17145] = 1
      "0000001" when "00100001011111010", -- t[17146] = 1
      "0000001" when "00100001011111011", -- t[17147] = 1
      "0000001" when "00100001011111100", -- t[17148] = 1
      "0000001" when "00100001011111101", -- t[17149] = 1
      "0000001" when "00100001011111110", -- t[17150] = 1
      "0000001" when "00100001011111111", -- t[17151] = 1
      "0000001" when "00100001100000000", -- t[17152] = 1
      "0000001" when "00100001100000001", -- t[17153] = 1
      "0000001" when "00100001100000010", -- t[17154] = 1
      "0000001" when "00100001100000011", -- t[17155] = 1
      "0000001" when "00100001100000100", -- t[17156] = 1
      "0000001" when "00100001100000101", -- t[17157] = 1
      "0000001" when "00100001100000110", -- t[17158] = 1
      "0000001" when "00100001100000111", -- t[17159] = 1
      "0000001" when "00100001100001000", -- t[17160] = 1
      "0000001" when "00100001100001001", -- t[17161] = 1
      "0000001" when "00100001100001010", -- t[17162] = 1
      "0000001" when "00100001100001011", -- t[17163] = 1
      "0000001" when "00100001100001100", -- t[17164] = 1
      "0000001" when "00100001100001101", -- t[17165] = 1
      "0000001" when "00100001100001110", -- t[17166] = 1
      "0000001" when "00100001100001111", -- t[17167] = 1
      "0000001" when "00100001100010000", -- t[17168] = 1
      "0000001" when "00100001100010001", -- t[17169] = 1
      "0000001" when "00100001100010010", -- t[17170] = 1
      "0000001" when "00100001100010011", -- t[17171] = 1
      "0000001" when "00100001100010100", -- t[17172] = 1
      "0000001" when "00100001100010101", -- t[17173] = 1
      "0000001" when "00100001100010110", -- t[17174] = 1
      "0000001" when "00100001100010111", -- t[17175] = 1
      "0000001" when "00100001100011000", -- t[17176] = 1
      "0000001" when "00100001100011001", -- t[17177] = 1
      "0000001" when "00100001100011010", -- t[17178] = 1
      "0000001" when "00100001100011011", -- t[17179] = 1
      "0000001" when "00100001100011100", -- t[17180] = 1
      "0000001" when "00100001100011101", -- t[17181] = 1
      "0000001" when "00100001100011110", -- t[17182] = 1
      "0000001" when "00100001100011111", -- t[17183] = 1
      "0000001" when "00100001100100000", -- t[17184] = 1
      "0000001" when "00100001100100001", -- t[17185] = 1
      "0000001" when "00100001100100010", -- t[17186] = 1
      "0000001" when "00100001100100011", -- t[17187] = 1
      "0000001" when "00100001100100100", -- t[17188] = 1
      "0000001" when "00100001100100101", -- t[17189] = 1
      "0000001" when "00100001100100110", -- t[17190] = 1
      "0000001" when "00100001100100111", -- t[17191] = 1
      "0000001" when "00100001100101000", -- t[17192] = 1
      "0000001" when "00100001100101001", -- t[17193] = 1
      "0000001" when "00100001100101010", -- t[17194] = 1
      "0000001" when "00100001100101011", -- t[17195] = 1
      "0000001" when "00100001100101100", -- t[17196] = 1
      "0000001" when "00100001100101101", -- t[17197] = 1
      "0000001" when "00100001100101110", -- t[17198] = 1
      "0000001" when "00100001100101111", -- t[17199] = 1
      "0000001" when "00100001100110000", -- t[17200] = 1
      "0000001" when "00100001100110001", -- t[17201] = 1
      "0000001" when "00100001100110010", -- t[17202] = 1
      "0000001" when "00100001100110011", -- t[17203] = 1
      "0000001" when "00100001100110100", -- t[17204] = 1
      "0000001" when "00100001100110101", -- t[17205] = 1
      "0000001" when "00100001100110110", -- t[17206] = 1
      "0000001" when "00100001100110111", -- t[17207] = 1
      "0000001" when "00100001100111000", -- t[17208] = 1
      "0000001" when "00100001100111001", -- t[17209] = 1
      "0000001" when "00100001100111010", -- t[17210] = 1
      "0000001" when "00100001100111011", -- t[17211] = 1
      "0000001" when "00100001100111100", -- t[17212] = 1
      "0000001" when "00100001100111101", -- t[17213] = 1
      "0000001" when "00100001100111110", -- t[17214] = 1
      "0000001" when "00100001100111111", -- t[17215] = 1
      "0000001" when "00100001101000000", -- t[17216] = 1
      "0000001" when "00100001101000001", -- t[17217] = 1
      "0000001" when "00100001101000010", -- t[17218] = 1
      "0000001" when "00100001101000011", -- t[17219] = 1
      "0000001" when "00100001101000100", -- t[17220] = 1
      "0000001" when "00100001101000101", -- t[17221] = 1
      "0000001" when "00100001101000110", -- t[17222] = 1
      "0000001" when "00100001101000111", -- t[17223] = 1
      "0000001" when "00100001101001000", -- t[17224] = 1
      "0000001" when "00100001101001001", -- t[17225] = 1
      "0000001" when "00100001101001010", -- t[17226] = 1
      "0000001" when "00100001101001011", -- t[17227] = 1
      "0000001" when "00100001101001100", -- t[17228] = 1
      "0000001" when "00100001101001101", -- t[17229] = 1
      "0000001" when "00100001101001110", -- t[17230] = 1
      "0000001" when "00100001101001111", -- t[17231] = 1
      "0000001" when "00100001101010000", -- t[17232] = 1
      "0000001" when "00100001101010001", -- t[17233] = 1
      "0000001" when "00100001101010010", -- t[17234] = 1
      "0000001" when "00100001101010011", -- t[17235] = 1
      "0000001" when "00100001101010100", -- t[17236] = 1
      "0000001" when "00100001101010101", -- t[17237] = 1
      "0000001" when "00100001101010110", -- t[17238] = 1
      "0000001" when "00100001101010111", -- t[17239] = 1
      "0000001" when "00100001101011000", -- t[17240] = 1
      "0000001" when "00100001101011001", -- t[17241] = 1
      "0000001" when "00100001101011010", -- t[17242] = 1
      "0000001" when "00100001101011011", -- t[17243] = 1
      "0000001" when "00100001101011100", -- t[17244] = 1
      "0000001" when "00100001101011101", -- t[17245] = 1
      "0000001" when "00100001101011110", -- t[17246] = 1
      "0000001" when "00100001101011111", -- t[17247] = 1
      "0000001" when "00100001101100000", -- t[17248] = 1
      "0000001" when "00100001101100001", -- t[17249] = 1
      "0000001" when "00100001101100010", -- t[17250] = 1
      "0000001" when "00100001101100011", -- t[17251] = 1
      "0000001" when "00100001101100100", -- t[17252] = 1
      "0000001" when "00100001101100101", -- t[17253] = 1
      "0000001" when "00100001101100110", -- t[17254] = 1
      "0000001" when "00100001101100111", -- t[17255] = 1
      "0000001" when "00100001101101000", -- t[17256] = 1
      "0000001" when "00100001101101001", -- t[17257] = 1
      "0000001" when "00100001101101010", -- t[17258] = 1
      "0000001" when "00100001101101011", -- t[17259] = 1
      "0000001" when "00100001101101100", -- t[17260] = 1
      "0000001" when "00100001101101101", -- t[17261] = 1
      "0000001" when "00100001101101110", -- t[17262] = 1
      "0000001" when "00100001101101111", -- t[17263] = 1
      "0000001" when "00100001101110000", -- t[17264] = 1
      "0000001" when "00100001101110001", -- t[17265] = 1
      "0000001" when "00100001101110010", -- t[17266] = 1
      "0000001" when "00100001101110011", -- t[17267] = 1
      "0000001" when "00100001101110100", -- t[17268] = 1
      "0000001" when "00100001101110101", -- t[17269] = 1
      "0000001" when "00100001101110110", -- t[17270] = 1
      "0000001" when "00100001101110111", -- t[17271] = 1
      "0000001" when "00100001101111000", -- t[17272] = 1
      "0000001" when "00100001101111001", -- t[17273] = 1
      "0000001" when "00100001101111010", -- t[17274] = 1
      "0000001" when "00100001101111011", -- t[17275] = 1
      "0000001" when "00100001101111100", -- t[17276] = 1
      "0000001" when "00100001101111101", -- t[17277] = 1
      "0000001" when "00100001101111110", -- t[17278] = 1
      "0000001" when "00100001101111111", -- t[17279] = 1
      "0000001" when "00100001110000000", -- t[17280] = 1
      "0000001" when "00100001110000001", -- t[17281] = 1
      "0000001" when "00100001110000010", -- t[17282] = 1
      "0000001" when "00100001110000011", -- t[17283] = 1
      "0000001" when "00100001110000100", -- t[17284] = 1
      "0000001" when "00100001110000101", -- t[17285] = 1
      "0000001" when "00100001110000110", -- t[17286] = 1
      "0000001" when "00100001110000111", -- t[17287] = 1
      "0000001" when "00100001110001000", -- t[17288] = 1
      "0000001" when "00100001110001001", -- t[17289] = 1
      "0000001" when "00100001110001010", -- t[17290] = 1
      "0000001" when "00100001110001011", -- t[17291] = 1
      "0000001" when "00100001110001100", -- t[17292] = 1
      "0000001" when "00100001110001101", -- t[17293] = 1
      "0000001" when "00100001110001110", -- t[17294] = 1
      "0000001" when "00100001110001111", -- t[17295] = 1
      "0000001" when "00100001110010000", -- t[17296] = 1
      "0000001" when "00100001110010001", -- t[17297] = 1
      "0000001" when "00100001110010010", -- t[17298] = 1
      "0000001" when "00100001110010011", -- t[17299] = 1
      "0000001" when "00100001110010100", -- t[17300] = 1
      "0000001" when "00100001110010101", -- t[17301] = 1
      "0000001" when "00100001110010110", -- t[17302] = 1
      "0000001" when "00100001110010111", -- t[17303] = 1
      "0000001" when "00100001110011000", -- t[17304] = 1
      "0000001" when "00100001110011001", -- t[17305] = 1
      "0000001" when "00100001110011010", -- t[17306] = 1
      "0000001" when "00100001110011011", -- t[17307] = 1
      "0000001" when "00100001110011100", -- t[17308] = 1
      "0000001" when "00100001110011101", -- t[17309] = 1
      "0000001" when "00100001110011110", -- t[17310] = 1
      "0000001" when "00100001110011111", -- t[17311] = 1
      "0000001" when "00100001110100000", -- t[17312] = 1
      "0000001" when "00100001110100001", -- t[17313] = 1
      "0000001" when "00100001110100010", -- t[17314] = 1
      "0000001" when "00100001110100011", -- t[17315] = 1
      "0000001" when "00100001110100100", -- t[17316] = 1
      "0000001" when "00100001110100101", -- t[17317] = 1
      "0000001" when "00100001110100110", -- t[17318] = 1
      "0000001" when "00100001110100111", -- t[17319] = 1
      "0000001" when "00100001110101000", -- t[17320] = 1
      "0000001" when "00100001110101001", -- t[17321] = 1
      "0000001" when "00100001110101010", -- t[17322] = 1
      "0000001" when "00100001110101011", -- t[17323] = 1
      "0000001" when "00100001110101100", -- t[17324] = 1
      "0000001" when "00100001110101101", -- t[17325] = 1
      "0000001" when "00100001110101110", -- t[17326] = 1
      "0000001" when "00100001110101111", -- t[17327] = 1
      "0000001" when "00100001110110000", -- t[17328] = 1
      "0000001" when "00100001110110001", -- t[17329] = 1
      "0000001" when "00100001110110010", -- t[17330] = 1
      "0000001" when "00100001110110011", -- t[17331] = 1
      "0000001" when "00100001110110100", -- t[17332] = 1
      "0000001" when "00100001110110101", -- t[17333] = 1
      "0000001" when "00100001110110110", -- t[17334] = 1
      "0000001" when "00100001110110111", -- t[17335] = 1
      "0000001" when "00100001110111000", -- t[17336] = 1
      "0000001" when "00100001110111001", -- t[17337] = 1
      "0000001" when "00100001110111010", -- t[17338] = 1
      "0000001" when "00100001110111011", -- t[17339] = 1
      "0000001" when "00100001110111100", -- t[17340] = 1
      "0000001" when "00100001110111101", -- t[17341] = 1
      "0000001" when "00100001110111110", -- t[17342] = 1
      "0000001" when "00100001110111111", -- t[17343] = 1
      "0000001" when "00100001111000000", -- t[17344] = 1
      "0000001" when "00100001111000001", -- t[17345] = 1
      "0000001" when "00100001111000010", -- t[17346] = 1
      "0000001" when "00100001111000011", -- t[17347] = 1
      "0000001" when "00100001111000100", -- t[17348] = 1
      "0000001" when "00100001111000101", -- t[17349] = 1
      "0000001" when "00100001111000110", -- t[17350] = 1
      "0000001" when "00100001111000111", -- t[17351] = 1
      "0000001" when "00100001111001000", -- t[17352] = 1
      "0000001" when "00100001111001001", -- t[17353] = 1
      "0000001" when "00100001111001010", -- t[17354] = 1
      "0000001" when "00100001111001011", -- t[17355] = 1
      "0000001" when "00100001111001100", -- t[17356] = 1
      "0000001" when "00100001111001101", -- t[17357] = 1
      "0000001" when "00100001111001110", -- t[17358] = 1
      "0000001" when "00100001111001111", -- t[17359] = 1
      "0000001" when "00100001111010000", -- t[17360] = 1
      "0000001" when "00100001111010001", -- t[17361] = 1
      "0000001" when "00100001111010010", -- t[17362] = 1
      "0000001" when "00100001111010011", -- t[17363] = 1
      "0000001" when "00100001111010100", -- t[17364] = 1
      "0000001" when "00100001111010101", -- t[17365] = 1
      "0000001" when "00100001111010110", -- t[17366] = 1
      "0000001" when "00100001111010111", -- t[17367] = 1
      "0000001" when "00100001111011000", -- t[17368] = 1
      "0000001" when "00100001111011001", -- t[17369] = 1
      "0000001" when "00100001111011010", -- t[17370] = 1
      "0000001" when "00100001111011011", -- t[17371] = 1
      "0000001" when "00100001111011100", -- t[17372] = 1
      "0000001" when "00100001111011101", -- t[17373] = 1
      "0000001" when "00100001111011110", -- t[17374] = 1
      "0000001" when "00100001111011111", -- t[17375] = 1
      "0000001" when "00100001111100000", -- t[17376] = 1
      "0000001" when "00100001111100001", -- t[17377] = 1
      "0000001" when "00100001111100010", -- t[17378] = 1
      "0000001" when "00100001111100011", -- t[17379] = 1
      "0000001" when "00100001111100100", -- t[17380] = 1
      "0000001" when "00100001111100101", -- t[17381] = 1
      "0000001" when "00100001111100110", -- t[17382] = 1
      "0000001" when "00100001111100111", -- t[17383] = 1
      "0000001" when "00100001111101000", -- t[17384] = 1
      "0000001" when "00100001111101001", -- t[17385] = 1
      "0000001" when "00100001111101010", -- t[17386] = 1
      "0000001" when "00100001111101011", -- t[17387] = 1
      "0000001" when "00100001111101100", -- t[17388] = 1
      "0000001" when "00100001111101101", -- t[17389] = 1
      "0000001" when "00100001111101110", -- t[17390] = 1
      "0000001" when "00100001111101111", -- t[17391] = 1
      "0000001" when "00100001111110000", -- t[17392] = 1
      "0000001" when "00100001111110001", -- t[17393] = 1
      "0000001" when "00100001111110010", -- t[17394] = 1
      "0000001" when "00100001111110011", -- t[17395] = 1
      "0000001" when "00100001111110100", -- t[17396] = 1
      "0000001" when "00100001111110101", -- t[17397] = 1
      "0000001" when "00100001111110110", -- t[17398] = 1
      "0000001" when "00100001111110111", -- t[17399] = 1
      "0000001" when "00100001111111000", -- t[17400] = 1
      "0000001" when "00100001111111001", -- t[17401] = 1
      "0000001" when "00100001111111010", -- t[17402] = 1
      "0000001" when "00100001111111011", -- t[17403] = 1
      "0000001" when "00100001111111100", -- t[17404] = 1
      "0000001" when "00100001111111101", -- t[17405] = 1
      "0000001" when "00100001111111110", -- t[17406] = 1
      "0000001" when "00100001111111111", -- t[17407] = 1
      "0000001" when "00100010000000000", -- t[17408] = 1
      "0000001" when "00100010000000001", -- t[17409] = 1
      "0000001" when "00100010000000010", -- t[17410] = 1
      "0000001" when "00100010000000011", -- t[17411] = 1
      "0000001" when "00100010000000100", -- t[17412] = 1
      "0000001" when "00100010000000101", -- t[17413] = 1
      "0000001" when "00100010000000110", -- t[17414] = 1
      "0000001" when "00100010000000111", -- t[17415] = 1
      "0000001" when "00100010000001000", -- t[17416] = 1
      "0000001" when "00100010000001001", -- t[17417] = 1
      "0000001" when "00100010000001010", -- t[17418] = 1
      "0000001" when "00100010000001011", -- t[17419] = 1
      "0000001" when "00100010000001100", -- t[17420] = 1
      "0000001" when "00100010000001101", -- t[17421] = 1
      "0000001" when "00100010000001110", -- t[17422] = 1
      "0000001" when "00100010000001111", -- t[17423] = 1
      "0000001" when "00100010000010000", -- t[17424] = 1
      "0000001" when "00100010000010001", -- t[17425] = 1
      "0000001" when "00100010000010010", -- t[17426] = 1
      "0000001" when "00100010000010011", -- t[17427] = 1
      "0000001" when "00100010000010100", -- t[17428] = 1
      "0000001" when "00100010000010101", -- t[17429] = 1
      "0000001" when "00100010000010110", -- t[17430] = 1
      "0000001" when "00100010000010111", -- t[17431] = 1
      "0000001" when "00100010000011000", -- t[17432] = 1
      "0000001" when "00100010000011001", -- t[17433] = 1
      "0000001" when "00100010000011010", -- t[17434] = 1
      "0000001" when "00100010000011011", -- t[17435] = 1
      "0000001" when "00100010000011100", -- t[17436] = 1
      "0000001" when "00100010000011101", -- t[17437] = 1
      "0000001" when "00100010000011110", -- t[17438] = 1
      "0000001" when "00100010000011111", -- t[17439] = 1
      "0000001" when "00100010000100000", -- t[17440] = 1
      "0000001" when "00100010000100001", -- t[17441] = 1
      "0000001" when "00100010000100010", -- t[17442] = 1
      "0000001" when "00100010000100011", -- t[17443] = 1
      "0000001" when "00100010000100100", -- t[17444] = 1
      "0000001" when "00100010000100101", -- t[17445] = 1
      "0000001" when "00100010000100110", -- t[17446] = 1
      "0000001" when "00100010000100111", -- t[17447] = 1
      "0000001" when "00100010000101000", -- t[17448] = 1
      "0000001" when "00100010000101001", -- t[17449] = 1
      "0000001" when "00100010000101010", -- t[17450] = 1
      "0000001" when "00100010000101011", -- t[17451] = 1
      "0000001" when "00100010000101100", -- t[17452] = 1
      "0000001" when "00100010000101101", -- t[17453] = 1
      "0000001" when "00100010000101110", -- t[17454] = 1
      "0000001" when "00100010000101111", -- t[17455] = 1
      "0000001" when "00100010000110000", -- t[17456] = 1
      "0000001" when "00100010000110001", -- t[17457] = 1
      "0000001" when "00100010000110010", -- t[17458] = 1
      "0000001" when "00100010000110011", -- t[17459] = 1
      "0000001" when "00100010000110100", -- t[17460] = 1
      "0000001" when "00100010000110101", -- t[17461] = 1
      "0000001" when "00100010000110110", -- t[17462] = 1
      "0000001" when "00100010000110111", -- t[17463] = 1
      "0000001" when "00100010000111000", -- t[17464] = 1
      "0000001" when "00100010000111001", -- t[17465] = 1
      "0000001" when "00100010000111010", -- t[17466] = 1
      "0000001" when "00100010000111011", -- t[17467] = 1
      "0000001" when "00100010000111100", -- t[17468] = 1
      "0000001" when "00100010000111101", -- t[17469] = 1
      "0000001" when "00100010000111110", -- t[17470] = 1
      "0000001" when "00100010000111111", -- t[17471] = 1
      "0000001" when "00100010001000000", -- t[17472] = 1
      "0000001" when "00100010001000001", -- t[17473] = 1
      "0000001" when "00100010001000010", -- t[17474] = 1
      "0000001" when "00100010001000011", -- t[17475] = 1
      "0000001" when "00100010001000100", -- t[17476] = 1
      "0000001" when "00100010001000101", -- t[17477] = 1
      "0000001" when "00100010001000110", -- t[17478] = 1
      "0000001" when "00100010001000111", -- t[17479] = 1
      "0000001" when "00100010001001000", -- t[17480] = 1
      "0000001" when "00100010001001001", -- t[17481] = 1
      "0000001" when "00100010001001010", -- t[17482] = 1
      "0000001" when "00100010001001011", -- t[17483] = 1
      "0000001" when "00100010001001100", -- t[17484] = 1
      "0000001" when "00100010001001101", -- t[17485] = 1
      "0000001" when "00100010001001110", -- t[17486] = 1
      "0000001" when "00100010001001111", -- t[17487] = 1
      "0000001" when "00100010001010000", -- t[17488] = 1
      "0000001" when "00100010001010001", -- t[17489] = 1
      "0000001" when "00100010001010010", -- t[17490] = 1
      "0000001" when "00100010001010011", -- t[17491] = 1
      "0000001" when "00100010001010100", -- t[17492] = 1
      "0000001" when "00100010001010101", -- t[17493] = 1
      "0000001" when "00100010001010110", -- t[17494] = 1
      "0000001" when "00100010001010111", -- t[17495] = 1
      "0000001" when "00100010001011000", -- t[17496] = 1
      "0000001" when "00100010001011001", -- t[17497] = 1
      "0000001" when "00100010001011010", -- t[17498] = 1
      "0000001" when "00100010001011011", -- t[17499] = 1
      "0000001" when "00100010001011100", -- t[17500] = 1
      "0000001" when "00100010001011101", -- t[17501] = 1
      "0000001" when "00100010001011110", -- t[17502] = 1
      "0000001" when "00100010001011111", -- t[17503] = 1
      "0000001" when "00100010001100000", -- t[17504] = 1
      "0000001" when "00100010001100001", -- t[17505] = 1
      "0000001" when "00100010001100010", -- t[17506] = 1
      "0000001" when "00100010001100011", -- t[17507] = 1
      "0000001" when "00100010001100100", -- t[17508] = 1
      "0000001" when "00100010001100101", -- t[17509] = 1
      "0000001" when "00100010001100110", -- t[17510] = 1
      "0000001" when "00100010001100111", -- t[17511] = 1
      "0000001" when "00100010001101000", -- t[17512] = 1
      "0000001" when "00100010001101001", -- t[17513] = 1
      "0000001" when "00100010001101010", -- t[17514] = 1
      "0000001" when "00100010001101011", -- t[17515] = 1
      "0000001" when "00100010001101100", -- t[17516] = 1
      "0000001" when "00100010001101101", -- t[17517] = 1
      "0000001" when "00100010001101110", -- t[17518] = 1
      "0000001" when "00100010001101111", -- t[17519] = 1
      "0000001" when "00100010001110000", -- t[17520] = 1
      "0000001" when "00100010001110001", -- t[17521] = 1
      "0000001" when "00100010001110010", -- t[17522] = 1
      "0000001" when "00100010001110011", -- t[17523] = 1
      "0000001" when "00100010001110100", -- t[17524] = 1
      "0000001" when "00100010001110101", -- t[17525] = 1
      "0000001" when "00100010001110110", -- t[17526] = 1
      "0000001" when "00100010001110111", -- t[17527] = 1
      "0000001" when "00100010001111000", -- t[17528] = 1
      "0000001" when "00100010001111001", -- t[17529] = 1
      "0000001" when "00100010001111010", -- t[17530] = 1
      "0000001" when "00100010001111011", -- t[17531] = 1
      "0000001" when "00100010001111100", -- t[17532] = 1
      "0000001" when "00100010001111101", -- t[17533] = 1
      "0000001" when "00100010001111110", -- t[17534] = 1
      "0000001" when "00100010001111111", -- t[17535] = 1
      "0000001" when "00100010010000000", -- t[17536] = 1
      "0000001" when "00100010010000001", -- t[17537] = 1
      "0000001" when "00100010010000010", -- t[17538] = 1
      "0000001" when "00100010010000011", -- t[17539] = 1
      "0000001" when "00100010010000100", -- t[17540] = 1
      "0000001" when "00100010010000101", -- t[17541] = 1
      "0000001" when "00100010010000110", -- t[17542] = 1
      "0000001" when "00100010010000111", -- t[17543] = 1
      "0000001" when "00100010010001000", -- t[17544] = 1
      "0000001" when "00100010010001001", -- t[17545] = 1
      "0000001" when "00100010010001010", -- t[17546] = 1
      "0000001" when "00100010010001011", -- t[17547] = 1
      "0000001" when "00100010010001100", -- t[17548] = 1
      "0000001" when "00100010010001101", -- t[17549] = 1
      "0000001" when "00100010010001110", -- t[17550] = 1
      "0000001" when "00100010010001111", -- t[17551] = 1
      "0000001" when "00100010010010000", -- t[17552] = 1
      "0000001" when "00100010010010001", -- t[17553] = 1
      "0000001" when "00100010010010010", -- t[17554] = 1
      "0000001" when "00100010010010011", -- t[17555] = 1
      "0000001" when "00100010010010100", -- t[17556] = 1
      "0000001" when "00100010010010101", -- t[17557] = 1
      "0000001" when "00100010010010110", -- t[17558] = 1
      "0000001" when "00100010010010111", -- t[17559] = 1
      "0000001" when "00100010010011000", -- t[17560] = 1
      "0000001" when "00100010010011001", -- t[17561] = 1
      "0000001" when "00100010010011010", -- t[17562] = 1
      "0000001" when "00100010010011011", -- t[17563] = 1
      "0000001" when "00100010010011100", -- t[17564] = 1
      "0000001" when "00100010010011101", -- t[17565] = 1
      "0000001" when "00100010010011110", -- t[17566] = 1
      "0000001" when "00100010010011111", -- t[17567] = 1
      "0000001" when "00100010010100000", -- t[17568] = 1
      "0000001" when "00100010010100001", -- t[17569] = 1
      "0000001" when "00100010010100010", -- t[17570] = 1
      "0000001" when "00100010010100011", -- t[17571] = 1
      "0000001" when "00100010010100100", -- t[17572] = 1
      "0000001" when "00100010010100101", -- t[17573] = 1
      "0000001" when "00100010010100110", -- t[17574] = 1
      "0000001" when "00100010010100111", -- t[17575] = 1
      "0000001" when "00100010010101000", -- t[17576] = 1
      "0000001" when "00100010010101001", -- t[17577] = 1
      "0000001" when "00100010010101010", -- t[17578] = 1
      "0000001" when "00100010010101011", -- t[17579] = 1
      "0000001" when "00100010010101100", -- t[17580] = 1
      "0000001" when "00100010010101101", -- t[17581] = 1
      "0000001" when "00100010010101110", -- t[17582] = 1
      "0000001" when "00100010010101111", -- t[17583] = 1
      "0000001" when "00100010010110000", -- t[17584] = 1
      "0000001" when "00100010010110001", -- t[17585] = 1
      "0000001" when "00100010010110010", -- t[17586] = 1
      "0000001" when "00100010010110011", -- t[17587] = 1
      "0000001" when "00100010010110100", -- t[17588] = 1
      "0000001" when "00100010010110101", -- t[17589] = 1
      "0000001" when "00100010010110110", -- t[17590] = 1
      "0000001" when "00100010010110111", -- t[17591] = 1
      "0000001" when "00100010010111000", -- t[17592] = 1
      "0000001" when "00100010010111001", -- t[17593] = 1
      "0000001" when "00100010010111010", -- t[17594] = 1
      "0000001" when "00100010010111011", -- t[17595] = 1
      "0000001" when "00100010010111100", -- t[17596] = 1
      "0000001" when "00100010010111101", -- t[17597] = 1
      "0000001" when "00100010010111110", -- t[17598] = 1
      "0000001" when "00100010010111111", -- t[17599] = 1
      "0000001" when "00100010011000000", -- t[17600] = 1
      "0000001" when "00100010011000001", -- t[17601] = 1
      "0000001" when "00100010011000010", -- t[17602] = 1
      "0000001" when "00100010011000011", -- t[17603] = 1
      "0000001" when "00100010011000100", -- t[17604] = 1
      "0000001" when "00100010011000101", -- t[17605] = 1
      "0000001" when "00100010011000110", -- t[17606] = 1
      "0000001" when "00100010011000111", -- t[17607] = 1
      "0000001" when "00100010011001000", -- t[17608] = 1
      "0000001" when "00100010011001001", -- t[17609] = 1
      "0000001" when "00100010011001010", -- t[17610] = 1
      "0000001" when "00100010011001011", -- t[17611] = 1
      "0000001" when "00100010011001100", -- t[17612] = 1
      "0000001" when "00100010011001101", -- t[17613] = 1
      "0000001" when "00100010011001110", -- t[17614] = 1
      "0000001" when "00100010011001111", -- t[17615] = 1
      "0000001" when "00100010011010000", -- t[17616] = 1
      "0000001" when "00100010011010001", -- t[17617] = 1
      "0000001" when "00100010011010010", -- t[17618] = 1
      "0000001" when "00100010011010011", -- t[17619] = 1
      "0000001" when "00100010011010100", -- t[17620] = 1
      "0000001" when "00100010011010101", -- t[17621] = 1
      "0000001" when "00100010011010110", -- t[17622] = 1
      "0000001" when "00100010011010111", -- t[17623] = 1
      "0000001" when "00100010011011000", -- t[17624] = 1
      "0000001" when "00100010011011001", -- t[17625] = 1
      "0000001" when "00100010011011010", -- t[17626] = 1
      "0000001" when "00100010011011011", -- t[17627] = 1
      "0000001" when "00100010011011100", -- t[17628] = 1
      "0000001" when "00100010011011101", -- t[17629] = 1
      "0000001" when "00100010011011110", -- t[17630] = 1
      "0000001" when "00100010011011111", -- t[17631] = 1
      "0000001" when "00100010011100000", -- t[17632] = 1
      "0000001" when "00100010011100001", -- t[17633] = 1
      "0000001" when "00100010011100010", -- t[17634] = 1
      "0000001" when "00100010011100011", -- t[17635] = 1
      "0000001" when "00100010011100100", -- t[17636] = 1
      "0000001" when "00100010011100101", -- t[17637] = 1
      "0000001" when "00100010011100110", -- t[17638] = 1
      "0000001" when "00100010011100111", -- t[17639] = 1
      "0000001" when "00100010011101000", -- t[17640] = 1
      "0000001" when "00100010011101001", -- t[17641] = 1
      "0000001" when "00100010011101010", -- t[17642] = 1
      "0000001" when "00100010011101011", -- t[17643] = 1
      "0000001" when "00100010011101100", -- t[17644] = 1
      "0000001" when "00100010011101101", -- t[17645] = 1
      "0000001" when "00100010011101110", -- t[17646] = 1
      "0000001" when "00100010011101111", -- t[17647] = 1
      "0000001" when "00100010011110000", -- t[17648] = 1
      "0000001" when "00100010011110001", -- t[17649] = 1
      "0000001" when "00100010011110010", -- t[17650] = 1
      "0000001" when "00100010011110011", -- t[17651] = 1
      "0000001" when "00100010011110100", -- t[17652] = 1
      "0000001" when "00100010011110101", -- t[17653] = 1
      "0000001" when "00100010011110110", -- t[17654] = 1
      "0000001" when "00100010011110111", -- t[17655] = 1
      "0000001" when "00100010011111000", -- t[17656] = 1
      "0000001" when "00100010011111001", -- t[17657] = 1
      "0000001" when "00100010011111010", -- t[17658] = 1
      "0000001" when "00100010011111011", -- t[17659] = 1
      "0000001" when "00100010011111100", -- t[17660] = 1
      "0000001" when "00100010011111101", -- t[17661] = 1
      "0000001" when "00100010011111110", -- t[17662] = 1
      "0000001" when "00100010011111111", -- t[17663] = 1
      "0000001" when "00100010100000000", -- t[17664] = 1
      "0000001" when "00100010100000001", -- t[17665] = 1
      "0000001" when "00100010100000010", -- t[17666] = 1
      "0000001" when "00100010100000011", -- t[17667] = 1
      "0000001" when "00100010100000100", -- t[17668] = 1
      "0000001" when "00100010100000101", -- t[17669] = 1
      "0000001" when "00100010100000110", -- t[17670] = 1
      "0000001" when "00100010100000111", -- t[17671] = 1
      "0000001" when "00100010100001000", -- t[17672] = 1
      "0000001" when "00100010100001001", -- t[17673] = 1
      "0000001" when "00100010100001010", -- t[17674] = 1
      "0000001" when "00100010100001011", -- t[17675] = 1
      "0000001" when "00100010100001100", -- t[17676] = 1
      "0000001" when "00100010100001101", -- t[17677] = 1
      "0000001" when "00100010100001110", -- t[17678] = 1
      "0000001" when "00100010100001111", -- t[17679] = 1
      "0000001" when "00100010100010000", -- t[17680] = 1
      "0000001" when "00100010100010001", -- t[17681] = 1
      "0000001" when "00100010100010010", -- t[17682] = 1
      "0000001" when "00100010100010011", -- t[17683] = 1
      "0000001" when "00100010100010100", -- t[17684] = 1
      "0000001" when "00100010100010101", -- t[17685] = 1
      "0000001" when "00100010100010110", -- t[17686] = 1
      "0000001" when "00100010100010111", -- t[17687] = 1
      "0000001" when "00100010100011000", -- t[17688] = 1
      "0000001" when "00100010100011001", -- t[17689] = 1
      "0000001" when "00100010100011010", -- t[17690] = 1
      "0000001" when "00100010100011011", -- t[17691] = 1
      "0000001" when "00100010100011100", -- t[17692] = 1
      "0000001" when "00100010100011101", -- t[17693] = 1
      "0000001" when "00100010100011110", -- t[17694] = 1
      "0000001" when "00100010100011111", -- t[17695] = 1
      "0000001" when "00100010100100000", -- t[17696] = 1
      "0000001" when "00100010100100001", -- t[17697] = 1
      "0000001" when "00100010100100010", -- t[17698] = 1
      "0000001" when "00100010100100011", -- t[17699] = 1
      "0000001" when "00100010100100100", -- t[17700] = 1
      "0000001" when "00100010100100101", -- t[17701] = 1
      "0000001" when "00100010100100110", -- t[17702] = 1
      "0000001" when "00100010100100111", -- t[17703] = 1
      "0000001" when "00100010100101000", -- t[17704] = 1
      "0000001" when "00100010100101001", -- t[17705] = 1
      "0000001" when "00100010100101010", -- t[17706] = 1
      "0000001" when "00100010100101011", -- t[17707] = 1
      "0000001" when "00100010100101100", -- t[17708] = 1
      "0000001" when "00100010100101101", -- t[17709] = 1
      "0000001" when "00100010100101110", -- t[17710] = 1
      "0000001" when "00100010100101111", -- t[17711] = 1
      "0000001" when "00100010100110000", -- t[17712] = 1
      "0000001" when "00100010100110001", -- t[17713] = 1
      "0000001" when "00100010100110010", -- t[17714] = 1
      "0000001" when "00100010100110011", -- t[17715] = 1
      "0000001" when "00100010100110100", -- t[17716] = 1
      "0000001" when "00100010100110101", -- t[17717] = 1
      "0000001" when "00100010100110110", -- t[17718] = 1
      "0000001" when "00100010100110111", -- t[17719] = 1
      "0000001" when "00100010100111000", -- t[17720] = 1
      "0000001" when "00100010100111001", -- t[17721] = 1
      "0000001" when "00100010100111010", -- t[17722] = 1
      "0000001" when "00100010100111011", -- t[17723] = 1
      "0000001" when "00100010100111100", -- t[17724] = 1
      "0000001" when "00100010100111101", -- t[17725] = 1
      "0000001" when "00100010100111110", -- t[17726] = 1
      "0000001" when "00100010100111111", -- t[17727] = 1
      "0000001" when "00100010101000000", -- t[17728] = 1
      "0000001" when "00100010101000001", -- t[17729] = 1
      "0000001" when "00100010101000010", -- t[17730] = 1
      "0000001" when "00100010101000011", -- t[17731] = 1
      "0000001" when "00100010101000100", -- t[17732] = 1
      "0000001" when "00100010101000101", -- t[17733] = 1
      "0000001" when "00100010101000110", -- t[17734] = 1
      "0000001" when "00100010101000111", -- t[17735] = 1
      "0000001" when "00100010101001000", -- t[17736] = 1
      "0000001" when "00100010101001001", -- t[17737] = 1
      "0000001" when "00100010101001010", -- t[17738] = 1
      "0000001" when "00100010101001011", -- t[17739] = 1
      "0000001" when "00100010101001100", -- t[17740] = 1
      "0000001" when "00100010101001101", -- t[17741] = 1
      "0000001" when "00100010101001110", -- t[17742] = 1
      "0000001" when "00100010101001111", -- t[17743] = 1
      "0000001" when "00100010101010000", -- t[17744] = 1
      "0000001" when "00100010101010001", -- t[17745] = 1
      "0000001" when "00100010101010010", -- t[17746] = 1
      "0000001" when "00100010101010011", -- t[17747] = 1
      "0000001" when "00100010101010100", -- t[17748] = 1
      "0000001" when "00100010101010101", -- t[17749] = 1
      "0000001" when "00100010101010110", -- t[17750] = 1
      "0000001" when "00100010101010111", -- t[17751] = 1
      "0000001" when "00100010101011000", -- t[17752] = 1
      "0000001" when "00100010101011001", -- t[17753] = 1
      "0000001" when "00100010101011010", -- t[17754] = 1
      "0000001" when "00100010101011011", -- t[17755] = 1
      "0000001" when "00100010101011100", -- t[17756] = 1
      "0000001" when "00100010101011101", -- t[17757] = 1
      "0000001" when "00100010101011110", -- t[17758] = 1
      "0000001" when "00100010101011111", -- t[17759] = 1
      "0000001" when "00100010101100000", -- t[17760] = 1
      "0000001" when "00100010101100001", -- t[17761] = 1
      "0000001" when "00100010101100010", -- t[17762] = 1
      "0000001" when "00100010101100011", -- t[17763] = 1
      "0000001" when "00100010101100100", -- t[17764] = 1
      "0000001" when "00100010101100101", -- t[17765] = 1
      "0000001" when "00100010101100110", -- t[17766] = 1
      "0000001" when "00100010101100111", -- t[17767] = 1
      "0000001" when "00100010101101000", -- t[17768] = 1
      "0000001" when "00100010101101001", -- t[17769] = 1
      "0000001" when "00100010101101010", -- t[17770] = 1
      "0000001" when "00100010101101011", -- t[17771] = 1
      "0000001" when "00100010101101100", -- t[17772] = 1
      "0000001" when "00100010101101101", -- t[17773] = 1
      "0000001" when "00100010101101110", -- t[17774] = 1
      "0000001" when "00100010101101111", -- t[17775] = 1
      "0000001" when "00100010101110000", -- t[17776] = 1
      "0000001" when "00100010101110001", -- t[17777] = 1
      "0000001" when "00100010101110010", -- t[17778] = 1
      "0000001" when "00100010101110011", -- t[17779] = 1
      "0000001" when "00100010101110100", -- t[17780] = 1
      "0000001" when "00100010101110101", -- t[17781] = 1
      "0000001" when "00100010101110110", -- t[17782] = 1
      "0000001" when "00100010101110111", -- t[17783] = 1
      "0000001" when "00100010101111000", -- t[17784] = 1
      "0000001" when "00100010101111001", -- t[17785] = 1
      "0000001" when "00100010101111010", -- t[17786] = 1
      "0000001" when "00100010101111011", -- t[17787] = 1
      "0000001" when "00100010101111100", -- t[17788] = 1
      "0000001" when "00100010101111101", -- t[17789] = 1
      "0000001" when "00100010101111110", -- t[17790] = 1
      "0000001" when "00100010101111111", -- t[17791] = 1
      "0000001" when "00100010110000000", -- t[17792] = 1
      "0000001" when "00100010110000001", -- t[17793] = 1
      "0000001" when "00100010110000010", -- t[17794] = 1
      "0000001" when "00100010110000011", -- t[17795] = 1
      "0000001" when "00100010110000100", -- t[17796] = 1
      "0000001" when "00100010110000101", -- t[17797] = 1
      "0000001" when "00100010110000110", -- t[17798] = 1
      "0000001" when "00100010110000111", -- t[17799] = 1
      "0000001" when "00100010110001000", -- t[17800] = 1
      "0000001" when "00100010110001001", -- t[17801] = 1
      "0000001" when "00100010110001010", -- t[17802] = 1
      "0000001" when "00100010110001011", -- t[17803] = 1
      "0000001" when "00100010110001100", -- t[17804] = 1
      "0000001" when "00100010110001101", -- t[17805] = 1
      "0000001" when "00100010110001110", -- t[17806] = 1
      "0000001" when "00100010110001111", -- t[17807] = 1
      "0000001" when "00100010110010000", -- t[17808] = 1
      "0000001" when "00100010110010001", -- t[17809] = 1
      "0000001" when "00100010110010010", -- t[17810] = 1
      "0000001" when "00100010110010011", -- t[17811] = 1
      "0000001" when "00100010110010100", -- t[17812] = 1
      "0000001" when "00100010110010101", -- t[17813] = 1
      "0000001" when "00100010110010110", -- t[17814] = 1
      "0000001" when "00100010110010111", -- t[17815] = 1
      "0000001" when "00100010110011000", -- t[17816] = 1
      "0000001" when "00100010110011001", -- t[17817] = 1
      "0000001" when "00100010110011010", -- t[17818] = 1
      "0000001" when "00100010110011011", -- t[17819] = 1
      "0000001" when "00100010110011100", -- t[17820] = 1
      "0000001" when "00100010110011101", -- t[17821] = 1
      "0000001" when "00100010110011110", -- t[17822] = 1
      "0000001" when "00100010110011111", -- t[17823] = 1
      "0000001" when "00100010110100000", -- t[17824] = 1
      "0000001" when "00100010110100001", -- t[17825] = 1
      "0000001" when "00100010110100010", -- t[17826] = 1
      "0000001" when "00100010110100011", -- t[17827] = 1
      "0000001" when "00100010110100100", -- t[17828] = 1
      "0000001" when "00100010110100101", -- t[17829] = 1
      "0000001" when "00100010110100110", -- t[17830] = 1
      "0000001" when "00100010110100111", -- t[17831] = 1
      "0000001" when "00100010110101000", -- t[17832] = 1
      "0000001" when "00100010110101001", -- t[17833] = 1
      "0000001" when "00100010110101010", -- t[17834] = 1
      "0000001" when "00100010110101011", -- t[17835] = 1
      "0000001" when "00100010110101100", -- t[17836] = 1
      "0000001" when "00100010110101101", -- t[17837] = 1
      "0000001" when "00100010110101110", -- t[17838] = 1
      "0000001" when "00100010110101111", -- t[17839] = 1
      "0000001" when "00100010110110000", -- t[17840] = 1
      "0000001" when "00100010110110001", -- t[17841] = 1
      "0000001" when "00100010110110010", -- t[17842] = 1
      "0000001" when "00100010110110011", -- t[17843] = 1
      "0000001" when "00100010110110100", -- t[17844] = 1
      "0000001" when "00100010110110101", -- t[17845] = 1
      "0000001" when "00100010110110110", -- t[17846] = 1
      "0000001" when "00100010110110111", -- t[17847] = 1
      "0000001" when "00100010110111000", -- t[17848] = 1
      "0000001" when "00100010110111001", -- t[17849] = 1
      "0000001" when "00100010110111010", -- t[17850] = 1
      "0000001" when "00100010110111011", -- t[17851] = 1
      "0000001" when "00100010110111100", -- t[17852] = 1
      "0000001" when "00100010110111101", -- t[17853] = 1
      "0000001" when "00100010110111110", -- t[17854] = 1
      "0000001" when "00100010110111111", -- t[17855] = 1
      "0000001" when "00100010111000000", -- t[17856] = 1
      "0000001" when "00100010111000001", -- t[17857] = 1
      "0000001" when "00100010111000010", -- t[17858] = 1
      "0000001" when "00100010111000011", -- t[17859] = 1
      "0000001" when "00100010111000100", -- t[17860] = 1
      "0000001" when "00100010111000101", -- t[17861] = 1
      "0000001" when "00100010111000110", -- t[17862] = 1
      "0000001" when "00100010111000111", -- t[17863] = 1
      "0000001" when "00100010111001000", -- t[17864] = 1
      "0000001" when "00100010111001001", -- t[17865] = 1
      "0000001" when "00100010111001010", -- t[17866] = 1
      "0000001" when "00100010111001011", -- t[17867] = 1
      "0000001" when "00100010111001100", -- t[17868] = 1
      "0000001" when "00100010111001101", -- t[17869] = 1
      "0000001" when "00100010111001110", -- t[17870] = 1
      "0000001" when "00100010111001111", -- t[17871] = 1
      "0000001" when "00100010111010000", -- t[17872] = 1
      "0000001" when "00100010111010001", -- t[17873] = 1
      "0000001" when "00100010111010010", -- t[17874] = 1
      "0000001" when "00100010111010011", -- t[17875] = 1
      "0000001" when "00100010111010100", -- t[17876] = 1
      "0000001" when "00100010111010101", -- t[17877] = 1
      "0000001" when "00100010111010110", -- t[17878] = 1
      "0000001" when "00100010111010111", -- t[17879] = 1
      "0000001" when "00100010111011000", -- t[17880] = 1
      "0000001" when "00100010111011001", -- t[17881] = 1
      "0000001" when "00100010111011010", -- t[17882] = 1
      "0000001" when "00100010111011011", -- t[17883] = 1
      "0000001" when "00100010111011100", -- t[17884] = 1
      "0000001" when "00100010111011101", -- t[17885] = 1
      "0000001" when "00100010111011110", -- t[17886] = 1
      "0000001" when "00100010111011111", -- t[17887] = 1
      "0000001" when "00100010111100000", -- t[17888] = 1
      "0000001" when "00100010111100001", -- t[17889] = 1
      "0000001" when "00100010111100010", -- t[17890] = 1
      "0000001" when "00100010111100011", -- t[17891] = 1
      "0000001" when "00100010111100100", -- t[17892] = 1
      "0000001" when "00100010111100101", -- t[17893] = 1
      "0000001" when "00100010111100110", -- t[17894] = 1
      "0000001" when "00100010111100111", -- t[17895] = 1
      "0000001" when "00100010111101000", -- t[17896] = 1
      "0000001" when "00100010111101001", -- t[17897] = 1
      "0000001" when "00100010111101010", -- t[17898] = 1
      "0000001" when "00100010111101011", -- t[17899] = 1
      "0000001" when "00100010111101100", -- t[17900] = 1
      "0000001" when "00100010111101101", -- t[17901] = 1
      "0000001" when "00100010111101110", -- t[17902] = 1
      "0000001" when "00100010111101111", -- t[17903] = 1
      "0000001" when "00100010111110000", -- t[17904] = 1
      "0000001" when "00100010111110001", -- t[17905] = 1
      "0000001" when "00100010111110010", -- t[17906] = 1
      "0000001" when "00100010111110011", -- t[17907] = 1
      "0000001" when "00100010111110100", -- t[17908] = 1
      "0000001" when "00100010111110101", -- t[17909] = 1
      "0000001" when "00100010111110110", -- t[17910] = 1
      "0000001" when "00100010111110111", -- t[17911] = 1
      "0000001" when "00100010111111000", -- t[17912] = 1
      "0000001" when "00100010111111001", -- t[17913] = 1
      "0000001" when "00100010111111010", -- t[17914] = 1
      "0000001" when "00100010111111011", -- t[17915] = 1
      "0000001" when "00100010111111100", -- t[17916] = 1
      "0000001" when "00100010111111101", -- t[17917] = 1
      "0000001" when "00100010111111110", -- t[17918] = 1
      "0000001" when "00100010111111111", -- t[17919] = 1
      "0000001" when "00100011000000000", -- t[17920] = 1
      "0000001" when "00100011000000001", -- t[17921] = 1
      "0000001" when "00100011000000010", -- t[17922] = 1
      "0000001" when "00100011000000011", -- t[17923] = 1
      "0000001" when "00100011000000100", -- t[17924] = 1
      "0000001" when "00100011000000101", -- t[17925] = 1
      "0000001" when "00100011000000110", -- t[17926] = 1
      "0000001" when "00100011000000111", -- t[17927] = 1
      "0000001" when "00100011000001000", -- t[17928] = 1
      "0000001" when "00100011000001001", -- t[17929] = 1
      "0000001" when "00100011000001010", -- t[17930] = 1
      "0000001" when "00100011000001011", -- t[17931] = 1
      "0000001" when "00100011000001100", -- t[17932] = 1
      "0000001" when "00100011000001101", -- t[17933] = 1
      "0000001" when "00100011000001110", -- t[17934] = 1
      "0000001" when "00100011000001111", -- t[17935] = 1
      "0000001" when "00100011000010000", -- t[17936] = 1
      "0000001" when "00100011000010001", -- t[17937] = 1
      "0000001" when "00100011000010010", -- t[17938] = 1
      "0000001" when "00100011000010011", -- t[17939] = 1
      "0000001" when "00100011000010100", -- t[17940] = 1
      "0000001" when "00100011000010101", -- t[17941] = 1
      "0000001" when "00100011000010110", -- t[17942] = 1
      "0000001" when "00100011000010111", -- t[17943] = 1
      "0000001" when "00100011000011000", -- t[17944] = 1
      "0000001" when "00100011000011001", -- t[17945] = 1
      "0000001" when "00100011000011010", -- t[17946] = 1
      "0000001" when "00100011000011011", -- t[17947] = 1
      "0000001" when "00100011000011100", -- t[17948] = 1
      "0000001" when "00100011000011101", -- t[17949] = 1
      "0000001" when "00100011000011110", -- t[17950] = 1
      "0000001" when "00100011000011111", -- t[17951] = 1
      "0000001" when "00100011000100000", -- t[17952] = 1
      "0000001" when "00100011000100001", -- t[17953] = 1
      "0000001" when "00100011000100010", -- t[17954] = 1
      "0000001" when "00100011000100011", -- t[17955] = 1
      "0000001" when "00100011000100100", -- t[17956] = 1
      "0000001" when "00100011000100101", -- t[17957] = 1
      "0000001" when "00100011000100110", -- t[17958] = 1
      "0000001" when "00100011000100111", -- t[17959] = 1
      "0000001" when "00100011000101000", -- t[17960] = 1
      "0000001" when "00100011000101001", -- t[17961] = 1
      "0000001" when "00100011000101010", -- t[17962] = 1
      "0000001" when "00100011000101011", -- t[17963] = 1
      "0000001" when "00100011000101100", -- t[17964] = 1
      "0000001" when "00100011000101101", -- t[17965] = 1
      "0000001" when "00100011000101110", -- t[17966] = 1
      "0000001" when "00100011000101111", -- t[17967] = 1
      "0000001" when "00100011000110000", -- t[17968] = 1
      "0000001" when "00100011000110001", -- t[17969] = 1
      "0000001" when "00100011000110010", -- t[17970] = 1
      "0000001" when "00100011000110011", -- t[17971] = 1
      "0000001" when "00100011000110100", -- t[17972] = 1
      "0000001" when "00100011000110101", -- t[17973] = 1
      "0000001" when "00100011000110110", -- t[17974] = 1
      "0000001" when "00100011000110111", -- t[17975] = 1
      "0000001" when "00100011000111000", -- t[17976] = 1
      "0000001" when "00100011000111001", -- t[17977] = 1
      "0000001" when "00100011000111010", -- t[17978] = 1
      "0000001" when "00100011000111011", -- t[17979] = 1
      "0000001" when "00100011000111100", -- t[17980] = 1
      "0000001" when "00100011000111101", -- t[17981] = 1
      "0000001" when "00100011000111110", -- t[17982] = 1
      "0000001" when "00100011000111111", -- t[17983] = 1
      "0000001" when "00100011001000000", -- t[17984] = 1
      "0000001" when "00100011001000001", -- t[17985] = 1
      "0000001" when "00100011001000010", -- t[17986] = 1
      "0000001" when "00100011001000011", -- t[17987] = 1
      "0000001" when "00100011001000100", -- t[17988] = 1
      "0000001" when "00100011001000101", -- t[17989] = 1
      "0000001" when "00100011001000110", -- t[17990] = 1
      "0000001" when "00100011001000111", -- t[17991] = 1
      "0000001" when "00100011001001000", -- t[17992] = 1
      "0000001" when "00100011001001001", -- t[17993] = 1
      "0000001" when "00100011001001010", -- t[17994] = 1
      "0000001" when "00100011001001011", -- t[17995] = 1
      "0000001" when "00100011001001100", -- t[17996] = 1
      "0000001" when "00100011001001101", -- t[17997] = 1
      "0000001" when "00100011001001110", -- t[17998] = 1
      "0000001" when "00100011001001111", -- t[17999] = 1
      "0000001" when "00100011001010000", -- t[18000] = 1
      "0000001" when "00100011001010001", -- t[18001] = 1
      "0000001" when "00100011001010010", -- t[18002] = 1
      "0000001" when "00100011001010011", -- t[18003] = 1
      "0000001" when "00100011001010100", -- t[18004] = 1
      "0000001" when "00100011001010101", -- t[18005] = 1
      "0000001" when "00100011001010110", -- t[18006] = 1
      "0000001" when "00100011001010111", -- t[18007] = 1
      "0000001" when "00100011001011000", -- t[18008] = 1
      "0000001" when "00100011001011001", -- t[18009] = 1
      "0000001" when "00100011001011010", -- t[18010] = 1
      "0000001" when "00100011001011011", -- t[18011] = 1
      "0000001" when "00100011001011100", -- t[18012] = 1
      "0000001" when "00100011001011101", -- t[18013] = 1
      "0000001" when "00100011001011110", -- t[18014] = 1
      "0000001" when "00100011001011111", -- t[18015] = 1
      "0000001" when "00100011001100000", -- t[18016] = 1
      "0000001" when "00100011001100001", -- t[18017] = 1
      "0000001" when "00100011001100010", -- t[18018] = 1
      "0000001" when "00100011001100011", -- t[18019] = 1
      "0000001" when "00100011001100100", -- t[18020] = 1
      "0000001" when "00100011001100101", -- t[18021] = 1
      "0000001" when "00100011001100110", -- t[18022] = 1
      "0000001" when "00100011001100111", -- t[18023] = 1
      "0000001" when "00100011001101000", -- t[18024] = 1
      "0000001" when "00100011001101001", -- t[18025] = 1
      "0000001" when "00100011001101010", -- t[18026] = 1
      "0000001" when "00100011001101011", -- t[18027] = 1
      "0000001" when "00100011001101100", -- t[18028] = 1
      "0000001" when "00100011001101101", -- t[18029] = 1
      "0000001" when "00100011001101110", -- t[18030] = 1
      "0000001" when "00100011001101111", -- t[18031] = 1
      "0000001" when "00100011001110000", -- t[18032] = 1
      "0000001" when "00100011001110001", -- t[18033] = 1
      "0000001" when "00100011001110010", -- t[18034] = 1
      "0000001" when "00100011001110011", -- t[18035] = 1
      "0000001" when "00100011001110100", -- t[18036] = 1
      "0000001" when "00100011001110101", -- t[18037] = 1
      "0000001" when "00100011001110110", -- t[18038] = 1
      "0000001" when "00100011001110111", -- t[18039] = 1
      "0000001" when "00100011001111000", -- t[18040] = 1
      "0000001" when "00100011001111001", -- t[18041] = 1
      "0000001" when "00100011001111010", -- t[18042] = 1
      "0000001" when "00100011001111011", -- t[18043] = 1
      "0000001" when "00100011001111100", -- t[18044] = 1
      "0000001" when "00100011001111101", -- t[18045] = 1
      "0000001" when "00100011001111110", -- t[18046] = 1
      "0000001" when "00100011001111111", -- t[18047] = 1
      "0000001" when "00100011010000000", -- t[18048] = 1
      "0000001" when "00100011010000001", -- t[18049] = 1
      "0000001" when "00100011010000010", -- t[18050] = 1
      "0000001" when "00100011010000011", -- t[18051] = 1
      "0000001" when "00100011010000100", -- t[18052] = 1
      "0000001" when "00100011010000101", -- t[18053] = 1
      "0000001" when "00100011010000110", -- t[18054] = 1
      "0000001" when "00100011010000111", -- t[18055] = 1
      "0000001" when "00100011010001000", -- t[18056] = 1
      "0000001" when "00100011010001001", -- t[18057] = 1
      "0000001" when "00100011010001010", -- t[18058] = 1
      "0000001" when "00100011010001011", -- t[18059] = 1
      "0000001" when "00100011010001100", -- t[18060] = 1
      "0000001" when "00100011010001101", -- t[18061] = 1
      "0000001" when "00100011010001110", -- t[18062] = 1
      "0000001" when "00100011010001111", -- t[18063] = 1
      "0000001" when "00100011010010000", -- t[18064] = 1
      "0000001" when "00100011010010001", -- t[18065] = 1
      "0000001" when "00100011010010010", -- t[18066] = 1
      "0000001" when "00100011010010011", -- t[18067] = 1
      "0000001" when "00100011010010100", -- t[18068] = 1
      "0000001" when "00100011010010101", -- t[18069] = 1
      "0000001" when "00100011010010110", -- t[18070] = 1
      "0000001" when "00100011010010111", -- t[18071] = 1
      "0000001" when "00100011010011000", -- t[18072] = 1
      "0000001" when "00100011010011001", -- t[18073] = 1
      "0000001" when "00100011010011010", -- t[18074] = 1
      "0000001" when "00100011010011011", -- t[18075] = 1
      "0000001" when "00100011010011100", -- t[18076] = 1
      "0000001" when "00100011010011101", -- t[18077] = 1
      "0000001" when "00100011010011110", -- t[18078] = 1
      "0000001" when "00100011010011111", -- t[18079] = 1
      "0000001" when "00100011010100000", -- t[18080] = 1
      "0000001" when "00100011010100001", -- t[18081] = 1
      "0000001" when "00100011010100010", -- t[18082] = 1
      "0000001" when "00100011010100011", -- t[18083] = 1
      "0000001" when "00100011010100100", -- t[18084] = 1
      "0000001" when "00100011010100101", -- t[18085] = 1
      "0000001" when "00100011010100110", -- t[18086] = 1
      "0000001" when "00100011010100111", -- t[18087] = 1
      "0000001" when "00100011010101000", -- t[18088] = 1
      "0000001" when "00100011010101001", -- t[18089] = 1
      "0000001" when "00100011010101010", -- t[18090] = 1
      "0000001" when "00100011010101011", -- t[18091] = 1
      "0000001" when "00100011010101100", -- t[18092] = 1
      "0000001" when "00100011010101101", -- t[18093] = 1
      "0000001" when "00100011010101110", -- t[18094] = 1
      "0000001" when "00100011010101111", -- t[18095] = 1
      "0000001" when "00100011010110000", -- t[18096] = 1
      "0000001" when "00100011010110001", -- t[18097] = 1
      "0000001" when "00100011010110010", -- t[18098] = 1
      "0000001" when "00100011010110011", -- t[18099] = 1
      "0000001" when "00100011010110100", -- t[18100] = 1
      "0000001" when "00100011010110101", -- t[18101] = 1
      "0000001" when "00100011010110110", -- t[18102] = 1
      "0000001" when "00100011010110111", -- t[18103] = 1
      "0000001" when "00100011010111000", -- t[18104] = 1
      "0000001" when "00100011010111001", -- t[18105] = 1
      "0000001" when "00100011010111010", -- t[18106] = 1
      "0000001" when "00100011010111011", -- t[18107] = 1
      "0000001" when "00100011010111100", -- t[18108] = 1
      "0000001" when "00100011010111101", -- t[18109] = 1
      "0000001" when "00100011010111110", -- t[18110] = 1
      "0000001" when "00100011010111111", -- t[18111] = 1
      "0000001" when "00100011011000000", -- t[18112] = 1
      "0000001" when "00100011011000001", -- t[18113] = 1
      "0000001" when "00100011011000010", -- t[18114] = 1
      "0000001" when "00100011011000011", -- t[18115] = 1
      "0000001" when "00100011011000100", -- t[18116] = 1
      "0000001" when "00100011011000101", -- t[18117] = 1
      "0000001" when "00100011011000110", -- t[18118] = 1
      "0000001" when "00100011011000111", -- t[18119] = 1
      "0000001" when "00100011011001000", -- t[18120] = 1
      "0000001" when "00100011011001001", -- t[18121] = 1
      "0000001" when "00100011011001010", -- t[18122] = 1
      "0000001" when "00100011011001011", -- t[18123] = 1
      "0000001" when "00100011011001100", -- t[18124] = 1
      "0000001" when "00100011011001101", -- t[18125] = 1
      "0000001" when "00100011011001110", -- t[18126] = 1
      "0000001" when "00100011011001111", -- t[18127] = 1
      "0000001" when "00100011011010000", -- t[18128] = 1
      "0000001" when "00100011011010001", -- t[18129] = 1
      "0000001" when "00100011011010010", -- t[18130] = 1
      "0000001" when "00100011011010011", -- t[18131] = 1
      "0000001" when "00100011011010100", -- t[18132] = 1
      "0000001" when "00100011011010101", -- t[18133] = 1
      "0000001" when "00100011011010110", -- t[18134] = 1
      "0000001" when "00100011011010111", -- t[18135] = 1
      "0000001" when "00100011011011000", -- t[18136] = 1
      "0000001" when "00100011011011001", -- t[18137] = 1
      "0000001" when "00100011011011010", -- t[18138] = 1
      "0000001" when "00100011011011011", -- t[18139] = 1
      "0000001" when "00100011011011100", -- t[18140] = 1
      "0000001" when "00100011011011101", -- t[18141] = 1
      "0000001" when "00100011011011110", -- t[18142] = 1
      "0000001" when "00100011011011111", -- t[18143] = 1
      "0000001" when "00100011011100000", -- t[18144] = 1
      "0000001" when "00100011011100001", -- t[18145] = 1
      "0000001" when "00100011011100010", -- t[18146] = 1
      "0000001" when "00100011011100011", -- t[18147] = 1
      "0000001" when "00100011011100100", -- t[18148] = 1
      "0000001" when "00100011011100101", -- t[18149] = 1
      "0000001" when "00100011011100110", -- t[18150] = 1
      "0000001" when "00100011011100111", -- t[18151] = 1
      "0000001" when "00100011011101000", -- t[18152] = 1
      "0000001" when "00100011011101001", -- t[18153] = 1
      "0000001" when "00100011011101010", -- t[18154] = 1
      "0000001" when "00100011011101011", -- t[18155] = 1
      "0000001" when "00100011011101100", -- t[18156] = 1
      "0000001" when "00100011011101101", -- t[18157] = 1
      "0000001" when "00100011011101110", -- t[18158] = 1
      "0000001" when "00100011011101111", -- t[18159] = 1
      "0000001" when "00100011011110000", -- t[18160] = 1
      "0000001" when "00100011011110001", -- t[18161] = 1
      "0000001" when "00100011011110010", -- t[18162] = 1
      "0000001" when "00100011011110011", -- t[18163] = 1
      "0000001" when "00100011011110100", -- t[18164] = 1
      "0000001" when "00100011011110101", -- t[18165] = 1
      "0000001" when "00100011011110110", -- t[18166] = 1
      "0000001" when "00100011011110111", -- t[18167] = 1
      "0000001" when "00100011011111000", -- t[18168] = 1
      "0000001" when "00100011011111001", -- t[18169] = 1
      "0000001" when "00100011011111010", -- t[18170] = 1
      "0000001" when "00100011011111011", -- t[18171] = 1
      "0000001" when "00100011011111100", -- t[18172] = 1
      "0000001" when "00100011011111101", -- t[18173] = 1
      "0000001" when "00100011011111110", -- t[18174] = 1
      "0000001" when "00100011011111111", -- t[18175] = 1
      "0000001" when "00100011100000000", -- t[18176] = 1
      "0000001" when "00100011100000001", -- t[18177] = 1
      "0000001" when "00100011100000010", -- t[18178] = 1
      "0000001" when "00100011100000011", -- t[18179] = 1
      "0000001" when "00100011100000100", -- t[18180] = 1
      "0000001" when "00100011100000101", -- t[18181] = 1
      "0000001" when "00100011100000110", -- t[18182] = 1
      "0000001" when "00100011100000111", -- t[18183] = 1
      "0000001" when "00100011100001000", -- t[18184] = 1
      "0000001" when "00100011100001001", -- t[18185] = 1
      "0000001" when "00100011100001010", -- t[18186] = 1
      "0000001" when "00100011100001011", -- t[18187] = 1
      "0000001" when "00100011100001100", -- t[18188] = 1
      "0000001" when "00100011100001101", -- t[18189] = 1
      "0000001" when "00100011100001110", -- t[18190] = 1
      "0000001" when "00100011100001111", -- t[18191] = 1
      "0000001" when "00100011100010000", -- t[18192] = 1
      "0000001" when "00100011100010001", -- t[18193] = 1
      "0000001" when "00100011100010010", -- t[18194] = 1
      "0000001" when "00100011100010011", -- t[18195] = 1
      "0000001" when "00100011100010100", -- t[18196] = 1
      "0000001" when "00100011100010101", -- t[18197] = 1
      "0000001" when "00100011100010110", -- t[18198] = 1
      "0000001" when "00100011100010111", -- t[18199] = 1
      "0000001" when "00100011100011000", -- t[18200] = 1
      "0000001" when "00100011100011001", -- t[18201] = 1
      "0000001" when "00100011100011010", -- t[18202] = 1
      "0000001" when "00100011100011011", -- t[18203] = 1
      "0000001" when "00100011100011100", -- t[18204] = 1
      "0000001" when "00100011100011101", -- t[18205] = 1
      "0000001" when "00100011100011110", -- t[18206] = 1
      "0000001" when "00100011100011111", -- t[18207] = 1
      "0000001" when "00100011100100000", -- t[18208] = 1
      "0000001" when "00100011100100001", -- t[18209] = 1
      "0000001" when "00100011100100010", -- t[18210] = 1
      "0000001" when "00100011100100011", -- t[18211] = 1
      "0000001" when "00100011100100100", -- t[18212] = 1
      "0000001" when "00100011100100101", -- t[18213] = 1
      "0000001" when "00100011100100110", -- t[18214] = 1
      "0000001" when "00100011100100111", -- t[18215] = 1
      "0000001" when "00100011100101000", -- t[18216] = 1
      "0000001" when "00100011100101001", -- t[18217] = 1
      "0000001" when "00100011100101010", -- t[18218] = 1
      "0000001" when "00100011100101011", -- t[18219] = 1
      "0000001" when "00100011100101100", -- t[18220] = 1
      "0000001" when "00100011100101101", -- t[18221] = 1
      "0000001" when "00100011100101110", -- t[18222] = 1
      "0000001" when "00100011100101111", -- t[18223] = 1
      "0000001" when "00100011100110000", -- t[18224] = 1
      "0000001" when "00100011100110001", -- t[18225] = 1
      "0000001" when "00100011100110010", -- t[18226] = 1
      "0000001" when "00100011100110011", -- t[18227] = 1
      "0000001" when "00100011100110100", -- t[18228] = 1
      "0000001" when "00100011100110101", -- t[18229] = 1
      "0000001" when "00100011100110110", -- t[18230] = 1
      "0000001" when "00100011100110111", -- t[18231] = 1
      "0000001" when "00100011100111000", -- t[18232] = 1
      "0000001" when "00100011100111001", -- t[18233] = 1
      "0000001" when "00100011100111010", -- t[18234] = 1
      "0000001" when "00100011100111011", -- t[18235] = 1
      "0000001" when "00100011100111100", -- t[18236] = 1
      "0000001" when "00100011100111101", -- t[18237] = 1
      "0000001" when "00100011100111110", -- t[18238] = 1
      "0000001" when "00100011100111111", -- t[18239] = 1
      "0000001" when "00100011101000000", -- t[18240] = 1
      "0000001" when "00100011101000001", -- t[18241] = 1
      "0000001" when "00100011101000010", -- t[18242] = 1
      "0000001" when "00100011101000011", -- t[18243] = 1
      "0000001" when "00100011101000100", -- t[18244] = 1
      "0000001" when "00100011101000101", -- t[18245] = 1
      "0000001" when "00100011101000110", -- t[18246] = 1
      "0000001" when "00100011101000111", -- t[18247] = 1
      "0000001" when "00100011101001000", -- t[18248] = 1
      "0000001" when "00100011101001001", -- t[18249] = 1
      "0000001" when "00100011101001010", -- t[18250] = 1
      "0000001" when "00100011101001011", -- t[18251] = 1
      "0000001" when "00100011101001100", -- t[18252] = 1
      "0000001" when "00100011101001101", -- t[18253] = 1
      "0000001" when "00100011101001110", -- t[18254] = 1
      "0000001" when "00100011101001111", -- t[18255] = 1
      "0000001" when "00100011101010000", -- t[18256] = 1
      "0000001" when "00100011101010001", -- t[18257] = 1
      "0000001" when "00100011101010010", -- t[18258] = 1
      "0000001" when "00100011101010011", -- t[18259] = 1
      "0000001" when "00100011101010100", -- t[18260] = 1
      "0000001" when "00100011101010101", -- t[18261] = 1
      "0000001" when "00100011101010110", -- t[18262] = 1
      "0000001" when "00100011101010111", -- t[18263] = 1
      "0000001" when "00100011101011000", -- t[18264] = 1
      "0000001" when "00100011101011001", -- t[18265] = 1
      "0000001" when "00100011101011010", -- t[18266] = 1
      "0000001" when "00100011101011011", -- t[18267] = 1
      "0000001" when "00100011101011100", -- t[18268] = 1
      "0000001" when "00100011101011101", -- t[18269] = 1
      "0000001" when "00100011101011110", -- t[18270] = 1
      "0000001" when "00100011101011111", -- t[18271] = 1
      "0000001" when "00100011101100000", -- t[18272] = 1
      "0000001" when "00100011101100001", -- t[18273] = 1
      "0000001" when "00100011101100010", -- t[18274] = 1
      "0000001" when "00100011101100011", -- t[18275] = 1
      "0000001" when "00100011101100100", -- t[18276] = 1
      "0000001" when "00100011101100101", -- t[18277] = 1
      "0000001" when "00100011101100110", -- t[18278] = 1
      "0000001" when "00100011101100111", -- t[18279] = 1
      "0000001" when "00100011101101000", -- t[18280] = 1
      "0000001" when "00100011101101001", -- t[18281] = 1
      "0000001" when "00100011101101010", -- t[18282] = 1
      "0000001" when "00100011101101011", -- t[18283] = 1
      "0000001" when "00100011101101100", -- t[18284] = 1
      "0000001" when "00100011101101101", -- t[18285] = 1
      "0000001" when "00100011101101110", -- t[18286] = 1
      "0000001" when "00100011101101111", -- t[18287] = 1
      "0000001" when "00100011101110000", -- t[18288] = 1
      "0000001" when "00100011101110001", -- t[18289] = 1
      "0000001" when "00100011101110010", -- t[18290] = 1
      "0000001" when "00100011101110011", -- t[18291] = 1
      "0000001" when "00100011101110100", -- t[18292] = 1
      "0000001" when "00100011101110101", -- t[18293] = 1
      "0000001" when "00100011101110110", -- t[18294] = 1
      "0000001" when "00100011101110111", -- t[18295] = 1
      "0000001" when "00100011101111000", -- t[18296] = 1
      "0000001" when "00100011101111001", -- t[18297] = 1
      "0000001" when "00100011101111010", -- t[18298] = 1
      "0000001" when "00100011101111011", -- t[18299] = 1
      "0000001" when "00100011101111100", -- t[18300] = 1
      "0000001" when "00100011101111101", -- t[18301] = 1
      "0000001" when "00100011101111110", -- t[18302] = 1
      "0000001" when "00100011101111111", -- t[18303] = 1
      "0000001" when "00100011110000000", -- t[18304] = 1
      "0000001" when "00100011110000001", -- t[18305] = 1
      "0000001" when "00100011110000010", -- t[18306] = 1
      "0000001" when "00100011110000011", -- t[18307] = 1
      "0000001" when "00100011110000100", -- t[18308] = 1
      "0000001" when "00100011110000101", -- t[18309] = 1
      "0000001" when "00100011110000110", -- t[18310] = 1
      "0000001" when "00100011110000111", -- t[18311] = 1
      "0000001" when "00100011110001000", -- t[18312] = 1
      "0000001" when "00100011110001001", -- t[18313] = 1
      "0000001" when "00100011110001010", -- t[18314] = 1
      "0000001" when "00100011110001011", -- t[18315] = 1
      "0000001" when "00100011110001100", -- t[18316] = 1
      "0000001" when "00100011110001101", -- t[18317] = 1
      "0000001" when "00100011110001110", -- t[18318] = 1
      "0000001" when "00100011110001111", -- t[18319] = 1
      "0000001" when "00100011110010000", -- t[18320] = 1
      "0000001" when "00100011110010001", -- t[18321] = 1
      "0000001" when "00100011110010010", -- t[18322] = 1
      "0000001" when "00100011110010011", -- t[18323] = 1
      "0000001" when "00100011110010100", -- t[18324] = 1
      "0000001" when "00100011110010101", -- t[18325] = 1
      "0000001" when "00100011110010110", -- t[18326] = 1
      "0000001" when "00100011110010111", -- t[18327] = 1
      "0000001" when "00100011110011000", -- t[18328] = 1
      "0000001" when "00100011110011001", -- t[18329] = 1
      "0000001" when "00100011110011010", -- t[18330] = 1
      "0000001" when "00100011110011011", -- t[18331] = 1
      "0000001" when "00100011110011100", -- t[18332] = 1
      "0000001" when "00100011110011101", -- t[18333] = 1
      "0000001" when "00100011110011110", -- t[18334] = 1
      "0000001" when "00100011110011111", -- t[18335] = 1
      "0000001" when "00100011110100000", -- t[18336] = 1
      "0000001" when "00100011110100001", -- t[18337] = 1
      "0000001" when "00100011110100010", -- t[18338] = 1
      "0000001" when "00100011110100011", -- t[18339] = 1
      "0000001" when "00100011110100100", -- t[18340] = 1
      "0000001" when "00100011110100101", -- t[18341] = 1
      "0000001" when "00100011110100110", -- t[18342] = 1
      "0000001" when "00100011110100111", -- t[18343] = 1
      "0000001" when "00100011110101000", -- t[18344] = 1
      "0000001" when "00100011110101001", -- t[18345] = 1
      "0000001" when "00100011110101010", -- t[18346] = 1
      "0000001" when "00100011110101011", -- t[18347] = 1
      "0000001" when "00100011110101100", -- t[18348] = 1
      "0000001" when "00100011110101101", -- t[18349] = 1
      "0000001" when "00100011110101110", -- t[18350] = 1
      "0000001" when "00100011110101111", -- t[18351] = 1
      "0000001" when "00100011110110000", -- t[18352] = 1
      "0000001" when "00100011110110001", -- t[18353] = 1
      "0000001" when "00100011110110010", -- t[18354] = 1
      "0000001" when "00100011110110011", -- t[18355] = 1
      "0000001" when "00100011110110100", -- t[18356] = 1
      "0000001" when "00100011110110101", -- t[18357] = 1
      "0000001" when "00100011110110110", -- t[18358] = 1
      "0000001" when "00100011110110111", -- t[18359] = 1
      "0000001" when "00100011110111000", -- t[18360] = 1
      "0000001" when "00100011110111001", -- t[18361] = 1
      "0000001" when "00100011110111010", -- t[18362] = 1
      "0000001" when "00100011110111011", -- t[18363] = 1
      "0000001" when "00100011110111100", -- t[18364] = 1
      "0000001" when "00100011110111101", -- t[18365] = 1
      "0000001" when "00100011110111110", -- t[18366] = 1
      "0000001" when "00100011110111111", -- t[18367] = 1
      "0000001" when "00100011111000000", -- t[18368] = 1
      "0000001" when "00100011111000001", -- t[18369] = 1
      "0000001" when "00100011111000010", -- t[18370] = 1
      "0000001" when "00100011111000011", -- t[18371] = 1
      "0000001" when "00100011111000100", -- t[18372] = 1
      "0000001" when "00100011111000101", -- t[18373] = 1
      "0000001" when "00100011111000110", -- t[18374] = 1
      "0000001" when "00100011111000111", -- t[18375] = 1
      "0000001" when "00100011111001000", -- t[18376] = 1
      "0000001" when "00100011111001001", -- t[18377] = 1
      "0000001" when "00100011111001010", -- t[18378] = 1
      "0000001" when "00100011111001011", -- t[18379] = 1
      "0000001" when "00100011111001100", -- t[18380] = 1
      "0000001" when "00100011111001101", -- t[18381] = 1
      "0000001" when "00100011111001110", -- t[18382] = 1
      "0000001" when "00100011111001111", -- t[18383] = 1
      "0000001" when "00100011111010000", -- t[18384] = 1
      "0000001" when "00100011111010001", -- t[18385] = 1
      "0000001" when "00100011111010010", -- t[18386] = 1
      "0000001" when "00100011111010011", -- t[18387] = 1
      "0000001" when "00100011111010100", -- t[18388] = 1
      "0000001" when "00100011111010101", -- t[18389] = 1
      "0000001" when "00100011111010110", -- t[18390] = 1
      "0000001" when "00100011111010111", -- t[18391] = 1
      "0000001" when "00100011111011000", -- t[18392] = 1
      "0000001" when "00100011111011001", -- t[18393] = 1
      "0000001" when "00100011111011010", -- t[18394] = 1
      "0000001" when "00100011111011011", -- t[18395] = 1
      "0000001" when "00100011111011100", -- t[18396] = 1
      "0000001" when "00100011111011101", -- t[18397] = 1
      "0000001" when "00100011111011110", -- t[18398] = 1
      "0000001" when "00100011111011111", -- t[18399] = 1
      "0000001" when "00100011111100000", -- t[18400] = 1
      "0000001" when "00100011111100001", -- t[18401] = 1
      "0000001" when "00100011111100010", -- t[18402] = 1
      "0000001" when "00100011111100011", -- t[18403] = 1
      "0000001" when "00100011111100100", -- t[18404] = 1
      "0000001" when "00100011111100101", -- t[18405] = 1
      "0000001" when "00100011111100110", -- t[18406] = 1
      "0000001" when "00100011111100111", -- t[18407] = 1
      "0000001" when "00100011111101000", -- t[18408] = 1
      "0000001" when "00100011111101001", -- t[18409] = 1
      "0000001" when "00100011111101010", -- t[18410] = 1
      "0000001" when "00100011111101011", -- t[18411] = 1
      "0000001" when "00100011111101100", -- t[18412] = 1
      "0000001" when "00100011111101101", -- t[18413] = 1
      "0000001" when "00100011111101110", -- t[18414] = 1
      "0000001" when "00100011111101111", -- t[18415] = 1
      "0000001" when "00100011111110000", -- t[18416] = 1
      "0000001" when "00100011111110001", -- t[18417] = 1
      "0000001" when "00100011111110010", -- t[18418] = 1
      "0000001" when "00100011111110011", -- t[18419] = 1
      "0000001" when "00100011111110100", -- t[18420] = 1
      "0000001" when "00100011111110101", -- t[18421] = 1
      "0000001" when "00100011111110110", -- t[18422] = 1
      "0000001" when "00100011111110111", -- t[18423] = 1
      "0000001" when "00100011111111000", -- t[18424] = 1
      "0000001" when "00100011111111001", -- t[18425] = 1
      "0000001" when "00100011111111010", -- t[18426] = 1
      "0000001" when "00100011111111011", -- t[18427] = 1
      "0000001" when "00100011111111100", -- t[18428] = 1
      "0000001" when "00100011111111101", -- t[18429] = 1
      "0000001" when "00100011111111110", -- t[18430] = 1
      "0000001" when "00100011111111111", -- t[18431] = 1
      "0000001" when "00100100000000000", -- t[18432] = 1
      "0000001" when "00100100000000001", -- t[18433] = 1
      "0000001" when "00100100000000010", -- t[18434] = 1
      "0000001" when "00100100000000011", -- t[18435] = 1
      "0000001" when "00100100000000100", -- t[18436] = 1
      "0000001" when "00100100000000101", -- t[18437] = 1
      "0000001" when "00100100000000110", -- t[18438] = 1
      "0000001" when "00100100000000111", -- t[18439] = 1
      "0000001" when "00100100000001000", -- t[18440] = 1
      "0000001" when "00100100000001001", -- t[18441] = 1
      "0000001" when "00100100000001010", -- t[18442] = 1
      "0000001" when "00100100000001011", -- t[18443] = 1
      "0000001" when "00100100000001100", -- t[18444] = 1
      "0000001" when "00100100000001101", -- t[18445] = 1
      "0000001" when "00100100000001110", -- t[18446] = 1
      "0000001" when "00100100000001111", -- t[18447] = 1
      "0000001" when "00100100000010000", -- t[18448] = 1
      "0000001" when "00100100000010001", -- t[18449] = 1
      "0000001" when "00100100000010010", -- t[18450] = 1
      "0000001" when "00100100000010011", -- t[18451] = 1
      "0000001" when "00100100000010100", -- t[18452] = 1
      "0000001" when "00100100000010101", -- t[18453] = 1
      "0000001" when "00100100000010110", -- t[18454] = 1
      "0000001" when "00100100000010111", -- t[18455] = 1
      "0000001" when "00100100000011000", -- t[18456] = 1
      "0000001" when "00100100000011001", -- t[18457] = 1
      "0000001" when "00100100000011010", -- t[18458] = 1
      "0000001" when "00100100000011011", -- t[18459] = 1
      "0000001" when "00100100000011100", -- t[18460] = 1
      "0000001" when "00100100000011101", -- t[18461] = 1
      "0000001" when "00100100000011110", -- t[18462] = 1
      "0000001" when "00100100000011111", -- t[18463] = 1
      "0000001" when "00100100000100000", -- t[18464] = 1
      "0000001" when "00100100000100001", -- t[18465] = 1
      "0000001" when "00100100000100010", -- t[18466] = 1
      "0000001" when "00100100000100011", -- t[18467] = 1
      "0000001" when "00100100000100100", -- t[18468] = 1
      "0000001" when "00100100000100101", -- t[18469] = 1
      "0000001" when "00100100000100110", -- t[18470] = 1
      "0000001" when "00100100000100111", -- t[18471] = 1
      "0000001" when "00100100000101000", -- t[18472] = 1
      "0000001" when "00100100000101001", -- t[18473] = 1
      "0000001" when "00100100000101010", -- t[18474] = 1
      "0000001" when "00100100000101011", -- t[18475] = 1
      "0000001" when "00100100000101100", -- t[18476] = 1
      "0000001" when "00100100000101101", -- t[18477] = 1
      "0000001" when "00100100000101110", -- t[18478] = 1
      "0000001" when "00100100000101111", -- t[18479] = 1
      "0000001" when "00100100000110000", -- t[18480] = 1
      "0000001" when "00100100000110001", -- t[18481] = 1
      "0000001" when "00100100000110010", -- t[18482] = 1
      "0000001" when "00100100000110011", -- t[18483] = 1
      "0000001" when "00100100000110100", -- t[18484] = 1
      "0000001" when "00100100000110101", -- t[18485] = 1
      "0000001" when "00100100000110110", -- t[18486] = 1
      "0000001" when "00100100000110111", -- t[18487] = 1
      "0000001" when "00100100000111000", -- t[18488] = 1
      "0000001" when "00100100000111001", -- t[18489] = 1
      "0000001" when "00100100000111010", -- t[18490] = 1
      "0000001" when "00100100000111011", -- t[18491] = 1
      "0000001" when "00100100000111100", -- t[18492] = 1
      "0000001" when "00100100000111101", -- t[18493] = 1
      "0000001" when "00100100000111110", -- t[18494] = 1
      "0000001" when "00100100000111111", -- t[18495] = 1
      "0000001" when "00100100001000000", -- t[18496] = 1
      "0000001" when "00100100001000001", -- t[18497] = 1
      "0000001" when "00100100001000010", -- t[18498] = 1
      "0000001" when "00100100001000011", -- t[18499] = 1
      "0000001" when "00100100001000100", -- t[18500] = 1
      "0000001" when "00100100001000101", -- t[18501] = 1
      "0000001" when "00100100001000110", -- t[18502] = 1
      "0000001" when "00100100001000111", -- t[18503] = 1
      "0000001" when "00100100001001000", -- t[18504] = 1
      "0000001" when "00100100001001001", -- t[18505] = 1
      "0000001" when "00100100001001010", -- t[18506] = 1
      "0000001" when "00100100001001011", -- t[18507] = 1
      "0000001" when "00100100001001100", -- t[18508] = 1
      "0000001" when "00100100001001101", -- t[18509] = 1
      "0000001" when "00100100001001110", -- t[18510] = 1
      "0000001" when "00100100001001111", -- t[18511] = 1
      "0000001" when "00100100001010000", -- t[18512] = 1
      "0000001" when "00100100001010001", -- t[18513] = 1
      "0000001" when "00100100001010010", -- t[18514] = 1
      "0000001" when "00100100001010011", -- t[18515] = 1
      "0000001" when "00100100001010100", -- t[18516] = 1
      "0000001" when "00100100001010101", -- t[18517] = 1
      "0000001" when "00100100001010110", -- t[18518] = 1
      "0000001" when "00100100001010111", -- t[18519] = 1
      "0000001" when "00100100001011000", -- t[18520] = 1
      "0000001" when "00100100001011001", -- t[18521] = 1
      "0000001" when "00100100001011010", -- t[18522] = 1
      "0000001" when "00100100001011011", -- t[18523] = 1
      "0000001" when "00100100001011100", -- t[18524] = 1
      "0000001" when "00100100001011101", -- t[18525] = 1
      "0000001" when "00100100001011110", -- t[18526] = 1
      "0000001" when "00100100001011111", -- t[18527] = 1
      "0000001" when "00100100001100000", -- t[18528] = 1
      "0000001" when "00100100001100001", -- t[18529] = 1
      "0000001" when "00100100001100010", -- t[18530] = 1
      "0000001" when "00100100001100011", -- t[18531] = 1
      "0000001" when "00100100001100100", -- t[18532] = 1
      "0000001" when "00100100001100101", -- t[18533] = 1
      "0000001" when "00100100001100110", -- t[18534] = 1
      "0000001" when "00100100001100111", -- t[18535] = 1
      "0000001" when "00100100001101000", -- t[18536] = 1
      "0000001" when "00100100001101001", -- t[18537] = 1
      "0000001" when "00100100001101010", -- t[18538] = 1
      "0000001" when "00100100001101011", -- t[18539] = 1
      "0000001" when "00100100001101100", -- t[18540] = 1
      "0000001" when "00100100001101101", -- t[18541] = 1
      "0000001" when "00100100001101110", -- t[18542] = 1
      "0000001" when "00100100001101111", -- t[18543] = 1
      "0000001" when "00100100001110000", -- t[18544] = 1
      "0000001" when "00100100001110001", -- t[18545] = 1
      "0000001" when "00100100001110010", -- t[18546] = 1
      "0000001" when "00100100001110011", -- t[18547] = 1
      "0000001" when "00100100001110100", -- t[18548] = 1
      "0000001" when "00100100001110101", -- t[18549] = 1
      "0000001" when "00100100001110110", -- t[18550] = 1
      "0000001" when "00100100001110111", -- t[18551] = 1
      "0000001" when "00100100001111000", -- t[18552] = 1
      "0000001" when "00100100001111001", -- t[18553] = 1
      "0000001" when "00100100001111010", -- t[18554] = 1
      "0000001" when "00100100001111011", -- t[18555] = 1
      "0000001" when "00100100001111100", -- t[18556] = 1
      "0000001" when "00100100001111101", -- t[18557] = 1
      "0000001" when "00100100001111110", -- t[18558] = 1
      "0000001" when "00100100001111111", -- t[18559] = 1
      "0000001" when "00100100010000000", -- t[18560] = 1
      "0000001" when "00100100010000001", -- t[18561] = 1
      "0000001" when "00100100010000010", -- t[18562] = 1
      "0000001" when "00100100010000011", -- t[18563] = 1
      "0000001" when "00100100010000100", -- t[18564] = 1
      "0000001" when "00100100010000101", -- t[18565] = 1
      "0000001" when "00100100010000110", -- t[18566] = 1
      "0000001" when "00100100010000111", -- t[18567] = 1
      "0000001" when "00100100010001000", -- t[18568] = 1
      "0000001" when "00100100010001001", -- t[18569] = 1
      "0000001" when "00100100010001010", -- t[18570] = 1
      "0000001" when "00100100010001011", -- t[18571] = 1
      "0000001" when "00100100010001100", -- t[18572] = 1
      "0000001" when "00100100010001101", -- t[18573] = 1
      "0000001" when "00100100010001110", -- t[18574] = 1
      "0000001" when "00100100010001111", -- t[18575] = 1
      "0000001" when "00100100010010000", -- t[18576] = 1
      "0000001" when "00100100010010001", -- t[18577] = 1
      "0000001" when "00100100010010010", -- t[18578] = 1
      "0000001" when "00100100010010011", -- t[18579] = 1
      "0000001" when "00100100010010100", -- t[18580] = 1
      "0000001" when "00100100010010101", -- t[18581] = 1
      "0000001" when "00100100010010110", -- t[18582] = 1
      "0000001" when "00100100010010111", -- t[18583] = 1
      "0000001" when "00100100010011000", -- t[18584] = 1
      "0000001" when "00100100010011001", -- t[18585] = 1
      "0000001" when "00100100010011010", -- t[18586] = 1
      "0000001" when "00100100010011011", -- t[18587] = 1
      "0000001" when "00100100010011100", -- t[18588] = 1
      "0000001" when "00100100010011101", -- t[18589] = 1
      "0000001" when "00100100010011110", -- t[18590] = 1
      "0000001" when "00100100010011111", -- t[18591] = 1
      "0000001" when "00100100010100000", -- t[18592] = 1
      "0000001" when "00100100010100001", -- t[18593] = 1
      "0000001" when "00100100010100010", -- t[18594] = 1
      "0000001" when "00100100010100011", -- t[18595] = 1
      "0000001" when "00100100010100100", -- t[18596] = 1
      "0000001" when "00100100010100101", -- t[18597] = 1
      "0000001" when "00100100010100110", -- t[18598] = 1
      "0000001" when "00100100010100111", -- t[18599] = 1
      "0000001" when "00100100010101000", -- t[18600] = 1
      "0000001" when "00100100010101001", -- t[18601] = 1
      "0000001" when "00100100010101010", -- t[18602] = 1
      "0000001" when "00100100010101011", -- t[18603] = 1
      "0000001" when "00100100010101100", -- t[18604] = 1
      "0000001" when "00100100010101101", -- t[18605] = 1
      "0000001" when "00100100010101110", -- t[18606] = 1
      "0000001" when "00100100010101111", -- t[18607] = 1
      "0000001" when "00100100010110000", -- t[18608] = 1
      "0000001" when "00100100010110001", -- t[18609] = 1
      "0000001" when "00100100010110010", -- t[18610] = 1
      "0000001" when "00100100010110011", -- t[18611] = 1
      "0000001" when "00100100010110100", -- t[18612] = 1
      "0000001" when "00100100010110101", -- t[18613] = 1
      "0000001" when "00100100010110110", -- t[18614] = 1
      "0000001" when "00100100010110111", -- t[18615] = 1
      "0000001" when "00100100010111000", -- t[18616] = 1
      "0000001" when "00100100010111001", -- t[18617] = 1
      "0000001" when "00100100010111010", -- t[18618] = 1
      "0000001" when "00100100010111011", -- t[18619] = 1
      "0000001" when "00100100010111100", -- t[18620] = 1
      "0000001" when "00100100010111101", -- t[18621] = 1
      "0000001" when "00100100010111110", -- t[18622] = 1
      "0000001" when "00100100010111111", -- t[18623] = 1
      "0000001" when "00100100011000000", -- t[18624] = 1
      "0000001" when "00100100011000001", -- t[18625] = 1
      "0000001" when "00100100011000010", -- t[18626] = 1
      "0000001" when "00100100011000011", -- t[18627] = 1
      "0000001" when "00100100011000100", -- t[18628] = 1
      "0000001" when "00100100011000101", -- t[18629] = 1
      "0000001" when "00100100011000110", -- t[18630] = 1
      "0000001" when "00100100011000111", -- t[18631] = 1
      "0000001" when "00100100011001000", -- t[18632] = 1
      "0000001" when "00100100011001001", -- t[18633] = 1
      "0000001" when "00100100011001010", -- t[18634] = 1
      "0000001" when "00100100011001011", -- t[18635] = 1
      "0000001" when "00100100011001100", -- t[18636] = 1
      "0000001" when "00100100011001101", -- t[18637] = 1
      "0000001" when "00100100011001110", -- t[18638] = 1
      "0000001" when "00100100011001111", -- t[18639] = 1
      "0000001" when "00100100011010000", -- t[18640] = 1
      "0000001" when "00100100011010001", -- t[18641] = 1
      "0000001" when "00100100011010010", -- t[18642] = 1
      "0000001" when "00100100011010011", -- t[18643] = 1
      "0000001" when "00100100011010100", -- t[18644] = 1
      "0000001" when "00100100011010101", -- t[18645] = 1
      "0000001" when "00100100011010110", -- t[18646] = 1
      "0000001" when "00100100011010111", -- t[18647] = 1
      "0000001" when "00100100011011000", -- t[18648] = 1
      "0000001" when "00100100011011001", -- t[18649] = 1
      "0000001" when "00100100011011010", -- t[18650] = 1
      "0000001" when "00100100011011011", -- t[18651] = 1
      "0000001" when "00100100011011100", -- t[18652] = 1
      "0000001" when "00100100011011101", -- t[18653] = 1
      "0000001" when "00100100011011110", -- t[18654] = 1
      "0000001" when "00100100011011111", -- t[18655] = 1
      "0000001" when "00100100011100000", -- t[18656] = 1
      "0000001" when "00100100011100001", -- t[18657] = 1
      "0000001" when "00100100011100010", -- t[18658] = 1
      "0000001" when "00100100011100011", -- t[18659] = 1
      "0000001" when "00100100011100100", -- t[18660] = 1
      "0000001" when "00100100011100101", -- t[18661] = 1
      "0000001" when "00100100011100110", -- t[18662] = 1
      "0000001" when "00100100011100111", -- t[18663] = 1
      "0000001" when "00100100011101000", -- t[18664] = 1
      "0000001" when "00100100011101001", -- t[18665] = 1
      "0000001" when "00100100011101010", -- t[18666] = 1
      "0000001" when "00100100011101011", -- t[18667] = 1
      "0000001" when "00100100011101100", -- t[18668] = 1
      "0000001" when "00100100011101101", -- t[18669] = 1
      "0000001" when "00100100011101110", -- t[18670] = 1
      "0000001" when "00100100011101111", -- t[18671] = 1
      "0000001" when "00100100011110000", -- t[18672] = 1
      "0000001" when "00100100011110001", -- t[18673] = 1
      "0000001" when "00100100011110010", -- t[18674] = 1
      "0000001" when "00100100011110011", -- t[18675] = 1
      "0000001" when "00100100011110100", -- t[18676] = 1
      "0000001" when "00100100011110101", -- t[18677] = 1
      "0000001" when "00100100011110110", -- t[18678] = 1
      "0000001" when "00100100011110111", -- t[18679] = 1
      "0000001" when "00100100011111000", -- t[18680] = 1
      "0000001" when "00100100011111001", -- t[18681] = 1
      "0000001" when "00100100011111010", -- t[18682] = 1
      "0000001" when "00100100011111011", -- t[18683] = 1
      "0000001" when "00100100011111100", -- t[18684] = 1
      "0000001" when "00100100011111101", -- t[18685] = 1
      "0000001" when "00100100011111110", -- t[18686] = 1
      "0000001" when "00100100011111111", -- t[18687] = 1
      "0000001" when "00100100100000000", -- t[18688] = 1
      "0000001" when "00100100100000001", -- t[18689] = 1
      "0000001" when "00100100100000010", -- t[18690] = 1
      "0000001" when "00100100100000011", -- t[18691] = 1
      "0000001" when "00100100100000100", -- t[18692] = 1
      "0000001" when "00100100100000101", -- t[18693] = 1
      "0000001" when "00100100100000110", -- t[18694] = 1
      "0000001" when "00100100100000111", -- t[18695] = 1
      "0000001" when "00100100100001000", -- t[18696] = 1
      "0000001" when "00100100100001001", -- t[18697] = 1
      "0000001" when "00100100100001010", -- t[18698] = 1
      "0000001" when "00100100100001011", -- t[18699] = 1
      "0000001" when "00100100100001100", -- t[18700] = 1
      "0000001" when "00100100100001101", -- t[18701] = 1
      "0000001" when "00100100100001110", -- t[18702] = 1
      "0000001" when "00100100100001111", -- t[18703] = 1
      "0000001" when "00100100100010000", -- t[18704] = 1
      "0000001" when "00100100100010001", -- t[18705] = 1
      "0000001" when "00100100100010010", -- t[18706] = 1
      "0000001" when "00100100100010011", -- t[18707] = 1
      "0000001" when "00100100100010100", -- t[18708] = 1
      "0000001" when "00100100100010101", -- t[18709] = 1
      "0000001" when "00100100100010110", -- t[18710] = 1
      "0000001" when "00100100100010111", -- t[18711] = 1
      "0000001" when "00100100100011000", -- t[18712] = 1
      "0000001" when "00100100100011001", -- t[18713] = 1
      "0000001" when "00100100100011010", -- t[18714] = 1
      "0000001" when "00100100100011011", -- t[18715] = 1
      "0000001" when "00100100100011100", -- t[18716] = 1
      "0000001" when "00100100100011101", -- t[18717] = 1
      "0000001" when "00100100100011110", -- t[18718] = 1
      "0000001" when "00100100100011111", -- t[18719] = 1
      "0000001" when "00100100100100000", -- t[18720] = 1
      "0000001" when "00100100100100001", -- t[18721] = 1
      "0000001" when "00100100100100010", -- t[18722] = 1
      "0000001" when "00100100100100011", -- t[18723] = 1
      "0000001" when "00100100100100100", -- t[18724] = 1
      "0000001" when "00100100100100101", -- t[18725] = 1
      "0000001" when "00100100100100110", -- t[18726] = 1
      "0000001" when "00100100100100111", -- t[18727] = 1
      "0000001" when "00100100100101000", -- t[18728] = 1
      "0000001" when "00100100100101001", -- t[18729] = 1
      "0000001" when "00100100100101010", -- t[18730] = 1
      "0000001" when "00100100100101011", -- t[18731] = 1
      "0000001" when "00100100100101100", -- t[18732] = 1
      "0000001" when "00100100100101101", -- t[18733] = 1
      "0000001" when "00100100100101110", -- t[18734] = 1
      "0000001" when "00100100100101111", -- t[18735] = 1
      "0000001" when "00100100100110000", -- t[18736] = 1
      "0000001" when "00100100100110001", -- t[18737] = 1
      "0000001" when "00100100100110010", -- t[18738] = 1
      "0000001" when "00100100100110011", -- t[18739] = 1
      "0000001" when "00100100100110100", -- t[18740] = 1
      "0000001" when "00100100100110101", -- t[18741] = 1
      "0000001" when "00100100100110110", -- t[18742] = 1
      "0000001" when "00100100100110111", -- t[18743] = 1
      "0000001" when "00100100100111000", -- t[18744] = 1
      "0000001" when "00100100100111001", -- t[18745] = 1
      "0000001" when "00100100100111010", -- t[18746] = 1
      "0000001" when "00100100100111011", -- t[18747] = 1
      "0000001" when "00100100100111100", -- t[18748] = 1
      "0000001" when "00100100100111101", -- t[18749] = 1
      "0000001" when "00100100100111110", -- t[18750] = 1
      "0000001" when "00100100100111111", -- t[18751] = 1
      "0000001" when "00100100101000000", -- t[18752] = 1
      "0000001" when "00100100101000001", -- t[18753] = 1
      "0000001" when "00100100101000010", -- t[18754] = 1
      "0000001" when "00100100101000011", -- t[18755] = 1
      "0000001" when "00100100101000100", -- t[18756] = 1
      "0000001" when "00100100101000101", -- t[18757] = 1
      "0000001" when "00100100101000110", -- t[18758] = 1
      "0000001" when "00100100101000111", -- t[18759] = 1
      "0000001" when "00100100101001000", -- t[18760] = 1
      "0000001" when "00100100101001001", -- t[18761] = 1
      "0000001" when "00100100101001010", -- t[18762] = 1
      "0000001" when "00100100101001011", -- t[18763] = 1
      "0000001" when "00100100101001100", -- t[18764] = 1
      "0000001" when "00100100101001101", -- t[18765] = 1
      "0000001" when "00100100101001110", -- t[18766] = 1
      "0000001" when "00100100101001111", -- t[18767] = 1
      "0000001" when "00100100101010000", -- t[18768] = 1
      "0000001" when "00100100101010001", -- t[18769] = 1
      "0000001" when "00100100101010010", -- t[18770] = 1
      "0000001" when "00100100101010011", -- t[18771] = 1
      "0000001" when "00100100101010100", -- t[18772] = 1
      "0000001" when "00100100101010101", -- t[18773] = 1
      "0000001" when "00100100101010110", -- t[18774] = 1
      "0000001" when "00100100101010111", -- t[18775] = 1
      "0000001" when "00100100101011000", -- t[18776] = 1
      "0000001" when "00100100101011001", -- t[18777] = 1
      "0000001" when "00100100101011010", -- t[18778] = 1
      "0000001" when "00100100101011011", -- t[18779] = 1
      "0000001" when "00100100101011100", -- t[18780] = 1
      "0000001" when "00100100101011101", -- t[18781] = 1
      "0000001" when "00100100101011110", -- t[18782] = 1
      "0000001" when "00100100101011111", -- t[18783] = 1
      "0000001" when "00100100101100000", -- t[18784] = 1
      "0000001" when "00100100101100001", -- t[18785] = 1
      "0000001" when "00100100101100010", -- t[18786] = 1
      "0000001" when "00100100101100011", -- t[18787] = 1
      "0000001" when "00100100101100100", -- t[18788] = 1
      "0000001" when "00100100101100101", -- t[18789] = 1
      "0000001" when "00100100101100110", -- t[18790] = 1
      "0000001" when "00100100101100111", -- t[18791] = 1
      "0000001" when "00100100101101000", -- t[18792] = 1
      "0000001" when "00100100101101001", -- t[18793] = 1
      "0000001" when "00100100101101010", -- t[18794] = 1
      "0000001" when "00100100101101011", -- t[18795] = 1
      "0000001" when "00100100101101100", -- t[18796] = 1
      "0000001" when "00100100101101101", -- t[18797] = 1
      "0000001" when "00100100101101110", -- t[18798] = 1
      "0000001" when "00100100101101111", -- t[18799] = 1
      "0000001" when "00100100101110000", -- t[18800] = 1
      "0000001" when "00100100101110001", -- t[18801] = 1
      "0000001" when "00100100101110010", -- t[18802] = 1
      "0000001" when "00100100101110011", -- t[18803] = 1
      "0000001" when "00100100101110100", -- t[18804] = 1
      "0000001" when "00100100101110101", -- t[18805] = 1
      "0000001" when "00100100101110110", -- t[18806] = 1
      "0000001" when "00100100101110111", -- t[18807] = 1
      "0000001" when "00100100101111000", -- t[18808] = 1
      "0000001" when "00100100101111001", -- t[18809] = 1
      "0000001" when "00100100101111010", -- t[18810] = 1
      "0000001" when "00100100101111011", -- t[18811] = 1
      "0000001" when "00100100101111100", -- t[18812] = 1
      "0000001" when "00100100101111101", -- t[18813] = 1
      "0000001" when "00100100101111110", -- t[18814] = 1
      "0000001" when "00100100101111111", -- t[18815] = 1
      "0000001" when "00100100110000000", -- t[18816] = 1
      "0000001" when "00100100110000001", -- t[18817] = 1
      "0000001" when "00100100110000010", -- t[18818] = 1
      "0000001" when "00100100110000011", -- t[18819] = 1
      "0000001" when "00100100110000100", -- t[18820] = 1
      "0000001" when "00100100110000101", -- t[18821] = 1
      "0000001" when "00100100110000110", -- t[18822] = 1
      "0000001" when "00100100110000111", -- t[18823] = 1
      "0000001" when "00100100110001000", -- t[18824] = 1
      "0000001" when "00100100110001001", -- t[18825] = 1
      "0000001" when "00100100110001010", -- t[18826] = 1
      "0000001" when "00100100110001011", -- t[18827] = 1
      "0000001" when "00100100110001100", -- t[18828] = 1
      "0000001" when "00100100110001101", -- t[18829] = 1
      "0000001" when "00100100110001110", -- t[18830] = 1
      "0000001" when "00100100110001111", -- t[18831] = 1
      "0000001" when "00100100110010000", -- t[18832] = 1
      "0000001" when "00100100110010001", -- t[18833] = 1
      "0000001" when "00100100110010010", -- t[18834] = 1
      "0000001" when "00100100110010011", -- t[18835] = 1
      "0000001" when "00100100110010100", -- t[18836] = 1
      "0000001" when "00100100110010101", -- t[18837] = 1
      "0000001" when "00100100110010110", -- t[18838] = 1
      "0000001" when "00100100110010111", -- t[18839] = 1
      "0000001" when "00100100110011000", -- t[18840] = 1
      "0000001" when "00100100110011001", -- t[18841] = 1
      "0000001" when "00100100110011010", -- t[18842] = 1
      "0000001" when "00100100110011011", -- t[18843] = 1
      "0000001" when "00100100110011100", -- t[18844] = 1
      "0000001" when "00100100110011101", -- t[18845] = 1
      "0000001" when "00100100110011110", -- t[18846] = 1
      "0000001" when "00100100110011111", -- t[18847] = 1
      "0000001" when "00100100110100000", -- t[18848] = 1
      "0000001" when "00100100110100001", -- t[18849] = 1
      "0000001" when "00100100110100010", -- t[18850] = 1
      "0000001" when "00100100110100011", -- t[18851] = 1
      "0000001" when "00100100110100100", -- t[18852] = 1
      "0000001" when "00100100110100101", -- t[18853] = 1
      "0000001" when "00100100110100110", -- t[18854] = 1
      "0000001" when "00100100110100111", -- t[18855] = 1
      "0000001" when "00100100110101000", -- t[18856] = 1
      "0000001" when "00100100110101001", -- t[18857] = 1
      "0000001" when "00100100110101010", -- t[18858] = 1
      "0000001" when "00100100110101011", -- t[18859] = 1
      "0000001" when "00100100110101100", -- t[18860] = 1
      "0000001" when "00100100110101101", -- t[18861] = 1
      "0000001" when "00100100110101110", -- t[18862] = 1
      "0000001" when "00100100110101111", -- t[18863] = 1
      "0000001" when "00100100110110000", -- t[18864] = 1
      "0000001" when "00100100110110001", -- t[18865] = 1
      "0000001" when "00100100110110010", -- t[18866] = 1
      "0000001" when "00100100110110011", -- t[18867] = 1
      "0000001" when "00100100110110100", -- t[18868] = 1
      "0000001" when "00100100110110101", -- t[18869] = 1
      "0000001" when "00100100110110110", -- t[18870] = 1
      "0000001" when "00100100110110111", -- t[18871] = 1
      "0000001" when "00100100110111000", -- t[18872] = 1
      "0000001" when "00100100110111001", -- t[18873] = 1
      "0000001" when "00100100110111010", -- t[18874] = 1
      "0000001" when "00100100110111011", -- t[18875] = 1
      "0000001" when "00100100110111100", -- t[18876] = 1
      "0000001" when "00100100110111101", -- t[18877] = 1
      "0000001" when "00100100110111110", -- t[18878] = 1
      "0000001" when "00100100110111111", -- t[18879] = 1
      "0000001" when "00100100111000000", -- t[18880] = 1
      "0000001" when "00100100111000001", -- t[18881] = 1
      "0000001" when "00100100111000010", -- t[18882] = 1
      "0000001" when "00100100111000011", -- t[18883] = 1
      "0000001" when "00100100111000100", -- t[18884] = 1
      "0000001" when "00100100111000101", -- t[18885] = 1
      "0000001" when "00100100111000110", -- t[18886] = 1
      "0000001" when "00100100111000111", -- t[18887] = 1
      "0000001" when "00100100111001000", -- t[18888] = 1
      "0000001" when "00100100111001001", -- t[18889] = 1
      "0000001" when "00100100111001010", -- t[18890] = 1
      "0000001" when "00100100111001011", -- t[18891] = 1
      "0000001" when "00100100111001100", -- t[18892] = 1
      "0000001" when "00100100111001101", -- t[18893] = 1
      "0000001" when "00100100111001110", -- t[18894] = 1
      "0000001" when "00100100111001111", -- t[18895] = 1
      "0000001" when "00100100111010000", -- t[18896] = 1
      "0000001" when "00100100111010001", -- t[18897] = 1
      "0000001" when "00100100111010010", -- t[18898] = 1
      "0000001" when "00100100111010011", -- t[18899] = 1
      "0000001" when "00100100111010100", -- t[18900] = 1
      "0000001" when "00100100111010101", -- t[18901] = 1
      "0000001" when "00100100111010110", -- t[18902] = 1
      "0000001" when "00100100111010111", -- t[18903] = 1
      "0000001" when "00100100111011000", -- t[18904] = 1
      "0000001" when "00100100111011001", -- t[18905] = 1
      "0000001" when "00100100111011010", -- t[18906] = 1
      "0000001" when "00100100111011011", -- t[18907] = 1
      "0000001" when "00100100111011100", -- t[18908] = 1
      "0000001" when "00100100111011101", -- t[18909] = 1
      "0000001" when "00100100111011110", -- t[18910] = 1
      "0000001" when "00100100111011111", -- t[18911] = 1
      "0000001" when "00100100111100000", -- t[18912] = 1
      "0000001" when "00100100111100001", -- t[18913] = 1
      "0000001" when "00100100111100010", -- t[18914] = 1
      "0000001" when "00100100111100011", -- t[18915] = 1
      "0000001" when "00100100111100100", -- t[18916] = 1
      "0000001" when "00100100111100101", -- t[18917] = 1
      "0000001" when "00100100111100110", -- t[18918] = 1
      "0000001" when "00100100111100111", -- t[18919] = 1
      "0000001" when "00100100111101000", -- t[18920] = 1
      "0000001" when "00100100111101001", -- t[18921] = 1
      "0000001" when "00100100111101010", -- t[18922] = 1
      "0000001" when "00100100111101011", -- t[18923] = 1
      "0000001" when "00100100111101100", -- t[18924] = 1
      "0000001" when "00100100111101101", -- t[18925] = 1
      "0000001" when "00100100111101110", -- t[18926] = 1
      "0000001" when "00100100111101111", -- t[18927] = 1
      "0000001" when "00100100111110000", -- t[18928] = 1
      "0000001" when "00100100111110001", -- t[18929] = 1
      "0000001" when "00100100111110010", -- t[18930] = 1
      "0000001" when "00100100111110011", -- t[18931] = 1
      "0000001" when "00100100111110100", -- t[18932] = 1
      "0000001" when "00100100111110101", -- t[18933] = 1
      "0000001" when "00100100111110110", -- t[18934] = 1
      "0000001" when "00100100111110111", -- t[18935] = 1
      "0000001" when "00100100111111000", -- t[18936] = 1
      "0000001" when "00100100111111001", -- t[18937] = 1
      "0000001" when "00100100111111010", -- t[18938] = 1
      "0000001" when "00100100111111011", -- t[18939] = 1
      "0000001" when "00100100111111100", -- t[18940] = 1
      "0000001" when "00100100111111101", -- t[18941] = 1
      "0000001" when "00100100111111110", -- t[18942] = 1
      "0000001" when "00100100111111111", -- t[18943] = 1
      "0000001" when "00100101000000000", -- t[18944] = 1
      "0000001" when "00100101000000001", -- t[18945] = 1
      "0000001" when "00100101000000010", -- t[18946] = 1
      "0000001" when "00100101000000011", -- t[18947] = 1
      "0000001" when "00100101000000100", -- t[18948] = 1
      "0000001" when "00100101000000101", -- t[18949] = 1
      "0000001" when "00100101000000110", -- t[18950] = 1
      "0000001" when "00100101000000111", -- t[18951] = 1
      "0000001" when "00100101000001000", -- t[18952] = 1
      "0000001" when "00100101000001001", -- t[18953] = 1
      "0000001" when "00100101000001010", -- t[18954] = 1
      "0000001" when "00100101000001011", -- t[18955] = 1
      "0000001" when "00100101000001100", -- t[18956] = 1
      "0000001" when "00100101000001101", -- t[18957] = 1
      "0000001" when "00100101000001110", -- t[18958] = 1
      "0000001" when "00100101000001111", -- t[18959] = 1
      "0000001" when "00100101000010000", -- t[18960] = 1
      "0000001" when "00100101000010001", -- t[18961] = 1
      "0000001" when "00100101000010010", -- t[18962] = 1
      "0000001" when "00100101000010011", -- t[18963] = 1
      "0000001" when "00100101000010100", -- t[18964] = 1
      "0000001" when "00100101000010101", -- t[18965] = 1
      "0000001" when "00100101000010110", -- t[18966] = 1
      "0000001" when "00100101000010111", -- t[18967] = 1
      "0000001" when "00100101000011000", -- t[18968] = 1
      "0000001" when "00100101000011001", -- t[18969] = 1
      "0000001" when "00100101000011010", -- t[18970] = 1
      "0000001" when "00100101000011011", -- t[18971] = 1
      "0000001" when "00100101000011100", -- t[18972] = 1
      "0000001" when "00100101000011101", -- t[18973] = 1
      "0000001" when "00100101000011110", -- t[18974] = 1
      "0000001" when "00100101000011111", -- t[18975] = 1
      "0000001" when "00100101000100000", -- t[18976] = 1
      "0000001" when "00100101000100001", -- t[18977] = 1
      "0000001" when "00100101000100010", -- t[18978] = 1
      "0000001" when "00100101000100011", -- t[18979] = 1
      "0000001" when "00100101000100100", -- t[18980] = 1
      "0000001" when "00100101000100101", -- t[18981] = 1
      "0000001" when "00100101000100110", -- t[18982] = 1
      "0000001" when "00100101000100111", -- t[18983] = 1
      "0000001" when "00100101000101000", -- t[18984] = 1
      "0000001" when "00100101000101001", -- t[18985] = 1
      "0000001" when "00100101000101010", -- t[18986] = 1
      "0000001" when "00100101000101011", -- t[18987] = 1
      "0000001" when "00100101000101100", -- t[18988] = 1
      "0000001" when "00100101000101101", -- t[18989] = 1
      "0000001" when "00100101000101110", -- t[18990] = 1
      "0000001" when "00100101000101111", -- t[18991] = 1
      "0000001" when "00100101000110000", -- t[18992] = 1
      "0000001" when "00100101000110001", -- t[18993] = 1
      "0000001" when "00100101000110010", -- t[18994] = 1
      "0000001" when "00100101000110011", -- t[18995] = 1
      "0000001" when "00100101000110100", -- t[18996] = 1
      "0000001" when "00100101000110101", -- t[18997] = 1
      "0000001" when "00100101000110110", -- t[18998] = 1
      "0000001" when "00100101000110111", -- t[18999] = 1
      "0000001" when "00100101000111000", -- t[19000] = 1
      "0000001" when "00100101000111001", -- t[19001] = 1
      "0000001" when "00100101000111010", -- t[19002] = 1
      "0000001" when "00100101000111011", -- t[19003] = 1
      "0000001" when "00100101000111100", -- t[19004] = 1
      "0000001" when "00100101000111101", -- t[19005] = 1
      "0000001" when "00100101000111110", -- t[19006] = 1
      "0000001" when "00100101000111111", -- t[19007] = 1
      "0000001" when "00100101001000000", -- t[19008] = 1
      "0000001" when "00100101001000001", -- t[19009] = 1
      "0000001" when "00100101001000010", -- t[19010] = 1
      "0000001" when "00100101001000011", -- t[19011] = 1
      "0000001" when "00100101001000100", -- t[19012] = 1
      "0000001" when "00100101001000101", -- t[19013] = 1
      "0000001" when "00100101001000110", -- t[19014] = 1
      "0000001" when "00100101001000111", -- t[19015] = 1
      "0000001" when "00100101001001000", -- t[19016] = 1
      "0000001" when "00100101001001001", -- t[19017] = 1
      "0000001" when "00100101001001010", -- t[19018] = 1
      "0000001" when "00100101001001011", -- t[19019] = 1
      "0000001" when "00100101001001100", -- t[19020] = 1
      "0000001" when "00100101001001101", -- t[19021] = 1
      "0000001" when "00100101001001110", -- t[19022] = 1
      "0000001" when "00100101001001111", -- t[19023] = 1
      "0000001" when "00100101001010000", -- t[19024] = 1
      "0000001" when "00100101001010001", -- t[19025] = 1
      "0000001" when "00100101001010010", -- t[19026] = 1
      "0000001" when "00100101001010011", -- t[19027] = 1
      "0000001" when "00100101001010100", -- t[19028] = 1
      "0000001" when "00100101001010101", -- t[19029] = 1
      "0000001" when "00100101001010110", -- t[19030] = 1
      "0000001" when "00100101001010111", -- t[19031] = 1
      "0000001" when "00100101001011000", -- t[19032] = 1
      "0000001" when "00100101001011001", -- t[19033] = 1
      "0000001" when "00100101001011010", -- t[19034] = 1
      "0000001" when "00100101001011011", -- t[19035] = 1
      "0000001" when "00100101001011100", -- t[19036] = 1
      "0000001" when "00100101001011101", -- t[19037] = 1
      "0000001" when "00100101001011110", -- t[19038] = 1
      "0000001" when "00100101001011111", -- t[19039] = 1
      "0000001" when "00100101001100000", -- t[19040] = 1
      "0000001" when "00100101001100001", -- t[19041] = 1
      "0000001" when "00100101001100010", -- t[19042] = 1
      "0000001" when "00100101001100011", -- t[19043] = 1
      "0000001" when "00100101001100100", -- t[19044] = 1
      "0000001" when "00100101001100101", -- t[19045] = 1
      "0000001" when "00100101001100110", -- t[19046] = 1
      "0000001" when "00100101001100111", -- t[19047] = 1
      "0000001" when "00100101001101000", -- t[19048] = 1
      "0000001" when "00100101001101001", -- t[19049] = 1
      "0000001" when "00100101001101010", -- t[19050] = 1
      "0000001" when "00100101001101011", -- t[19051] = 1
      "0000001" when "00100101001101100", -- t[19052] = 1
      "0000001" when "00100101001101101", -- t[19053] = 1
      "0000001" when "00100101001101110", -- t[19054] = 1
      "0000001" when "00100101001101111", -- t[19055] = 1
      "0000001" when "00100101001110000", -- t[19056] = 1
      "0000001" when "00100101001110001", -- t[19057] = 1
      "0000001" when "00100101001110010", -- t[19058] = 1
      "0000001" when "00100101001110011", -- t[19059] = 1
      "0000001" when "00100101001110100", -- t[19060] = 1
      "0000001" when "00100101001110101", -- t[19061] = 1
      "0000001" when "00100101001110110", -- t[19062] = 1
      "0000001" when "00100101001110111", -- t[19063] = 1
      "0000001" when "00100101001111000", -- t[19064] = 1
      "0000001" when "00100101001111001", -- t[19065] = 1
      "0000001" when "00100101001111010", -- t[19066] = 1
      "0000001" when "00100101001111011", -- t[19067] = 1
      "0000001" when "00100101001111100", -- t[19068] = 1
      "0000001" when "00100101001111101", -- t[19069] = 1
      "0000001" when "00100101001111110", -- t[19070] = 1
      "0000001" when "00100101001111111", -- t[19071] = 1
      "0000001" when "00100101010000000", -- t[19072] = 1
      "0000001" when "00100101010000001", -- t[19073] = 1
      "0000001" when "00100101010000010", -- t[19074] = 1
      "0000001" when "00100101010000011", -- t[19075] = 1
      "0000001" when "00100101010000100", -- t[19076] = 1
      "0000001" when "00100101010000101", -- t[19077] = 1
      "0000001" when "00100101010000110", -- t[19078] = 1
      "0000001" when "00100101010000111", -- t[19079] = 1
      "0000001" when "00100101010001000", -- t[19080] = 1
      "0000001" when "00100101010001001", -- t[19081] = 1
      "0000001" when "00100101010001010", -- t[19082] = 1
      "0000001" when "00100101010001011", -- t[19083] = 1
      "0000001" when "00100101010001100", -- t[19084] = 1
      "0000001" when "00100101010001101", -- t[19085] = 1
      "0000001" when "00100101010001110", -- t[19086] = 1
      "0000001" when "00100101010001111", -- t[19087] = 1
      "0000001" when "00100101010010000", -- t[19088] = 1
      "0000001" when "00100101010010001", -- t[19089] = 1
      "0000001" when "00100101010010010", -- t[19090] = 1
      "0000001" when "00100101010010011", -- t[19091] = 1
      "0000001" when "00100101010010100", -- t[19092] = 1
      "0000001" when "00100101010010101", -- t[19093] = 1
      "0000001" when "00100101010010110", -- t[19094] = 1
      "0000001" when "00100101010010111", -- t[19095] = 1
      "0000001" when "00100101010011000", -- t[19096] = 1
      "0000001" when "00100101010011001", -- t[19097] = 1
      "0000001" when "00100101010011010", -- t[19098] = 1
      "0000001" when "00100101010011011", -- t[19099] = 1
      "0000001" when "00100101010011100", -- t[19100] = 1
      "0000001" when "00100101010011101", -- t[19101] = 1
      "0000001" when "00100101010011110", -- t[19102] = 1
      "0000001" when "00100101010011111", -- t[19103] = 1
      "0000001" when "00100101010100000", -- t[19104] = 1
      "0000001" when "00100101010100001", -- t[19105] = 1
      "0000001" when "00100101010100010", -- t[19106] = 1
      "0000001" when "00100101010100011", -- t[19107] = 1
      "0000001" when "00100101010100100", -- t[19108] = 1
      "0000001" when "00100101010100101", -- t[19109] = 1
      "0000001" when "00100101010100110", -- t[19110] = 1
      "0000001" when "00100101010100111", -- t[19111] = 1
      "0000001" when "00100101010101000", -- t[19112] = 1
      "0000001" when "00100101010101001", -- t[19113] = 1
      "0000001" when "00100101010101010", -- t[19114] = 1
      "0000001" when "00100101010101011", -- t[19115] = 1
      "0000001" when "00100101010101100", -- t[19116] = 1
      "0000001" when "00100101010101101", -- t[19117] = 1
      "0000001" when "00100101010101110", -- t[19118] = 1
      "0000001" when "00100101010101111", -- t[19119] = 1
      "0000001" when "00100101010110000", -- t[19120] = 1
      "0000001" when "00100101010110001", -- t[19121] = 1
      "0000001" when "00100101010110010", -- t[19122] = 1
      "0000001" when "00100101010110011", -- t[19123] = 1
      "0000001" when "00100101010110100", -- t[19124] = 1
      "0000001" when "00100101010110101", -- t[19125] = 1
      "0000001" when "00100101010110110", -- t[19126] = 1
      "0000001" when "00100101010110111", -- t[19127] = 1
      "0000001" when "00100101010111000", -- t[19128] = 1
      "0000001" when "00100101010111001", -- t[19129] = 1
      "0000001" when "00100101010111010", -- t[19130] = 1
      "0000001" when "00100101010111011", -- t[19131] = 1
      "0000001" when "00100101010111100", -- t[19132] = 1
      "0000001" when "00100101010111101", -- t[19133] = 1
      "0000001" when "00100101010111110", -- t[19134] = 1
      "0000001" when "00100101010111111", -- t[19135] = 1
      "0000001" when "00100101011000000", -- t[19136] = 1
      "0000001" when "00100101011000001", -- t[19137] = 1
      "0000001" when "00100101011000010", -- t[19138] = 1
      "0000001" when "00100101011000011", -- t[19139] = 1
      "0000001" when "00100101011000100", -- t[19140] = 1
      "0000001" when "00100101011000101", -- t[19141] = 1
      "0000001" when "00100101011000110", -- t[19142] = 1
      "0000001" when "00100101011000111", -- t[19143] = 1
      "0000001" when "00100101011001000", -- t[19144] = 1
      "0000001" when "00100101011001001", -- t[19145] = 1
      "0000001" when "00100101011001010", -- t[19146] = 1
      "0000001" when "00100101011001011", -- t[19147] = 1
      "0000001" when "00100101011001100", -- t[19148] = 1
      "0000001" when "00100101011001101", -- t[19149] = 1
      "0000001" when "00100101011001110", -- t[19150] = 1
      "0000001" when "00100101011001111", -- t[19151] = 1
      "0000001" when "00100101011010000", -- t[19152] = 1
      "0000001" when "00100101011010001", -- t[19153] = 1
      "0000001" when "00100101011010010", -- t[19154] = 1
      "0000001" when "00100101011010011", -- t[19155] = 1
      "0000001" when "00100101011010100", -- t[19156] = 1
      "0000001" when "00100101011010101", -- t[19157] = 1
      "0000001" when "00100101011010110", -- t[19158] = 1
      "0000001" when "00100101011010111", -- t[19159] = 1
      "0000001" when "00100101011011000", -- t[19160] = 1
      "0000001" when "00100101011011001", -- t[19161] = 1
      "0000001" when "00100101011011010", -- t[19162] = 1
      "0000001" when "00100101011011011", -- t[19163] = 1
      "0000001" when "00100101011011100", -- t[19164] = 1
      "0000001" when "00100101011011101", -- t[19165] = 1
      "0000001" when "00100101011011110", -- t[19166] = 1
      "0000001" when "00100101011011111", -- t[19167] = 1
      "0000001" when "00100101011100000", -- t[19168] = 1
      "0000001" when "00100101011100001", -- t[19169] = 1
      "0000001" when "00100101011100010", -- t[19170] = 1
      "0000001" when "00100101011100011", -- t[19171] = 1
      "0000001" when "00100101011100100", -- t[19172] = 1
      "0000001" when "00100101011100101", -- t[19173] = 1
      "0000001" when "00100101011100110", -- t[19174] = 1
      "0000001" when "00100101011100111", -- t[19175] = 1
      "0000001" when "00100101011101000", -- t[19176] = 1
      "0000001" when "00100101011101001", -- t[19177] = 1
      "0000001" when "00100101011101010", -- t[19178] = 1
      "0000001" when "00100101011101011", -- t[19179] = 1
      "0000001" when "00100101011101100", -- t[19180] = 1
      "0000001" when "00100101011101101", -- t[19181] = 1
      "0000001" when "00100101011101110", -- t[19182] = 1
      "0000001" when "00100101011101111", -- t[19183] = 1
      "0000001" when "00100101011110000", -- t[19184] = 1
      "0000001" when "00100101011110001", -- t[19185] = 1
      "0000001" when "00100101011110010", -- t[19186] = 1
      "0000001" when "00100101011110011", -- t[19187] = 1
      "0000001" when "00100101011110100", -- t[19188] = 1
      "0000001" when "00100101011110101", -- t[19189] = 1
      "0000001" when "00100101011110110", -- t[19190] = 1
      "0000001" when "00100101011110111", -- t[19191] = 1
      "0000001" when "00100101011111000", -- t[19192] = 1
      "0000001" when "00100101011111001", -- t[19193] = 1
      "0000001" when "00100101011111010", -- t[19194] = 1
      "0000001" when "00100101011111011", -- t[19195] = 1
      "0000001" when "00100101011111100", -- t[19196] = 1
      "0000001" when "00100101011111101", -- t[19197] = 1
      "0000001" when "00100101011111110", -- t[19198] = 1
      "0000001" when "00100101011111111", -- t[19199] = 1
      "0000001" when "00100101100000000", -- t[19200] = 1
      "0000001" when "00100101100000001", -- t[19201] = 1
      "0000001" when "00100101100000010", -- t[19202] = 1
      "0000001" when "00100101100000011", -- t[19203] = 1
      "0000001" when "00100101100000100", -- t[19204] = 1
      "0000001" when "00100101100000101", -- t[19205] = 1
      "0000001" when "00100101100000110", -- t[19206] = 1
      "0000001" when "00100101100000111", -- t[19207] = 1
      "0000001" when "00100101100001000", -- t[19208] = 1
      "0000001" when "00100101100001001", -- t[19209] = 1
      "0000001" when "00100101100001010", -- t[19210] = 1
      "0000001" when "00100101100001011", -- t[19211] = 1
      "0000001" when "00100101100001100", -- t[19212] = 1
      "0000001" when "00100101100001101", -- t[19213] = 1
      "0000001" when "00100101100001110", -- t[19214] = 1
      "0000001" when "00100101100001111", -- t[19215] = 1
      "0000001" when "00100101100010000", -- t[19216] = 1
      "0000001" when "00100101100010001", -- t[19217] = 1
      "0000001" when "00100101100010010", -- t[19218] = 1
      "0000001" when "00100101100010011", -- t[19219] = 1
      "0000001" when "00100101100010100", -- t[19220] = 1
      "0000001" when "00100101100010101", -- t[19221] = 1
      "0000001" when "00100101100010110", -- t[19222] = 1
      "0000001" when "00100101100010111", -- t[19223] = 1
      "0000001" when "00100101100011000", -- t[19224] = 1
      "0000001" when "00100101100011001", -- t[19225] = 1
      "0000001" when "00100101100011010", -- t[19226] = 1
      "0000001" when "00100101100011011", -- t[19227] = 1
      "0000001" when "00100101100011100", -- t[19228] = 1
      "0000001" when "00100101100011101", -- t[19229] = 1
      "0000001" when "00100101100011110", -- t[19230] = 1
      "0000001" when "00100101100011111", -- t[19231] = 1
      "0000001" when "00100101100100000", -- t[19232] = 1
      "0000001" when "00100101100100001", -- t[19233] = 1
      "0000001" when "00100101100100010", -- t[19234] = 1
      "0000001" when "00100101100100011", -- t[19235] = 1
      "0000001" when "00100101100100100", -- t[19236] = 1
      "0000001" when "00100101100100101", -- t[19237] = 1
      "0000001" when "00100101100100110", -- t[19238] = 1
      "0000001" when "00100101100100111", -- t[19239] = 1
      "0000001" when "00100101100101000", -- t[19240] = 1
      "0000001" when "00100101100101001", -- t[19241] = 1
      "0000001" when "00100101100101010", -- t[19242] = 1
      "0000001" when "00100101100101011", -- t[19243] = 1
      "0000001" when "00100101100101100", -- t[19244] = 1
      "0000001" when "00100101100101101", -- t[19245] = 1
      "0000001" when "00100101100101110", -- t[19246] = 1
      "0000001" when "00100101100101111", -- t[19247] = 1
      "0000001" when "00100101100110000", -- t[19248] = 1
      "0000001" when "00100101100110001", -- t[19249] = 1
      "0000001" when "00100101100110010", -- t[19250] = 1
      "0000001" when "00100101100110011", -- t[19251] = 1
      "0000001" when "00100101100110100", -- t[19252] = 1
      "0000001" when "00100101100110101", -- t[19253] = 1
      "0000001" when "00100101100110110", -- t[19254] = 1
      "0000001" when "00100101100110111", -- t[19255] = 1
      "0000001" when "00100101100111000", -- t[19256] = 1
      "0000001" when "00100101100111001", -- t[19257] = 1
      "0000001" when "00100101100111010", -- t[19258] = 1
      "0000001" when "00100101100111011", -- t[19259] = 1
      "0000001" when "00100101100111100", -- t[19260] = 1
      "0000001" when "00100101100111101", -- t[19261] = 1
      "0000001" when "00100101100111110", -- t[19262] = 1
      "0000001" when "00100101100111111", -- t[19263] = 1
      "0000001" when "00100101101000000", -- t[19264] = 1
      "0000001" when "00100101101000001", -- t[19265] = 1
      "0000001" when "00100101101000010", -- t[19266] = 1
      "0000001" when "00100101101000011", -- t[19267] = 1
      "0000001" when "00100101101000100", -- t[19268] = 1
      "0000001" when "00100101101000101", -- t[19269] = 1
      "0000001" when "00100101101000110", -- t[19270] = 1
      "0000001" when "00100101101000111", -- t[19271] = 1
      "0000001" when "00100101101001000", -- t[19272] = 1
      "0000001" when "00100101101001001", -- t[19273] = 1
      "0000001" when "00100101101001010", -- t[19274] = 1
      "0000001" when "00100101101001011", -- t[19275] = 1
      "0000001" when "00100101101001100", -- t[19276] = 1
      "0000001" when "00100101101001101", -- t[19277] = 1
      "0000001" when "00100101101001110", -- t[19278] = 1
      "0000001" when "00100101101001111", -- t[19279] = 1
      "0000001" when "00100101101010000", -- t[19280] = 1
      "0000001" when "00100101101010001", -- t[19281] = 1
      "0000001" when "00100101101010010", -- t[19282] = 1
      "0000001" when "00100101101010011", -- t[19283] = 1
      "0000001" when "00100101101010100", -- t[19284] = 1
      "0000001" when "00100101101010101", -- t[19285] = 1
      "0000001" when "00100101101010110", -- t[19286] = 1
      "0000001" when "00100101101010111", -- t[19287] = 1
      "0000001" when "00100101101011000", -- t[19288] = 1
      "0000001" when "00100101101011001", -- t[19289] = 1
      "0000001" when "00100101101011010", -- t[19290] = 1
      "0000001" when "00100101101011011", -- t[19291] = 1
      "0000001" when "00100101101011100", -- t[19292] = 1
      "0000001" when "00100101101011101", -- t[19293] = 1
      "0000001" when "00100101101011110", -- t[19294] = 1
      "0000001" when "00100101101011111", -- t[19295] = 1
      "0000001" when "00100101101100000", -- t[19296] = 1
      "0000001" when "00100101101100001", -- t[19297] = 1
      "0000001" when "00100101101100010", -- t[19298] = 1
      "0000001" when "00100101101100011", -- t[19299] = 1
      "0000001" when "00100101101100100", -- t[19300] = 1
      "0000001" when "00100101101100101", -- t[19301] = 1
      "0000001" when "00100101101100110", -- t[19302] = 1
      "0000001" when "00100101101100111", -- t[19303] = 1
      "0000001" when "00100101101101000", -- t[19304] = 1
      "0000001" when "00100101101101001", -- t[19305] = 1
      "0000001" when "00100101101101010", -- t[19306] = 1
      "0000001" when "00100101101101011", -- t[19307] = 1
      "0000001" when "00100101101101100", -- t[19308] = 1
      "0000001" when "00100101101101101", -- t[19309] = 1
      "0000001" when "00100101101101110", -- t[19310] = 1
      "0000001" when "00100101101101111", -- t[19311] = 1
      "0000001" when "00100101101110000", -- t[19312] = 1
      "0000001" when "00100101101110001", -- t[19313] = 1
      "0000001" when "00100101101110010", -- t[19314] = 1
      "0000001" when "00100101101110011", -- t[19315] = 1
      "0000001" when "00100101101110100", -- t[19316] = 1
      "0000001" when "00100101101110101", -- t[19317] = 1
      "0000001" when "00100101101110110", -- t[19318] = 1
      "0000001" when "00100101101110111", -- t[19319] = 1
      "0000001" when "00100101101111000", -- t[19320] = 1
      "0000001" when "00100101101111001", -- t[19321] = 1
      "0000001" when "00100101101111010", -- t[19322] = 1
      "0000001" when "00100101101111011", -- t[19323] = 1
      "0000001" when "00100101101111100", -- t[19324] = 1
      "0000001" when "00100101101111101", -- t[19325] = 1
      "0000001" when "00100101101111110", -- t[19326] = 1
      "0000001" when "00100101101111111", -- t[19327] = 1
      "0000001" when "00100101110000000", -- t[19328] = 1
      "0000001" when "00100101110000001", -- t[19329] = 1
      "0000001" when "00100101110000010", -- t[19330] = 1
      "0000001" when "00100101110000011", -- t[19331] = 1
      "0000001" when "00100101110000100", -- t[19332] = 1
      "0000001" when "00100101110000101", -- t[19333] = 1
      "0000001" when "00100101110000110", -- t[19334] = 1
      "0000001" when "00100101110000111", -- t[19335] = 1
      "0000001" when "00100101110001000", -- t[19336] = 1
      "0000001" when "00100101110001001", -- t[19337] = 1
      "0000001" when "00100101110001010", -- t[19338] = 1
      "0000001" when "00100101110001011", -- t[19339] = 1
      "0000001" when "00100101110001100", -- t[19340] = 1
      "0000001" when "00100101110001101", -- t[19341] = 1
      "0000001" when "00100101110001110", -- t[19342] = 1
      "0000001" when "00100101110001111", -- t[19343] = 1
      "0000001" when "00100101110010000", -- t[19344] = 1
      "0000001" when "00100101110010001", -- t[19345] = 1
      "0000001" when "00100101110010010", -- t[19346] = 1
      "0000001" when "00100101110010011", -- t[19347] = 1
      "0000001" when "00100101110010100", -- t[19348] = 1
      "0000001" when "00100101110010101", -- t[19349] = 1
      "0000001" when "00100101110010110", -- t[19350] = 1
      "0000001" when "00100101110010111", -- t[19351] = 1
      "0000001" when "00100101110011000", -- t[19352] = 1
      "0000001" when "00100101110011001", -- t[19353] = 1
      "0000001" when "00100101110011010", -- t[19354] = 1
      "0000001" when "00100101110011011", -- t[19355] = 1
      "0000001" when "00100101110011100", -- t[19356] = 1
      "0000001" when "00100101110011101", -- t[19357] = 1
      "0000001" when "00100101110011110", -- t[19358] = 1
      "0000001" when "00100101110011111", -- t[19359] = 1
      "0000001" when "00100101110100000", -- t[19360] = 1
      "0000001" when "00100101110100001", -- t[19361] = 1
      "0000001" when "00100101110100010", -- t[19362] = 1
      "0000001" when "00100101110100011", -- t[19363] = 1
      "0000001" when "00100101110100100", -- t[19364] = 1
      "0000001" when "00100101110100101", -- t[19365] = 1
      "0000001" when "00100101110100110", -- t[19366] = 1
      "0000001" when "00100101110100111", -- t[19367] = 1
      "0000001" when "00100101110101000", -- t[19368] = 1
      "0000001" when "00100101110101001", -- t[19369] = 1
      "0000001" when "00100101110101010", -- t[19370] = 1
      "0000001" when "00100101110101011", -- t[19371] = 1
      "0000001" when "00100101110101100", -- t[19372] = 1
      "0000001" when "00100101110101101", -- t[19373] = 1
      "0000001" when "00100101110101110", -- t[19374] = 1
      "0000001" when "00100101110101111", -- t[19375] = 1
      "0000001" when "00100101110110000", -- t[19376] = 1
      "0000001" when "00100101110110001", -- t[19377] = 1
      "0000001" when "00100101110110010", -- t[19378] = 1
      "0000001" when "00100101110110011", -- t[19379] = 1
      "0000001" when "00100101110110100", -- t[19380] = 1
      "0000001" when "00100101110110101", -- t[19381] = 1
      "0000001" when "00100101110110110", -- t[19382] = 1
      "0000001" when "00100101110110111", -- t[19383] = 1
      "0000001" when "00100101110111000", -- t[19384] = 1
      "0000001" when "00100101110111001", -- t[19385] = 1
      "0000001" when "00100101110111010", -- t[19386] = 1
      "0000001" when "00100101110111011", -- t[19387] = 1
      "0000001" when "00100101110111100", -- t[19388] = 1
      "0000001" when "00100101110111101", -- t[19389] = 1
      "0000001" when "00100101110111110", -- t[19390] = 1
      "0000001" when "00100101110111111", -- t[19391] = 1
      "0000001" when "00100101111000000", -- t[19392] = 1
      "0000001" when "00100101111000001", -- t[19393] = 1
      "0000001" when "00100101111000010", -- t[19394] = 1
      "0000001" when "00100101111000011", -- t[19395] = 1
      "0000001" when "00100101111000100", -- t[19396] = 1
      "0000001" when "00100101111000101", -- t[19397] = 1
      "0000001" when "00100101111000110", -- t[19398] = 1
      "0000001" when "00100101111000111", -- t[19399] = 1
      "0000001" when "00100101111001000", -- t[19400] = 1
      "0000001" when "00100101111001001", -- t[19401] = 1
      "0000001" when "00100101111001010", -- t[19402] = 1
      "0000001" when "00100101111001011", -- t[19403] = 1
      "0000001" when "00100101111001100", -- t[19404] = 1
      "0000001" when "00100101111001101", -- t[19405] = 1
      "0000001" when "00100101111001110", -- t[19406] = 1
      "0000001" when "00100101111001111", -- t[19407] = 1
      "0000001" when "00100101111010000", -- t[19408] = 1
      "0000001" when "00100101111010001", -- t[19409] = 1
      "0000001" when "00100101111010010", -- t[19410] = 1
      "0000001" when "00100101111010011", -- t[19411] = 1
      "0000001" when "00100101111010100", -- t[19412] = 1
      "0000001" when "00100101111010101", -- t[19413] = 1
      "0000001" when "00100101111010110", -- t[19414] = 1
      "0000001" when "00100101111010111", -- t[19415] = 1
      "0000001" when "00100101111011000", -- t[19416] = 1
      "0000001" when "00100101111011001", -- t[19417] = 1
      "0000001" when "00100101111011010", -- t[19418] = 1
      "0000001" when "00100101111011011", -- t[19419] = 1
      "0000001" when "00100101111011100", -- t[19420] = 1
      "0000001" when "00100101111011101", -- t[19421] = 1
      "0000001" when "00100101111011110", -- t[19422] = 1
      "0000001" when "00100101111011111", -- t[19423] = 1
      "0000001" when "00100101111100000", -- t[19424] = 1
      "0000001" when "00100101111100001", -- t[19425] = 1
      "0000001" when "00100101111100010", -- t[19426] = 1
      "0000001" when "00100101111100011", -- t[19427] = 1
      "0000001" when "00100101111100100", -- t[19428] = 1
      "0000001" when "00100101111100101", -- t[19429] = 1
      "0000001" when "00100101111100110", -- t[19430] = 1
      "0000001" when "00100101111100111", -- t[19431] = 1
      "0000001" when "00100101111101000", -- t[19432] = 1
      "0000001" when "00100101111101001", -- t[19433] = 1
      "0000001" when "00100101111101010", -- t[19434] = 1
      "0000001" when "00100101111101011", -- t[19435] = 1
      "0000001" when "00100101111101100", -- t[19436] = 1
      "0000001" when "00100101111101101", -- t[19437] = 1
      "0000001" when "00100101111101110", -- t[19438] = 1
      "0000001" when "00100101111101111", -- t[19439] = 1
      "0000001" when "00100101111110000", -- t[19440] = 1
      "0000001" when "00100101111110001", -- t[19441] = 1
      "0000001" when "00100101111110010", -- t[19442] = 1
      "0000001" when "00100101111110011", -- t[19443] = 1
      "0000001" when "00100101111110100", -- t[19444] = 1
      "0000001" when "00100101111110101", -- t[19445] = 1
      "0000001" when "00100101111110110", -- t[19446] = 1
      "0000001" when "00100101111110111", -- t[19447] = 1
      "0000001" when "00100101111111000", -- t[19448] = 1
      "0000001" when "00100101111111001", -- t[19449] = 1
      "0000001" when "00100101111111010", -- t[19450] = 1
      "0000001" when "00100101111111011", -- t[19451] = 1
      "0000001" when "00100101111111100", -- t[19452] = 1
      "0000001" when "00100101111111101", -- t[19453] = 1
      "0000001" when "00100101111111110", -- t[19454] = 1
      "0000001" when "00100101111111111", -- t[19455] = 1
      "0000001" when "00100110000000000", -- t[19456] = 1
      "0000001" when "00100110000000001", -- t[19457] = 1
      "0000001" when "00100110000000010", -- t[19458] = 1
      "0000001" when "00100110000000011", -- t[19459] = 1
      "0000001" when "00100110000000100", -- t[19460] = 1
      "0000001" when "00100110000000101", -- t[19461] = 1
      "0000001" when "00100110000000110", -- t[19462] = 1
      "0000001" when "00100110000000111", -- t[19463] = 1
      "0000001" when "00100110000001000", -- t[19464] = 1
      "0000001" when "00100110000001001", -- t[19465] = 1
      "0000001" when "00100110000001010", -- t[19466] = 1
      "0000001" when "00100110000001011", -- t[19467] = 1
      "0000001" when "00100110000001100", -- t[19468] = 1
      "0000001" when "00100110000001101", -- t[19469] = 1
      "0000001" when "00100110000001110", -- t[19470] = 1
      "0000001" when "00100110000001111", -- t[19471] = 1
      "0000001" when "00100110000010000", -- t[19472] = 1
      "0000001" when "00100110000010001", -- t[19473] = 1
      "0000001" when "00100110000010010", -- t[19474] = 1
      "0000001" when "00100110000010011", -- t[19475] = 1
      "0000001" when "00100110000010100", -- t[19476] = 1
      "0000001" when "00100110000010101", -- t[19477] = 1
      "0000001" when "00100110000010110", -- t[19478] = 1
      "0000001" when "00100110000010111", -- t[19479] = 1
      "0000001" when "00100110000011000", -- t[19480] = 1
      "0000001" when "00100110000011001", -- t[19481] = 1
      "0000001" when "00100110000011010", -- t[19482] = 1
      "0000001" when "00100110000011011", -- t[19483] = 1
      "0000001" when "00100110000011100", -- t[19484] = 1
      "0000001" when "00100110000011101", -- t[19485] = 1
      "0000001" when "00100110000011110", -- t[19486] = 1
      "0000001" when "00100110000011111", -- t[19487] = 1
      "0000001" when "00100110000100000", -- t[19488] = 1
      "0000001" when "00100110000100001", -- t[19489] = 1
      "0000001" when "00100110000100010", -- t[19490] = 1
      "0000001" when "00100110000100011", -- t[19491] = 1
      "0000001" when "00100110000100100", -- t[19492] = 1
      "0000001" when "00100110000100101", -- t[19493] = 1
      "0000001" when "00100110000100110", -- t[19494] = 1
      "0000001" when "00100110000100111", -- t[19495] = 1
      "0000001" when "00100110000101000", -- t[19496] = 1
      "0000001" when "00100110000101001", -- t[19497] = 1
      "0000001" when "00100110000101010", -- t[19498] = 1
      "0000001" when "00100110000101011", -- t[19499] = 1
      "0000001" when "00100110000101100", -- t[19500] = 1
      "0000001" when "00100110000101101", -- t[19501] = 1
      "0000001" when "00100110000101110", -- t[19502] = 1
      "0000001" when "00100110000101111", -- t[19503] = 1
      "0000001" when "00100110000110000", -- t[19504] = 1
      "0000001" when "00100110000110001", -- t[19505] = 1
      "0000001" when "00100110000110010", -- t[19506] = 1
      "0000001" when "00100110000110011", -- t[19507] = 1
      "0000001" when "00100110000110100", -- t[19508] = 1
      "0000001" when "00100110000110101", -- t[19509] = 1
      "0000001" when "00100110000110110", -- t[19510] = 1
      "0000001" when "00100110000110111", -- t[19511] = 1
      "0000001" when "00100110000111000", -- t[19512] = 1
      "0000001" when "00100110000111001", -- t[19513] = 1
      "0000001" when "00100110000111010", -- t[19514] = 1
      "0000001" when "00100110000111011", -- t[19515] = 1
      "0000001" when "00100110000111100", -- t[19516] = 1
      "0000001" when "00100110000111101", -- t[19517] = 1
      "0000001" when "00100110000111110", -- t[19518] = 1
      "0000001" when "00100110000111111", -- t[19519] = 1
      "0000001" when "00100110001000000", -- t[19520] = 1
      "0000001" when "00100110001000001", -- t[19521] = 1
      "0000001" when "00100110001000010", -- t[19522] = 1
      "0000001" when "00100110001000011", -- t[19523] = 1
      "0000001" when "00100110001000100", -- t[19524] = 1
      "0000001" when "00100110001000101", -- t[19525] = 1
      "0000001" when "00100110001000110", -- t[19526] = 1
      "0000001" when "00100110001000111", -- t[19527] = 1
      "0000001" when "00100110001001000", -- t[19528] = 1
      "0000001" when "00100110001001001", -- t[19529] = 1
      "0000001" when "00100110001001010", -- t[19530] = 1
      "0000001" when "00100110001001011", -- t[19531] = 1
      "0000001" when "00100110001001100", -- t[19532] = 1
      "0000001" when "00100110001001101", -- t[19533] = 1
      "0000001" when "00100110001001110", -- t[19534] = 1
      "0000001" when "00100110001001111", -- t[19535] = 1
      "0000001" when "00100110001010000", -- t[19536] = 1
      "0000001" when "00100110001010001", -- t[19537] = 1
      "0000001" when "00100110001010010", -- t[19538] = 1
      "0000001" when "00100110001010011", -- t[19539] = 1
      "0000001" when "00100110001010100", -- t[19540] = 1
      "0000001" when "00100110001010101", -- t[19541] = 1
      "0000001" when "00100110001010110", -- t[19542] = 1
      "0000001" when "00100110001010111", -- t[19543] = 1
      "0000001" when "00100110001011000", -- t[19544] = 1
      "0000001" when "00100110001011001", -- t[19545] = 1
      "0000001" when "00100110001011010", -- t[19546] = 1
      "0000001" when "00100110001011011", -- t[19547] = 1
      "0000001" when "00100110001011100", -- t[19548] = 1
      "0000001" when "00100110001011101", -- t[19549] = 1
      "0000001" when "00100110001011110", -- t[19550] = 1
      "0000001" when "00100110001011111", -- t[19551] = 1
      "0000001" when "00100110001100000", -- t[19552] = 1
      "0000001" when "00100110001100001", -- t[19553] = 1
      "0000001" when "00100110001100010", -- t[19554] = 1
      "0000001" when "00100110001100011", -- t[19555] = 1
      "0000001" when "00100110001100100", -- t[19556] = 1
      "0000001" when "00100110001100101", -- t[19557] = 1
      "0000001" when "00100110001100110", -- t[19558] = 1
      "0000001" when "00100110001100111", -- t[19559] = 1
      "0000001" when "00100110001101000", -- t[19560] = 1
      "0000001" when "00100110001101001", -- t[19561] = 1
      "0000001" when "00100110001101010", -- t[19562] = 1
      "0000001" when "00100110001101011", -- t[19563] = 1
      "0000001" when "00100110001101100", -- t[19564] = 1
      "0000001" when "00100110001101101", -- t[19565] = 1
      "0000001" when "00100110001101110", -- t[19566] = 1
      "0000001" when "00100110001101111", -- t[19567] = 1
      "0000001" when "00100110001110000", -- t[19568] = 1
      "0000001" when "00100110001110001", -- t[19569] = 1
      "0000001" when "00100110001110010", -- t[19570] = 1
      "0000001" when "00100110001110011", -- t[19571] = 1
      "0000001" when "00100110001110100", -- t[19572] = 1
      "0000001" when "00100110001110101", -- t[19573] = 1
      "0000001" when "00100110001110110", -- t[19574] = 1
      "0000001" when "00100110001110111", -- t[19575] = 1
      "0000001" when "00100110001111000", -- t[19576] = 1
      "0000001" when "00100110001111001", -- t[19577] = 1
      "0000001" when "00100110001111010", -- t[19578] = 1
      "0000001" when "00100110001111011", -- t[19579] = 1
      "0000001" when "00100110001111100", -- t[19580] = 1
      "0000001" when "00100110001111101", -- t[19581] = 1
      "0000001" when "00100110001111110", -- t[19582] = 1
      "0000001" when "00100110001111111", -- t[19583] = 1
      "0000001" when "00100110010000000", -- t[19584] = 1
      "0000001" when "00100110010000001", -- t[19585] = 1
      "0000001" when "00100110010000010", -- t[19586] = 1
      "0000001" when "00100110010000011", -- t[19587] = 1
      "0000001" when "00100110010000100", -- t[19588] = 1
      "0000001" when "00100110010000101", -- t[19589] = 1
      "0000001" when "00100110010000110", -- t[19590] = 1
      "0000001" when "00100110010000111", -- t[19591] = 1
      "0000001" when "00100110010001000", -- t[19592] = 1
      "0000001" when "00100110010001001", -- t[19593] = 1
      "0000001" when "00100110010001010", -- t[19594] = 1
      "0000001" when "00100110010001011", -- t[19595] = 1
      "0000001" when "00100110010001100", -- t[19596] = 1
      "0000001" when "00100110010001101", -- t[19597] = 1
      "0000001" when "00100110010001110", -- t[19598] = 1
      "0000001" when "00100110010001111", -- t[19599] = 1
      "0000001" when "00100110010010000", -- t[19600] = 1
      "0000001" when "00100110010010001", -- t[19601] = 1
      "0000001" when "00100110010010010", -- t[19602] = 1
      "0000001" when "00100110010010011", -- t[19603] = 1
      "0000001" when "00100110010010100", -- t[19604] = 1
      "0000001" when "00100110010010101", -- t[19605] = 1
      "0000001" when "00100110010010110", -- t[19606] = 1
      "0000001" when "00100110010010111", -- t[19607] = 1
      "0000001" when "00100110010011000", -- t[19608] = 1
      "0000001" when "00100110010011001", -- t[19609] = 1
      "0000001" when "00100110010011010", -- t[19610] = 1
      "0000001" when "00100110010011011", -- t[19611] = 1
      "0000001" when "00100110010011100", -- t[19612] = 1
      "0000001" when "00100110010011101", -- t[19613] = 1
      "0000001" when "00100110010011110", -- t[19614] = 1
      "0000001" when "00100110010011111", -- t[19615] = 1
      "0000001" when "00100110010100000", -- t[19616] = 1
      "0000001" when "00100110010100001", -- t[19617] = 1
      "0000001" when "00100110010100010", -- t[19618] = 1
      "0000001" when "00100110010100011", -- t[19619] = 1
      "0000001" when "00100110010100100", -- t[19620] = 1
      "0000001" when "00100110010100101", -- t[19621] = 1
      "0000001" when "00100110010100110", -- t[19622] = 1
      "0000001" when "00100110010100111", -- t[19623] = 1
      "0000001" when "00100110010101000", -- t[19624] = 1
      "0000001" when "00100110010101001", -- t[19625] = 1
      "0000001" when "00100110010101010", -- t[19626] = 1
      "0000001" when "00100110010101011", -- t[19627] = 1
      "0000001" when "00100110010101100", -- t[19628] = 1
      "0000001" when "00100110010101101", -- t[19629] = 1
      "0000001" when "00100110010101110", -- t[19630] = 1
      "0000001" when "00100110010101111", -- t[19631] = 1
      "0000001" when "00100110010110000", -- t[19632] = 1
      "0000001" when "00100110010110001", -- t[19633] = 1
      "0000001" when "00100110010110010", -- t[19634] = 1
      "0000001" when "00100110010110011", -- t[19635] = 1
      "0000001" when "00100110010110100", -- t[19636] = 1
      "0000001" when "00100110010110101", -- t[19637] = 1
      "0000001" when "00100110010110110", -- t[19638] = 1
      "0000001" when "00100110010110111", -- t[19639] = 1
      "0000001" when "00100110010111000", -- t[19640] = 1
      "0000001" when "00100110010111001", -- t[19641] = 1
      "0000001" when "00100110010111010", -- t[19642] = 1
      "0000001" when "00100110010111011", -- t[19643] = 1
      "0000001" when "00100110010111100", -- t[19644] = 1
      "0000001" when "00100110010111101", -- t[19645] = 1
      "0000001" when "00100110010111110", -- t[19646] = 1
      "0000001" when "00100110010111111", -- t[19647] = 1
      "0000001" when "00100110011000000", -- t[19648] = 1
      "0000001" when "00100110011000001", -- t[19649] = 1
      "0000001" when "00100110011000010", -- t[19650] = 1
      "0000001" when "00100110011000011", -- t[19651] = 1
      "0000001" when "00100110011000100", -- t[19652] = 1
      "0000001" when "00100110011000101", -- t[19653] = 1
      "0000001" when "00100110011000110", -- t[19654] = 1
      "0000001" when "00100110011000111", -- t[19655] = 1
      "0000001" when "00100110011001000", -- t[19656] = 1
      "0000001" when "00100110011001001", -- t[19657] = 1
      "0000001" when "00100110011001010", -- t[19658] = 1
      "0000001" when "00100110011001011", -- t[19659] = 1
      "0000001" when "00100110011001100", -- t[19660] = 1
      "0000001" when "00100110011001101", -- t[19661] = 1
      "0000001" when "00100110011001110", -- t[19662] = 1
      "0000001" when "00100110011001111", -- t[19663] = 1
      "0000001" when "00100110011010000", -- t[19664] = 1
      "0000001" when "00100110011010001", -- t[19665] = 1
      "0000001" when "00100110011010010", -- t[19666] = 1
      "0000001" when "00100110011010011", -- t[19667] = 1
      "0000001" when "00100110011010100", -- t[19668] = 1
      "0000001" when "00100110011010101", -- t[19669] = 1
      "0000001" when "00100110011010110", -- t[19670] = 1
      "0000001" when "00100110011010111", -- t[19671] = 1
      "0000001" when "00100110011011000", -- t[19672] = 1
      "0000001" when "00100110011011001", -- t[19673] = 1
      "0000001" when "00100110011011010", -- t[19674] = 1
      "0000001" when "00100110011011011", -- t[19675] = 1
      "0000001" when "00100110011011100", -- t[19676] = 1
      "0000001" when "00100110011011101", -- t[19677] = 1
      "0000001" when "00100110011011110", -- t[19678] = 1
      "0000001" when "00100110011011111", -- t[19679] = 1
      "0000001" when "00100110011100000", -- t[19680] = 1
      "0000001" when "00100110011100001", -- t[19681] = 1
      "0000001" when "00100110011100010", -- t[19682] = 1
      "0000001" when "00100110011100011", -- t[19683] = 1
      "0000001" when "00100110011100100", -- t[19684] = 1
      "0000001" when "00100110011100101", -- t[19685] = 1
      "0000001" when "00100110011100110", -- t[19686] = 1
      "0000001" when "00100110011100111", -- t[19687] = 1
      "0000001" when "00100110011101000", -- t[19688] = 1
      "0000001" when "00100110011101001", -- t[19689] = 1
      "0000001" when "00100110011101010", -- t[19690] = 1
      "0000001" when "00100110011101011", -- t[19691] = 1
      "0000001" when "00100110011101100", -- t[19692] = 1
      "0000001" when "00100110011101101", -- t[19693] = 1
      "0000001" when "00100110011101110", -- t[19694] = 1
      "0000001" when "00100110011101111", -- t[19695] = 1
      "0000001" when "00100110011110000", -- t[19696] = 1
      "0000001" when "00100110011110001", -- t[19697] = 1
      "0000001" when "00100110011110010", -- t[19698] = 1
      "0000001" when "00100110011110011", -- t[19699] = 1
      "0000001" when "00100110011110100", -- t[19700] = 1
      "0000001" when "00100110011110101", -- t[19701] = 1
      "0000001" when "00100110011110110", -- t[19702] = 1
      "0000001" when "00100110011110111", -- t[19703] = 1
      "0000001" when "00100110011111000", -- t[19704] = 1
      "0000001" when "00100110011111001", -- t[19705] = 1
      "0000001" when "00100110011111010", -- t[19706] = 1
      "0000001" when "00100110011111011", -- t[19707] = 1
      "0000001" when "00100110011111100", -- t[19708] = 1
      "0000001" when "00100110011111101", -- t[19709] = 1
      "0000001" when "00100110011111110", -- t[19710] = 1
      "0000001" when "00100110011111111", -- t[19711] = 1
      "0000001" when "00100110100000000", -- t[19712] = 1
      "0000001" when "00100110100000001", -- t[19713] = 1
      "0000001" when "00100110100000010", -- t[19714] = 1
      "0000001" when "00100110100000011", -- t[19715] = 1
      "0000001" when "00100110100000100", -- t[19716] = 1
      "0000001" when "00100110100000101", -- t[19717] = 1
      "0000001" when "00100110100000110", -- t[19718] = 1
      "0000001" when "00100110100000111", -- t[19719] = 1
      "0000001" when "00100110100001000", -- t[19720] = 1
      "0000001" when "00100110100001001", -- t[19721] = 1
      "0000001" when "00100110100001010", -- t[19722] = 1
      "0000001" when "00100110100001011", -- t[19723] = 1
      "0000001" when "00100110100001100", -- t[19724] = 1
      "0000001" when "00100110100001101", -- t[19725] = 1
      "0000001" when "00100110100001110", -- t[19726] = 1
      "0000001" when "00100110100001111", -- t[19727] = 1
      "0000001" when "00100110100010000", -- t[19728] = 1
      "0000001" when "00100110100010001", -- t[19729] = 1
      "0000001" when "00100110100010010", -- t[19730] = 1
      "0000001" when "00100110100010011", -- t[19731] = 1
      "0000001" when "00100110100010100", -- t[19732] = 1
      "0000001" when "00100110100010101", -- t[19733] = 1
      "0000001" when "00100110100010110", -- t[19734] = 1
      "0000001" when "00100110100010111", -- t[19735] = 1
      "0000001" when "00100110100011000", -- t[19736] = 1
      "0000001" when "00100110100011001", -- t[19737] = 1
      "0000001" when "00100110100011010", -- t[19738] = 1
      "0000001" when "00100110100011011", -- t[19739] = 1
      "0000001" when "00100110100011100", -- t[19740] = 1
      "0000001" when "00100110100011101", -- t[19741] = 1
      "0000001" when "00100110100011110", -- t[19742] = 1
      "0000001" when "00100110100011111", -- t[19743] = 1
      "0000001" when "00100110100100000", -- t[19744] = 1
      "0000001" when "00100110100100001", -- t[19745] = 1
      "0000001" when "00100110100100010", -- t[19746] = 1
      "0000001" when "00100110100100011", -- t[19747] = 1
      "0000001" when "00100110100100100", -- t[19748] = 1
      "0000001" when "00100110100100101", -- t[19749] = 1
      "0000001" when "00100110100100110", -- t[19750] = 1
      "0000001" when "00100110100100111", -- t[19751] = 1
      "0000001" when "00100110100101000", -- t[19752] = 1
      "0000001" when "00100110100101001", -- t[19753] = 1
      "0000001" when "00100110100101010", -- t[19754] = 1
      "0000001" when "00100110100101011", -- t[19755] = 1
      "0000001" when "00100110100101100", -- t[19756] = 1
      "0000001" when "00100110100101101", -- t[19757] = 1
      "0000001" when "00100110100101110", -- t[19758] = 1
      "0000001" when "00100110100101111", -- t[19759] = 1
      "0000001" when "00100110100110000", -- t[19760] = 1
      "0000001" when "00100110100110001", -- t[19761] = 1
      "0000001" when "00100110100110010", -- t[19762] = 1
      "0000001" when "00100110100110011", -- t[19763] = 1
      "0000001" when "00100110100110100", -- t[19764] = 1
      "0000001" when "00100110100110101", -- t[19765] = 1
      "0000001" when "00100110100110110", -- t[19766] = 1
      "0000001" when "00100110100110111", -- t[19767] = 1
      "0000001" when "00100110100111000", -- t[19768] = 1
      "0000001" when "00100110100111001", -- t[19769] = 1
      "0000001" when "00100110100111010", -- t[19770] = 1
      "0000001" when "00100110100111011", -- t[19771] = 1
      "0000001" when "00100110100111100", -- t[19772] = 1
      "0000001" when "00100110100111101", -- t[19773] = 1
      "0000001" when "00100110100111110", -- t[19774] = 1
      "0000001" when "00100110100111111", -- t[19775] = 1
      "0000001" when "00100110101000000", -- t[19776] = 1
      "0000001" when "00100110101000001", -- t[19777] = 1
      "0000001" when "00100110101000010", -- t[19778] = 1
      "0000001" when "00100110101000011", -- t[19779] = 1
      "0000001" when "00100110101000100", -- t[19780] = 1
      "0000001" when "00100110101000101", -- t[19781] = 1
      "0000001" when "00100110101000110", -- t[19782] = 1
      "0000001" when "00100110101000111", -- t[19783] = 1
      "0000001" when "00100110101001000", -- t[19784] = 1
      "0000001" when "00100110101001001", -- t[19785] = 1
      "0000001" when "00100110101001010", -- t[19786] = 1
      "0000001" when "00100110101001011", -- t[19787] = 1
      "0000001" when "00100110101001100", -- t[19788] = 1
      "0000001" when "00100110101001101", -- t[19789] = 1
      "0000001" when "00100110101001110", -- t[19790] = 1
      "0000001" when "00100110101001111", -- t[19791] = 1
      "0000001" when "00100110101010000", -- t[19792] = 1
      "0000001" when "00100110101010001", -- t[19793] = 1
      "0000001" when "00100110101010010", -- t[19794] = 1
      "0000001" when "00100110101010011", -- t[19795] = 1
      "0000001" when "00100110101010100", -- t[19796] = 1
      "0000001" when "00100110101010101", -- t[19797] = 1
      "0000001" when "00100110101010110", -- t[19798] = 1
      "0000001" when "00100110101010111", -- t[19799] = 1
      "0000001" when "00100110101011000", -- t[19800] = 1
      "0000001" when "00100110101011001", -- t[19801] = 1
      "0000001" when "00100110101011010", -- t[19802] = 1
      "0000001" when "00100110101011011", -- t[19803] = 1
      "0000001" when "00100110101011100", -- t[19804] = 1
      "0000001" when "00100110101011101", -- t[19805] = 1
      "0000001" when "00100110101011110", -- t[19806] = 1
      "0000001" when "00100110101011111", -- t[19807] = 1
      "0000001" when "00100110101100000", -- t[19808] = 1
      "0000001" when "00100110101100001", -- t[19809] = 1
      "0000001" when "00100110101100010", -- t[19810] = 1
      "0000001" when "00100110101100011", -- t[19811] = 1
      "0000001" when "00100110101100100", -- t[19812] = 1
      "0000001" when "00100110101100101", -- t[19813] = 1
      "0000001" when "00100110101100110", -- t[19814] = 1
      "0000001" when "00100110101100111", -- t[19815] = 1
      "0000001" when "00100110101101000", -- t[19816] = 1
      "0000001" when "00100110101101001", -- t[19817] = 1
      "0000001" when "00100110101101010", -- t[19818] = 1
      "0000001" when "00100110101101011", -- t[19819] = 1
      "0000001" when "00100110101101100", -- t[19820] = 1
      "0000001" when "00100110101101101", -- t[19821] = 1
      "0000001" when "00100110101101110", -- t[19822] = 1
      "0000001" when "00100110101101111", -- t[19823] = 1
      "0000001" when "00100110101110000", -- t[19824] = 1
      "0000001" when "00100110101110001", -- t[19825] = 1
      "0000001" when "00100110101110010", -- t[19826] = 1
      "0000001" when "00100110101110011", -- t[19827] = 1
      "0000001" when "00100110101110100", -- t[19828] = 1
      "0000001" when "00100110101110101", -- t[19829] = 1
      "0000001" when "00100110101110110", -- t[19830] = 1
      "0000001" when "00100110101110111", -- t[19831] = 1
      "0000001" when "00100110101111000", -- t[19832] = 1
      "0000001" when "00100110101111001", -- t[19833] = 1
      "0000001" when "00100110101111010", -- t[19834] = 1
      "0000001" when "00100110101111011", -- t[19835] = 1
      "0000001" when "00100110101111100", -- t[19836] = 1
      "0000001" when "00100110101111101", -- t[19837] = 1
      "0000001" when "00100110101111110", -- t[19838] = 1
      "0000001" when "00100110101111111", -- t[19839] = 1
      "0000001" when "00100110110000000", -- t[19840] = 1
      "0000001" when "00100110110000001", -- t[19841] = 1
      "0000001" when "00100110110000010", -- t[19842] = 1
      "0000001" when "00100110110000011", -- t[19843] = 1
      "0000001" when "00100110110000100", -- t[19844] = 1
      "0000001" when "00100110110000101", -- t[19845] = 1
      "0000001" when "00100110110000110", -- t[19846] = 1
      "0000001" when "00100110110000111", -- t[19847] = 1
      "0000001" when "00100110110001000", -- t[19848] = 1
      "0000001" when "00100110110001001", -- t[19849] = 1
      "0000001" when "00100110110001010", -- t[19850] = 1
      "0000001" when "00100110110001011", -- t[19851] = 1
      "0000001" when "00100110110001100", -- t[19852] = 1
      "0000001" when "00100110110001101", -- t[19853] = 1
      "0000001" when "00100110110001110", -- t[19854] = 1
      "0000001" when "00100110110001111", -- t[19855] = 1
      "0000001" when "00100110110010000", -- t[19856] = 1
      "0000001" when "00100110110010001", -- t[19857] = 1
      "0000001" when "00100110110010010", -- t[19858] = 1
      "0000001" when "00100110110010011", -- t[19859] = 1
      "0000001" when "00100110110010100", -- t[19860] = 1
      "0000001" when "00100110110010101", -- t[19861] = 1
      "0000001" when "00100110110010110", -- t[19862] = 1
      "0000001" when "00100110110010111", -- t[19863] = 1
      "0000001" when "00100110110011000", -- t[19864] = 1
      "0000001" when "00100110110011001", -- t[19865] = 1
      "0000001" when "00100110110011010", -- t[19866] = 1
      "0000001" when "00100110110011011", -- t[19867] = 1
      "0000001" when "00100110110011100", -- t[19868] = 1
      "0000001" when "00100110110011101", -- t[19869] = 1
      "0000001" when "00100110110011110", -- t[19870] = 1
      "0000001" when "00100110110011111", -- t[19871] = 1
      "0000001" when "00100110110100000", -- t[19872] = 1
      "0000001" when "00100110110100001", -- t[19873] = 1
      "0000001" when "00100110110100010", -- t[19874] = 1
      "0000001" when "00100110110100011", -- t[19875] = 1
      "0000001" when "00100110110100100", -- t[19876] = 1
      "0000001" when "00100110110100101", -- t[19877] = 1
      "0000001" when "00100110110100110", -- t[19878] = 1
      "0000001" when "00100110110100111", -- t[19879] = 1
      "0000001" when "00100110110101000", -- t[19880] = 1
      "0000001" when "00100110110101001", -- t[19881] = 1
      "0000001" when "00100110110101010", -- t[19882] = 1
      "0000001" when "00100110110101011", -- t[19883] = 1
      "0000001" when "00100110110101100", -- t[19884] = 1
      "0000001" when "00100110110101101", -- t[19885] = 1
      "0000001" when "00100110110101110", -- t[19886] = 1
      "0000001" when "00100110110101111", -- t[19887] = 1
      "0000001" when "00100110110110000", -- t[19888] = 1
      "0000001" when "00100110110110001", -- t[19889] = 1
      "0000001" when "00100110110110010", -- t[19890] = 1
      "0000001" when "00100110110110011", -- t[19891] = 1
      "0000001" when "00100110110110100", -- t[19892] = 1
      "0000001" when "00100110110110101", -- t[19893] = 1
      "0000001" when "00100110110110110", -- t[19894] = 1
      "0000001" when "00100110110110111", -- t[19895] = 1
      "0000001" when "00100110110111000", -- t[19896] = 1
      "0000001" when "00100110110111001", -- t[19897] = 1
      "0000001" when "00100110110111010", -- t[19898] = 1
      "0000001" when "00100110110111011", -- t[19899] = 1
      "0000001" when "00100110110111100", -- t[19900] = 1
      "0000001" when "00100110110111101", -- t[19901] = 1
      "0000001" when "00100110110111110", -- t[19902] = 1
      "0000001" when "00100110110111111", -- t[19903] = 1
      "0000001" when "00100110111000000", -- t[19904] = 1
      "0000001" when "00100110111000001", -- t[19905] = 1
      "0000001" when "00100110111000010", -- t[19906] = 1
      "0000001" when "00100110111000011", -- t[19907] = 1
      "0000001" when "00100110111000100", -- t[19908] = 1
      "0000001" when "00100110111000101", -- t[19909] = 1
      "0000001" when "00100110111000110", -- t[19910] = 1
      "0000001" when "00100110111000111", -- t[19911] = 1
      "0000001" when "00100110111001000", -- t[19912] = 1
      "0000001" when "00100110111001001", -- t[19913] = 1
      "0000001" when "00100110111001010", -- t[19914] = 1
      "0000001" when "00100110111001011", -- t[19915] = 1
      "0000001" when "00100110111001100", -- t[19916] = 1
      "0000001" when "00100110111001101", -- t[19917] = 1
      "0000001" when "00100110111001110", -- t[19918] = 1
      "0000001" when "00100110111001111", -- t[19919] = 1
      "0000001" when "00100110111010000", -- t[19920] = 1
      "0000001" when "00100110111010001", -- t[19921] = 1
      "0000001" when "00100110111010010", -- t[19922] = 1
      "0000001" when "00100110111010011", -- t[19923] = 1
      "0000001" when "00100110111010100", -- t[19924] = 1
      "0000001" when "00100110111010101", -- t[19925] = 1
      "0000001" when "00100110111010110", -- t[19926] = 1
      "0000001" when "00100110111010111", -- t[19927] = 1
      "0000001" when "00100110111011000", -- t[19928] = 1
      "0000001" when "00100110111011001", -- t[19929] = 1
      "0000001" when "00100110111011010", -- t[19930] = 1
      "0000001" when "00100110111011011", -- t[19931] = 1
      "0000001" when "00100110111011100", -- t[19932] = 1
      "0000001" when "00100110111011101", -- t[19933] = 1
      "0000001" when "00100110111011110", -- t[19934] = 1
      "0000001" when "00100110111011111", -- t[19935] = 1
      "0000001" when "00100110111100000", -- t[19936] = 1
      "0000001" when "00100110111100001", -- t[19937] = 1
      "0000001" when "00100110111100010", -- t[19938] = 1
      "0000001" when "00100110111100011", -- t[19939] = 1
      "0000001" when "00100110111100100", -- t[19940] = 1
      "0000001" when "00100110111100101", -- t[19941] = 1
      "0000001" when "00100110111100110", -- t[19942] = 1
      "0000001" when "00100110111100111", -- t[19943] = 1
      "0000001" when "00100110111101000", -- t[19944] = 1
      "0000001" when "00100110111101001", -- t[19945] = 1
      "0000001" when "00100110111101010", -- t[19946] = 1
      "0000001" when "00100110111101011", -- t[19947] = 1
      "0000001" when "00100110111101100", -- t[19948] = 1
      "0000001" when "00100110111101101", -- t[19949] = 1
      "0000001" when "00100110111101110", -- t[19950] = 1
      "0000001" when "00100110111101111", -- t[19951] = 1
      "0000001" when "00100110111110000", -- t[19952] = 1
      "0000001" when "00100110111110001", -- t[19953] = 1
      "0000001" when "00100110111110010", -- t[19954] = 1
      "0000001" when "00100110111110011", -- t[19955] = 1
      "0000001" when "00100110111110100", -- t[19956] = 1
      "0000001" when "00100110111110101", -- t[19957] = 1
      "0000001" when "00100110111110110", -- t[19958] = 1
      "0000001" when "00100110111110111", -- t[19959] = 1
      "0000001" when "00100110111111000", -- t[19960] = 1
      "0000001" when "00100110111111001", -- t[19961] = 1
      "0000001" when "00100110111111010", -- t[19962] = 1
      "0000001" when "00100110111111011", -- t[19963] = 1
      "0000001" when "00100110111111100", -- t[19964] = 1
      "0000001" when "00100110111111101", -- t[19965] = 1
      "0000001" when "00100110111111110", -- t[19966] = 1
      "0000001" when "00100110111111111", -- t[19967] = 1
      "0000001" when "00100111000000000", -- t[19968] = 1
      "0000001" when "00100111000000001", -- t[19969] = 1
      "0000001" when "00100111000000010", -- t[19970] = 1
      "0000001" when "00100111000000011", -- t[19971] = 1
      "0000001" when "00100111000000100", -- t[19972] = 1
      "0000001" when "00100111000000101", -- t[19973] = 1
      "0000001" when "00100111000000110", -- t[19974] = 1
      "0000001" when "00100111000000111", -- t[19975] = 1
      "0000001" when "00100111000001000", -- t[19976] = 1
      "0000001" when "00100111000001001", -- t[19977] = 1
      "0000001" when "00100111000001010", -- t[19978] = 1
      "0000001" when "00100111000001011", -- t[19979] = 1
      "0000001" when "00100111000001100", -- t[19980] = 1
      "0000001" when "00100111000001101", -- t[19981] = 1
      "0000001" when "00100111000001110", -- t[19982] = 1
      "0000001" when "00100111000001111", -- t[19983] = 1
      "0000001" when "00100111000010000", -- t[19984] = 1
      "0000001" when "00100111000010001", -- t[19985] = 1
      "0000001" when "00100111000010010", -- t[19986] = 1
      "0000001" when "00100111000010011", -- t[19987] = 1
      "0000001" when "00100111000010100", -- t[19988] = 1
      "0000001" when "00100111000010101", -- t[19989] = 1
      "0000001" when "00100111000010110", -- t[19990] = 1
      "0000001" when "00100111000010111", -- t[19991] = 1
      "0000001" when "00100111000011000", -- t[19992] = 1
      "0000001" when "00100111000011001", -- t[19993] = 1
      "0000001" when "00100111000011010", -- t[19994] = 1
      "0000001" when "00100111000011011", -- t[19995] = 1
      "0000001" when "00100111000011100", -- t[19996] = 1
      "0000001" when "00100111000011101", -- t[19997] = 1
      "0000001" when "00100111000011110", -- t[19998] = 1
      "0000001" when "00100111000011111", -- t[19999] = 1
      "0000001" when "00100111000100000", -- t[20000] = 1
      "0000001" when "00100111000100001", -- t[20001] = 1
      "0000001" when "00100111000100010", -- t[20002] = 1
      "0000001" when "00100111000100011", -- t[20003] = 1
      "0000001" when "00100111000100100", -- t[20004] = 1
      "0000001" when "00100111000100101", -- t[20005] = 1
      "0000001" when "00100111000100110", -- t[20006] = 1
      "0000001" when "00100111000100111", -- t[20007] = 1
      "0000001" when "00100111000101000", -- t[20008] = 1
      "0000001" when "00100111000101001", -- t[20009] = 1
      "0000001" when "00100111000101010", -- t[20010] = 1
      "0000001" when "00100111000101011", -- t[20011] = 1
      "0000001" when "00100111000101100", -- t[20012] = 1
      "0000001" when "00100111000101101", -- t[20013] = 1
      "0000001" when "00100111000101110", -- t[20014] = 1
      "0000001" when "00100111000101111", -- t[20015] = 1
      "0000001" when "00100111000110000", -- t[20016] = 1
      "0000001" when "00100111000110001", -- t[20017] = 1
      "0000001" when "00100111000110010", -- t[20018] = 1
      "0000001" when "00100111000110011", -- t[20019] = 1
      "0000001" when "00100111000110100", -- t[20020] = 1
      "0000001" when "00100111000110101", -- t[20021] = 1
      "0000001" when "00100111000110110", -- t[20022] = 1
      "0000001" when "00100111000110111", -- t[20023] = 1
      "0000001" when "00100111000111000", -- t[20024] = 1
      "0000001" when "00100111000111001", -- t[20025] = 1
      "0000001" when "00100111000111010", -- t[20026] = 1
      "0000001" when "00100111000111011", -- t[20027] = 1
      "0000001" when "00100111000111100", -- t[20028] = 1
      "0000001" when "00100111000111101", -- t[20029] = 1
      "0000001" when "00100111000111110", -- t[20030] = 1
      "0000001" when "00100111000111111", -- t[20031] = 1
      "0000001" when "00100111001000000", -- t[20032] = 1
      "0000001" when "00100111001000001", -- t[20033] = 1
      "0000001" when "00100111001000010", -- t[20034] = 1
      "0000001" when "00100111001000011", -- t[20035] = 1
      "0000001" when "00100111001000100", -- t[20036] = 1
      "0000001" when "00100111001000101", -- t[20037] = 1
      "0000001" when "00100111001000110", -- t[20038] = 1
      "0000001" when "00100111001000111", -- t[20039] = 1
      "0000001" when "00100111001001000", -- t[20040] = 1
      "0000001" when "00100111001001001", -- t[20041] = 1
      "0000001" when "00100111001001010", -- t[20042] = 1
      "0000001" when "00100111001001011", -- t[20043] = 1
      "0000001" when "00100111001001100", -- t[20044] = 1
      "0000001" when "00100111001001101", -- t[20045] = 1
      "0000001" when "00100111001001110", -- t[20046] = 1
      "0000001" when "00100111001001111", -- t[20047] = 1
      "0000001" when "00100111001010000", -- t[20048] = 1
      "0000001" when "00100111001010001", -- t[20049] = 1
      "0000001" when "00100111001010010", -- t[20050] = 1
      "0000001" when "00100111001010011", -- t[20051] = 1
      "0000001" when "00100111001010100", -- t[20052] = 1
      "0000001" when "00100111001010101", -- t[20053] = 1
      "0000001" when "00100111001010110", -- t[20054] = 1
      "0000001" when "00100111001010111", -- t[20055] = 1
      "0000001" when "00100111001011000", -- t[20056] = 1
      "0000001" when "00100111001011001", -- t[20057] = 1
      "0000001" when "00100111001011010", -- t[20058] = 1
      "0000001" when "00100111001011011", -- t[20059] = 1
      "0000001" when "00100111001011100", -- t[20060] = 1
      "0000001" when "00100111001011101", -- t[20061] = 1
      "0000001" when "00100111001011110", -- t[20062] = 1
      "0000001" when "00100111001011111", -- t[20063] = 1
      "0000001" when "00100111001100000", -- t[20064] = 1
      "0000001" when "00100111001100001", -- t[20065] = 1
      "0000001" when "00100111001100010", -- t[20066] = 1
      "0000001" when "00100111001100011", -- t[20067] = 1
      "0000001" when "00100111001100100", -- t[20068] = 1
      "0000001" when "00100111001100101", -- t[20069] = 1
      "0000001" when "00100111001100110", -- t[20070] = 1
      "0000001" when "00100111001100111", -- t[20071] = 1
      "0000001" when "00100111001101000", -- t[20072] = 1
      "0000001" when "00100111001101001", -- t[20073] = 1
      "0000001" when "00100111001101010", -- t[20074] = 1
      "0000001" when "00100111001101011", -- t[20075] = 1
      "0000001" when "00100111001101100", -- t[20076] = 1
      "0000001" when "00100111001101101", -- t[20077] = 1
      "0000001" when "00100111001101110", -- t[20078] = 1
      "0000001" when "00100111001101111", -- t[20079] = 1
      "0000001" when "00100111001110000", -- t[20080] = 1
      "0000001" when "00100111001110001", -- t[20081] = 1
      "0000001" when "00100111001110010", -- t[20082] = 1
      "0000001" when "00100111001110011", -- t[20083] = 1
      "0000001" when "00100111001110100", -- t[20084] = 1
      "0000001" when "00100111001110101", -- t[20085] = 1
      "0000001" when "00100111001110110", -- t[20086] = 1
      "0000001" when "00100111001110111", -- t[20087] = 1
      "0000001" when "00100111001111000", -- t[20088] = 1
      "0000001" when "00100111001111001", -- t[20089] = 1
      "0000001" when "00100111001111010", -- t[20090] = 1
      "0000001" when "00100111001111011", -- t[20091] = 1
      "0000001" when "00100111001111100", -- t[20092] = 1
      "0000001" when "00100111001111101", -- t[20093] = 1
      "0000001" when "00100111001111110", -- t[20094] = 1
      "0000001" when "00100111001111111", -- t[20095] = 1
      "0000001" when "00100111010000000", -- t[20096] = 1
      "0000001" when "00100111010000001", -- t[20097] = 1
      "0000001" when "00100111010000010", -- t[20098] = 1
      "0000001" when "00100111010000011", -- t[20099] = 1
      "0000001" when "00100111010000100", -- t[20100] = 1
      "0000001" when "00100111010000101", -- t[20101] = 1
      "0000001" when "00100111010000110", -- t[20102] = 1
      "0000001" when "00100111010000111", -- t[20103] = 1
      "0000001" when "00100111010001000", -- t[20104] = 1
      "0000001" when "00100111010001001", -- t[20105] = 1
      "0000001" when "00100111010001010", -- t[20106] = 1
      "0000001" when "00100111010001011", -- t[20107] = 1
      "0000001" when "00100111010001100", -- t[20108] = 1
      "0000001" when "00100111010001101", -- t[20109] = 1
      "0000001" when "00100111010001110", -- t[20110] = 1
      "0000001" when "00100111010001111", -- t[20111] = 1
      "0000001" when "00100111010010000", -- t[20112] = 1
      "0000001" when "00100111010010001", -- t[20113] = 1
      "0000001" when "00100111010010010", -- t[20114] = 1
      "0000001" when "00100111010010011", -- t[20115] = 1
      "0000001" when "00100111010010100", -- t[20116] = 1
      "0000001" when "00100111010010101", -- t[20117] = 1
      "0000001" when "00100111010010110", -- t[20118] = 1
      "0000001" when "00100111010010111", -- t[20119] = 1
      "0000001" when "00100111010011000", -- t[20120] = 1
      "0000001" when "00100111010011001", -- t[20121] = 1
      "0000001" when "00100111010011010", -- t[20122] = 1
      "0000001" when "00100111010011011", -- t[20123] = 1
      "0000001" when "00100111010011100", -- t[20124] = 1
      "0000001" when "00100111010011101", -- t[20125] = 1
      "0000001" when "00100111010011110", -- t[20126] = 1
      "0000001" when "00100111010011111", -- t[20127] = 1
      "0000001" when "00100111010100000", -- t[20128] = 1
      "0000001" when "00100111010100001", -- t[20129] = 1
      "0000001" when "00100111010100010", -- t[20130] = 1
      "0000001" when "00100111010100011", -- t[20131] = 1
      "0000001" when "00100111010100100", -- t[20132] = 1
      "0000001" when "00100111010100101", -- t[20133] = 1
      "0000001" when "00100111010100110", -- t[20134] = 1
      "0000001" when "00100111010100111", -- t[20135] = 1
      "0000001" when "00100111010101000", -- t[20136] = 1
      "0000001" when "00100111010101001", -- t[20137] = 1
      "0000001" when "00100111010101010", -- t[20138] = 1
      "0000001" when "00100111010101011", -- t[20139] = 1
      "0000001" when "00100111010101100", -- t[20140] = 1
      "0000001" when "00100111010101101", -- t[20141] = 1
      "0000001" when "00100111010101110", -- t[20142] = 1
      "0000001" when "00100111010101111", -- t[20143] = 1
      "0000001" when "00100111010110000", -- t[20144] = 1
      "0000001" when "00100111010110001", -- t[20145] = 1
      "0000001" when "00100111010110010", -- t[20146] = 1
      "0000001" when "00100111010110011", -- t[20147] = 1
      "0000001" when "00100111010110100", -- t[20148] = 1
      "0000001" when "00100111010110101", -- t[20149] = 1
      "0000001" when "00100111010110110", -- t[20150] = 1
      "0000001" when "00100111010110111", -- t[20151] = 1
      "0000001" when "00100111010111000", -- t[20152] = 1
      "0000001" when "00100111010111001", -- t[20153] = 1
      "0000001" when "00100111010111010", -- t[20154] = 1
      "0000001" when "00100111010111011", -- t[20155] = 1
      "0000001" when "00100111010111100", -- t[20156] = 1
      "0000001" when "00100111010111101", -- t[20157] = 1
      "0000001" when "00100111010111110", -- t[20158] = 1
      "0000001" when "00100111010111111", -- t[20159] = 1
      "0000001" when "00100111011000000", -- t[20160] = 1
      "0000001" when "00100111011000001", -- t[20161] = 1
      "0000001" when "00100111011000010", -- t[20162] = 1
      "0000001" when "00100111011000011", -- t[20163] = 1
      "0000001" when "00100111011000100", -- t[20164] = 1
      "0000001" when "00100111011000101", -- t[20165] = 1
      "0000001" when "00100111011000110", -- t[20166] = 1
      "0000001" when "00100111011000111", -- t[20167] = 1
      "0000001" when "00100111011001000", -- t[20168] = 1
      "0000001" when "00100111011001001", -- t[20169] = 1
      "0000001" when "00100111011001010", -- t[20170] = 1
      "0000001" when "00100111011001011", -- t[20171] = 1
      "0000001" when "00100111011001100", -- t[20172] = 1
      "0000001" when "00100111011001101", -- t[20173] = 1
      "0000001" when "00100111011001110", -- t[20174] = 1
      "0000001" when "00100111011001111", -- t[20175] = 1
      "0000001" when "00100111011010000", -- t[20176] = 1
      "0000001" when "00100111011010001", -- t[20177] = 1
      "0000001" when "00100111011010010", -- t[20178] = 1
      "0000001" when "00100111011010011", -- t[20179] = 1
      "0000001" when "00100111011010100", -- t[20180] = 1
      "0000001" when "00100111011010101", -- t[20181] = 1
      "0000001" when "00100111011010110", -- t[20182] = 1
      "0000001" when "00100111011010111", -- t[20183] = 1
      "0000001" when "00100111011011000", -- t[20184] = 1
      "0000001" when "00100111011011001", -- t[20185] = 1
      "0000001" when "00100111011011010", -- t[20186] = 1
      "0000001" when "00100111011011011", -- t[20187] = 1
      "0000001" when "00100111011011100", -- t[20188] = 1
      "0000001" when "00100111011011101", -- t[20189] = 1
      "0000001" when "00100111011011110", -- t[20190] = 1
      "0000001" when "00100111011011111", -- t[20191] = 1
      "0000001" when "00100111011100000", -- t[20192] = 1
      "0000001" when "00100111011100001", -- t[20193] = 1
      "0000001" when "00100111011100010", -- t[20194] = 1
      "0000001" when "00100111011100011", -- t[20195] = 1
      "0000001" when "00100111011100100", -- t[20196] = 1
      "0000001" when "00100111011100101", -- t[20197] = 1
      "0000001" when "00100111011100110", -- t[20198] = 1
      "0000001" when "00100111011100111", -- t[20199] = 1
      "0000001" when "00100111011101000", -- t[20200] = 1
      "0000001" when "00100111011101001", -- t[20201] = 1
      "0000001" when "00100111011101010", -- t[20202] = 1
      "0000001" when "00100111011101011", -- t[20203] = 1
      "0000001" when "00100111011101100", -- t[20204] = 1
      "0000001" when "00100111011101101", -- t[20205] = 1
      "0000001" when "00100111011101110", -- t[20206] = 1
      "0000001" when "00100111011101111", -- t[20207] = 1
      "0000001" when "00100111011110000", -- t[20208] = 1
      "0000001" when "00100111011110001", -- t[20209] = 1
      "0000001" when "00100111011110010", -- t[20210] = 1
      "0000001" when "00100111011110011", -- t[20211] = 1
      "0000001" when "00100111011110100", -- t[20212] = 1
      "0000001" when "00100111011110101", -- t[20213] = 1
      "0000001" when "00100111011110110", -- t[20214] = 1
      "0000001" when "00100111011110111", -- t[20215] = 1
      "0000001" when "00100111011111000", -- t[20216] = 1
      "0000001" when "00100111011111001", -- t[20217] = 1
      "0000001" when "00100111011111010", -- t[20218] = 1
      "0000001" when "00100111011111011", -- t[20219] = 1
      "0000001" when "00100111011111100", -- t[20220] = 1
      "0000001" when "00100111011111101", -- t[20221] = 1
      "0000001" when "00100111011111110", -- t[20222] = 1
      "0000001" when "00100111011111111", -- t[20223] = 1
      "0000001" when "00100111100000000", -- t[20224] = 1
      "0000001" when "00100111100000001", -- t[20225] = 1
      "0000001" when "00100111100000010", -- t[20226] = 1
      "0000001" when "00100111100000011", -- t[20227] = 1
      "0000001" when "00100111100000100", -- t[20228] = 1
      "0000001" when "00100111100000101", -- t[20229] = 1
      "0000001" when "00100111100000110", -- t[20230] = 1
      "0000001" when "00100111100000111", -- t[20231] = 1
      "0000001" when "00100111100001000", -- t[20232] = 1
      "0000001" when "00100111100001001", -- t[20233] = 1
      "0000001" when "00100111100001010", -- t[20234] = 1
      "0000001" when "00100111100001011", -- t[20235] = 1
      "0000001" when "00100111100001100", -- t[20236] = 1
      "0000001" when "00100111100001101", -- t[20237] = 1
      "0000001" when "00100111100001110", -- t[20238] = 1
      "0000001" when "00100111100001111", -- t[20239] = 1
      "0000001" when "00100111100010000", -- t[20240] = 1
      "0000001" when "00100111100010001", -- t[20241] = 1
      "0000001" when "00100111100010010", -- t[20242] = 1
      "0000001" when "00100111100010011", -- t[20243] = 1
      "0000001" when "00100111100010100", -- t[20244] = 1
      "0000001" when "00100111100010101", -- t[20245] = 1
      "0000001" when "00100111100010110", -- t[20246] = 1
      "0000001" when "00100111100010111", -- t[20247] = 1
      "0000001" when "00100111100011000", -- t[20248] = 1
      "0000001" when "00100111100011001", -- t[20249] = 1
      "0000001" when "00100111100011010", -- t[20250] = 1
      "0000001" when "00100111100011011", -- t[20251] = 1
      "0000001" when "00100111100011100", -- t[20252] = 1
      "0000001" when "00100111100011101", -- t[20253] = 1
      "0000001" when "00100111100011110", -- t[20254] = 1
      "0000001" when "00100111100011111", -- t[20255] = 1
      "0000001" when "00100111100100000", -- t[20256] = 1
      "0000001" when "00100111100100001", -- t[20257] = 1
      "0000001" when "00100111100100010", -- t[20258] = 1
      "0000001" when "00100111100100011", -- t[20259] = 1
      "0000001" when "00100111100100100", -- t[20260] = 1
      "0000001" when "00100111100100101", -- t[20261] = 1
      "0000001" when "00100111100100110", -- t[20262] = 1
      "0000001" when "00100111100100111", -- t[20263] = 1
      "0000001" when "00100111100101000", -- t[20264] = 1
      "0000001" when "00100111100101001", -- t[20265] = 1
      "0000001" when "00100111100101010", -- t[20266] = 1
      "0000001" when "00100111100101011", -- t[20267] = 1
      "0000001" when "00100111100101100", -- t[20268] = 1
      "0000001" when "00100111100101101", -- t[20269] = 1
      "0000001" when "00100111100101110", -- t[20270] = 1
      "0000001" when "00100111100101111", -- t[20271] = 1
      "0000001" when "00100111100110000", -- t[20272] = 1
      "0000001" when "00100111100110001", -- t[20273] = 1
      "0000001" when "00100111100110010", -- t[20274] = 1
      "0000001" when "00100111100110011", -- t[20275] = 1
      "0000001" when "00100111100110100", -- t[20276] = 1
      "0000001" when "00100111100110101", -- t[20277] = 1
      "0000001" when "00100111100110110", -- t[20278] = 1
      "0000001" when "00100111100110111", -- t[20279] = 1
      "0000001" when "00100111100111000", -- t[20280] = 1
      "0000001" when "00100111100111001", -- t[20281] = 1
      "0000001" when "00100111100111010", -- t[20282] = 1
      "0000001" when "00100111100111011", -- t[20283] = 1
      "0000001" when "00100111100111100", -- t[20284] = 1
      "0000001" when "00100111100111101", -- t[20285] = 1
      "0000001" when "00100111100111110", -- t[20286] = 1
      "0000001" when "00100111100111111", -- t[20287] = 1
      "0000001" when "00100111101000000", -- t[20288] = 1
      "0000001" when "00100111101000001", -- t[20289] = 1
      "0000001" when "00100111101000010", -- t[20290] = 1
      "0000001" when "00100111101000011", -- t[20291] = 1
      "0000001" when "00100111101000100", -- t[20292] = 1
      "0000001" when "00100111101000101", -- t[20293] = 1
      "0000001" when "00100111101000110", -- t[20294] = 1
      "0000001" when "00100111101000111", -- t[20295] = 1
      "0000001" when "00100111101001000", -- t[20296] = 1
      "0000001" when "00100111101001001", -- t[20297] = 1
      "0000001" when "00100111101001010", -- t[20298] = 1
      "0000001" when "00100111101001011", -- t[20299] = 1
      "0000001" when "00100111101001100", -- t[20300] = 1
      "0000001" when "00100111101001101", -- t[20301] = 1
      "0000001" when "00100111101001110", -- t[20302] = 1
      "0000001" when "00100111101001111", -- t[20303] = 1
      "0000001" when "00100111101010000", -- t[20304] = 1
      "0000001" when "00100111101010001", -- t[20305] = 1
      "0000001" when "00100111101010010", -- t[20306] = 1
      "0000001" when "00100111101010011", -- t[20307] = 1
      "0000001" when "00100111101010100", -- t[20308] = 1
      "0000001" when "00100111101010101", -- t[20309] = 1
      "0000001" when "00100111101010110", -- t[20310] = 1
      "0000001" when "00100111101010111", -- t[20311] = 1
      "0000001" when "00100111101011000", -- t[20312] = 1
      "0000001" when "00100111101011001", -- t[20313] = 1
      "0000001" when "00100111101011010", -- t[20314] = 1
      "0000001" when "00100111101011011", -- t[20315] = 1
      "0000001" when "00100111101011100", -- t[20316] = 1
      "0000001" when "00100111101011101", -- t[20317] = 1
      "0000001" when "00100111101011110", -- t[20318] = 1
      "0000001" when "00100111101011111", -- t[20319] = 1
      "0000001" when "00100111101100000", -- t[20320] = 1
      "0000001" when "00100111101100001", -- t[20321] = 1
      "0000001" when "00100111101100010", -- t[20322] = 1
      "0000001" when "00100111101100011", -- t[20323] = 1
      "0000001" when "00100111101100100", -- t[20324] = 1
      "0000001" when "00100111101100101", -- t[20325] = 1
      "0000001" when "00100111101100110", -- t[20326] = 1
      "0000001" when "00100111101100111", -- t[20327] = 1
      "0000001" when "00100111101101000", -- t[20328] = 1
      "0000001" when "00100111101101001", -- t[20329] = 1
      "0000001" when "00100111101101010", -- t[20330] = 1
      "0000001" when "00100111101101011", -- t[20331] = 1
      "0000001" when "00100111101101100", -- t[20332] = 1
      "0000001" when "00100111101101101", -- t[20333] = 1
      "0000001" when "00100111101101110", -- t[20334] = 1
      "0000001" when "00100111101101111", -- t[20335] = 1
      "0000001" when "00100111101110000", -- t[20336] = 1
      "0000001" when "00100111101110001", -- t[20337] = 1
      "0000001" when "00100111101110010", -- t[20338] = 1
      "0000001" when "00100111101110011", -- t[20339] = 1
      "0000001" when "00100111101110100", -- t[20340] = 1
      "0000001" when "00100111101110101", -- t[20341] = 1
      "0000001" when "00100111101110110", -- t[20342] = 1
      "0000001" when "00100111101110111", -- t[20343] = 1
      "0000001" when "00100111101111000", -- t[20344] = 1
      "0000001" when "00100111101111001", -- t[20345] = 1
      "0000001" when "00100111101111010", -- t[20346] = 1
      "0000001" when "00100111101111011", -- t[20347] = 1
      "0000001" when "00100111101111100", -- t[20348] = 1
      "0000001" when "00100111101111101", -- t[20349] = 1
      "0000001" when "00100111101111110", -- t[20350] = 1
      "0000001" when "00100111101111111", -- t[20351] = 1
      "0000001" when "00100111110000000", -- t[20352] = 1
      "0000001" when "00100111110000001", -- t[20353] = 1
      "0000001" when "00100111110000010", -- t[20354] = 1
      "0000001" when "00100111110000011", -- t[20355] = 1
      "0000001" when "00100111110000100", -- t[20356] = 1
      "0000001" when "00100111110000101", -- t[20357] = 1
      "0000001" when "00100111110000110", -- t[20358] = 1
      "0000001" when "00100111110000111", -- t[20359] = 1
      "0000001" when "00100111110001000", -- t[20360] = 1
      "0000001" when "00100111110001001", -- t[20361] = 1
      "0000001" when "00100111110001010", -- t[20362] = 1
      "0000001" when "00100111110001011", -- t[20363] = 1
      "0000001" when "00100111110001100", -- t[20364] = 1
      "0000001" when "00100111110001101", -- t[20365] = 1
      "0000001" when "00100111110001110", -- t[20366] = 1
      "0000001" when "00100111110001111", -- t[20367] = 1
      "0000001" when "00100111110010000", -- t[20368] = 1
      "0000001" when "00100111110010001", -- t[20369] = 1
      "0000001" when "00100111110010010", -- t[20370] = 1
      "0000001" when "00100111110010011", -- t[20371] = 1
      "0000001" when "00100111110010100", -- t[20372] = 1
      "0000001" when "00100111110010101", -- t[20373] = 1
      "0000001" when "00100111110010110", -- t[20374] = 1
      "0000001" when "00100111110010111", -- t[20375] = 1
      "0000001" when "00100111110011000", -- t[20376] = 1
      "0000001" when "00100111110011001", -- t[20377] = 1
      "0000001" when "00100111110011010", -- t[20378] = 1
      "0000001" when "00100111110011011", -- t[20379] = 1
      "0000001" when "00100111110011100", -- t[20380] = 1
      "0000001" when "00100111110011101", -- t[20381] = 1
      "0000001" when "00100111110011110", -- t[20382] = 1
      "0000001" when "00100111110011111", -- t[20383] = 1
      "0000001" when "00100111110100000", -- t[20384] = 1
      "0000001" when "00100111110100001", -- t[20385] = 1
      "0000001" when "00100111110100010", -- t[20386] = 1
      "0000001" when "00100111110100011", -- t[20387] = 1
      "0000001" when "00100111110100100", -- t[20388] = 1
      "0000001" when "00100111110100101", -- t[20389] = 1
      "0000001" when "00100111110100110", -- t[20390] = 1
      "0000001" when "00100111110100111", -- t[20391] = 1
      "0000001" when "00100111110101000", -- t[20392] = 1
      "0000001" when "00100111110101001", -- t[20393] = 1
      "0000001" when "00100111110101010", -- t[20394] = 1
      "0000001" when "00100111110101011", -- t[20395] = 1
      "0000001" when "00100111110101100", -- t[20396] = 1
      "0000001" when "00100111110101101", -- t[20397] = 1
      "0000001" when "00100111110101110", -- t[20398] = 1
      "0000001" when "00100111110101111", -- t[20399] = 1
      "0000001" when "00100111110110000", -- t[20400] = 1
      "0000001" when "00100111110110001", -- t[20401] = 1
      "0000001" when "00100111110110010", -- t[20402] = 1
      "0000001" when "00100111110110011", -- t[20403] = 1
      "0000001" when "00100111110110100", -- t[20404] = 1
      "0000001" when "00100111110110101", -- t[20405] = 1
      "0000001" when "00100111110110110", -- t[20406] = 1
      "0000001" when "00100111110110111", -- t[20407] = 1
      "0000001" when "00100111110111000", -- t[20408] = 1
      "0000001" when "00100111110111001", -- t[20409] = 1
      "0000001" when "00100111110111010", -- t[20410] = 1
      "0000001" when "00100111110111011", -- t[20411] = 1
      "0000001" when "00100111110111100", -- t[20412] = 1
      "0000001" when "00100111110111101", -- t[20413] = 1
      "0000001" when "00100111110111110", -- t[20414] = 1
      "0000001" when "00100111110111111", -- t[20415] = 1
      "0000001" when "00100111111000000", -- t[20416] = 1
      "0000001" when "00100111111000001", -- t[20417] = 1
      "0000001" when "00100111111000010", -- t[20418] = 1
      "0000001" when "00100111111000011", -- t[20419] = 1
      "0000001" when "00100111111000100", -- t[20420] = 1
      "0000001" when "00100111111000101", -- t[20421] = 1
      "0000001" when "00100111111000110", -- t[20422] = 1
      "0000001" when "00100111111000111", -- t[20423] = 1
      "0000001" when "00100111111001000", -- t[20424] = 1
      "0000001" when "00100111111001001", -- t[20425] = 1
      "0000001" when "00100111111001010", -- t[20426] = 1
      "0000001" when "00100111111001011", -- t[20427] = 1
      "0000001" when "00100111111001100", -- t[20428] = 1
      "0000001" when "00100111111001101", -- t[20429] = 1
      "0000001" when "00100111111001110", -- t[20430] = 1
      "0000001" when "00100111111001111", -- t[20431] = 1
      "0000001" when "00100111111010000", -- t[20432] = 1
      "0000001" when "00100111111010001", -- t[20433] = 1
      "0000001" when "00100111111010010", -- t[20434] = 1
      "0000001" when "00100111111010011", -- t[20435] = 1
      "0000001" when "00100111111010100", -- t[20436] = 1
      "0000001" when "00100111111010101", -- t[20437] = 1
      "0000001" when "00100111111010110", -- t[20438] = 1
      "0000001" when "00100111111010111", -- t[20439] = 1
      "0000001" when "00100111111011000", -- t[20440] = 1
      "0000001" when "00100111111011001", -- t[20441] = 1
      "0000001" when "00100111111011010", -- t[20442] = 1
      "0000001" when "00100111111011011", -- t[20443] = 1
      "0000001" when "00100111111011100", -- t[20444] = 1
      "0000001" when "00100111111011101", -- t[20445] = 1
      "0000001" when "00100111111011110", -- t[20446] = 1
      "0000001" when "00100111111011111", -- t[20447] = 1
      "0000001" when "00100111111100000", -- t[20448] = 1
      "0000001" when "00100111111100001", -- t[20449] = 1
      "0000001" when "00100111111100010", -- t[20450] = 1
      "0000001" when "00100111111100011", -- t[20451] = 1
      "0000001" when "00100111111100100", -- t[20452] = 1
      "0000001" when "00100111111100101", -- t[20453] = 1
      "0000001" when "00100111111100110", -- t[20454] = 1
      "0000001" when "00100111111100111", -- t[20455] = 1
      "0000001" when "00100111111101000", -- t[20456] = 1
      "0000001" when "00100111111101001", -- t[20457] = 1
      "0000001" when "00100111111101010", -- t[20458] = 1
      "0000001" when "00100111111101011", -- t[20459] = 1
      "0000001" when "00100111111101100", -- t[20460] = 1
      "0000001" when "00100111111101101", -- t[20461] = 1
      "0000001" when "00100111111101110", -- t[20462] = 1
      "0000001" when "00100111111101111", -- t[20463] = 1
      "0000001" when "00100111111110000", -- t[20464] = 1
      "0000001" when "00100111111110001", -- t[20465] = 1
      "0000001" when "00100111111110010", -- t[20466] = 1
      "0000001" when "00100111111110011", -- t[20467] = 1
      "0000001" when "00100111111110100", -- t[20468] = 1
      "0000001" when "00100111111110101", -- t[20469] = 1
      "0000001" when "00100111111110110", -- t[20470] = 1
      "0000001" when "00100111111110111", -- t[20471] = 1
      "0000001" when "00100111111111000", -- t[20472] = 1
      "0000001" when "00100111111111001", -- t[20473] = 1
      "0000001" when "00100111111111010", -- t[20474] = 1
      "0000001" when "00100111111111011", -- t[20475] = 1
      "0000001" when "00100111111111100", -- t[20476] = 1
      "0000001" when "00100111111111101", -- t[20477] = 1
      "0000001" when "00100111111111110", -- t[20478] = 1
      "0000001" when "00100111111111111", -- t[20479] = 1
      "0000001" when "00101000000000000", -- t[20480] = 1
      "0000001" when "00101000000000001", -- t[20481] = 1
      "0000001" when "00101000000000010", -- t[20482] = 1
      "0000001" when "00101000000000011", -- t[20483] = 1
      "0000001" when "00101000000000100", -- t[20484] = 1
      "0000001" when "00101000000000101", -- t[20485] = 1
      "0000001" when "00101000000000110", -- t[20486] = 1
      "0000001" when "00101000000000111", -- t[20487] = 1
      "0000001" when "00101000000001000", -- t[20488] = 1
      "0000001" when "00101000000001001", -- t[20489] = 1
      "0000001" when "00101000000001010", -- t[20490] = 1
      "0000001" when "00101000000001011", -- t[20491] = 1
      "0000001" when "00101000000001100", -- t[20492] = 1
      "0000001" when "00101000000001101", -- t[20493] = 1
      "0000001" when "00101000000001110", -- t[20494] = 1
      "0000001" when "00101000000001111", -- t[20495] = 1
      "0000001" when "00101000000010000", -- t[20496] = 1
      "0000001" when "00101000000010001", -- t[20497] = 1
      "0000001" when "00101000000010010", -- t[20498] = 1
      "0000001" when "00101000000010011", -- t[20499] = 1
      "0000001" when "00101000000010100", -- t[20500] = 1
      "0000001" when "00101000000010101", -- t[20501] = 1
      "0000001" when "00101000000010110", -- t[20502] = 1
      "0000001" when "00101000000010111", -- t[20503] = 1
      "0000001" when "00101000000011000", -- t[20504] = 1
      "0000001" when "00101000000011001", -- t[20505] = 1
      "0000001" when "00101000000011010", -- t[20506] = 1
      "0000001" when "00101000000011011", -- t[20507] = 1
      "0000001" when "00101000000011100", -- t[20508] = 1
      "0000001" when "00101000000011101", -- t[20509] = 1
      "0000001" when "00101000000011110", -- t[20510] = 1
      "0000001" when "00101000000011111", -- t[20511] = 1
      "0000001" when "00101000000100000", -- t[20512] = 1
      "0000001" when "00101000000100001", -- t[20513] = 1
      "0000001" when "00101000000100010", -- t[20514] = 1
      "0000001" when "00101000000100011", -- t[20515] = 1
      "0000001" when "00101000000100100", -- t[20516] = 1
      "0000001" when "00101000000100101", -- t[20517] = 1
      "0000001" when "00101000000100110", -- t[20518] = 1
      "0000001" when "00101000000100111", -- t[20519] = 1
      "0000001" when "00101000000101000", -- t[20520] = 1
      "0000001" when "00101000000101001", -- t[20521] = 1
      "0000001" when "00101000000101010", -- t[20522] = 1
      "0000001" when "00101000000101011", -- t[20523] = 1
      "0000001" when "00101000000101100", -- t[20524] = 1
      "0000001" when "00101000000101101", -- t[20525] = 1
      "0000001" when "00101000000101110", -- t[20526] = 1
      "0000001" when "00101000000101111", -- t[20527] = 1
      "0000001" when "00101000000110000", -- t[20528] = 1
      "0000001" when "00101000000110001", -- t[20529] = 1
      "0000001" when "00101000000110010", -- t[20530] = 1
      "0000001" when "00101000000110011", -- t[20531] = 1
      "0000001" when "00101000000110100", -- t[20532] = 1
      "0000001" when "00101000000110101", -- t[20533] = 1
      "0000001" when "00101000000110110", -- t[20534] = 1
      "0000001" when "00101000000110111", -- t[20535] = 1
      "0000001" when "00101000000111000", -- t[20536] = 1
      "0000001" when "00101000000111001", -- t[20537] = 1
      "0000001" when "00101000000111010", -- t[20538] = 1
      "0000001" when "00101000000111011", -- t[20539] = 1
      "0000001" when "00101000000111100", -- t[20540] = 1
      "0000001" when "00101000000111101", -- t[20541] = 1
      "0000001" when "00101000000111110", -- t[20542] = 1
      "0000001" when "00101000000111111", -- t[20543] = 1
      "0000001" when "00101000001000000", -- t[20544] = 1
      "0000001" when "00101000001000001", -- t[20545] = 1
      "0000001" when "00101000001000010", -- t[20546] = 1
      "0000001" when "00101000001000011", -- t[20547] = 1
      "0000001" when "00101000001000100", -- t[20548] = 1
      "0000001" when "00101000001000101", -- t[20549] = 1
      "0000001" when "00101000001000110", -- t[20550] = 1
      "0000001" when "00101000001000111", -- t[20551] = 1
      "0000001" when "00101000001001000", -- t[20552] = 1
      "0000001" when "00101000001001001", -- t[20553] = 1
      "0000001" when "00101000001001010", -- t[20554] = 1
      "0000001" when "00101000001001011", -- t[20555] = 1
      "0000001" when "00101000001001100", -- t[20556] = 1
      "0000001" when "00101000001001101", -- t[20557] = 1
      "0000001" when "00101000001001110", -- t[20558] = 1
      "0000001" when "00101000001001111", -- t[20559] = 1
      "0000001" when "00101000001010000", -- t[20560] = 1
      "0000001" when "00101000001010001", -- t[20561] = 1
      "0000001" when "00101000001010010", -- t[20562] = 1
      "0000001" when "00101000001010011", -- t[20563] = 1
      "0000001" when "00101000001010100", -- t[20564] = 1
      "0000001" when "00101000001010101", -- t[20565] = 1
      "0000001" when "00101000001010110", -- t[20566] = 1
      "0000001" when "00101000001010111", -- t[20567] = 1
      "0000001" when "00101000001011000", -- t[20568] = 1
      "0000001" when "00101000001011001", -- t[20569] = 1
      "0000001" when "00101000001011010", -- t[20570] = 1
      "0000001" when "00101000001011011", -- t[20571] = 1
      "0000001" when "00101000001011100", -- t[20572] = 1
      "0000001" when "00101000001011101", -- t[20573] = 1
      "0000001" when "00101000001011110", -- t[20574] = 1
      "0000001" when "00101000001011111", -- t[20575] = 1
      "0000001" when "00101000001100000", -- t[20576] = 1
      "0000001" when "00101000001100001", -- t[20577] = 1
      "0000001" when "00101000001100010", -- t[20578] = 1
      "0000001" when "00101000001100011", -- t[20579] = 1
      "0000001" when "00101000001100100", -- t[20580] = 1
      "0000001" when "00101000001100101", -- t[20581] = 1
      "0000001" when "00101000001100110", -- t[20582] = 1
      "0000001" when "00101000001100111", -- t[20583] = 1
      "0000001" when "00101000001101000", -- t[20584] = 1
      "0000001" when "00101000001101001", -- t[20585] = 1
      "0000001" when "00101000001101010", -- t[20586] = 1
      "0000001" when "00101000001101011", -- t[20587] = 1
      "0000001" when "00101000001101100", -- t[20588] = 1
      "0000001" when "00101000001101101", -- t[20589] = 1
      "0000001" when "00101000001101110", -- t[20590] = 1
      "0000001" when "00101000001101111", -- t[20591] = 1
      "0000001" when "00101000001110000", -- t[20592] = 1
      "0000001" when "00101000001110001", -- t[20593] = 1
      "0000001" when "00101000001110010", -- t[20594] = 1
      "0000001" when "00101000001110011", -- t[20595] = 1
      "0000001" when "00101000001110100", -- t[20596] = 1
      "0000001" when "00101000001110101", -- t[20597] = 1
      "0000001" when "00101000001110110", -- t[20598] = 1
      "0000001" when "00101000001110111", -- t[20599] = 1
      "0000001" when "00101000001111000", -- t[20600] = 1
      "0000001" when "00101000001111001", -- t[20601] = 1
      "0000001" when "00101000001111010", -- t[20602] = 1
      "0000001" when "00101000001111011", -- t[20603] = 1
      "0000001" when "00101000001111100", -- t[20604] = 1
      "0000001" when "00101000001111101", -- t[20605] = 1
      "0000001" when "00101000001111110", -- t[20606] = 1
      "0000001" when "00101000001111111", -- t[20607] = 1
      "0000001" when "00101000010000000", -- t[20608] = 1
      "0000001" when "00101000010000001", -- t[20609] = 1
      "0000001" when "00101000010000010", -- t[20610] = 1
      "0000001" when "00101000010000011", -- t[20611] = 1
      "0000001" when "00101000010000100", -- t[20612] = 1
      "0000001" when "00101000010000101", -- t[20613] = 1
      "0000001" when "00101000010000110", -- t[20614] = 1
      "0000001" when "00101000010000111", -- t[20615] = 1
      "0000001" when "00101000010001000", -- t[20616] = 1
      "0000001" when "00101000010001001", -- t[20617] = 1
      "0000001" when "00101000010001010", -- t[20618] = 1
      "0000001" when "00101000010001011", -- t[20619] = 1
      "0000001" when "00101000010001100", -- t[20620] = 1
      "0000001" when "00101000010001101", -- t[20621] = 1
      "0000001" when "00101000010001110", -- t[20622] = 1
      "0000001" when "00101000010001111", -- t[20623] = 1
      "0000001" when "00101000010010000", -- t[20624] = 1
      "0000001" when "00101000010010001", -- t[20625] = 1
      "0000001" when "00101000010010010", -- t[20626] = 1
      "0000001" when "00101000010010011", -- t[20627] = 1
      "0000001" when "00101000010010100", -- t[20628] = 1
      "0000001" when "00101000010010101", -- t[20629] = 1
      "0000001" when "00101000010010110", -- t[20630] = 1
      "0000001" when "00101000010010111", -- t[20631] = 1
      "0000001" when "00101000010011000", -- t[20632] = 1
      "0000001" when "00101000010011001", -- t[20633] = 1
      "0000001" when "00101000010011010", -- t[20634] = 1
      "0000001" when "00101000010011011", -- t[20635] = 1
      "0000001" when "00101000010011100", -- t[20636] = 1
      "0000001" when "00101000010011101", -- t[20637] = 1
      "0000001" when "00101000010011110", -- t[20638] = 1
      "0000001" when "00101000010011111", -- t[20639] = 1
      "0000001" when "00101000010100000", -- t[20640] = 1
      "0000001" when "00101000010100001", -- t[20641] = 1
      "0000001" when "00101000010100010", -- t[20642] = 1
      "0000001" when "00101000010100011", -- t[20643] = 1
      "0000001" when "00101000010100100", -- t[20644] = 1
      "0000001" when "00101000010100101", -- t[20645] = 1
      "0000001" when "00101000010100110", -- t[20646] = 1
      "0000001" when "00101000010100111", -- t[20647] = 1
      "0000001" when "00101000010101000", -- t[20648] = 1
      "0000001" when "00101000010101001", -- t[20649] = 1
      "0000001" when "00101000010101010", -- t[20650] = 1
      "0000001" when "00101000010101011", -- t[20651] = 1
      "0000001" when "00101000010101100", -- t[20652] = 1
      "0000001" when "00101000010101101", -- t[20653] = 1
      "0000001" when "00101000010101110", -- t[20654] = 1
      "0000001" when "00101000010101111", -- t[20655] = 1
      "0000001" when "00101000010110000", -- t[20656] = 1
      "0000001" when "00101000010110001", -- t[20657] = 1
      "0000001" when "00101000010110010", -- t[20658] = 1
      "0000001" when "00101000010110011", -- t[20659] = 1
      "0000001" when "00101000010110100", -- t[20660] = 1
      "0000001" when "00101000010110101", -- t[20661] = 1
      "0000001" when "00101000010110110", -- t[20662] = 1
      "0000001" when "00101000010110111", -- t[20663] = 1
      "0000001" when "00101000010111000", -- t[20664] = 1
      "0000001" when "00101000010111001", -- t[20665] = 1
      "0000001" when "00101000010111010", -- t[20666] = 1
      "0000001" when "00101000010111011", -- t[20667] = 1
      "0000001" when "00101000010111100", -- t[20668] = 1
      "0000001" when "00101000010111101", -- t[20669] = 1
      "0000001" when "00101000010111110", -- t[20670] = 1
      "0000001" when "00101000010111111", -- t[20671] = 1
      "0000001" when "00101000011000000", -- t[20672] = 1
      "0000001" when "00101000011000001", -- t[20673] = 1
      "0000001" when "00101000011000010", -- t[20674] = 1
      "0000001" when "00101000011000011", -- t[20675] = 1
      "0000001" when "00101000011000100", -- t[20676] = 1
      "0000001" when "00101000011000101", -- t[20677] = 1
      "0000001" when "00101000011000110", -- t[20678] = 1
      "0000001" when "00101000011000111", -- t[20679] = 1
      "0000001" when "00101000011001000", -- t[20680] = 1
      "0000001" when "00101000011001001", -- t[20681] = 1
      "0000001" when "00101000011001010", -- t[20682] = 1
      "0000001" when "00101000011001011", -- t[20683] = 1
      "0000001" when "00101000011001100", -- t[20684] = 1
      "0000001" when "00101000011001101", -- t[20685] = 1
      "0000001" when "00101000011001110", -- t[20686] = 1
      "0000001" when "00101000011001111", -- t[20687] = 1
      "0000001" when "00101000011010000", -- t[20688] = 1
      "0000001" when "00101000011010001", -- t[20689] = 1
      "0000001" when "00101000011010010", -- t[20690] = 1
      "0000001" when "00101000011010011", -- t[20691] = 1
      "0000001" when "00101000011010100", -- t[20692] = 1
      "0000001" when "00101000011010101", -- t[20693] = 1
      "0000001" when "00101000011010110", -- t[20694] = 1
      "0000001" when "00101000011010111", -- t[20695] = 1
      "0000001" when "00101000011011000", -- t[20696] = 1
      "0000001" when "00101000011011001", -- t[20697] = 1
      "0000001" when "00101000011011010", -- t[20698] = 1
      "0000001" when "00101000011011011", -- t[20699] = 1
      "0000001" when "00101000011011100", -- t[20700] = 1
      "0000001" when "00101000011011101", -- t[20701] = 1
      "0000001" when "00101000011011110", -- t[20702] = 1
      "0000001" when "00101000011011111", -- t[20703] = 1
      "0000001" when "00101000011100000", -- t[20704] = 1
      "0000001" when "00101000011100001", -- t[20705] = 1
      "0000001" when "00101000011100010", -- t[20706] = 1
      "0000001" when "00101000011100011", -- t[20707] = 1
      "0000001" when "00101000011100100", -- t[20708] = 1
      "0000001" when "00101000011100101", -- t[20709] = 1
      "0000001" when "00101000011100110", -- t[20710] = 1
      "0000001" when "00101000011100111", -- t[20711] = 1
      "0000001" when "00101000011101000", -- t[20712] = 1
      "0000001" when "00101000011101001", -- t[20713] = 1
      "0000001" when "00101000011101010", -- t[20714] = 1
      "0000001" when "00101000011101011", -- t[20715] = 1
      "0000001" when "00101000011101100", -- t[20716] = 1
      "0000001" when "00101000011101101", -- t[20717] = 1
      "0000001" when "00101000011101110", -- t[20718] = 1
      "0000001" when "00101000011101111", -- t[20719] = 1
      "0000001" when "00101000011110000", -- t[20720] = 1
      "0000001" when "00101000011110001", -- t[20721] = 1
      "0000001" when "00101000011110010", -- t[20722] = 1
      "0000001" when "00101000011110011", -- t[20723] = 1
      "0000001" when "00101000011110100", -- t[20724] = 1
      "0000001" when "00101000011110101", -- t[20725] = 1
      "0000001" when "00101000011110110", -- t[20726] = 1
      "0000001" when "00101000011110111", -- t[20727] = 1
      "0000001" when "00101000011111000", -- t[20728] = 1
      "0000001" when "00101000011111001", -- t[20729] = 1
      "0000001" when "00101000011111010", -- t[20730] = 1
      "0000001" when "00101000011111011", -- t[20731] = 1
      "0000001" when "00101000011111100", -- t[20732] = 1
      "0000001" when "00101000011111101", -- t[20733] = 1
      "0000001" when "00101000011111110", -- t[20734] = 1
      "0000001" when "00101000011111111", -- t[20735] = 1
      "0000001" when "00101000100000000", -- t[20736] = 1
      "0000001" when "00101000100000001", -- t[20737] = 1
      "0000001" when "00101000100000010", -- t[20738] = 1
      "0000001" when "00101000100000011", -- t[20739] = 1
      "0000001" when "00101000100000100", -- t[20740] = 1
      "0000001" when "00101000100000101", -- t[20741] = 1
      "0000001" when "00101000100000110", -- t[20742] = 1
      "0000001" when "00101000100000111", -- t[20743] = 1
      "0000001" when "00101000100001000", -- t[20744] = 1
      "0000001" when "00101000100001001", -- t[20745] = 1
      "0000001" when "00101000100001010", -- t[20746] = 1
      "0000001" when "00101000100001011", -- t[20747] = 1
      "0000001" when "00101000100001100", -- t[20748] = 1
      "0000001" when "00101000100001101", -- t[20749] = 1
      "0000001" when "00101000100001110", -- t[20750] = 1
      "0000001" when "00101000100001111", -- t[20751] = 1
      "0000001" when "00101000100010000", -- t[20752] = 1
      "0000001" when "00101000100010001", -- t[20753] = 1
      "0000001" when "00101000100010010", -- t[20754] = 1
      "0000001" when "00101000100010011", -- t[20755] = 1
      "0000001" when "00101000100010100", -- t[20756] = 1
      "0000001" when "00101000100010101", -- t[20757] = 1
      "0000001" when "00101000100010110", -- t[20758] = 1
      "0000001" when "00101000100010111", -- t[20759] = 1
      "0000001" when "00101000100011000", -- t[20760] = 1
      "0000001" when "00101000100011001", -- t[20761] = 1
      "0000001" when "00101000100011010", -- t[20762] = 1
      "0000001" when "00101000100011011", -- t[20763] = 1
      "0000001" when "00101000100011100", -- t[20764] = 1
      "0000001" when "00101000100011101", -- t[20765] = 1
      "0000001" when "00101000100011110", -- t[20766] = 1
      "0000001" when "00101000100011111", -- t[20767] = 1
      "0000001" when "00101000100100000", -- t[20768] = 1
      "0000001" when "00101000100100001", -- t[20769] = 1
      "0000001" when "00101000100100010", -- t[20770] = 1
      "0000001" when "00101000100100011", -- t[20771] = 1
      "0000001" when "00101000100100100", -- t[20772] = 1
      "0000001" when "00101000100100101", -- t[20773] = 1
      "0000001" when "00101000100100110", -- t[20774] = 1
      "0000001" when "00101000100100111", -- t[20775] = 1
      "0000001" when "00101000100101000", -- t[20776] = 1
      "0000001" when "00101000100101001", -- t[20777] = 1
      "0000001" when "00101000100101010", -- t[20778] = 1
      "0000001" when "00101000100101011", -- t[20779] = 1
      "0000001" when "00101000100101100", -- t[20780] = 1
      "0000001" when "00101000100101101", -- t[20781] = 1
      "0000001" when "00101000100101110", -- t[20782] = 1
      "0000001" when "00101000100101111", -- t[20783] = 1
      "0000001" when "00101000100110000", -- t[20784] = 1
      "0000001" when "00101000100110001", -- t[20785] = 1
      "0000001" when "00101000100110010", -- t[20786] = 1
      "0000001" when "00101000100110011", -- t[20787] = 1
      "0000001" when "00101000100110100", -- t[20788] = 1
      "0000001" when "00101000100110101", -- t[20789] = 1
      "0000001" when "00101000100110110", -- t[20790] = 1
      "0000001" when "00101000100110111", -- t[20791] = 1
      "0000001" when "00101000100111000", -- t[20792] = 1
      "0000001" when "00101000100111001", -- t[20793] = 1
      "0000001" when "00101000100111010", -- t[20794] = 1
      "0000001" when "00101000100111011", -- t[20795] = 1
      "0000001" when "00101000100111100", -- t[20796] = 1
      "0000001" when "00101000100111101", -- t[20797] = 1
      "0000001" when "00101000100111110", -- t[20798] = 1
      "0000001" when "00101000100111111", -- t[20799] = 1
      "0000001" when "00101000101000000", -- t[20800] = 1
      "0000001" when "00101000101000001", -- t[20801] = 1
      "0000001" when "00101000101000010", -- t[20802] = 1
      "0000001" when "00101000101000011", -- t[20803] = 1
      "0000001" when "00101000101000100", -- t[20804] = 1
      "0000001" when "00101000101000101", -- t[20805] = 1
      "0000001" when "00101000101000110", -- t[20806] = 1
      "0000001" when "00101000101000111", -- t[20807] = 1
      "0000001" when "00101000101001000", -- t[20808] = 1
      "0000001" when "00101000101001001", -- t[20809] = 1
      "0000001" when "00101000101001010", -- t[20810] = 1
      "0000001" when "00101000101001011", -- t[20811] = 1
      "0000001" when "00101000101001100", -- t[20812] = 1
      "0000001" when "00101000101001101", -- t[20813] = 1
      "0000001" when "00101000101001110", -- t[20814] = 1
      "0000001" when "00101000101001111", -- t[20815] = 1
      "0000001" when "00101000101010000", -- t[20816] = 1
      "0000001" when "00101000101010001", -- t[20817] = 1
      "0000001" when "00101000101010010", -- t[20818] = 1
      "0000001" when "00101000101010011", -- t[20819] = 1
      "0000001" when "00101000101010100", -- t[20820] = 1
      "0000001" when "00101000101010101", -- t[20821] = 1
      "0000001" when "00101000101010110", -- t[20822] = 1
      "0000001" when "00101000101010111", -- t[20823] = 1
      "0000001" when "00101000101011000", -- t[20824] = 1
      "0000001" when "00101000101011001", -- t[20825] = 1
      "0000001" when "00101000101011010", -- t[20826] = 1
      "0000001" when "00101000101011011", -- t[20827] = 1
      "0000001" when "00101000101011100", -- t[20828] = 1
      "0000001" when "00101000101011101", -- t[20829] = 1
      "0000001" when "00101000101011110", -- t[20830] = 1
      "0000001" when "00101000101011111", -- t[20831] = 1
      "0000001" when "00101000101100000", -- t[20832] = 1
      "0000001" when "00101000101100001", -- t[20833] = 1
      "0000001" when "00101000101100010", -- t[20834] = 1
      "0000001" when "00101000101100011", -- t[20835] = 1
      "0000001" when "00101000101100100", -- t[20836] = 1
      "0000001" when "00101000101100101", -- t[20837] = 1
      "0000001" when "00101000101100110", -- t[20838] = 1
      "0000001" when "00101000101100111", -- t[20839] = 1
      "0000001" when "00101000101101000", -- t[20840] = 1
      "0000001" when "00101000101101001", -- t[20841] = 1
      "0000001" when "00101000101101010", -- t[20842] = 1
      "0000001" when "00101000101101011", -- t[20843] = 1
      "0000001" when "00101000101101100", -- t[20844] = 1
      "0000001" when "00101000101101101", -- t[20845] = 1
      "0000001" when "00101000101101110", -- t[20846] = 1
      "0000001" when "00101000101101111", -- t[20847] = 1
      "0000001" when "00101000101110000", -- t[20848] = 1
      "0000001" when "00101000101110001", -- t[20849] = 1
      "0000001" when "00101000101110010", -- t[20850] = 1
      "0000001" when "00101000101110011", -- t[20851] = 1
      "0000001" when "00101000101110100", -- t[20852] = 1
      "0000001" when "00101000101110101", -- t[20853] = 1
      "0000001" when "00101000101110110", -- t[20854] = 1
      "0000001" when "00101000101110111", -- t[20855] = 1
      "0000001" when "00101000101111000", -- t[20856] = 1
      "0000001" when "00101000101111001", -- t[20857] = 1
      "0000001" when "00101000101111010", -- t[20858] = 1
      "0000001" when "00101000101111011", -- t[20859] = 1
      "0000001" when "00101000101111100", -- t[20860] = 1
      "0000001" when "00101000101111101", -- t[20861] = 1
      "0000001" when "00101000101111110", -- t[20862] = 1
      "0000001" when "00101000101111111", -- t[20863] = 1
      "0000001" when "00101000110000000", -- t[20864] = 1
      "0000001" when "00101000110000001", -- t[20865] = 1
      "0000001" when "00101000110000010", -- t[20866] = 1
      "0000001" when "00101000110000011", -- t[20867] = 1
      "0000001" when "00101000110000100", -- t[20868] = 1
      "0000001" when "00101000110000101", -- t[20869] = 1
      "0000001" when "00101000110000110", -- t[20870] = 1
      "0000001" when "00101000110000111", -- t[20871] = 1
      "0000001" when "00101000110001000", -- t[20872] = 1
      "0000001" when "00101000110001001", -- t[20873] = 1
      "0000001" when "00101000110001010", -- t[20874] = 1
      "0000001" when "00101000110001011", -- t[20875] = 1
      "0000001" when "00101000110001100", -- t[20876] = 1
      "0000001" when "00101000110001101", -- t[20877] = 1
      "0000001" when "00101000110001110", -- t[20878] = 1
      "0000001" when "00101000110001111", -- t[20879] = 1
      "0000001" when "00101000110010000", -- t[20880] = 1
      "0000001" when "00101000110010001", -- t[20881] = 1
      "0000001" when "00101000110010010", -- t[20882] = 1
      "0000001" when "00101000110010011", -- t[20883] = 1
      "0000001" when "00101000110010100", -- t[20884] = 1
      "0000001" when "00101000110010101", -- t[20885] = 1
      "0000001" when "00101000110010110", -- t[20886] = 1
      "0000001" when "00101000110010111", -- t[20887] = 1
      "0000001" when "00101000110011000", -- t[20888] = 1
      "0000001" when "00101000110011001", -- t[20889] = 1
      "0000001" when "00101000110011010", -- t[20890] = 1
      "0000001" when "00101000110011011", -- t[20891] = 1
      "0000001" when "00101000110011100", -- t[20892] = 1
      "0000001" when "00101000110011101", -- t[20893] = 1
      "0000001" when "00101000110011110", -- t[20894] = 1
      "0000001" when "00101000110011111", -- t[20895] = 1
      "0000001" when "00101000110100000", -- t[20896] = 1
      "0000001" when "00101000110100001", -- t[20897] = 1
      "0000001" when "00101000110100010", -- t[20898] = 1
      "0000001" when "00101000110100011", -- t[20899] = 1
      "0000001" when "00101000110100100", -- t[20900] = 1
      "0000001" when "00101000110100101", -- t[20901] = 1
      "0000001" when "00101000110100110", -- t[20902] = 1
      "0000001" when "00101000110100111", -- t[20903] = 1
      "0000001" when "00101000110101000", -- t[20904] = 1
      "0000001" when "00101000110101001", -- t[20905] = 1
      "0000001" when "00101000110101010", -- t[20906] = 1
      "0000001" when "00101000110101011", -- t[20907] = 1
      "0000001" when "00101000110101100", -- t[20908] = 1
      "0000001" when "00101000110101101", -- t[20909] = 1
      "0000001" when "00101000110101110", -- t[20910] = 1
      "0000001" when "00101000110101111", -- t[20911] = 1
      "0000001" when "00101000110110000", -- t[20912] = 1
      "0000001" when "00101000110110001", -- t[20913] = 1
      "0000001" when "00101000110110010", -- t[20914] = 1
      "0000001" when "00101000110110011", -- t[20915] = 1
      "0000001" when "00101000110110100", -- t[20916] = 1
      "0000001" when "00101000110110101", -- t[20917] = 1
      "0000001" when "00101000110110110", -- t[20918] = 1
      "0000001" when "00101000110110111", -- t[20919] = 1
      "0000001" when "00101000110111000", -- t[20920] = 1
      "0000001" when "00101000110111001", -- t[20921] = 1
      "0000001" when "00101000110111010", -- t[20922] = 1
      "0000001" when "00101000110111011", -- t[20923] = 1
      "0000001" when "00101000110111100", -- t[20924] = 1
      "0000001" when "00101000110111101", -- t[20925] = 1
      "0000001" when "00101000110111110", -- t[20926] = 1
      "0000001" when "00101000110111111", -- t[20927] = 1
      "0000001" when "00101000111000000", -- t[20928] = 1
      "0000001" when "00101000111000001", -- t[20929] = 1
      "0000001" when "00101000111000010", -- t[20930] = 1
      "0000001" when "00101000111000011", -- t[20931] = 1
      "0000001" when "00101000111000100", -- t[20932] = 1
      "0000001" when "00101000111000101", -- t[20933] = 1
      "0000001" when "00101000111000110", -- t[20934] = 1
      "0000001" when "00101000111000111", -- t[20935] = 1
      "0000001" when "00101000111001000", -- t[20936] = 1
      "0000001" when "00101000111001001", -- t[20937] = 1
      "0000001" when "00101000111001010", -- t[20938] = 1
      "0000001" when "00101000111001011", -- t[20939] = 1
      "0000001" when "00101000111001100", -- t[20940] = 1
      "0000001" when "00101000111001101", -- t[20941] = 1
      "0000001" when "00101000111001110", -- t[20942] = 1
      "0000001" when "00101000111001111", -- t[20943] = 1
      "0000001" when "00101000111010000", -- t[20944] = 1
      "0000001" when "00101000111010001", -- t[20945] = 1
      "0000001" when "00101000111010010", -- t[20946] = 1
      "0000001" when "00101000111010011", -- t[20947] = 1
      "0000001" when "00101000111010100", -- t[20948] = 1
      "0000001" when "00101000111010101", -- t[20949] = 1
      "0000001" when "00101000111010110", -- t[20950] = 1
      "0000001" when "00101000111010111", -- t[20951] = 1
      "0000001" when "00101000111011000", -- t[20952] = 1
      "0000001" when "00101000111011001", -- t[20953] = 1
      "0000001" when "00101000111011010", -- t[20954] = 1
      "0000001" when "00101000111011011", -- t[20955] = 1
      "0000001" when "00101000111011100", -- t[20956] = 1
      "0000001" when "00101000111011101", -- t[20957] = 1
      "0000001" when "00101000111011110", -- t[20958] = 1
      "0000001" when "00101000111011111", -- t[20959] = 1
      "0000001" when "00101000111100000", -- t[20960] = 1
      "0000001" when "00101000111100001", -- t[20961] = 1
      "0000001" when "00101000111100010", -- t[20962] = 1
      "0000001" when "00101000111100011", -- t[20963] = 1
      "0000001" when "00101000111100100", -- t[20964] = 1
      "0000001" when "00101000111100101", -- t[20965] = 1
      "0000001" when "00101000111100110", -- t[20966] = 1
      "0000001" when "00101000111100111", -- t[20967] = 1
      "0000001" when "00101000111101000", -- t[20968] = 1
      "0000001" when "00101000111101001", -- t[20969] = 1
      "0000001" when "00101000111101010", -- t[20970] = 1
      "0000001" when "00101000111101011", -- t[20971] = 1
      "0000001" when "00101000111101100", -- t[20972] = 1
      "0000001" when "00101000111101101", -- t[20973] = 1
      "0000001" when "00101000111101110", -- t[20974] = 1
      "0000001" when "00101000111101111", -- t[20975] = 1
      "0000001" when "00101000111110000", -- t[20976] = 1
      "0000001" when "00101000111110001", -- t[20977] = 1
      "0000001" when "00101000111110010", -- t[20978] = 1
      "0000001" when "00101000111110011", -- t[20979] = 1
      "0000001" when "00101000111110100", -- t[20980] = 1
      "0000001" when "00101000111110101", -- t[20981] = 1
      "0000001" when "00101000111110110", -- t[20982] = 1
      "0000001" when "00101000111110111", -- t[20983] = 1
      "0000001" when "00101000111111000", -- t[20984] = 1
      "0000001" when "00101000111111001", -- t[20985] = 1
      "0000001" when "00101000111111010", -- t[20986] = 1
      "0000001" when "00101000111111011", -- t[20987] = 1
      "0000001" when "00101000111111100", -- t[20988] = 1
      "0000001" when "00101000111111101", -- t[20989] = 1
      "0000001" when "00101000111111110", -- t[20990] = 1
      "0000001" when "00101000111111111", -- t[20991] = 1
      "0000001" when "00101001000000000", -- t[20992] = 1
      "0000001" when "00101001000000001", -- t[20993] = 1
      "0000001" when "00101001000000010", -- t[20994] = 1
      "0000001" when "00101001000000011", -- t[20995] = 1
      "0000001" when "00101001000000100", -- t[20996] = 1
      "0000001" when "00101001000000101", -- t[20997] = 1
      "0000001" when "00101001000000110", -- t[20998] = 1
      "0000001" when "00101001000000111", -- t[20999] = 1
      "0000001" when "00101001000001000", -- t[21000] = 1
      "0000001" when "00101001000001001", -- t[21001] = 1
      "0000001" when "00101001000001010", -- t[21002] = 1
      "0000001" when "00101001000001011", -- t[21003] = 1
      "0000001" when "00101001000001100", -- t[21004] = 1
      "0000001" when "00101001000001101", -- t[21005] = 1
      "0000001" when "00101001000001110", -- t[21006] = 1
      "0000001" when "00101001000001111", -- t[21007] = 1
      "0000001" when "00101001000010000", -- t[21008] = 1
      "0000001" when "00101001000010001", -- t[21009] = 1
      "0000001" when "00101001000010010", -- t[21010] = 1
      "0000001" when "00101001000010011", -- t[21011] = 1
      "0000001" when "00101001000010100", -- t[21012] = 1
      "0000001" when "00101001000010101", -- t[21013] = 1
      "0000001" when "00101001000010110", -- t[21014] = 1
      "0000001" when "00101001000010111", -- t[21015] = 1
      "0000001" when "00101001000011000", -- t[21016] = 1
      "0000001" when "00101001000011001", -- t[21017] = 1
      "0000001" when "00101001000011010", -- t[21018] = 1
      "0000001" when "00101001000011011", -- t[21019] = 1
      "0000001" when "00101001000011100", -- t[21020] = 1
      "0000001" when "00101001000011101", -- t[21021] = 1
      "0000001" when "00101001000011110", -- t[21022] = 1
      "0000001" when "00101001000011111", -- t[21023] = 1
      "0000001" when "00101001000100000", -- t[21024] = 1
      "0000001" when "00101001000100001", -- t[21025] = 1
      "0000001" when "00101001000100010", -- t[21026] = 1
      "0000001" when "00101001000100011", -- t[21027] = 1
      "0000001" when "00101001000100100", -- t[21028] = 1
      "0000001" when "00101001000100101", -- t[21029] = 1
      "0000001" when "00101001000100110", -- t[21030] = 1
      "0000001" when "00101001000100111", -- t[21031] = 1
      "0000001" when "00101001000101000", -- t[21032] = 1
      "0000001" when "00101001000101001", -- t[21033] = 1
      "0000001" when "00101001000101010", -- t[21034] = 1
      "0000001" when "00101001000101011", -- t[21035] = 1
      "0000001" when "00101001000101100", -- t[21036] = 1
      "0000001" when "00101001000101101", -- t[21037] = 1
      "0000001" when "00101001000101110", -- t[21038] = 1
      "0000001" when "00101001000101111", -- t[21039] = 1
      "0000001" when "00101001000110000", -- t[21040] = 1
      "0000001" when "00101001000110001", -- t[21041] = 1
      "0000001" when "00101001000110010", -- t[21042] = 1
      "0000001" when "00101001000110011", -- t[21043] = 1
      "0000001" when "00101001000110100", -- t[21044] = 1
      "0000001" when "00101001000110101", -- t[21045] = 1
      "0000001" when "00101001000110110", -- t[21046] = 1
      "0000001" when "00101001000110111", -- t[21047] = 1
      "0000001" when "00101001000111000", -- t[21048] = 1
      "0000001" when "00101001000111001", -- t[21049] = 1
      "0000001" when "00101001000111010", -- t[21050] = 1
      "0000001" when "00101001000111011", -- t[21051] = 1
      "0000001" when "00101001000111100", -- t[21052] = 1
      "0000001" when "00101001000111101", -- t[21053] = 1
      "0000001" when "00101001000111110", -- t[21054] = 1
      "0000001" when "00101001000111111", -- t[21055] = 1
      "0000001" when "00101001001000000", -- t[21056] = 1
      "0000001" when "00101001001000001", -- t[21057] = 1
      "0000001" when "00101001001000010", -- t[21058] = 1
      "0000001" when "00101001001000011", -- t[21059] = 1
      "0000001" when "00101001001000100", -- t[21060] = 1
      "0000001" when "00101001001000101", -- t[21061] = 1
      "0000001" when "00101001001000110", -- t[21062] = 1
      "0000001" when "00101001001000111", -- t[21063] = 1
      "0000001" when "00101001001001000", -- t[21064] = 1
      "0000001" when "00101001001001001", -- t[21065] = 1
      "0000001" when "00101001001001010", -- t[21066] = 1
      "0000001" when "00101001001001011", -- t[21067] = 1
      "0000001" when "00101001001001100", -- t[21068] = 1
      "0000001" when "00101001001001101", -- t[21069] = 1
      "0000001" when "00101001001001110", -- t[21070] = 1
      "0000001" when "00101001001001111", -- t[21071] = 1
      "0000001" when "00101001001010000", -- t[21072] = 1
      "0000001" when "00101001001010001", -- t[21073] = 1
      "0000001" when "00101001001010010", -- t[21074] = 1
      "0000001" when "00101001001010011", -- t[21075] = 1
      "0000001" when "00101001001010100", -- t[21076] = 1
      "0000001" when "00101001001010101", -- t[21077] = 1
      "0000001" when "00101001001010110", -- t[21078] = 1
      "0000001" when "00101001001010111", -- t[21079] = 1
      "0000001" when "00101001001011000", -- t[21080] = 1
      "0000001" when "00101001001011001", -- t[21081] = 1
      "0000001" when "00101001001011010", -- t[21082] = 1
      "0000001" when "00101001001011011", -- t[21083] = 1
      "0000001" when "00101001001011100", -- t[21084] = 1
      "0000001" when "00101001001011101", -- t[21085] = 1
      "0000001" when "00101001001011110", -- t[21086] = 1
      "0000001" when "00101001001011111", -- t[21087] = 1
      "0000001" when "00101001001100000", -- t[21088] = 1
      "0000001" when "00101001001100001", -- t[21089] = 1
      "0000001" when "00101001001100010", -- t[21090] = 1
      "0000001" when "00101001001100011", -- t[21091] = 1
      "0000001" when "00101001001100100", -- t[21092] = 1
      "0000001" when "00101001001100101", -- t[21093] = 1
      "0000001" when "00101001001100110", -- t[21094] = 1
      "0000001" when "00101001001100111", -- t[21095] = 1
      "0000001" when "00101001001101000", -- t[21096] = 1
      "0000001" when "00101001001101001", -- t[21097] = 1
      "0000001" when "00101001001101010", -- t[21098] = 1
      "0000001" when "00101001001101011", -- t[21099] = 1
      "0000001" when "00101001001101100", -- t[21100] = 1
      "0000001" when "00101001001101101", -- t[21101] = 1
      "0000001" when "00101001001101110", -- t[21102] = 1
      "0000001" when "00101001001101111", -- t[21103] = 1
      "0000001" when "00101001001110000", -- t[21104] = 1
      "0000001" when "00101001001110001", -- t[21105] = 1
      "0000001" when "00101001001110010", -- t[21106] = 1
      "0000001" when "00101001001110011", -- t[21107] = 1
      "0000001" when "00101001001110100", -- t[21108] = 1
      "0000001" when "00101001001110101", -- t[21109] = 1
      "0000001" when "00101001001110110", -- t[21110] = 1
      "0000001" when "00101001001110111", -- t[21111] = 1
      "0000001" when "00101001001111000", -- t[21112] = 1
      "0000001" when "00101001001111001", -- t[21113] = 1
      "0000001" when "00101001001111010", -- t[21114] = 1
      "0000001" when "00101001001111011", -- t[21115] = 1
      "0000001" when "00101001001111100", -- t[21116] = 1
      "0000001" when "00101001001111101", -- t[21117] = 1
      "0000001" when "00101001001111110", -- t[21118] = 1
      "0000001" when "00101001001111111", -- t[21119] = 1
      "0000001" when "00101001010000000", -- t[21120] = 1
      "0000001" when "00101001010000001", -- t[21121] = 1
      "0000001" when "00101001010000010", -- t[21122] = 1
      "0000001" when "00101001010000011", -- t[21123] = 1
      "0000001" when "00101001010000100", -- t[21124] = 1
      "0000001" when "00101001010000101", -- t[21125] = 1
      "0000001" when "00101001010000110", -- t[21126] = 1
      "0000001" when "00101001010000111", -- t[21127] = 1
      "0000001" when "00101001010001000", -- t[21128] = 1
      "0000001" when "00101001010001001", -- t[21129] = 1
      "0000001" when "00101001010001010", -- t[21130] = 1
      "0000001" when "00101001010001011", -- t[21131] = 1
      "0000001" when "00101001010001100", -- t[21132] = 1
      "0000001" when "00101001010001101", -- t[21133] = 1
      "0000001" when "00101001010001110", -- t[21134] = 1
      "0000001" when "00101001010001111", -- t[21135] = 1
      "0000001" when "00101001010010000", -- t[21136] = 1
      "0000001" when "00101001010010001", -- t[21137] = 1
      "0000001" when "00101001010010010", -- t[21138] = 1
      "0000001" when "00101001010010011", -- t[21139] = 1
      "0000001" when "00101001010010100", -- t[21140] = 1
      "0000001" when "00101001010010101", -- t[21141] = 1
      "0000001" when "00101001010010110", -- t[21142] = 1
      "0000001" when "00101001010010111", -- t[21143] = 1
      "0000001" when "00101001010011000", -- t[21144] = 1
      "0000001" when "00101001010011001", -- t[21145] = 1
      "0000001" when "00101001010011010", -- t[21146] = 1
      "0000001" when "00101001010011011", -- t[21147] = 1
      "0000001" when "00101001010011100", -- t[21148] = 1
      "0000001" when "00101001010011101", -- t[21149] = 1
      "0000001" when "00101001010011110", -- t[21150] = 1
      "0000001" when "00101001010011111", -- t[21151] = 1
      "0000001" when "00101001010100000", -- t[21152] = 1
      "0000001" when "00101001010100001", -- t[21153] = 1
      "0000001" when "00101001010100010", -- t[21154] = 1
      "0000001" when "00101001010100011", -- t[21155] = 1
      "0000001" when "00101001010100100", -- t[21156] = 1
      "0000001" when "00101001010100101", -- t[21157] = 1
      "0000001" when "00101001010100110", -- t[21158] = 1
      "0000001" when "00101001010100111", -- t[21159] = 1
      "0000001" when "00101001010101000", -- t[21160] = 1
      "0000001" when "00101001010101001", -- t[21161] = 1
      "0000001" when "00101001010101010", -- t[21162] = 1
      "0000001" when "00101001010101011", -- t[21163] = 1
      "0000001" when "00101001010101100", -- t[21164] = 1
      "0000001" when "00101001010101101", -- t[21165] = 1
      "0000001" when "00101001010101110", -- t[21166] = 1
      "0000001" when "00101001010101111", -- t[21167] = 1
      "0000001" when "00101001010110000", -- t[21168] = 1
      "0000001" when "00101001010110001", -- t[21169] = 1
      "0000001" when "00101001010110010", -- t[21170] = 1
      "0000001" when "00101001010110011", -- t[21171] = 1
      "0000001" when "00101001010110100", -- t[21172] = 1
      "0000001" when "00101001010110101", -- t[21173] = 1
      "0000001" when "00101001010110110", -- t[21174] = 1
      "0000001" when "00101001010110111", -- t[21175] = 1
      "0000001" when "00101001010111000", -- t[21176] = 1
      "0000001" when "00101001010111001", -- t[21177] = 1
      "0000001" when "00101001010111010", -- t[21178] = 1
      "0000001" when "00101001010111011", -- t[21179] = 1
      "0000001" when "00101001010111100", -- t[21180] = 1
      "0000001" when "00101001010111101", -- t[21181] = 1
      "0000001" when "00101001010111110", -- t[21182] = 1
      "0000001" when "00101001010111111", -- t[21183] = 1
      "0000001" when "00101001011000000", -- t[21184] = 1
      "0000001" when "00101001011000001", -- t[21185] = 1
      "0000001" when "00101001011000010", -- t[21186] = 1
      "0000001" when "00101001011000011", -- t[21187] = 1
      "0000001" when "00101001011000100", -- t[21188] = 1
      "0000001" when "00101001011000101", -- t[21189] = 1
      "0000001" when "00101001011000110", -- t[21190] = 1
      "0000001" when "00101001011000111", -- t[21191] = 1
      "0000001" when "00101001011001000", -- t[21192] = 1
      "0000001" when "00101001011001001", -- t[21193] = 1
      "0000001" when "00101001011001010", -- t[21194] = 1
      "0000001" when "00101001011001011", -- t[21195] = 1
      "0000001" when "00101001011001100", -- t[21196] = 1
      "0000001" when "00101001011001101", -- t[21197] = 1
      "0000001" when "00101001011001110", -- t[21198] = 1
      "0000001" when "00101001011001111", -- t[21199] = 1
      "0000001" when "00101001011010000", -- t[21200] = 1
      "0000001" when "00101001011010001", -- t[21201] = 1
      "0000001" when "00101001011010010", -- t[21202] = 1
      "0000001" when "00101001011010011", -- t[21203] = 1
      "0000001" when "00101001011010100", -- t[21204] = 1
      "0000001" when "00101001011010101", -- t[21205] = 1
      "0000001" when "00101001011010110", -- t[21206] = 1
      "0000001" when "00101001011010111", -- t[21207] = 1
      "0000001" when "00101001011011000", -- t[21208] = 1
      "0000001" when "00101001011011001", -- t[21209] = 1
      "0000001" when "00101001011011010", -- t[21210] = 1
      "0000001" when "00101001011011011", -- t[21211] = 1
      "0000001" when "00101001011011100", -- t[21212] = 1
      "0000001" when "00101001011011101", -- t[21213] = 1
      "0000001" when "00101001011011110", -- t[21214] = 1
      "0000001" when "00101001011011111", -- t[21215] = 1
      "0000001" when "00101001011100000", -- t[21216] = 1
      "0000001" when "00101001011100001", -- t[21217] = 1
      "0000001" when "00101001011100010", -- t[21218] = 1
      "0000001" when "00101001011100011", -- t[21219] = 1
      "0000001" when "00101001011100100", -- t[21220] = 1
      "0000001" when "00101001011100101", -- t[21221] = 1
      "0000001" when "00101001011100110", -- t[21222] = 1
      "0000001" when "00101001011100111", -- t[21223] = 1
      "0000001" when "00101001011101000", -- t[21224] = 1
      "0000001" when "00101001011101001", -- t[21225] = 1
      "0000001" when "00101001011101010", -- t[21226] = 1
      "0000001" when "00101001011101011", -- t[21227] = 1
      "0000001" when "00101001011101100", -- t[21228] = 1
      "0000001" when "00101001011101101", -- t[21229] = 1
      "0000001" when "00101001011101110", -- t[21230] = 1
      "0000001" when "00101001011101111", -- t[21231] = 1
      "0000001" when "00101001011110000", -- t[21232] = 1
      "0000001" when "00101001011110001", -- t[21233] = 1
      "0000001" when "00101001011110010", -- t[21234] = 1
      "0000001" when "00101001011110011", -- t[21235] = 1
      "0000001" when "00101001011110100", -- t[21236] = 1
      "0000001" when "00101001011110101", -- t[21237] = 1
      "0000001" when "00101001011110110", -- t[21238] = 1
      "0000001" when "00101001011110111", -- t[21239] = 1
      "0000001" when "00101001011111000", -- t[21240] = 1
      "0000001" when "00101001011111001", -- t[21241] = 1
      "0000001" when "00101001011111010", -- t[21242] = 1
      "0000001" when "00101001011111011", -- t[21243] = 1
      "0000001" when "00101001011111100", -- t[21244] = 1
      "0000001" when "00101001011111101", -- t[21245] = 1
      "0000001" when "00101001011111110", -- t[21246] = 1
      "0000001" when "00101001011111111", -- t[21247] = 1
      "0000001" when "00101001100000000", -- t[21248] = 1
      "0000001" when "00101001100000001", -- t[21249] = 1
      "0000001" when "00101001100000010", -- t[21250] = 1
      "0000001" when "00101001100000011", -- t[21251] = 1
      "0000001" when "00101001100000100", -- t[21252] = 1
      "0000001" when "00101001100000101", -- t[21253] = 1
      "0000001" when "00101001100000110", -- t[21254] = 1
      "0000001" when "00101001100000111", -- t[21255] = 1
      "0000001" when "00101001100001000", -- t[21256] = 1
      "0000001" when "00101001100001001", -- t[21257] = 1
      "0000001" when "00101001100001010", -- t[21258] = 1
      "0000001" when "00101001100001011", -- t[21259] = 1
      "0000001" when "00101001100001100", -- t[21260] = 1
      "0000001" when "00101001100001101", -- t[21261] = 1
      "0000001" when "00101001100001110", -- t[21262] = 1
      "0000001" when "00101001100001111", -- t[21263] = 1
      "0000001" when "00101001100010000", -- t[21264] = 1
      "0000001" when "00101001100010001", -- t[21265] = 1
      "0000001" when "00101001100010010", -- t[21266] = 1
      "0000001" when "00101001100010011", -- t[21267] = 1
      "0000001" when "00101001100010100", -- t[21268] = 1
      "0000001" when "00101001100010101", -- t[21269] = 1
      "0000001" when "00101001100010110", -- t[21270] = 1
      "0000001" when "00101001100010111", -- t[21271] = 1
      "0000001" when "00101001100011000", -- t[21272] = 1
      "0000001" when "00101001100011001", -- t[21273] = 1
      "0000001" when "00101001100011010", -- t[21274] = 1
      "0000001" when "00101001100011011", -- t[21275] = 1
      "0000001" when "00101001100011100", -- t[21276] = 1
      "0000001" when "00101001100011101", -- t[21277] = 1
      "0000001" when "00101001100011110", -- t[21278] = 1
      "0000001" when "00101001100011111", -- t[21279] = 1
      "0000001" when "00101001100100000", -- t[21280] = 1
      "0000001" when "00101001100100001", -- t[21281] = 1
      "0000001" when "00101001100100010", -- t[21282] = 1
      "0000001" when "00101001100100011", -- t[21283] = 1
      "0000001" when "00101001100100100", -- t[21284] = 1
      "0000001" when "00101001100100101", -- t[21285] = 1
      "0000001" when "00101001100100110", -- t[21286] = 1
      "0000001" when "00101001100100111", -- t[21287] = 1
      "0000001" when "00101001100101000", -- t[21288] = 1
      "0000001" when "00101001100101001", -- t[21289] = 1
      "0000001" when "00101001100101010", -- t[21290] = 1
      "0000001" when "00101001100101011", -- t[21291] = 1
      "0000001" when "00101001100101100", -- t[21292] = 1
      "0000001" when "00101001100101101", -- t[21293] = 1
      "0000001" when "00101001100101110", -- t[21294] = 1
      "0000001" when "00101001100101111", -- t[21295] = 1
      "0000001" when "00101001100110000", -- t[21296] = 1
      "0000001" when "00101001100110001", -- t[21297] = 1
      "0000001" when "00101001100110010", -- t[21298] = 1
      "0000001" when "00101001100110011", -- t[21299] = 1
      "0000001" when "00101001100110100", -- t[21300] = 1
      "0000001" when "00101001100110101", -- t[21301] = 1
      "0000001" when "00101001100110110", -- t[21302] = 1
      "0000001" when "00101001100110111", -- t[21303] = 1
      "0000001" when "00101001100111000", -- t[21304] = 1
      "0000001" when "00101001100111001", -- t[21305] = 1
      "0000001" when "00101001100111010", -- t[21306] = 1
      "0000001" when "00101001100111011", -- t[21307] = 1
      "0000001" when "00101001100111100", -- t[21308] = 1
      "0000001" when "00101001100111101", -- t[21309] = 1
      "0000001" when "00101001100111110", -- t[21310] = 1
      "0000001" when "00101001100111111", -- t[21311] = 1
      "0000001" when "00101001101000000", -- t[21312] = 1
      "0000001" when "00101001101000001", -- t[21313] = 1
      "0000001" when "00101001101000010", -- t[21314] = 1
      "0000001" when "00101001101000011", -- t[21315] = 1
      "0000001" when "00101001101000100", -- t[21316] = 1
      "0000001" when "00101001101000101", -- t[21317] = 1
      "0000001" when "00101001101000110", -- t[21318] = 1
      "0000001" when "00101001101000111", -- t[21319] = 1
      "0000001" when "00101001101001000", -- t[21320] = 1
      "0000001" when "00101001101001001", -- t[21321] = 1
      "0000001" when "00101001101001010", -- t[21322] = 1
      "0000001" when "00101001101001011", -- t[21323] = 1
      "0000001" when "00101001101001100", -- t[21324] = 1
      "0000001" when "00101001101001101", -- t[21325] = 1
      "0000001" when "00101001101001110", -- t[21326] = 1
      "0000001" when "00101001101001111", -- t[21327] = 1
      "0000001" when "00101001101010000", -- t[21328] = 1
      "0000001" when "00101001101010001", -- t[21329] = 1
      "0000001" when "00101001101010010", -- t[21330] = 1
      "0000001" when "00101001101010011", -- t[21331] = 1
      "0000001" when "00101001101010100", -- t[21332] = 1
      "0000001" when "00101001101010101", -- t[21333] = 1
      "0000001" when "00101001101010110", -- t[21334] = 1
      "0000001" when "00101001101010111", -- t[21335] = 1
      "0000001" when "00101001101011000", -- t[21336] = 1
      "0000001" when "00101001101011001", -- t[21337] = 1
      "0000001" when "00101001101011010", -- t[21338] = 1
      "0000001" when "00101001101011011", -- t[21339] = 1
      "0000001" when "00101001101011100", -- t[21340] = 1
      "0000001" when "00101001101011101", -- t[21341] = 1
      "0000001" when "00101001101011110", -- t[21342] = 1
      "0000001" when "00101001101011111", -- t[21343] = 1
      "0000001" when "00101001101100000", -- t[21344] = 1
      "0000001" when "00101001101100001", -- t[21345] = 1
      "0000001" when "00101001101100010", -- t[21346] = 1
      "0000001" when "00101001101100011", -- t[21347] = 1
      "0000001" when "00101001101100100", -- t[21348] = 1
      "0000001" when "00101001101100101", -- t[21349] = 1
      "0000001" when "00101001101100110", -- t[21350] = 1
      "0000001" when "00101001101100111", -- t[21351] = 1
      "0000001" when "00101001101101000", -- t[21352] = 1
      "0000001" when "00101001101101001", -- t[21353] = 1
      "0000001" when "00101001101101010", -- t[21354] = 1
      "0000001" when "00101001101101011", -- t[21355] = 1
      "0000001" when "00101001101101100", -- t[21356] = 1
      "0000001" when "00101001101101101", -- t[21357] = 1
      "0000001" when "00101001101101110", -- t[21358] = 1
      "0000001" when "00101001101101111", -- t[21359] = 1
      "0000001" when "00101001101110000", -- t[21360] = 1
      "0000001" when "00101001101110001", -- t[21361] = 1
      "0000001" when "00101001101110010", -- t[21362] = 1
      "0000001" when "00101001101110011", -- t[21363] = 1
      "0000001" when "00101001101110100", -- t[21364] = 1
      "0000001" when "00101001101110101", -- t[21365] = 1
      "0000001" when "00101001101110110", -- t[21366] = 1
      "0000001" when "00101001101110111", -- t[21367] = 1
      "0000001" when "00101001101111000", -- t[21368] = 1
      "0000001" when "00101001101111001", -- t[21369] = 1
      "0000001" when "00101001101111010", -- t[21370] = 1
      "0000001" when "00101001101111011", -- t[21371] = 1
      "0000001" when "00101001101111100", -- t[21372] = 1
      "0000001" when "00101001101111101", -- t[21373] = 1
      "0000001" when "00101001101111110", -- t[21374] = 1
      "0000001" when "00101001101111111", -- t[21375] = 1
      "0000001" when "00101001110000000", -- t[21376] = 1
      "0000001" when "00101001110000001", -- t[21377] = 1
      "0000001" when "00101001110000010", -- t[21378] = 1
      "0000001" when "00101001110000011", -- t[21379] = 1
      "0000001" when "00101001110000100", -- t[21380] = 1
      "0000001" when "00101001110000101", -- t[21381] = 1
      "0000001" when "00101001110000110", -- t[21382] = 1
      "0000001" when "00101001110000111", -- t[21383] = 1
      "0000001" when "00101001110001000", -- t[21384] = 1
      "0000001" when "00101001110001001", -- t[21385] = 1
      "0000001" when "00101001110001010", -- t[21386] = 1
      "0000001" when "00101001110001011", -- t[21387] = 1
      "0000001" when "00101001110001100", -- t[21388] = 1
      "0000001" when "00101001110001101", -- t[21389] = 1
      "0000001" when "00101001110001110", -- t[21390] = 1
      "0000001" when "00101001110001111", -- t[21391] = 1
      "0000001" when "00101001110010000", -- t[21392] = 1
      "0000001" when "00101001110010001", -- t[21393] = 1
      "0000001" when "00101001110010010", -- t[21394] = 1
      "0000001" when "00101001110010011", -- t[21395] = 1
      "0000001" when "00101001110010100", -- t[21396] = 1
      "0000001" when "00101001110010101", -- t[21397] = 1
      "0000001" when "00101001110010110", -- t[21398] = 1
      "0000001" when "00101001110010111", -- t[21399] = 1
      "0000001" when "00101001110011000", -- t[21400] = 1
      "0000001" when "00101001110011001", -- t[21401] = 1
      "0000001" when "00101001110011010", -- t[21402] = 1
      "0000001" when "00101001110011011", -- t[21403] = 1
      "0000001" when "00101001110011100", -- t[21404] = 1
      "0000001" when "00101001110011101", -- t[21405] = 1
      "0000001" when "00101001110011110", -- t[21406] = 1
      "0000001" when "00101001110011111", -- t[21407] = 1
      "0000001" when "00101001110100000", -- t[21408] = 1
      "0000001" when "00101001110100001", -- t[21409] = 1
      "0000001" when "00101001110100010", -- t[21410] = 1
      "0000001" when "00101001110100011", -- t[21411] = 1
      "0000001" when "00101001110100100", -- t[21412] = 1
      "0000001" when "00101001110100101", -- t[21413] = 1
      "0000001" when "00101001110100110", -- t[21414] = 1
      "0000001" when "00101001110100111", -- t[21415] = 1
      "0000001" when "00101001110101000", -- t[21416] = 1
      "0000001" when "00101001110101001", -- t[21417] = 1
      "0000001" when "00101001110101010", -- t[21418] = 1
      "0000001" when "00101001110101011", -- t[21419] = 1
      "0000001" when "00101001110101100", -- t[21420] = 1
      "0000001" when "00101001110101101", -- t[21421] = 1
      "0000001" when "00101001110101110", -- t[21422] = 1
      "0000001" when "00101001110101111", -- t[21423] = 1
      "0000001" when "00101001110110000", -- t[21424] = 1
      "0000001" when "00101001110110001", -- t[21425] = 1
      "0000001" when "00101001110110010", -- t[21426] = 1
      "0000001" when "00101001110110011", -- t[21427] = 1
      "0000001" when "00101001110110100", -- t[21428] = 1
      "0000001" when "00101001110110101", -- t[21429] = 1
      "0000001" when "00101001110110110", -- t[21430] = 1
      "0000001" when "00101001110110111", -- t[21431] = 1
      "0000001" when "00101001110111000", -- t[21432] = 1
      "0000001" when "00101001110111001", -- t[21433] = 1
      "0000001" when "00101001110111010", -- t[21434] = 1
      "0000001" when "00101001110111011", -- t[21435] = 1
      "0000001" when "00101001110111100", -- t[21436] = 1
      "0000001" when "00101001110111101", -- t[21437] = 1
      "0000001" when "00101001110111110", -- t[21438] = 1
      "0000001" when "00101001110111111", -- t[21439] = 1
      "0000001" when "00101001111000000", -- t[21440] = 1
      "0000001" when "00101001111000001", -- t[21441] = 1
      "0000001" when "00101001111000010", -- t[21442] = 1
      "0000001" when "00101001111000011", -- t[21443] = 1
      "0000001" when "00101001111000100", -- t[21444] = 1
      "0000001" when "00101001111000101", -- t[21445] = 1
      "0000001" when "00101001111000110", -- t[21446] = 1
      "0000001" when "00101001111000111", -- t[21447] = 1
      "0000001" when "00101001111001000", -- t[21448] = 1
      "0000001" when "00101001111001001", -- t[21449] = 1
      "0000001" when "00101001111001010", -- t[21450] = 1
      "0000001" when "00101001111001011", -- t[21451] = 1
      "0000001" when "00101001111001100", -- t[21452] = 1
      "0000001" when "00101001111001101", -- t[21453] = 1
      "0000001" when "00101001111001110", -- t[21454] = 1
      "0000001" when "00101001111001111", -- t[21455] = 1
      "0000001" when "00101001111010000", -- t[21456] = 1
      "0000001" when "00101001111010001", -- t[21457] = 1
      "0000001" when "00101001111010010", -- t[21458] = 1
      "0000001" when "00101001111010011", -- t[21459] = 1
      "0000001" when "00101001111010100", -- t[21460] = 1
      "0000001" when "00101001111010101", -- t[21461] = 1
      "0000001" when "00101001111010110", -- t[21462] = 1
      "0000001" when "00101001111010111", -- t[21463] = 1
      "0000001" when "00101001111011000", -- t[21464] = 1
      "0000001" when "00101001111011001", -- t[21465] = 1
      "0000001" when "00101001111011010", -- t[21466] = 1
      "0000001" when "00101001111011011", -- t[21467] = 1
      "0000001" when "00101001111011100", -- t[21468] = 1
      "0000001" when "00101001111011101", -- t[21469] = 1
      "0000001" when "00101001111011110", -- t[21470] = 1
      "0000001" when "00101001111011111", -- t[21471] = 1
      "0000001" when "00101001111100000", -- t[21472] = 1
      "0000001" when "00101001111100001", -- t[21473] = 1
      "0000001" when "00101001111100010", -- t[21474] = 1
      "0000001" when "00101001111100011", -- t[21475] = 1
      "0000001" when "00101001111100100", -- t[21476] = 1
      "0000001" when "00101001111100101", -- t[21477] = 1
      "0000001" when "00101001111100110", -- t[21478] = 1
      "0000001" when "00101001111100111", -- t[21479] = 1
      "0000001" when "00101001111101000", -- t[21480] = 1
      "0000001" when "00101001111101001", -- t[21481] = 1
      "0000001" when "00101001111101010", -- t[21482] = 1
      "0000001" when "00101001111101011", -- t[21483] = 1
      "0000001" when "00101001111101100", -- t[21484] = 1
      "0000001" when "00101001111101101", -- t[21485] = 1
      "0000001" when "00101001111101110", -- t[21486] = 1
      "0000001" when "00101001111101111", -- t[21487] = 1
      "0000001" when "00101001111110000", -- t[21488] = 1
      "0000001" when "00101001111110001", -- t[21489] = 1
      "0000001" when "00101001111110010", -- t[21490] = 1
      "0000001" when "00101001111110011", -- t[21491] = 1
      "0000001" when "00101001111110100", -- t[21492] = 1
      "0000001" when "00101001111110101", -- t[21493] = 1
      "0000001" when "00101001111110110", -- t[21494] = 1
      "0000001" when "00101001111110111", -- t[21495] = 1
      "0000001" when "00101001111111000", -- t[21496] = 1
      "0000001" when "00101001111111001", -- t[21497] = 1
      "0000001" when "00101001111111010", -- t[21498] = 1
      "0000001" when "00101001111111011", -- t[21499] = 1
      "0000001" when "00101001111111100", -- t[21500] = 1
      "0000001" when "00101001111111101", -- t[21501] = 1
      "0000001" when "00101001111111110", -- t[21502] = 1
      "0000001" when "00101001111111111", -- t[21503] = 1
      "0000001" when "00101010000000000", -- t[21504] = 1
      "0000001" when "00101010000000001", -- t[21505] = 1
      "0000001" when "00101010000000010", -- t[21506] = 1
      "0000001" when "00101010000000011", -- t[21507] = 1
      "0000001" when "00101010000000100", -- t[21508] = 1
      "0000001" when "00101010000000101", -- t[21509] = 1
      "0000001" when "00101010000000110", -- t[21510] = 1
      "0000001" when "00101010000000111", -- t[21511] = 1
      "0000001" when "00101010000001000", -- t[21512] = 1
      "0000001" when "00101010000001001", -- t[21513] = 1
      "0000001" when "00101010000001010", -- t[21514] = 1
      "0000001" when "00101010000001011", -- t[21515] = 1
      "0000001" when "00101010000001100", -- t[21516] = 1
      "0000001" when "00101010000001101", -- t[21517] = 1
      "0000001" when "00101010000001110", -- t[21518] = 1
      "0000001" when "00101010000001111", -- t[21519] = 1
      "0000001" when "00101010000010000", -- t[21520] = 1
      "0000001" when "00101010000010001", -- t[21521] = 1
      "0000001" when "00101010000010010", -- t[21522] = 1
      "0000001" when "00101010000010011", -- t[21523] = 1
      "0000001" when "00101010000010100", -- t[21524] = 1
      "0000001" when "00101010000010101", -- t[21525] = 1
      "0000001" when "00101010000010110", -- t[21526] = 1
      "0000001" when "00101010000010111", -- t[21527] = 1
      "0000001" when "00101010000011000", -- t[21528] = 1
      "0000001" when "00101010000011001", -- t[21529] = 1
      "0000001" when "00101010000011010", -- t[21530] = 1
      "0000001" when "00101010000011011", -- t[21531] = 1
      "0000001" when "00101010000011100", -- t[21532] = 1
      "0000001" when "00101010000011101", -- t[21533] = 1
      "0000001" when "00101010000011110", -- t[21534] = 1
      "0000001" when "00101010000011111", -- t[21535] = 1
      "0000001" when "00101010000100000", -- t[21536] = 1
      "0000001" when "00101010000100001", -- t[21537] = 1
      "0000001" when "00101010000100010", -- t[21538] = 1
      "0000001" when "00101010000100011", -- t[21539] = 1
      "0000001" when "00101010000100100", -- t[21540] = 1
      "0000001" when "00101010000100101", -- t[21541] = 1
      "0000001" when "00101010000100110", -- t[21542] = 1
      "0000001" when "00101010000100111", -- t[21543] = 1
      "0000001" when "00101010000101000", -- t[21544] = 1
      "0000001" when "00101010000101001", -- t[21545] = 1
      "0000001" when "00101010000101010", -- t[21546] = 1
      "0000001" when "00101010000101011", -- t[21547] = 1
      "0000001" when "00101010000101100", -- t[21548] = 1
      "0000001" when "00101010000101101", -- t[21549] = 1
      "0000001" when "00101010000101110", -- t[21550] = 1
      "0000001" when "00101010000101111", -- t[21551] = 1
      "0000001" when "00101010000110000", -- t[21552] = 1
      "0000001" when "00101010000110001", -- t[21553] = 1
      "0000001" when "00101010000110010", -- t[21554] = 1
      "0000001" when "00101010000110011", -- t[21555] = 1
      "0000001" when "00101010000110100", -- t[21556] = 1
      "0000001" when "00101010000110101", -- t[21557] = 1
      "0000001" when "00101010000110110", -- t[21558] = 1
      "0000001" when "00101010000110111", -- t[21559] = 1
      "0000001" when "00101010000111000", -- t[21560] = 1
      "0000001" when "00101010000111001", -- t[21561] = 1
      "0000001" when "00101010000111010", -- t[21562] = 1
      "0000001" when "00101010000111011", -- t[21563] = 1
      "0000001" when "00101010000111100", -- t[21564] = 1
      "0000001" when "00101010000111101", -- t[21565] = 1
      "0000001" when "00101010000111110", -- t[21566] = 1
      "0000001" when "00101010000111111", -- t[21567] = 1
      "0000001" when "00101010001000000", -- t[21568] = 1
      "0000001" when "00101010001000001", -- t[21569] = 1
      "0000001" when "00101010001000010", -- t[21570] = 1
      "0000001" when "00101010001000011", -- t[21571] = 1
      "0000001" when "00101010001000100", -- t[21572] = 1
      "0000001" when "00101010001000101", -- t[21573] = 1
      "0000001" when "00101010001000110", -- t[21574] = 1
      "0000001" when "00101010001000111", -- t[21575] = 1
      "0000001" when "00101010001001000", -- t[21576] = 1
      "0000001" when "00101010001001001", -- t[21577] = 1
      "0000001" when "00101010001001010", -- t[21578] = 1
      "0000001" when "00101010001001011", -- t[21579] = 1
      "0000001" when "00101010001001100", -- t[21580] = 1
      "0000001" when "00101010001001101", -- t[21581] = 1
      "0000001" when "00101010001001110", -- t[21582] = 1
      "0000001" when "00101010001001111", -- t[21583] = 1
      "0000001" when "00101010001010000", -- t[21584] = 1
      "0000001" when "00101010001010001", -- t[21585] = 1
      "0000001" when "00101010001010010", -- t[21586] = 1
      "0000001" when "00101010001010011", -- t[21587] = 1
      "0000001" when "00101010001010100", -- t[21588] = 1
      "0000001" when "00101010001010101", -- t[21589] = 1
      "0000001" when "00101010001010110", -- t[21590] = 1
      "0000001" when "00101010001010111", -- t[21591] = 1
      "0000001" when "00101010001011000", -- t[21592] = 1
      "0000001" when "00101010001011001", -- t[21593] = 1
      "0000001" when "00101010001011010", -- t[21594] = 1
      "0000001" when "00101010001011011", -- t[21595] = 1
      "0000001" when "00101010001011100", -- t[21596] = 1
      "0000001" when "00101010001011101", -- t[21597] = 1
      "0000001" when "00101010001011110", -- t[21598] = 1
      "0000001" when "00101010001011111", -- t[21599] = 1
      "0000001" when "00101010001100000", -- t[21600] = 1
      "0000001" when "00101010001100001", -- t[21601] = 1
      "0000001" when "00101010001100010", -- t[21602] = 1
      "0000001" when "00101010001100011", -- t[21603] = 1
      "0000001" when "00101010001100100", -- t[21604] = 1
      "0000001" when "00101010001100101", -- t[21605] = 1
      "0000001" when "00101010001100110", -- t[21606] = 1
      "0000001" when "00101010001100111", -- t[21607] = 1
      "0000001" when "00101010001101000", -- t[21608] = 1
      "0000001" when "00101010001101001", -- t[21609] = 1
      "0000001" when "00101010001101010", -- t[21610] = 1
      "0000001" when "00101010001101011", -- t[21611] = 1
      "0000001" when "00101010001101100", -- t[21612] = 1
      "0000001" when "00101010001101101", -- t[21613] = 1
      "0000001" when "00101010001101110", -- t[21614] = 1
      "0000001" when "00101010001101111", -- t[21615] = 1
      "0000001" when "00101010001110000", -- t[21616] = 1
      "0000001" when "00101010001110001", -- t[21617] = 1
      "0000001" when "00101010001110010", -- t[21618] = 1
      "0000001" when "00101010001110011", -- t[21619] = 1
      "0000001" when "00101010001110100", -- t[21620] = 1
      "0000001" when "00101010001110101", -- t[21621] = 1
      "0000001" when "00101010001110110", -- t[21622] = 1
      "0000001" when "00101010001110111", -- t[21623] = 1
      "0000001" when "00101010001111000", -- t[21624] = 1
      "0000001" when "00101010001111001", -- t[21625] = 1
      "0000001" when "00101010001111010", -- t[21626] = 1
      "0000001" when "00101010001111011", -- t[21627] = 1
      "0000001" when "00101010001111100", -- t[21628] = 1
      "0000001" when "00101010001111101", -- t[21629] = 1
      "0000001" when "00101010001111110", -- t[21630] = 1
      "0000001" when "00101010001111111", -- t[21631] = 1
      "0000001" when "00101010010000000", -- t[21632] = 1
      "0000001" when "00101010010000001", -- t[21633] = 1
      "0000001" when "00101010010000010", -- t[21634] = 1
      "0000001" when "00101010010000011", -- t[21635] = 1
      "0000001" when "00101010010000100", -- t[21636] = 1
      "0000001" when "00101010010000101", -- t[21637] = 1
      "0000001" when "00101010010000110", -- t[21638] = 1
      "0000001" when "00101010010000111", -- t[21639] = 1
      "0000001" when "00101010010001000", -- t[21640] = 1
      "0000001" when "00101010010001001", -- t[21641] = 1
      "0000001" when "00101010010001010", -- t[21642] = 1
      "0000001" when "00101010010001011", -- t[21643] = 1
      "0000001" when "00101010010001100", -- t[21644] = 1
      "0000001" when "00101010010001101", -- t[21645] = 1
      "0000001" when "00101010010001110", -- t[21646] = 1
      "0000001" when "00101010010001111", -- t[21647] = 1
      "0000001" when "00101010010010000", -- t[21648] = 1
      "0000001" when "00101010010010001", -- t[21649] = 1
      "0000001" when "00101010010010010", -- t[21650] = 1
      "0000001" when "00101010010010011", -- t[21651] = 1
      "0000001" when "00101010010010100", -- t[21652] = 1
      "0000001" when "00101010010010101", -- t[21653] = 1
      "0000001" when "00101010010010110", -- t[21654] = 1
      "0000001" when "00101010010010111", -- t[21655] = 1
      "0000001" when "00101010010011000", -- t[21656] = 1
      "0000001" when "00101010010011001", -- t[21657] = 1
      "0000001" when "00101010010011010", -- t[21658] = 1
      "0000001" when "00101010010011011", -- t[21659] = 1
      "0000001" when "00101010010011100", -- t[21660] = 1
      "0000001" when "00101010010011101", -- t[21661] = 1
      "0000001" when "00101010010011110", -- t[21662] = 1
      "0000001" when "00101010010011111", -- t[21663] = 1
      "0000001" when "00101010010100000", -- t[21664] = 1
      "0000001" when "00101010010100001", -- t[21665] = 1
      "0000001" when "00101010010100010", -- t[21666] = 1
      "0000001" when "00101010010100011", -- t[21667] = 1
      "0000001" when "00101010010100100", -- t[21668] = 1
      "0000001" when "00101010010100101", -- t[21669] = 1
      "0000001" when "00101010010100110", -- t[21670] = 1
      "0000001" when "00101010010100111", -- t[21671] = 1
      "0000001" when "00101010010101000", -- t[21672] = 1
      "0000001" when "00101010010101001", -- t[21673] = 1
      "0000001" when "00101010010101010", -- t[21674] = 1
      "0000001" when "00101010010101011", -- t[21675] = 1
      "0000001" when "00101010010101100", -- t[21676] = 1
      "0000001" when "00101010010101101", -- t[21677] = 1
      "0000001" when "00101010010101110", -- t[21678] = 1
      "0000001" when "00101010010101111", -- t[21679] = 1
      "0000001" when "00101010010110000", -- t[21680] = 1
      "0000001" when "00101010010110001", -- t[21681] = 1
      "0000001" when "00101010010110010", -- t[21682] = 1
      "0000001" when "00101010010110011", -- t[21683] = 1
      "0000001" when "00101010010110100", -- t[21684] = 1
      "0000001" when "00101010010110101", -- t[21685] = 1
      "0000001" when "00101010010110110", -- t[21686] = 1
      "0000001" when "00101010010110111", -- t[21687] = 1
      "0000001" when "00101010010111000", -- t[21688] = 1
      "0000001" when "00101010010111001", -- t[21689] = 1
      "0000001" when "00101010010111010", -- t[21690] = 1
      "0000001" when "00101010010111011", -- t[21691] = 1
      "0000001" when "00101010010111100", -- t[21692] = 1
      "0000001" when "00101010010111101", -- t[21693] = 1
      "0000001" when "00101010010111110", -- t[21694] = 1
      "0000001" when "00101010010111111", -- t[21695] = 1
      "0000001" when "00101010011000000", -- t[21696] = 1
      "0000001" when "00101010011000001", -- t[21697] = 1
      "0000001" when "00101010011000010", -- t[21698] = 1
      "0000001" when "00101010011000011", -- t[21699] = 1
      "0000001" when "00101010011000100", -- t[21700] = 1
      "0000001" when "00101010011000101", -- t[21701] = 1
      "0000001" when "00101010011000110", -- t[21702] = 1
      "0000001" when "00101010011000111", -- t[21703] = 1
      "0000001" when "00101010011001000", -- t[21704] = 1
      "0000001" when "00101010011001001", -- t[21705] = 1
      "0000001" when "00101010011001010", -- t[21706] = 1
      "0000001" when "00101010011001011", -- t[21707] = 1
      "0000001" when "00101010011001100", -- t[21708] = 1
      "0000001" when "00101010011001101", -- t[21709] = 1
      "0000001" when "00101010011001110", -- t[21710] = 1
      "0000001" when "00101010011001111", -- t[21711] = 1
      "0000001" when "00101010011010000", -- t[21712] = 1
      "0000001" when "00101010011010001", -- t[21713] = 1
      "0000001" when "00101010011010010", -- t[21714] = 1
      "0000001" when "00101010011010011", -- t[21715] = 1
      "0000001" when "00101010011010100", -- t[21716] = 1
      "0000001" when "00101010011010101", -- t[21717] = 1
      "0000001" when "00101010011010110", -- t[21718] = 1
      "0000001" when "00101010011010111", -- t[21719] = 1
      "0000001" when "00101010011011000", -- t[21720] = 1
      "0000001" when "00101010011011001", -- t[21721] = 1
      "0000001" when "00101010011011010", -- t[21722] = 1
      "0000001" when "00101010011011011", -- t[21723] = 1
      "0000001" when "00101010011011100", -- t[21724] = 1
      "0000001" when "00101010011011101", -- t[21725] = 1
      "0000001" when "00101010011011110", -- t[21726] = 1
      "0000001" when "00101010011011111", -- t[21727] = 1
      "0000001" when "00101010011100000", -- t[21728] = 1
      "0000001" when "00101010011100001", -- t[21729] = 1
      "0000001" when "00101010011100010", -- t[21730] = 1
      "0000001" when "00101010011100011", -- t[21731] = 1
      "0000001" when "00101010011100100", -- t[21732] = 1
      "0000001" when "00101010011100101", -- t[21733] = 1
      "0000001" when "00101010011100110", -- t[21734] = 1
      "0000001" when "00101010011100111", -- t[21735] = 1
      "0000001" when "00101010011101000", -- t[21736] = 1
      "0000001" when "00101010011101001", -- t[21737] = 1
      "0000001" when "00101010011101010", -- t[21738] = 1
      "0000001" when "00101010011101011", -- t[21739] = 1
      "0000001" when "00101010011101100", -- t[21740] = 1
      "0000001" when "00101010011101101", -- t[21741] = 1
      "0000001" when "00101010011101110", -- t[21742] = 1
      "0000001" when "00101010011101111", -- t[21743] = 1
      "0000001" when "00101010011110000", -- t[21744] = 1
      "0000001" when "00101010011110001", -- t[21745] = 1
      "0000001" when "00101010011110010", -- t[21746] = 1
      "0000001" when "00101010011110011", -- t[21747] = 1
      "0000001" when "00101010011110100", -- t[21748] = 1
      "0000001" when "00101010011110101", -- t[21749] = 1
      "0000001" when "00101010011110110", -- t[21750] = 1
      "0000001" when "00101010011110111", -- t[21751] = 1
      "0000001" when "00101010011111000", -- t[21752] = 1
      "0000001" when "00101010011111001", -- t[21753] = 1
      "0000001" when "00101010011111010", -- t[21754] = 1
      "0000001" when "00101010011111011", -- t[21755] = 1
      "0000001" when "00101010011111100", -- t[21756] = 1
      "0000001" when "00101010011111101", -- t[21757] = 1
      "0000001" when "00101010011111110", -- t[21758] = 1
      "0000001" when "00101010011111111", -- t[21759] = 1
      "0000001" when "00101010100000000", -- t[21760] = 1
      "0000001" when "00101010100000001", -- t[21761] = 1
      "0000001" when "00101010100000010", -- t[21762] = 1
      "0000001" when "00101010100000011", -- t[21763] = 1
      "0000001" when "00101010100000100", -- t[21764] = 1
      "0000001" when "00101010100000101", -- t[21765] = 1
      "0000001" when "00101010100000110", -- t[21766] = 1
      "0000001" when "00101010100000111", -- t[21767] = 1
      "0000001" when "00101010100001000", -- t[21768] = 1
      "0000001" when "00101010100001001", -- t[21769] = 1
      "0000001" when "00101010100001010", -- t[21770] = 1
      "0000001" when "00101010100001011", -- t[21771] = 1
      "0000001" when "00101010100001100", -- t[21772] = 1
      "0000001" when "00101010100001101", -- t[21773] = 1
      "0000001" when "00101010100001110", -- t[21774] = 1
      "0000001" when "00101010100001111", -- t[21775] = 1
      "0000001" when "00101010100010000", -- t[21776] = 1
      "0000001" when "00101010100010001", -- t[21777] = 1
      "0000001" when "00101010100010010", -- t[21778] = 1
      "0000001" when "00101010100010011", -- t[21779] = 1
      "0000001" when "00101010100010100", -- t[21780] = 1
      "0000001" when "00101010100010101", -- t[21781] = 1
      "0000001" when "00101010100010110", -- t[21782] = 1
      "0000001" when "00101010100010111", -- t[21783] = 1
      "0000001" when "00101010100011000", -- t[21784] = 1
      "0000001" when "00101010100011001", -- t[21785] = 1
      "0000001" when "00101010100011010", -- t[21786] = 1
      "0000001" when "00101010100011011", -- t[21787] = 1
      "0000001" when "00101010100011100", -- t[21788] = 1
      "0000001" when "00101010100011101", -- t[21789] = 1
      "0000001" when "00101010100011110", -- t[21790] = 1
      "0000001" when "00101010100011111", -- t[21791] = 1
      "0000001" when "00101010100100000", -- t[21792] = 1
      "0000001" when "00101010100100001", -- t[21793] = 1
      "0000001" when "00101010100100010", -- t[21794] = 1
      "0000001" when "00101010100100011", -- t[21795] = 1
      "0000001" when "00101010100100100", -- t[21796] = 1
      "0000001" when "00101010100100101", -- t[21797] = 1
      "0000001" when "00101010100100110", -- t[21798] = 1
      "0000001" when "00101010100100111", -- t[21799] = 1
      "0000001" when "00101010100101000", -- t[21800] = 1
      "0000001" when "00101010100101001", -- t[21801] = 1
      "0000001" when "00101010100101010", -- t[21802] = 1
      "0000001" when "00101010100101011", -- t[21803] = 1
      "0000001" when "00101010100101100", -- t[21804] = 1
      "0000001" when "00101010100101101", -- t[21805] = 1
      "0000001" when "00101010100101110", -- t[21806] = 1
      "0000001" when "00101010100101111", -- t[21807] = 1
      "0000001" when "00101010100110000", -- t[21808] = 1
      "0000001" when "00101010100110001", -- t[21809] = 1
      "0000001" when "00101010100110010", -- t[21810] = 1
      "0000001" when "00101010100110011", -- t[21811] = 1
      "0000001" when "00101010100110100", -- t[21812] = 1
      "0000001" when "00101010100110101", -- t[21813] = 1
      "0000001" when "00101010100110110", -- t[21814] = 1
      "0000001" when "00101010100110111", -- t[21815] = 1
      "0000001" when "00101010100111000", -- t[21816] = 1
      "0000001" when "00101010100111001", -- t[21817] = 1
      "0000001" when "00101010100111010", -- t[21818] = 1
      "0000001" when "00101010100111011", -- t[21819] = 1
      "0000001" when "00101010100111100", -- t[21820] = 1
      "0000001" when "00101010100111101", -- t[21821] = 1
      "0000001" when "00101010100111110", -- t[21822] = 1
      "0000001" when "00101010100111111", -- t[21823] = 1
      "0000001" when "00101010101000000", -- t[21824] = 1
      "0000001" when "00101010101000001", -- t[21825] = 1
      "0000001" when "00101010101000010", -- t[21826] = 1
      "0000001" when "00101010101000011", -- t[21827] = 1
      "0000001" when "00101010101000100", -- t[21828] = 1
      "0000001" when "00101010101000101", -- t[21829] = 1
      "0000001" when "00101010101000110", -- t[21830] = 1
      "0000001" when "00101010101000111", -- t[21831] = 1
      "0000001" when "00101010101001000", -- t[21832] = 1
      "0000001" when "00101010101001001", -- t[21833] = 1
      "0000001" when "00101010101001010", -- t[21834] = 1
      "0000001" when "00101010101001011", -- t[21835] = 1
      "0000001" when "00101010101001100", -- t[21836] = 1
      "0000001" when "00101010101001101", -- t[21837] = 1
      "0000001" when "00101010101001110", -- t[21838] = 1
      "0000001" when "00101010101001111", -- t[21839] = 1
      "0000001" when "00101010101010000", -- t[21840] = 1
      "0000001" when "00101010101010001", -- t[21841] = 1
      "0000001" when "00101010101010010", -- t[21842] = 1
      "0000001" when "00101010101010011", -- t[21843] = 1
      "0000001" when "00101010101010100", -- t[21844] = 1
      "0000001" when "00101010101010101", -- t[21845] = 1
      "0000001" when "00101010101010110", -- t[21846] = 1
      "0000001" when "00101010101010111", -- t[21847] = 1
      "0000001" when "00101010101011000", -- t[21848] = 1
      "0000001" when "00101010101011001", -- t[21849] = 1
      "0000001" when "00101010101011010", -- t[21850] = 1
      "0000001" when "00101010101011011", -- t[21851] = 1
      "0000001" when "00101010101011100", -- t[21852] = 1
      "0000001" when "00101010101011101", -- t[21853] = 1
      "0000001" when "00101010101011110", -- t[21854] = 1
      "0000001" when "00101010101011111", -- t[21855] = 1
      "0000001" when "00101010101100000", -- t[21856] = 1
      "0000001" when "00101010101100001", -- t[21857] = 1
      "0000001" when "00101010101100010", -- t[21858] = 1
      "0000001" when "00101010101100011", -- t[21859] = 1
      "0000001" when "00101010101100100", -- t[21860] = 1
      "0000001" when "00101010101100101", -- t[21861] = 1
      "0000001" when "00101010101100110", -- t[21862] = 1
      "0000001" when "00101010101100111", -- t[21863] = 1
      "0000001" when "00101010101101000", -- t[21864] = 1
      "0000001" when "00101010101101001", -- t[21865] = 1
      "0000001" when "00101010101101010", -- t[21866] = 1
      "0000001" when "00101010101101011", -- t[21867] = 1
      "0000001" when "00101010101101100", -- t[21868] = 1
      "0000001" when "00101010101101101", -- t[21869] = 1
      "0000001" when "00101010101101110", -- t[21870] = 1
      "0000001" when "00101010101101111", -- t[21871] = 1
      "0000001" when "00101010101110000", -- t[21872] = 1
      "0000001" when "00101010101110001", -- t[21873] = 1
      "0000001" when "00101010101110010", -- t[21874] = 1
      "0000001" when "00101010101110011", -- t[21875] = 1
      "0000001" when "00101010101110100", -- t[21876] = 1
      "0000001" when "00101010101110101", -- t[21877] = 1
      "0000001" when "00101010101110110", -- t[21878] = 1
      "0000001" when "00101010101110111", -- t[21879] = 1
      "0000001" when "00101010101111000", -- t[21880] = 1
      "0000001" when "00101010101111001", -- t[21881] = 1
      "0000001" when "00101010101111010", -- t[21882] = 1
      "0000001" when "00101010101111011", -- t[21883] = 1
      "0000001" when "00101010101111100", -- t[21884] = 1
      "0000001" when "00101010101111101", -- t[21885] = 1
      "0000001" when "00101010101111110", -- t[21886] = 1
      "0000001" when "00101010101111111", -- t[21887] = 1
      "0000001" when "00101010110000000", -- t[21888] = 1
      "0000001" when "00101010110000001", -- t[21889] = 1
      "0000001" when "00101010110000010", -- t[21890] = 1
      "0000001" when "00101010110000011", -- t[21891] = 1
      "0000001" when "00101010110000100", -- t[21892] = 1
      "0000001" when "00101010110000101", -- t[21893] = 1
      "0000001" when "00101010110000110", -- t[21894] = 1
      "0000001" when "00101010110000111", -- t[21895] = 1
      "0000001" when "00101010110001000", -- t[21896] = 1
      "0000001" when "00101010110001001", -- t[21897] = 1
      "0000001" when "00101010110001010", -- t[21898] = 1
      "0000001" when "00101010110001011", -- t[21899] = 1
      "0000001" when "00101010110001100", -- t[21900] = 1
      "0000001" when "00101010110001101", -- t[21901] = 1
      "0000001" when "00101010110001110", -- t[21902] = 1
      "0000001" when "00101010110001111", -- t[21903] = 1
      "0000001" when "00101010110010000", -- t[21904] = 1
      "0000001" when "00101010110010001", -- t[21905] = 1
      "0000001" when "00101010110010010", -- t[21906] = 1
      "0000001" when "00101010110010011", -- t[21907] = 1
      "0000001" when "00101010110010100", -- t[21908] = 1
      "0000001" when "00101010110010101", -- t[21909] = 1
      "0000001" when "00101010110010110", -- t[21910] = 1
      "0000001" when "00101010110010111", -- t[21911] = 1
      "0000001" when "00101010110011000", -- t[21912] = 1
      "0000001" when "00101010110011001", -- t[21913] = 1
      "0000001" when "00101010110011010", -- t[21914] = 1
      "0000001" when "00101010110011011", -- t[21915] = 1
      "0000001" when "00101010110011100", -- t[21916] = 1
      "0000001" when "00101010110011101", -- t[21917] = 1
      "0000001" when "00101010110011110", -- t[21918] = 1
      "0000001" when "00101010110011111", -- t[21919] = 1
      "0000001" when "00101010110100000", -- t[21920] = 1
      "0000001" when "00101010110100001", -- t[21921] = 1
      "0000001" when "00101010110100010", -- t[21922] = 1
      "0000001" when "00101010110100011", -- t[21923] = 1
      "0000001" when "00101010110100100", -- t[21924] = 1
      "0000001" when "00101010110100101", -- t[21925] = 1
      "0000001" when "00101010110100110", -- t[21926] = 1
      "0000001" when "00101010110100111", -- t[21927] = 1
      "0000001" when "00101010110101000", -- t[21928] = 1
      "0000001" when "00101010110101001", -- t[21929] = 1
      "0000001" when "00101010110101010", -- t[21930] = 1
      "0000001" when "00101010110101011", -- t[21931] = 1
      "0000001" when "00101010110101100", -- t[21932] = 1
      "0000001" when "00101010110101101", -- t[21933] = 1
      "0000001" when "00101010110101110", -- t[21934] = 1
      "0000001" when "00101010110101111", -- t[21935] = 1
      "0000001" when "00101010110110000", -- t[21936] = 1
      "0000001" when "00101010110110001", -- t[21937] = 1
      "0000001" when "00101010110110010", -- t[21938] = 1
      "0000001" when "00101010110110011", -- t[21939] = 1
      "0000001" when "00101010110110100", -- t[21940] = 1
      "0000001" when "00101010110110101", -- t[21941] = 1
      "0000001" when "00101010110110110", -- t[21942] = 1
      "0000001" when "00101010110110111", -- t[21943] = 1
      "0000001" when "00101010110111000", -- t[21944] = 1
      "0000001" when "00101010110111001", -- t[21945] = 1
      "0000001" when "00101010110111010", -- t[21946] = 1
      "0000001" when "00101010110111011", -- t[21947] = 1
      "0000001" when "00101010110111100", -- t[21948] = 1
      "0000001" when "00101010110111101", -- t[21949] = 1
      "0000001" when "00101010110111110", -- t[21950] = 1
      "0000001" when "00101010110111111", -- t[21951] = 1
      "0000001" when "00101010111000000", -- t[21952] = 1
      "0000001" when "00101010111000001", -- t[21953] = 1
      "0000001" when "00101010111000010", -- t[21954] = 1
      "0000001" when "00101010111000011", -- t[21955] = 1
      "0000001" when "00101010111000100", -- t[21956] = 1
      "0000001" when "00101010111000101", -- t[21957] = 1
      "0000001" when "00101010111000110", -- t[21958] = 1
      "0000001" when "00101010111000111", -- t[21959] = 1
      "0000001" when "00101010111001000", -- t[21960] = 1
      "0000001" when "00101010111001001", -- t[21961] = 1
      "0000001" when "00101010111001010", -- t[21962] = 1
      "0000001" when "00101010111001011", -- t[21963] = 1
      "0000001" when "00101010111001100", -- t[21964] = 1
      "0000001" when "00101010111001101", -- t[21965] = 1
      "0000001" when "00101010111001110", -- t[21966] = 1
      "0000001" when "00101010111001111", -- t[21967] = 1
      "0000001" when "00101010111010000", -- t[21968] = 1
      "0000001" when "00101010111010001", -- t[21969] = 1
      "0000001" when "00101010111010010", -- t[21970] = 1
      "0000001" when "00101010111010011", -- t[21971] = 1
      "0000001" when "00101010111010100", -- t[21972] = 1
      "0000001" when "00101010111010101", -- t[21973] = 1
      "0000001" when "00101010111010110", -- t[21974] = 1
      "0000001" when "00101010111010111", -- t[21975] = 1
      "0000001" when "00101010111011000", -- t[21976] = 1
      "0000001" when "00101010111011001", -- t[21977] = 1
      "0000001" when "00101010111011010", -- t[21978] = 1
      "0000001" when "00101010111011011", -- t[21979] = 1
      "0000001" when "00101010111011100", -- t[21980] = 1
      "0000001" when "00101010111011101", -- t[21981] = 1
      "0000001" when "00101010111011110", -- t[21982] = 1
      "0000001" when "00101010111011111", -- t[21983] = 1
      "0000001" when "00101010111100000", -- t[21984] = 1
      "0000001" when "00101010111100001", -- t[21985] = 1
      "0000001" when "00101010111100010", -- t[21986] = 1
      "0000001" when "00101010111100011", -- t[21987] = 1
      "0000001" when "00101010111100100", -- t[21988] = 1
      "0000001" when "00101010111100101", -- t[21989] = 1
      "0000001" when "00101010111100110", -- t[21990] = 1
      "0000001" when "00101010111100111", -- t[21991] = 1
      "0000001" when "00101010111101000", -- t[21992] = 1
      "0000001" when "00101010111101001", -- t[21993] = 1
      "0000001" when "00101010111101010", -- t[21994] = 1
      "0000001" when "00101010111101011", -- t[21995] = 1
      "0000001" when "00101010111101100", -- t[21996] = 1
      "0000001" when "00101010111101101", -- t[21997] = 1
      "0000001" when "00101010111101110", -- t[21998] = 1
      "0000001" when "00101010111101111", -- t[21999] = 1
      "0000001" when "00101010111110000", -- t[22000] = 1
      "0000001" when "00101010111110001", -- t[22001] = 1
      "0000001" when "00101010111110010", -- t[22002] = 1
      "0000001" when "00101010111110011", -- t[22003] = 1
      "0000001" when "00101010111110100", -- t[22004] = 1
      "0000001" when "00101010111110101", -- t[22005] = 1
      "0000001" when "00101010111110110", -- t[22006] = 1
      "0000001" when "00101010111110111", -- t[22007] = 1
      "0000001" when "00101010111111000", -- t[22008] = 1
      "0000001" when "00101010111111001", -- t[22009] = 1
      "0000001" when "00101010111111010", -- t[22010] = 1
      "0000001" when "00101010111111011", -- t[22011] = 1
      "0000001" when "00101010111111100", -- t[22012] = 1
      "0000001" when "00101010111111101", -- t[22013] = 1
      "0000001" when "00101010111111110", -- t[22014] = 1
      "0000001" when "00101010111111111", -- t[22015] = 1
      "0000001" when "00101011000000000", -- t[22016] = 1
      "0000001" when "00101011000000001", -- t[22017] = 1
      "0000001" when "00101011000000010", -- t[22018] = 1
      "0000001" when "00101011000000011", -- t[22019] = 1
      "0000001" when "00101011000000100", -- t[22020] = 1
      "0000001" when "00101011000000101", -- t[22021] = 1
      "0000001" when "00101011000000110", -- t[22022] = 1
      "0000001" when "00101011000000111", -- t[22023] = 1
      "0000001" when "00101011000001000", -- t[22024] = 1
      "0000001" when "00101011000001001", -- t[22025] = 1
      "0000001" when "00101011000001010", -- t[22026] = 1
      "0000001" when "00101011000001011", -- t[22027] = 1
      "0000001" when "00101011000001100", -- t[22028] = 1
      "0000001" when "00101011000001101", -- t[22029] = 1
      "0000001" when "00101011000001110", -- t[22030] = 1
      "0000001" when "00101011000001111", -- t[22031] = 1
      "0000001" when "00101011000010000", -- t[22032] = 1
      "0000001" when "00101011000010001", -- t[22033] = 1
      "0000001" when "00101011000010010", -- t[22034] = 1
      "0000001" when "00101011000010011", -- t[22035] = 1
      "0000001" when "00101011000010100", -- t[22036] = 1
      "0000001" when "00101011000010101", -- t[22037] = 1
      "0000001" when "00101011000010110", -- t[22038] = 1
      "0000001" when "00101011000010111", -- t[22039] = 1
      "0000001" when "00101011000011000", -- t[22040] = 1
      "0000001" when "00101011000011001", -- t[22041] = 1
      "0000001" when "00101011000011010", -- t[22042] = 1
      "0000001" when "00101011000011011", -- t[22043] = 1
      "0000001" when "00101011000011100", -- t[22044] = 1
      "0000001" when "00101011000011101", -- t[22045] = 1
      "0000001" when "00101011000011110", -- t[22046] = 1
      "0000001" when "00101011000011111", -- t[22047] = 1
      "0000001" when "00101011000100000", -- t[22048] = 1
      "0000001" when "00101011000100001", -- t[22049] = 1
      "0000001" when "00101011000100010", -- t[22050] = 1
      "0000001" when "00101011000100011", -- t[22051] = 1
      "0000001" when "00101011000100100", -- t[22052] = 1
      "0000001" when "00101011000100101", -- t[22053] = 1
      "0000001" when "00101011000100110", -- t[22054] = 1
      "0000001" when "00101011000100111", -- t[22055] = 1
      "0000001" when "00101011000101000", -- t[22056] = 1
      "0000001" when "00101011000101001", -- t[22057] = 1
      "0000001" when "00101011000101010", -- t[22058] = 1
      "0000001" when "00101011000101011", -- t[22059] = 1
      "0000001" when "00101011000101100", -- t[22060] = 1
      "0000001" when "00101011000101101", -- t[22061] = 1
      "0000001" when "00101011000101110", -- t[22062] = 1
      "0000001" when "00101011000101111", -- t[22063] = 1
      "0000001" when "00101011000110000", -- t[22064] = 1
      "0000001" when "00101011000110001", -- t[22065] = 1
      "0000001" when "00101011000110010", -- t[22066] = 1
      "0000001" when "00101011000110011", -- t[22067] = 1
      "0000001" when "00101011000110100", -- t[22068] = 1
      "0000001" when "00101011000110101", -- t[22069] = 1
      "0000001" when "00101011000110110", -- t[22070] = 1
      "0000001" when "00101011000110111", -- t[22071] = 1
      "0000001" when "00101011000111000", -- t[22072] = 1
      "0000001" when "00101011000111001", -- t[22073] = 1
      "0000001" when "00101011000111010", -- t[22074] = 1
      "0000001" when "00101011000111011", -- t[22075] = 1
      "0000001" when "00101011000111100", -- t[22076] = 1
      "0000001" when "00101011000111101", -- t[22077] = 1
      "0000001" when "00101011000111110", -- t[22078] = 1
      "0000001" when "00101011000111111", -- t[22079] = 1
      "0000001" when "00101011001000000", -- t[22080] = 1
      "0000001" when "00101011001000001", -- t[22081] = 1
      "0000001" when "00101011001000010", -- t[22082] = 1
      "0000001" when "00101011001000011", -- t[22083] = 1
      "0000001" when "00101011001000100", -- t[22084] = 1
      "0000001" when "00101011001000101", -- t[22085] = 1
      "0000001" when "00101011001000110", -- t[22086] = 1
      "0000001" when "00101011001000111", -- t[22087] = 1
      "0000001" when "00101011001001000", -- t[22088] = 1
      "0000001" when "00101011001001001", -- t[22089] = 1
      "0000001" when "00101011001001010", -- t[22090] = 1
      "0000001" when "00101011001001011", -- t[22091] = 1
      "0000001" when "00101011001001100", -- t[22092] = 1
      "0000001" when "00101011001001101", -- t[22093] = 1
      "0000001" when "00101011001001110", -- t[22094] = 1
      "0000001" when "00101011001001111", -- t[22095] = 1
      "0000001" when "00101011001010000", -- t[22096] = 1
      "0000001" when "00101011001010001", -- t[22097] = 1
      "0000001" when "00101011001010010", -- t[22098] = 1
      "0000001" when "00101011001010011", -- t[22099] = 1
      "0000001" when "00101011001010100", -- t[22100] = 1
      "0000001" when "00101011001010101", -- t[22101] = 1
      "0000001" when "00101011001010110", -- t[22102] = 1
      "0000001" when "00101011001010111", -- t[22103] = 1
      "0000001" when "00101011001011000", -- t[22104] = 1
      "0000001" when "00101011001011001", -- t[22105] = 1
      "0000001" when "00101011001011010", -- t[22106] = 1
      "0000001" when "00101011001011011", -- t[22107] = 1
      "0000001" when "00101011001011100", -- t[22108] = 1
      "0000001" when "00101011001011101", -- t[22109] = 1
      "0000001" when "00101011001011110", -- t[22110] = 1
      "0000001" when "00101011001011111", -- t[22111] = 1
      "0000001" when "00101011001100000", -- t[22112] = 1
      "0000001" when "00101011001100001", -- t[22113] = 1
      "0000001" when "00101011001100010", -- t[22114] = 1
      "0000001" when "00101011001100011", -- t[22115] = 1
      "0000001" when "00101011001100100", -- t[22116] = 1
      "0000001" when "00101011001100101", -- t[22117] = 1
      "0000001" when "00101011001100110", -- t[22118] = 1
      "0000001" when "00101011001100111", -- t[22119] = 1
      "0000001" when "00101011001101000", -- t[22120] = 1
      "0000001" when "00101011001101001", -- t[22121] = 1
      "0000001" when "00101011001101010", -- t[22122] = 1
      "0000001" when "00101011001101011", -- t[22123] = 1
      "0000001" when "00101011001101100", -- t[22124] = 1
      "0000001" when "00101011001101101", -- t[22125] = 1
      "0000001" when "00101011001101110", -- t[22126] = 1
      "0000001" when "00101011001101111", -- t[22127] = 1
      "0000001" when "00101011001110000", -- t[22128] = 1
      "0000001" when "00101011001110001", -- t[22129] = 1
      "0000001" when "00101011001110010", -- t[22130] = 1
      "0000001" when "00101011001110011", -- t[22131] = 1
      "0000001" when "00101011001110100", -- t[22132] = 1
      "0000001" when "00101011001110101", -- t[22133] = 1
      "0000001" when "00101011001110110", -- t[22134] = 1
      "0000001" when "00101011001110111", -- t[22135] = 1
      "0000001" when "00101011001111000", -- t[22136] = 1
      "0000001" when "00101011001111001", -- t[22137] = 1
      "0000001" when "00101011001111010", -- t[22138] = 1
      "0000001" when "00101011001111011", -- t[22139] = 1
      "0000001" when "00101011001111100", -- t[22140] = 1
      "0000001" when "00101011001111101", -- t[22141] = 1
      "0000001" when "00101011001111110", -- t[22142] = 1
      "0000001" when "00101011001111111", -- t[22143] = 1
      "0000001" when "00101011010000000", -- t[22144] = 1
      "0000001" when "00101011010000001", -- t[22145] = 1
      "0000001" when "00101011010000010", -- t[22146] = 1
      "0000001" when "00101011010000011", -- t[22147] = 1
      "0000001" when "00101011010000100", -- t[22148] = 1
      "0000001" when "00101011010000101", -- t[22149] = 1
      "0000001" when "00101011010000110", -- t[22150] = 1
      "0000001" when "00101011010000111", -- t[22151] = 1
      "0000001" when "00101011010001000", -- t[22152] = 1
      "0000001" when "00101011010001001", -- t[22153] = 1
      "0000001" when "00101011010001010", -- t[22154] = 1
      "0000001" when "00101011010001011", -- t[22155] = 1
      "0000001" when "00101011010001100", -- t[22156] = 1
      "0000001" when "00101011010001101", -- t[22157] = 1
      "0000001" when "00101011010001110", -- t[22158] = 1
      "0000001" when "00101011010001111", -- t[22159] = 1
      "0000001" when "00101011010010000", -- t[22160] = 1
      "0000001" when "00101011010010001", -- t[22161] = 1
      "0000001" when "00101011010010010", -- t[22162] = 1
      "0000001" when "00101011010010011", -- t[22163] = 1
      "0000001" when "00101011010010100", -- t[22164] = 1
      "0000001" when "00101011010010101", -- t[22165] = 1
      "0000001" when "00101011010010110", -- t[22166] = 1
      "0000001" when "00101011010010111", -- t[22167] = 1
      "0000001" when "00101011010011000", -- t[22168] = 1
      "0000001" when "00101011010011001", -- t[22169] = 1
      "0000001" when "00101011010011010", -- t[22170] = 1
      "0000001" when "00101011010011011", -- t[22171] = 1
      "0000001" when "00101011010011100", -- t[22172] = 1
      "0000001" when "00101011010011101", -- t[22173] = 1
      "0000001" when "00101011010011110", -- t[22174] = 1
      "0000001" when "00101011010011111", -- t[22175] = 1
      "0000001" when "00101011010100000", -- t[22176] = 1
      "0000001" when "00101011010100001", -- t[22177] = 1
      "0000001" when "00101011010100010", -- t[22178] = 1
      "0000001" when "00101011010100011", -- t[22179] = 1
      "0000001" when "00101011010100100", -- t[22180] = 1
      "0000001" when "00101011010100101", -- t[22181] = 1
      "0000001" when "00101011010100110", -- t[22182] = 1
      "0000001" when "00101011010100111", -- t[22183] = 1
      "0000001" when "00101011010101000", -- t[22184] = 1
      "0000001" when "00101011010101001", -- t[22185] = 1
      "0000001" when "00101011010101010", -- t[22186] = 1
      "0000001" when "00101011010101011", -- t[22187] = 1
      "0000001" when "00101011010101100", -- t[22188] = 1
      "0000001" when "00101011010101101", -- t[22189] = 1
      "0000001" when "00101011010101110", -- t[22190] = 1
      "0000001" when "00101011010101111", -- t[22191] = 1
      "0000001" when "00101011010110000", -- t[22192] = 1
      "0000001" when "00101011010110001", -- t[22193] = 1
      "0000001" when "00101011010110010", -- t[22194] = 1
      "0000001" when "00101011010110011", -- t[22195] = 1
      "0000001" when "00101011010110100", -- t[22196] = 1
      "0000001" when "00101011010110101", -- t[22197] = 1
      "0000001" when "00101011010110110", -- t[22198] = 1
      "0000001" when "00101011010110111", -- t[22199] = 1
      "0000001" when "00101011010111000", -- t[22200] = 1
      "0000001" when "00101011010111001", -- t[22201] = 1
      "0000001" when "00101011010111010", -- t[22202] = 1
      "0000001" when "00101011010111011", -- t[22203] = 1
      "0000001" when "00101011010111100", -- t[22204] = 1
      "0000001" when "00101011010111101", -- t[22205] = 1
      "0000001" when "00101011010111110", -- t[22206] = 1
      "0000001" when "00101011010111111", -- t[22207] = 1
      "0000001" when "00101011011000000", -- t[22208] = 1
      "0000001" when "00101011011000001", -- t[22209] = 1
      "0000001" when "00101011011000010", -- t[22210] = 1
      "0000001" when "00101011011000011", -- t[22211] = 1
      "0000001" when "00101011011000100", -- t[22212] = 1
      "0000001" when "00101011011000101", -- t[22213] = 1
      "0000001" when "00101011011000110", -- t[22214] = 1
      "0000001" when "00101011011000111", -- t[22215] = 1
      "0000001" when "00101011011001000", -- t[22216] = 1
      "0000001" when "00101011011001001", -- t[22217] = 1
      "0000001" when "00101011011001010", -- t[22218] = 1
      "0000001" when "00101011011001011", -- t[22219] = 1
      "0000001" when "00101011011001100", -- t[22220] = 1
      "0000001" when "00101011011001101", -- t[22221] = 1
      "0000001" when "00101011011001110", -- t[22222] = 1
      "0000001" when "00101011011001111", -- t[22223] = 1
      "0000001" when "00101011011010000", -- t[22224] = 1
      "0000001" when "00101011011010001", -- t[22225] = 1
      "0000001" when "00101011011010010", -- t[22226] = 1
      "0000001" when "00101011011010011", -- t[22227] = 1
      "0000001" when "00101011011010100", -- t[22228] = 1
      "0000001" when "00101011011010101", -- t[22229] = 1
      "0000001" when "00101011011010110", -- t[22230] = 1
      "0000001" when "00101011011010111", -- t[22231] = 1
      "0000001" when "00101011011011000", -- t[22232] = 1
      "0000001" when "00101011011011001", -- t[22233] = 1
      "0000001" when "00101011011011010", -- t[22234] = 1
      "0000001" when "00101011011011011", -- t[22235] = 1
      "0000001" when "00101011011011100", -- t[22236] = 1
      "0000001" when "00101011011011101", -- t[22237] = 1
      "0000001" when "00101011011011110", -- t[22238] = 1
      "0000001" when "00101011011011111", -- t[22239] = 1
      "0000001" when "00101011011100000", -- t[22240] = 1
      "0000001" when "00101011011100001", -- t[22241] = 1
      "0000001" when "00101011011100010", -- t[22242] = 1
      "0000001" when "00101011011100011", -- t[22243] = 1
      "0000001" when "00101011011100100", -- t[22244] = 1
      "0000001" when "00101011011100101", -- t[22245] = 1
      "0000001" when "00101011011100110", -- t[22246] = 1
      "0000001" when "00101011011100111", -- t[22247] = 1
      "0000001" when "00101011011101000", -- t[22248] = 1
      "0000001" when "00101011011101001", -- t[22249] = 1
      "0000001" when "00101011011101010", -- t[22250] = 1
      "0000001" when "00101011011101011", -- t[22251] = 1
      "0000001" when "00101011011101100", -- t[22252] = 1
      "0000001" when "00101011011101101", -- t[22253] = 1
      "0000001" when "00101011011101110", -- t[22254] = 1
      "0000001" when "00101011011101111", -- t[22255] = 1
      "0000001" when "00101011011110000", -- t[22256] = 1
      "0000001" when "00101011011110001", -- t[22257] = 1
      "0000001" when "00101011011110010", -- t[22258] = 1
      "0000001" when "00101011011110011", -- t[22259] = 1
      "0000001" when "00101011011110100", -- t[22260] = 1
      "0000001" when "00101011011110101", -- t[22261] = 1
      "0000001" when "00101011011110110", -- t[22262] = 1
      "0000001" when "00101011011110111", -- t[22263] = 1
      "0000001" when "00101011011111000", -- t[22264] = 1
      "0000001" when "00101011011111001", -- t[22265] = 1
      "0000001" when "00101011011111010", -- t[22266] = 1
      "0000001" when "00101011011111011", -- t[22267] = 1
      "0000001" when "00101011011111100", -- t[22268] = 1
      "0000001" when "00101011011111101", -- t[22269] = 1
      "0000001" when "00101011011111110", -- t[22270] = 1
      "0000001" when "00101011011111111", -- t[22271] = 1
      "0000001" when "00101011100000000", -- t[22272] = 1
      "0000001" when "00101011100000001", -- t[22273] = 1
      "0000001" when "00101011100000010", -- t[22274] = 1
      "0000001" when "00101011100000011", -- t[22275] = 1
      "0000001" when "00101011100000100", -- t[22276] = 1
      "0000001" when "00101011100000101", -- t[22277] = 1
      "0000001" when "00101011100000110", -- t[22278] = 1
      "0000001" when "00101011100000111", -- t[22279] = 1
      "0000001" when "00101011100001000", -- t[22280] = 1
      "0000001" when "00101011100001001", -- t[22281] = 1
      "0000001" when "00101011100001010", -- t[22282] = 1
      "0000001" when "00101011100001011", -- t[22283] = 1
      "0000001" when "00101011100001100", -- t[22284] = 1
      "0000001" when "00101011100001101", -- t[22285] = 1
      "0000001" when "00101011100001110", -- t[22286] = 1
      "0000001" when "00101011100001111", -- t[22287] = 1
      "0000001" when "00101011100010000", -- t[22288] = 1
      "0000001" when "00101011100010001", -- t[22289] = 1
      "0000001" when "00101011100010010", -- t[22290] = 1
      "0000001" when "00101011100010011", -- t[22291] = 1
      "0000001" when "00101011100010100", -- t[22292] = 1
      "0000001" when "00101011100010101", -- t[22293] = 1
      "0000001" when "00101011100010110", -- t[22294] = 1
      "0000001" when "00101011100010111", -- t[22295] = 1
      "0000001" when "00101011100011000", -- t[22296] = 1
      "0000001" when "00101011100011001", -- t[22297] = 1
      "0000001" when "00101011100011010", -- t[22298] = 1
      "0000001" when "00101011100011011", -- t[22299] = 1
      "0000001" when "00101011100011100", -- t[22300] = 1
      "0000001" when "00101011100011101", -- t[22301] = 1
      "0000001" when "00101011100011110", -- t[22302] = 1
      "0000001" when "00101011100011111", -- t[22303] = 1
      "0000001" when "00101011100100000", -- t[22304] = 1
      "0000001" when "00101011100100001", -- t[22305] = 1
      "0000001" when "00101011100100010", -- t[22306] = 1
      "0000001" when "00101011100100011", -- t[22307] = 1
      "0000001" when "00101011100100100", -- t[22308] = 1
      "0000001" when "00101011100100101", -- t[22309] = 1
      "0000001" when "00101011100100110", -- t[22310] = 1
      "0000001" when "00101011100100111", -- t[22311] = 1
      "0000001" when "00101011100101000", -- t[22312] = 1
      "0000001" when "00101011100101001", -- t[22313] = 1
      "0000001" when "00101011100101010", -- t[22314] = 1
      "0000001" when "00101011100101011", -- t[22315] = 1
      "0000001" when "00101011100101100", -- t[22316] = 1
      "0000001" when "00101011100101101", -- t[22317] = 1
      "0000001" when "00101011100101110", -- t[22318] = 1
      "0000001" when "00101011100101111", -- t[22319] = 1
      "0000001" when "00101011100110000", -- t[22320] = 1
      "0000001" when "00101011100110001", -- t[22321] = 1
      "0000001" when "00101011100110010", -- t[22322] = 1
      "0000001" when "00101011100110011", -- t[22323] = 1
      "0000001" when "00101011100110100", -- t[22324] = 1
      "0000001" when "00101011100110101", -- t[22325] = 1
      "0000001" when "00101011100110110", -- t[22326] = 1
      "0000001" when "00101011100110111", -- t[22327] = 1
      "0000001" when "00101011100111000", -- t[22328] = 1
      "0000001" when "00101011100111001", -- t[22329] = 1
      "0000001" when "00101011100111010", -- t[22330] = 1
      "0000001" when "00101011100111011", -- t[22331] = 1
      "0000001" when "00101011100111100", -- t[22332] = 1
      "0000001" when "00101011100111101", -- t[22333] = 1
      "0000001" when "00101011100111110", -- t[22334] = 1
      "0000001" when "00101011100111111", -- t[22335] = 1
      "0000001" when "00101011101000000", -- t[22336] = 1
      "0000001" when "00101011101000001", -- t[22337] = 1
      "0000001" when "00101011101000010", -- t[22338] = 1
      "0000001" when "00101011101000011", -- t[22339] = 1
      "0000001" when "00101011101000100", -- t[22340] = 1
      "0000001" when "00101011101000101", -- t[22341] = 1
      "0000001" when "00101011101000110", -- t[22342] = 1
      "0000001" when "00101011101000111", -- t[22343] = 1
      "0000001" when "00101011101001000", -- t[22344] = 1
      "0000001" when "00101011101001001", -- t[22345] = 1
      "0000001" when "00101011101001010", -- t[22346] = 1
      "0000001" when "00101011101001011", -- t[22347] = 1
      "0000001" when "00101011101001100", -- t[22348] = 1
      "0000001" when "00101011101001101", -- t[22349] = 1
      "0000001" when "00101011101001110", -- t[22350] = 1
      "0000001" when "00101011101001111", -- t[22351] = 1
      "0000001" when "00101011101010000", -- t[22352] = 1
      "0000001" when "00101011101010001", -- t[22353] = 1
      "0000001" when "00101011101010010", -- t[22354] = 1
      "0000001" when "00101011101010011", -- t[22355] = 1
      "0000001" when "00101011101010100", -- t[22356] = 1
      "0000001" when "00101011101010101", -- t[22357] = 1
      "0000001" when "00101011101010110", -- t[22358] = 1
      "0000001" when "00101011101010111", -- t[22359] = 1
      "0000001" when "00101011101011000", -- t[22360] = 1
      "0000001" when "00101011101011001", -- t[22361] = 1
      "0000001" when "00101011101011010", -- t[22362] = 1
      "0000001" when "00101011101011011", -- t[22363] = 1
      "0000001" when "00101011101011100", -- t[22364] = 1
      "0000001" when "00101011101011101", -- t[22365] = 1
      "0000001" when "00101011101011110", -- t[22366] = 1
      "0000001" when "00101011101011111", -- t[22367] = 1
      "0000001" when "00101011101100000", -- t[22368] = 1
      "0000001" when "00101011101100001", -- t[22369] = 1
      "0000001" when "00101011101100010", -- t[22370] = 1
      "0000001" when "00101011101100011", -- t[22371] = 1
      "0000001" when "00101011101100100", -- t[22372] = 1
      "0000001" when "00101011101100101", -- t[22373] = 1
      "0000001" when "00101011101100110", -- t[22374] = 1
      "0000001" when "00101011101100111", -- t[22375] = 1
      "0000001" when "00101011101101000", -- t[22376] = 1
      "0000001" when "00101011101101001", -- t[22377] = 1
      "0000001" when "00101011101101010", -- t[22378] = 1
      "0000001" when "00101011101101011", -- t[22379] = 1
      "0000001" when "00101011101101100", -- t[22380] = 1
      "0000001" when "00101011101101101", -- t[22381] = 1
      "0000001" when "00101011101101110", -- t[22382] = 1
      "0000001" when "00101011101101111", -- t[22383] = 1
      "0000001" when "00101011101110000", -- t[22384] = 1
      "0000001" when "00101011101110001", -- t[22385] = 1
      "0000001" when "00101011101110010", -- t[22386] = 1
      "0000001" when "00101011101110011", -- t[22387] = 1
      "0000001" when "00101011101110100", -- t[22388] = 1
      "0000001" when "00101011101110101", -- t[22389] = 1
      "0000001" when "00101011101110110", -- t[22390] = 1
      "0000001" when "00101011101110111", -- t[22391] = 1
      "0000001" when "00101011101111000", -- t[22392] = 1
      "0000001" when "00101011101111001", -- t[22393] = 1
      "0000001" when "00101011101111010", -- t[22394] = 1
      "0000001" when "00101011101111011", -- t[22395] = 1
      "0000001" when "00101011101111100", -- t[22396] = 1
      "0000001" when "00101011101111101", -- t[22397] = 1
      "0000001" when "00101011101111110", -- t[22398] = 1
      "0000001" when "00101011101111111", -- t[22399] = 1
      "0000001" when "00101011110000000", -- t[22400] = 1
      "0000001" when "00101011110000001", -- t[22401] = 1
      "0000001" when "00101011110000010", -- t[22402] = 1
      "0000001" when "00101011110000011", -- t[22403] = 1
      "0000001" when "00101011110000100", -- t[22404] = 1
      "0000001" when "00101011110000101", -- t[22405] = 1
      "0000001" when "00101011110000110", -- t[22406] = 1
      "0000001" when "00101011110000111", -- t[22407] = 1
      "0000001" when "00101011110001000", -- t[22408] = 1
      "0000001" when "00101011110001001", -- t[22409] = 1
      "0000001" when "00101011110001010", -- t[22410] = 1
      "0000001" when "00101011110001011", -- t[22411] = 1
      "0000001" when "00101011110001100", -- t[22412] = 1
      "0000001" when "00101011110001101", -- t[22413] = 1
      "0000001" when "00101011110001110", -- t[22414] = 1
      "0000001" when "00101011110001111", -- t[22415] = 1
      "0000001" when "00101011110010000", -- t[22416] = 1
      "0000001" when "00101011110010001", -- t[22417] = 1
      "0000001" when "00101011110010010", -- t[22418] = 1
      "0000001" when "00101011110010011", -- t[22419] = 1
      "0000001" when "00101011110010100", -- t[22420] = 1
      "0000001" when "00101011110010101", -- t[22421] = 1
      "0000001" when "00101011110010110", -- t[22422] = 1
      "0000001" when "00101011110010111", -- t[22423] = 1
      "0000001" when "00101011110011000", -- t[22424] = 1
      "0000001" when "00101011110011001", -- t[22425] = 1
      "0000001" when "00101011110011010", -- t[22426] = 1
      "0000001" when "00101011110011011", -- t[22427] = 1
      "0000001" when "00101011110011100", -- t[22428] = 1
      "0000001" when "00101011110011101", -- t[22429] = 1
      "0000001" when "00101011110011110", -- t[22430] = 1
      "0000001" when "00101011110011111", -- t[22431] = 1
      "0000001" when "00101011110100000", -- t[22432] = 1
      "0000001" when "00101011110100001", -- t[22433] = 1
      "0000001" when "00101011110100010", -- t[22434] = 1
      "0000001" when "00101011110100011", -- t[22435] = 1
      "0000001" when "00101011110100100", -- t[22436] = 1
      "0000001" when "00101011110100101", -- t[22437] = 1
      "0000001" when "00101011110100110", -- t[22438] = 1
      "0000001" when "00101011110100111", -- t[22439] = 1
      "0000001" when "00101011110101000", -- t[22440] = 1
      "0000001" when "00101011110101001", -- t[22441] = 1
      "0000001" when "00101011110101010", -- t[22442] = 1
      "0000001" when "00101011110101011", -- t[22443] = 1
      "0000001" when "00101011110101100", -- t[22444] = 1
      "0000001" when "00101011110101101", -- t[22445] = 1
      "0000001" when "00101011110101110", -- t[22446] = 1
      "0000001" when "00101011110101111", -- t[22447] = 1
      "0000001" when "00101011110110000", -- t[22448] = 1
      "0000001" when "00101011110110001", -- t[22449] = 1
      "0000001" when "00101011110110010", -- t[22450] = 1
      "0000001" when "00101011110110011", -- t[22451] = 1
      "0000001" when "00101011110110100", -- t[22452] = 1
      "0000001" when "00101011110110101", -- t[22453] = 1
      "0000001" when "00101011110110110", -- t[22454] = 1
      "0000001" when "00101011110110111", -- t[22455] = 1
      "0000001" when "00101011110111000", -- t[22456] = 1
      "0000001" when "00101011110111001", -- t[22457] = 1
      "0000001" when "00101011110111010", -- t[22458] = 1
      "0000001" when "00101011110111011", -- t[22459] = 1
      "0000001" when "00101011110111100", -- t[22460] = 1
      "0000001" when "00101011110111101", -- t[22461] = 1
      "0000001" when "00101011110111110", -- t[22462] = 1
      "0000001" when "00101011110111111", -- t[22463] = 1
      "0000001" when "00101011111000000", -- t[22464] = 1
      "0000001" when "00101011111000001", -- t[22465] = 1
      "0000001" when "00101011111000010", -- t[22466] = 1
      "0000001" when "00101011111000011", -- t[22467] = 1
      "0000001" when "00101011111000100", -- t[22468] = 1
      "0000001" when "00101011111000101", -- t[22469] = 1
      "0000001" when "00101011111000110", -- t[22470] = 1
      "0000001" when "00101011111000111", -- t[22471] = 1
      "0000001" when "00101011111001000", -- t[22472] = 1
      "0000001" when "00101011111001001", -- t[22473] = 1
      "0000001" when "00101011111001010", -- t[22474] = 1
      "0000001" when "00101011111001011", -- t[22475] = 1
      "0000001" when "00101011111001100", -- t[22476] = 1
      "0000001" when "00101011111001101", -- t[22477] = 1
      "0000001" when "00101011111001110", -- t[22478] = 1
      "0000001" when "00101011111001111", -- t[22479] = 1
      "0000001" when "00101011111010000", -- t[22480] = 1
      "0000001" when "00101011111010001", -- t[22481] = 1
      "0000001" when "00101011111010010", -- t[22482] = 1
      "0000001" when "00101011111010011", -- t[22483] = 1
      "0000001" when "00101011111010100", -- t[22484] = 1
      "0000001" when "00101011111010101", -- t[22485] = 1
      "0000001" when "00101011111010110", -- t[22486] = 1
      "0000001" when "00101011111010111", -- t[22487] = 1
      "0000001" when "00101011111011000", -- t[22488] = 1
      "0000001" when "00101011111011001", -- t[22489] = 1
      "0000001" when "00101011111011010", -- t[22490] = 1
      "0000001" when "00101011111011011", -- t[22491] = 1
      "0000001" when "00101011111011100", -- t[22492] = 1
      "0000001" when "00101011111011101", -- t[22493] = 1
      "0000001" when "00101011111011110", -- t[22494] = 1
      "0000001" when "00101011111011111", -- t[22495] = 1
      "0000001" when "00101011111100000", -- t[22496] = 1
      "0000001" when "00101011111100001", -- t[22497] = 1
      "0000001" when "00101011111100010", -- t[22498] = 1
      "0000001" when "00101011111100011", -- t[22499] = 1
      "0000001" when "00101011111100100", -- t[22500] = 1
      "0000001" when "00101011111100101", -- t[22501] = 1
      "0000001" when "00101011111100110", -- t[22502] = 1
      "0000001" when "00101011111100111", -- t[22503] = 1
      "0000001" when "00101011111101000", -- t[22504] = 1
      "0000001" when "00101011111101001", -- t[22505] = 1
      "0000001" when "00101011111101010", -- t[22506] = 1
      "0000001" when "00101011111101011", -- t[22507] = 1
      "0000001" when "00101011111101100", -- t[22508] = 1
      "0000001" when "00101011111101101", -- t[22509] = 1
      "0000001" when "00101011111101110", -- t[22510] = 1
      "0000001" when "00101011111101111", -- t[22511] = 1
      "0000001" when "00101011111110000", -- t[22512] = 1
      "0000001" when "00101011111110001", -- t[22513] = 1
      "0000001" when "00101011111110010", -- t[22514] = 1
      "0000001" when "00101011111110011", -- t[22515] = 1
      "0000001" when "00101011111110100", -- t[22516] = 1
      "0000001" when "00101011111110101", -- t[22517] = 1
      "0000001" when "00101011111110110", -- t[22518] = 1
      "0000001" when "00101011111110111", -- t[22519] = 1
      "0000001" when "00101011111111000", -- t[22520] = 1
      "0000001" when "00101011111111001", -- t[22521] = 1
      "0000001" when "00101011111111010", -- t[22522] = 1
      "0000001" when "00101011111111011", -- t[22523] = 1
      "0000001" when "00101011111111100", -- t[22524] = 1
      "0000001" when "00101011111111101", -- t[22525] = 1
      "0000001" when "00101011111111110", -- t[22526] = 1
      "0000001" when "00101011111111111", -- t[22527] = 1
      "0000001" when "00101100000000000", -- t[22528] = 1
      "0000001" when "00101100000000001", -- t[22529] = 1
      "0000001" when "00101100000000010", -- t[22530] = 1
      "0000001" when "00101100000000011", -- t[22531] = 1
      "0000001" when "00101100000000100", -- t[22532] = 1
      "0000001" when "00101100000000101", -- t[22533] = 1
      "0000001" when "00101100000000110", -- t[22534] = 1
      "0000001" when "00101100000000111", -- t[22535] = 1
      "0000001" when "00101100000001000", -- t[22536] = 1
      "0000001" when "00101100000001001", -- t[22537] = 1
      "0000001" when "00101100000001010", -- t[22538] = 1
      "0000001" when "00101100000001011", -- t[22539] = 1
      "0000001" when "00101100000001100", -- t[22540] = 1
      "0000001" when "00101100000001101", -- t[22541] = 1
      "0000001" when "00101100000001110", -- t[22542] = 1
      "0000001" when "00101100000001111", -- t[22543] = 1
      "0000001" when "00101100000010000", -- t[22544] = 1
      "0000001" when "00101100000010001", -- t[22545] = 1
      "0000001" when "00101100000010010", -- t[22546] = 1
      "0000001" when "00101100000010011", -- t[22547] = 1
      "0000001" when "00101100000010100", -- t[22548] = 1
      "0000001" when "00101100000010101", -- t[22549] = 1
      "0000001" when "00101100000010110", -- t[22550] = 1
      "0000001" when "00101100000010111", -- t[22551] = 1
      "0000001" when "00101100000011000", -- t[22552] = 1
      "0000001" when "00101100000011001", -- t[22553] = 1
      "0000001" when "00101100000011010", -- t[22554] = 1
      "0000001" when "00101100000011011", -- t[22555] = 1
      "0000001" when "00101100000011100", -- t[22556] = 1
      "0000001" when "00101100000011101", -- t[22557] = 1
      "0000001" when "00101100000011110", -- t[22558] = 1
      "0000001" when "00101100000011111", -- t[22559] = 1
      "0000001" when "00101100000100000", -- t[22560] = 1
      "0000001" when "00101100000100001", -- t[22561] = 1
      "0000001" when "00101100000100010", -- t[22562] = 1
      "0000001" when "00101100000100011", -- t[22563] = 1
      "0000001" when "00101100000100100", -- t[22564] = 1
      "0000001" when "00101100000100101", -- t[22565] = 1
      "0000001" when "00101100000100110", -- t[22566] = 1
      "0000001" when "00101100000100111", -- t[22567] = 1
      "0000001" when "00101100000101000", -- t[22568] = 1
      "0000001" when "00101100000101001", -- t[22569] = 1
      "0000001" when "00101100000101010", -- t[22570] = 1
      "0000001" when "00101100000101011", -- t[22571] = 1
      "0000001" when "00101100000101100", -- t[22572] = 1
      "0000001" when "00101100000101101", -- t[22573] = 1
      "0000001" when "00101100000101110", -- t[22574] = 1
      "0000001" when "00101100000101111", -- t[22575] = 1
      "0000001" when "00101100000110000", -- t[22576] = 1
      "0000001" when "00101100000110001", -- t[22577] = 1
      "0000001" when "00101100000110010", -- t[22578] = 1
      "0000001" when "00101100000110011", -- t[22579] = 1
      "0000001" when "00101100000110100", -- t[22580] = 1
      "0000001" when "00101100000110101", -- t[22581] = 1
      "0000001" when "00101100000110110", -- t[22582] = 1
      "0000001" when "00101100000110111", -- t[22583] = 1
      "0000001" when "00101100000111000", -- t[22584] = 1
      "0000001" when "00101100000111001", -- t[22585] = 1
      "0000001" when "00101100000111010", -- t[22586] = 1
      "0000001" when "00101100000111011", -- t[22587] = 1
      "0000001" when "00101100000111100", -- t[22588] = 1
      "0000001" when "00101100000111101", -- t[22589] = 1
      "0000001" when "00101100000111110", -- t[22590] = 1
      "0000001" when "00101100000111111", -- t[22591] = 1
      "0000001" when "00101100001000000", -- t[22592] = 1
      "0000001" when "00101100001000001", -- t[22593] = 1
      "0000001" when "00101100001000010", -- t[22594] = 1
      "0000001" when "00101100001000011", -- t[22595] = 1
      "0000001" when "00101100001000100", -- t[22596] = 1
      "0000001" when "00101100001000101", -- t[22597] = 1
      "0000001" when "00101100001000110", -- t[22598] = 1
      "0000001" when "00101100001000111", -- t[22599] = 1
      "0000001" when "00101100001001000", -- t[22600] = 1
      "0000001" when "00101100001001001", -- t[22601] = 1
      "0000001" when "00101100001001010", -- t[22602] = 1
      "0000001" when "00101100001001011", -- t[22603] = 1
      "0000001" when "00101100001001100", -- t[22604] = 1
      "0000001" when "00101100001001101", -- t[22605] = 1
      "0000001" when "00101100001001110", -- t[22606] = 1
      "0000001" when "00101100001001111", -- t[22607] = 1
      "0000001" when "00101100001010000", -- t[22608] = 1
      "0000001" when "00101100001010001", -- t[22609] = 1
      "0000001" when "00101100001010010", -- t[22610] = 1
      "0000001" when "00101100001010011", -- t[22611] = 1
      "0000001" when "00101100001010100", -- t[22612] = 1
      "0000001" when "00101100001010101", -- t[22613] = 1
      "0000001" when "00101100001010110", -- t[22614] = 1
      "0000001" when "00101100001010111", -- t[22615] = 1
      "0000001" when "00101100001011000", -- t[22616] = 1
      "0000001" when "00101100001011001", -- t[22617] = 1
      "0000001" when "00101100001011010", -- t[22618] = 1
      "0000001" when "00101100001011011", -- t[22619] = 1
      "0000001" when "00101100001011100", -- t[22620] = 1
      "0000001" when "00101100001011101", -- t[22621] = 1
      "0000001" when "00101100001011110", -- t[22622] = 1
      "0000001" when "00101100001011111", -- t[22623] = 1
      "0000001" when "00101100001100000", -- t[22624] = 1
      "0000001" when "00101100001100001", -- t[22625] = 1
      "0000001" when "00101100001100010", -- t[22626] = 1
      "0000001" when "00101100001100011", -- t[22627] = 1
      "0000001" when "00101100001100100", -- t[22628] = 1
      "0000001" when "00101100001100101", -- t[22629] = 1
      "0000001" when "00101100001100110", -- t[22630] = 1
      "0000001" when "00101100001100111", -- t[22631] = 1
      "0000001" when "00101100001101000", -- t[22632] = 1
      "0000001" when "00101100001101001", -- t[22633] = 1
      "0000001" when "00101100001101010", -- t[22634] = 1
      "0000001" when "00101100001101011", -- t[22635] = 1
      "0000001" when "00101100001101100", -- t[22636] = 1
      "0000001" when "00101100001101101", -- t[22637] = 1
      "0000001" when "00101100001101110", -- t[22638] = 1
      "0000001" when "00101100001101111", -- t[22639] = 1
      "0000001" when "00101100001110000", -- t[22640] = 1
      "0000001" when "00101100001110001", -- t[22641] = 1
      "0000001" when "00101100001110010", -- t[22642] = 1
      "0000001" when "00101100001110011", -- t[22643] = 1
      "0000001" when "00101100001110100", -- t[22644] = 1
      "0000001" when "00101100001110101", -- t[22645] = 1
      "0000001" when "00101100001110110", -- t[22646] = 1
      "0000001" when "00101100001110111", -- t[22647] = 1
      "0000001" when "00101100001111000", -- t[22648] = 1
      "0000001" when "00101100001111001", -- t[22649] = 1
      "0000001" when "00101100001111010", -- t[22650] = 1
      "0000001" when "00101100001111011", -- t[22651] = 1
      "0000001" when "00101100001111100", -- t[22652] = 1
      "0000001" when "00101100001111101", -- t[22653] = 1
      "0000001" when "00101100001111110", -- t[22654] = 1
      "0000001" when "00101100001111111", -- t[22655] = 1
      "0000001" when "00101100010000000", -- t[22656] = 1
      "0000001" when "00101100010000001", -- t[22657] = 1
      "0000001" when "00101100010000010", -- t[22658] = 1
      "0000001" when "00101100010000011", -- t[22659] = 1
      "0000001" when "00101100010000100", -- t[22660] = 1
      "0000001" when "00101100010000101", -- t[22661] = 1
      "0000001" when "00101100010000110", -- t[22662] = 1
      "0000001" when "00101100010000111", -- t[22663] = 1
      "0000001" when "00101100010001000", -- t[22664] = 1
      "0000001" when "00101100010001001", -- t[22665] = 1
      "0000001" when "00101100010001010", -- t[22666] = 1
      "0000001" when "00101100010001011", -- t[22667] = 1
      "0000001" when "00101100010001100", -- t[22668] = 1
      "0000001" when "00101100010001101", -- t[22669] = 1
      "0000001" when "00101100010001110", -- t[22670] = 1
      "0000001" when "00101100010001111", -- t[22671] = 1
      "0000001" when "00101100010010000", -- t[22672] = 1
      "0000001" when "00101100010010001", -- t[22673] = 1
      "0000001" when "00101100010010010", -- t[22674] = 1
      "0000001" when "00101100010010011", -- t[22675] = 1
      "0000001" when "00101100010010100", -- t[22676] = 1
      "0000001" when "00101100010010101", -- t[22677] = 1
      "0000001" when "00101100010010110", -- t[22678] = 1
      "0000001" when "00101100010010111", -- t[22679] = 1
      "0000001" when "00101100010011000", -- t[22680] = 1
      "0000001" when "00101100010011001", -- t[22681] = 1
      "0000001" when "00101100010011010", -- t[22682] = 1
      "0000001" when "00101100010011011", -- t[22683] = 1
      "0000001" when "00101100010011100", -- t[22684] = 1
      "0000001" when "00101100010011101", -- t[22685] = 1
      "0000001" when "00101100010011110", -- t[22686] = 1
      "0000001" when "00101100010011111", -- t[22687] = 1
      "0000001" when "00101100010100000", -- t[22688] = 1
      "0000001" when "00101100010100001", -- t[22689] = 1
      "0000001" when "00101100010100010", -- t[22690] = 1
      "0000001" when "00101100010100011", -- t[22691] = 1
      "0000001" when "00101100010100100", -- t[22692] = 1
      "0000001" when "00101100010100101", -- t[22693] = 1
      "0000001" when "00101100010100110", -- t[22694] = 1
      "0000001" when "00101100010100111", -- t[22695] = 1
      "0000001" when "00101100010101000", -- t[22696] = 1
      "0000001" when "00101100010101001", -- t[22697] = 1
      "0000001" when "00101100010101010", -- t[22698] = 1
      "0000001" when "00101100010101011", -- t[22699] = 1
      "0000001" when "00101100010101100", -- t[22700] = 1
      "0000001" when "00101100010101101", -- t[22701] = 1
      "0000001" when "00101100010101110", -- t[22702] = 1
      "0000001" when "00101100010101111", -- t[22703] = 1
      "0000001" when "00101100010110000", -- t[22704] = 1
      "0000001" when "00101100010110001", -- t[22705] = 1
      "0000001" when "00101100010110010", -- t[22706] = 1
      "0000001" when "00101100010110011", -- t[22707] = 1
      "0000001" when "00101100010110100", -- t[22708] = 1
      "0000001" when "00101100010110101", -- t[22709] = 1
      "0000001" when "00101100010110110", -- t[22710] = 1
      "0000001" when "00101100010110111", -- t[22711] = 1
      "0000001" when "00101100010111000", -- t[22712] = 1
      "0000001" when "00101100010111001", -- t[22713] = 1
      "0000001" when "00101100010111010", -- t[22714] = 1
      "0000001" when "00101100010111011", -- t[22715] = 1
      "0000001" when "00101100010111100", -- t[22716] = 1
      "0000001" when "00101100010111101", -- t[22717] = 1
      "0000001" when "00101100010111110", -- t[22718] = 1
      "0000001" when "00101100010111111", -- t[22719] = 1
      "0000001" when "00101100011000000", -- t[22720] = 1
      "0000001" when "00101100011000001", -- t[22721] = 1
      "0000001" when "00101100011000010", -- t[22722] = 1
      "0000001" when "00101100011000011", -- t[22723] = 1
      "0000001" when "00101100011000100", -- t[22724] = 1
      "0000001" when "00101100011000101", -- t[22725] = 1
      "0000001" when "00101100011000110", -- t[22726] = 1
      "0000001" when "00101100011000111", -- t[22727] = 1
      "0000001" when "00101100011001000", -- t[22728] = 1
      "0000001" when "00101100011001001", -- t[22729] = 1
      "0000001" when "00101100011001010", -- t[22730] = 1
      "0000001" when "00101100011001011", -- t[22731] = 1
      "0000001" when "00101100011001100", -- t[22732] = 1
      "0000001" when "00101100011001101", -- t[22733] = 1
      "0000001" when "00101100011001110", -- t[22734] = 1
      "0000001" when "00101100011001111", -- t[22735] = 1
      "0000001" when "00101100011010000", -- t[22736] = 1
      "0000001" when "00101100011010001", -- t[22737] = 1
      "0000001" when "00101100011010010", -- t[22738] = 1
      "0000001" when "00101100011010011", -- t[22739] = 1
      "0000001" when "00101100011010100", -- t[22740] = 1
      "0000001" when "00101100011010101", -- t[22741] = 1
      "0000001" when "00101100011010110", -- t[22742] = 1
      "0000001" when "00101100011010111", -- t[22743] = 1
      "0000001" when "00101100011011000", -- t[22744] = 1
      "0000001" when "00101100011011001", -- t[22745] = 1
      "0000001" when "00101100011011010", -- t[22746] = 1
      "0000001" when "00101100011011011", -- t[22747] = 1
      "0000001" when "00101100011011100", -- t[22748] = 1
      "0000001" when "00101100011011101", -- t[22749] = 1
      "0000001" when "00101100011011110", -- t[22750] = 1
      "0000001" when "00101100011011111", -- t[22751] = 1
      "0000001" when "00101100011100000", -- t[22752] = 1
      "0000001" when "00101100011100001", -- t[22753] = 1
      "0000001" when "00101100011100010", -- t[22754] = 1
      "0000001" when "00101100011100011", -- t[22755] = 1
      "0000001" when "00101100011100100", -- t[22756] = 1
      "0000001" when "00101100011100101", -- t[22757] = 1
      "0000001" when "00101100011100110", -- t[22758] = 1
      "0000001" when "00101100011100111", -- t[22759] = 1
      "0000001" when "00101100011101000", -- t[22760] = 1
      "0000001" when "00101100011101001", -- t[22761] = 1
      "0000001" when "00101100011101010", -- t[22762] = 1
      "0000001" when "00101100011101011", -- t[22763] = 1
      "0000001" when "00101100011101100", -- t[22764] = 1
      "0000001" when "00101100011101101", -- t[22765] = 1
      "0000001" when "00101100011101110", -- t[22766] = 1
      "0000001" when "00101100011101111", -- t[22767] = 1
      "0000001" when "00101100011110000", -- t[22768] = 1
      "0000001" when "00101100011110001", -- t[22769] = 1
      "0000001" when "00101100011110010", -- t[22770] = 1
      "0000001" when "00101100011110011", -- t[22771] = 1
      "0000001" when "00101100011110100", -- t[22772] = 1
      "0000001" when "00101100011110101", -- t[22773] = 1
      "0000001" when "00101100011110110", -- t[22774] = 1
      "0000001" when "00101100011110111", -- t[22775] = 1
      "0000001" when "00101100011111000", -- t[22776] = 1
      "0000001" when "00101100011111001", -- t[22777] = 1
      "0000001" when "00101100011111010", -- t[22778] = 1
      "0000001" when "00101100011111011", -- t[22779] = 1
      "0000001" when "00101100011111100", -- t[22780] = 1
      "0000001" when "00101100011111101", -- t[22781] = 1
      "0000001" when "00101100011111110", -- t[22782] = 1
      "0000001" when "00101100011111111", -- t[22783] = 1
      "0000001" when "00101100100000000", -- t[22784] = 1
      "0000001" when "00101100100000001", -- t[22785] = 1
      "0000001" when "00101100100000010", -- t[22786] = 1
      "0000001" when "00101100100000011", -- t[22787] = 1
      "0000001" when "00101100100000100", -- t[22788] = 1
      "0000001" when "00101100100000101", -- t[22789] = 1
      "0000001" when "00101100100000110", -- t[22790] = 1
      "0000001" when "00101100100000111", -- t[22791] = 1
      "0000001" when "00101100100001000", -- t[22792] = 1
      "0000001" when "00101100100001001", -- t[22793] = 1
      "0000001" when "00101100100001010", -- t[22794] = 1
      "0000001" when "00101100100001011", -- t[22795] = 1
      "0000001" when "00101100100001100", -- t[22796] = 1
      "0000001" when "00101100100001101", -- t[22797] = 1
      "0000001" when "00101100100001110", -- t[22798] = 1
      "0000001" when "00101100100001111", -- t[22799] = 1
      "0000001" when "00101100100010000", -- t[22800] = 1
      "0000001" when "00101100100010001", -- t[22801] = 1
      "0000001" when "00101100100010010", -- t[22802] = 1
      "0000001" when "00101100100010011", -- t[22803] = 1
      "0000001" when "00101100100010100", -- t[22804] = 1
      "0000001" when "00101100100010101", -- t[22805] = 1
      "0000001" when "00101100100010110", -- t[22806] = 1
      "0000001" when "00101100100010111", -- t[22807] = 1
      "0000001" when "00101100100011000", -- t[22808] = 1
      "0000001" when "00101100100011001", -- t[22809] = 1
      "0000001" when "00101100100011010", -- t[22810] = 1
      "0000001" when "00101100100011011", -- t[22811] = 1
      "0000001" when "00101100100011100", -- t[22812] = 1
      "0000001" when "00101100100011101", -- t[22813] = 1
      "0000001" when "00101100100011110", -- t[22814] = 1
      "0000001" when "00101100100011111", -- t[22815] = 1
      "0000001" when "00101100100100000", -- t[22816] = 1
      "0000001" when "00101100100100001", -- t[22817] = 1
      "0000001" when "00101100100100010", -- t[22818] = 1
      "0000001" when "00101100100100011", -- t[22819] = 1
      "0000001" when "00101100100100100", -- t[22820] = 1
      "0000001" when "00101100100100101", -- t[22821] = 1
      "0000001" when "00101100100100110", -- t[22822] = 1
      "0000001" when "00101100100100111", -- t[22823] = 1
      "0000001" when "00101100100101000", -- t[22824] = 1
      "0000001" when "00101100100101001", -- t[22825] = 1
      "0000001" when "00101100100101010", -- t[22826] = 1
      "0000001" when "00101100100101011", -- t[22827] = 1
      "0000001" when "00101100100101100", -- t[22828] = 1
      "0000001" when "00101100100101101", -- t[22829] = 1
      "0000001" when "00101100100101110", -- t[22830] = 1
      "0000001" when "00101100100101111", -- t[22831] = 1
      "0000001" when "00101100100110000", -- t[22832] = 1
      "0000001" when "00101100100110001", -- t[22833] = 1
      "0000001" when "00101100100110010", -- t[22834] = 1
      "0000001" when "00101100100110011", -- t[22835] = 1
      "0000001" when "00101100100110100", -- t[22836] = 1
      "0000001" when "00101100100110101", -- t[22837] = 1
      "0000001" when "00101100100110110", -- t[22838] = 1
      "0000001" when "00101100100110111", -- t[22839] = 1
      "0000001" when "00101100100111000", -- t[22840] = 1
      "0000001" when "00101100100111001", -- t[22841] = 1
      "0000001" when "00101100100111010", -- t[22842] = 1
      "0000001" when "00101100100111011", -- t[22843] = 1
      "0000001" when "00101100100111100", -- t[22844] = 1
      "0000001" when "00101100100111101", -- t[22845] = 1
      "0000001" when "00101100100111110", -- t[22846] = 1
      "0000001" when "00101100100111111", -- t[22847] = 1
      "0000001" when "00101100101000000", -- t[22848] = 1
      "0000001" when "00101100101000001", -- t[22849] = 1
      "0000001" when "00101100101000010", -- t[22850] = 1
      "0000001" when "00101100101000011", -- t[22851] = 1
      "0000001" when "00101100101000100", -- t[22852] = 1
      "0000001" when "00101100101000101", -- t[22853] = 1
      "0000001" when "00101100101000110", -- t[22854] = 1
      "0000001" when "00101100101000111", -- t[22855] = 1
      "0000001" when "00101100101001000", -- t[22856] = 1
      "0000001" when "00101100101001001", -- t[22857] = 1
      "0000001" when "00101100101001010", -- t[22858] = 1
      "0000001" when "00101100101001011", -- t[22859] = 1
      "0000001" when "00101100101001100", -- t[22860] = 1
      "0000001" when "00101100101001101", -- t[22861] = 1
      "0000001" when "00101100101001110", -- t[22862] = 1
      "0000001" when "00101100101001111", -- t[22863] = 1
      "0000001" when "00101100101010000", -- t[22864] = 1
      "0000001" when "00101100101010001", -- t[22865] = 1
      "0000001" when "00101100101010010", -- t[22866] = 1
      "0000001" when "00101100101010011", -- t[22867] = 1
      "0000001" when "00101100101010100", -- t[22868] = 1
      "0000001" when "00101100101010101", -- t[22869] = 1
      "0000001" when "00101100101010110", -- t[22870] = 1
      "0000001" when "00101100101010111", -- t[22871] = 1
      "0000001" when "00101100101011000", -- t[22872] = 1
      "0000001" when "00101100101011001", -- t[22873] = 1
      "0000001" when "00101100101011010", -- t[22874] = 1
      "0000001" when "00101100101011011", -- t[22875] = 1
      "0000001" when "00101100101011100", -- t[22876] = 1
      "0000001" when "00101100101011101", -- t[22877] = 1
      "0000001" when "00101100101011110", -- t[22878] = 1
      "0000001" when "00101100101011111", -- t[22879] = 1
      "0000001" when "00101100101100000", -- t[22880] = 1
      "0000001" when "00101100101100001", -- t[22881] = 1
      "0000001" when "00101100101100010", -- t[22882] = 1
      "0000001" when "00101100101100011", -- t[22883] = 1
      "0000001" when "00101100101100100", -- t[22884] = 1
      "0000001" when "00101100101100101", -- t[22885] = 1
      "0000001" when "00101100101100110", -- t[22886] = 1
      "0000001" when "00101100101100111", -- t[22887] = 1
      "0000001" when "00101100101101000", -- t[22888] = 1
      "0000001" when "00101100101101001", -- t[22889] = 1
      "0000001" when "00101100101101010", -- t[22890] = 1
      "0000001" when "00101100101101011", -- t[22891] = 1
      "0000001" when "00101100101101100", -- t[22892] = 1
      "0000001" when "00101100101101101", -- t[22893] = 1
      "0000001" when "00101100101101110", -- t[22894] = 1
      "0000001" when "00101100101101111", -- t[22895] = 1
      "0000001" when "00101100101110000", -- t[22896] = 1
      "0000001" when "00101100101110001", -- t[22897] = 1
      "0000001" when "00101100101110010", -- t[22898] = 1
      "0000001" when "00101100101110011", -- t[22899] = 1
      "0000001" when "00101100101110100", -- t[22900] = 1
      "0000001" when "00101100101110101", -- t[22901] = 1
      "0000001" when "00101100101110110", -- t[22902] = 1
      "0000001" when "00101100101110111", -- t[22903] = 1
      "0000001" when "00101100101111000", -- t[22904] = 1
      "0000001" when "00101100101111001", -- t[22905] = 1
      "0000001" when "00101100101111010", -- t[22906] = 1
      "0000001" when "00101100101111011", -- t[22907] = 1
      "0000001" when "00101100101111100", -- t[22908] = 1
      "0000001" when "00101100101111101", -- t[22909] = 1
      "0000001" when "00101100101111110", -- t[22910] = 1
      "0000001" when "00101100101111111", -- t[22911] = 1
      "0000001" when "00101100110000000", -- t[22912] = 1
      "0000001" when "00101100110000001", -- t[22913] = 1
      "0000001" when "00101100110000010", -- t[22914] = 1
      "0000001" when "00101100110000011", -- t[22915] = 1
      "0000001" when "00101100110000100", -- t[22916] = 1
      "0000001" when "00101100110000101", -- t[22917] = 1
      "0000001" when "00101100110000110", -- t[22918] = 1
      "0000001" when "00101100110000111", -- t[22919] = 1
      "0000001" when "00101100110001000", -- t[22920] = 1
      "0000001" when "00101100110001001", -- t[22921] = 1
      "0000001" when "00101100110001010", -- t[22922] = 1
      "0000001" when "00101100110001011", -- t[22923] = 1
      "0000001" when "00101100110001100", -- t[22924] = 1
      "0000001" when "00101100110001101", -- t[22925] = 1
      "0000001" when "00101100110001110", -- t[22926] = 1
      "0000001" when "00101100110001111", -- t[22927] = 1
      "0000001" when "00101100110010000", -- t[22928] = 1
      "0000001" when "00101100110010001", -- t[22929] = 1
      "0000001" when "00101100110010010", -- t[22930] = 1
      "0000001" when "00101100110010011", -- t[22931] = 1
      "0000001" when "00101100110010100", -- t[22932] = 1
      "0000001" when "00101100110010101", -- t[22933] = 1
      "0000001" when "00101100110010110", -- t[22934] = 1
      "0000001" when "00101100110010111", -- t[22935] = 1
      "0000001" when "00101100110011000", -- t[22936] = 1
      "0000001" when "00101100110011001", -- t[22937] = 1
      "0000001" when "00101100110011010", -- t[22938] = 1
      "0000001" when "00101100110011011", -- t[22939] = 1
      "0000001" when "00101100110011100", -- t[22940] = 1
      "0000001" when "00101100110011101", -- t[22941] = 1
      "0000001" when "00101100110011110", -- t[22942] = 1
      "0000001" when "00101100110011111", -- t[22943] = 1
      "0000001" when "00101100110100000", -- t[22944] = 1
      "0000001" when "00101100110100001", -- t[22945] = 1
      "0000001" when "00101100110100010", -- t[22946] = 1
      "0000001" when "00101100110100011", -- t[22947] = 1
      "0000001" when "00101100110100100", -- t[22948] = 1
      "0000001" when "00101100110100101", -- t[22949] = 1
      "0000001" when "00101100110100110", -- t[22950] = 1
      "0000001" when "00101100110100111", -- t[22951] = 1
      "0000001" when "00101100110101000", -- t[22952] = 1
      "0000001" when "00101100110101001", -- t[22953] = 1
      "0000001" when "00101100110101010", -- t[22954] = 1
      "0000001" when "00101100110101011", -- t[22955] = 1
      "0000001" when "00101100110101100", -- t[22956] = 1
      "0000001" when "00101100110101101", -- t[22957] = 1
      "0000001" when "00101100110101110", -- t[22958] = 1
      "0000001" when "00101100110101111", -- t[22959] = 1
      "0000001" when "00101100110110000", -- t[22960] = 1
      "0000001" when "00101100110110001", -- t[22961] = 1
      "0000001" when "00101100110110010", -- t[22962] = 1
      "0000001" when "00101100110110011", -- t[22963] = 1
      "0000001" when "00101100110110100", -- t[22964] = 1
      "0000001" when "00101100110110101", -- t[22965] = 1
      "0000001" when "00101100110110110", -- t[22966] = 1
      "0000001" when "00101100110110111", -- t[22967] = 1
      "0000001" when "00101100110111000", -- t[22968] = 1
      "0000001" when "00101100110111001", -- t[22969] = 1
      "0000001" when "00101100110111010", -- t[22970] = 1
      "0000001" when "00101100110111011", -- t[22971] = 1
      "0000001" when "00101100110111100", -- t[22972] = 1
      "0000001" when "00101100110111101", -- t[22973] = 1
      "0000001" when "00101100110111110", -- t[22974] = 1
      "0000001" when "00101100110111111", -- t[22975] = 1
      "0000001" when "00101100111000000", -- t[22976] = 1
      "0000001" when "00101100111000001", -- t[22977] = 1
      "0000001" when "00101100111000010", -- t[22978] = 1
      "0000001" when "00101100111000011", -- t[22979] = 1
      "0000001" when "00101100111000100", -- t[22980] = 1
      "0000001" when "00101100111000101", -- t[22981] = 1
      "0000001" when "00101100111000110", -- t[22982] = 1
      "0000001" when "00101100111000111", -- t[22983] = 1
      "0000001" when "00101100111001000", -- t[22984] = 1
      "0000001" when "00101100111001001", -- t[22985] = 1
      "0000001" when "00101100111001010", -- t[22986] = 1
      "0000001" when "00101100111001011", -- t[22987] = 1
      "0000001" when "00101100111001100", -- t[22988] = 1
      "0000001" when "00101100111001101", -- t[22989] = 1
      "0000001" when "00101100111001110", -- t[22990] = 1
      "0000001" when "00101100111001111", -- t[22991] = 1
      "0000001" when "00101100111010000", -- t[22992] = 1
      "0000001" when "00101100111010001", -- t[22993] = 1
      "0000001" when "00101100111010010", -- t[22994] = 1
      "0000001" when "00101100111010011", -- t[22995] = 1
      "0000001" when "00101100111010100", -- t[22996] = 1
      "0000001" when "00101100111010101", -- t[22997] = 1
      "0000001" when "00101100111010110", -- t[22998] = 1
      "0000001" when "00101100111010111", -- t[22999] = 1
      "0000001" when "00101100111011000", -- t[23000] = 1
      "0000001" when "00101100111011001", -- t[23001] = 1
      "0000001" when "00101100111011010", -- t[23002] = 1
      "0000001" when "00101100111011011", -- t[23003] = 1
      "0000001" when "00101100111011100", -- t[23004] = 1
      "0000001" when "00101100111011101", -- t[23005] = 1
      "0000001" when "00101100111011110", -- t[23006] = 1
      "0000001" when "00101100111011111", -- t[23007] = 1
      "0000001" when "00101100111100000", -- t[23008] = 1
      "0000001" when "00101100111100001", -- t[23009] = 1
      "0000001" when "00101100111100010", -- t[23010] = 1
      "0000001" when "00101100111100011", -- t[23011] = 1
      "0000001" when "00101100111100100", -- t[23012] = 1
      "0000001" when "00101100111100101", -- t[23013] = 1
      "0000001" when "00101100111100110", -- t[23014] = 1
      "0000001" when "00101100111100111", -- t[23015] = 1
      "0000001" when "00101100111101000", -- t[23016] = 1
      "0000001" when "00101100111101001", -- t[23017] = 1
      "0000001" when "00101100111101010", -- t[23018] = 1
      "0000001" when "00101100111101011", -- t[23019] = 1
      "0000001" when "00101100111101100", -- t[23020] = 1
      "0000001" when "00101100111101101", -- t[23021] = 1
      "0000001" when "00101100111101110", -- t[23022] = 1
      "0000001" when "00101100111101111", -- t[23023] = 1
      "0000001" when "00101100111110000", -- t[23024] = 1
      "0000001" when "00101100111110001", -- t[23025] = 1
      "0000001" when "00101100111110010", -- t[23026] = 1
      "0000001" when "00101100111110011", -- t[23027] = 1
      "0000001" when "00101100111110100", -- t[23028] = 1
      "0000001" when "00101100111110101", -- t[23029] = 1
      "0000001" when "00101100111110110", -- t[23030] = 1
      "0000001" when "00101100111110111", -- t[23031] = 1
      "0000001" when "00101100111111000", -- t[23032] = 1
      "0000001" when "00101100111111001", -- t[23033] = 1
      "0000001" when "00101100111111010", -- t[23034] = 1
      "0000001" when "00101100111111011", -- t[23035] = 1
      "0000001" when "00101100111111100", -- t[23036] = 1
      "0000001" when "00101100111111101", -- t[23037] = 1
      "0000001" when "00101100111111110", -- t[23038] = 1
      "0000001" when "00101100111111111", -- t[23039] = 1
      "0000001" when "00101101000000000", -- t[23040] = 1
      "0000001" when "00101101000000001", -- t[23041] = 1
      "0000001" when "00101101000000010", -- t[23042] = 1
      "0000001" when "00101101000000011", -- t[23043] = 1
      "0000001" when "00101101000000100", -- t[23044] = 1
      "0000001" when "00101101000000101", -- t[23045] = 1
      "0000001" when "00101101000000110", -- t[23046] = 1
      "0000001" when "00101101000000111", -- t[23047] = 1
      "0000001" when "00101101000001000", -- t[23048] = 1
      "0000001" when "00101101000001001", -- t[23049] = 1
      "0000001" when "00101101000001010", -- t[23050] = 1
      "0000001" when "00101101000001011", -- t[23051] = 1
      "0000001" when "00101101000001100", -- t[23052] = 1
      "0000001" when "00101101000001101", -- t[23053] = 1
      "0000001" when "00101101000001110", -- t[23054] = 1
      "0000001" when "00101101000001111", -- t[23055] = 1
      "0000001" when "00101101000010000", -- t[23056] = 1
      "0000001" when "00101101000010001", -- t[23057] = 1
      "0000001" when "00101101000010010", -- t[23058] = 1
      "0000001" when "00101101000010011", -- t[23059] = 1
      "0000001" when "00101101000010100", -- t[23060] = 1
      "0000001" when "00101101000010101", -- t[23061] = 1
      "0000001" when "00101101000010110", -- t[23062] = 1
      "0000001" when "00101101000010111", -- t[23063] = 1
      "0000001" when "00101101000011000", -- t[23064] = 1
      "0000001" when "00101101000011001", -- t[23065] = 1
      "0000001" when "00101101000011010", -- t[23066] = 1
      "0000001" when "00101101000011011", -- t[23067] = 1
      "0000001" when "00101101000011100", -- t[23068] = 1
      "0000001" when "00101101000011101", -- t[23069] = 1
      "0000001" when "00101101000011110", -- t[23070] = 1
      "0000001" when "00101101000011111", -- t[23071] = 1
      "0000001" when "00101101000100000", -- t[23072] = 1
      "0000001" when "00101101000100001", -- t[23073] = 1
      "0000001" when "00101101000100010", -- t[23074] = 1
      "0000001" when "00101101000100011", -- t[23075] = 1
      "0000001" when "00101101000100100", -- t[23076] = 1
      "0000001" when "00101101000100101", -- t[23077] = 1
      "0000001" when "00101101000100110", -- t[23078] = 1
      "0000001" when "00101101000100111", -- t[23079] = 1
      "0000001" when "00101101000101000", -- t[23080] = 1
      "0000001" when "00101101000101001", -- t[23081] = 1
      "0000001" when "00101101000101010", -- t[23082] = 1
      "0000001" when "00101101000101011", -- t[23083] = 1
      "0000001" when "00101101000101100", -- t[23084] = 1
      "0000001" when "00101101000101101", -- t[23085] = 1
      "0000001" when "00101101000101110", -- t[23086] = 1
      "0000001" when "00101101000101111", -- t[23087] = 1
      "0000001" when "00101101000110000", -- t[23088] = 1
      "0000001" when "00101101000110001", -- t[23089] = 1
      "0000001" when "00101101000110010", -- t[23090] = 1
      "0000001" when "00101101000110011", -- t[23091] = 1
      "0000001" when "00101101000110100", -- t[23092] = 1
      "0000001" when "00101101000110101", -- t[23093] = 1
      "0000001" when "00101101000110110", -- t[23094] = 1
      "0000001" when "00101101000110111", -- t[23095] = 1
      "0000001" when "00101101000111000", -- t[23096] = 1
      "0000001" when "00101101000111001", -- t[23097] = 1
      "0000001" when "00101101000111010", -- t[23098] = 1
      "0000001" when "00101101000111011", -- t[23099] = 1
      "0000001" when "00101101000111100", -- t[23100] = 1
      "0000001" when "00101101000111101", -- t[23101] = 1
      "0000001" when "00101101000111110", -- t[23102] = 1
      "0000001" when "00101101000111111", -- t[23103] = 1
      "0000001" when "00101101001000000", -- t[23104] = 1
      "0000001" when "00101101001000001", -- t[23105] = 1
      "0000001" when "00101101001000010", -- t[23106] = 1
      "0000001" when "00101101001000011", -- t[23107] = 1
      "0000001" when "00101101001000100", -- t[23108] = 1
      "0000001" when "00101101001000101", -- t[23109] = 1
      "0000001" when "00101101001000110", -- t[23110] = 1
      "0000001" when "00101101001000111", -- t[23111] = 1
      "0000001" when "00101101001001000", -- t[23112] = 1
      "0000001" when "00101101001001001", -- t[23113] = 1
      "0000001" when "00101101001001010", -- t[23114] = 1
      "0000001" when "00101101001001011", -- t[23115] = 1
      "0000001" when "00101101001001100", -- t[23116] = 1
      "0000001" when "00101101001001101", -- t[23117] = 1
      "0000001" when "00101101001001110", -- t[23118] = 1
      "0000001" when "00101101001001111", -- t[23119] = 1
      "0000001" when "00101101001010000", -- t[23120] = 1
      "0000001" when "00101101001010001", -- t[23121] = 1
      "0000001" when "00101101001010010", -- t[23122] = 1
      "0000001" when "00101101001010011", -- t[23123] = 1
      "0000001" when "00101101001010100", -- t[23124] = 1
      "0000001" when "00101101001010101", -- t[23125] = 1
      "0000001" when "00101101001010110", -- t[23126] = 1
      "0000001" when "00101101001010111", -- t[23127] = 1
      "0000001" when "00101101001011000", -- t[23128] = 1
      "0000001" when "00101101001011001", -- t[23129] = 1
      "0000001" when "00101101001011010", -- t[23130] = 1
      "0000001" when "00101101001011011", -- t[23131] = 1
      "0000001" when "00101101001011100", -- t[23132] = 1
      "0000001" when "00101101001011101", -- t[23133] = 1
      "0000001" when "00101101001011110", -- t[23134] = 1
      "0000001" when "00101101001011111", -- t[23135] = 1
      "0000001" when "00101101001100000", -- t[23136] = 1
      "0000001" when "00101101001100001", -- t[23137] = 1
      "0000001" when "00101101001100010", -- t[23138] = 1
      "0000001" when "00101101001100011", -- t[23139] = 1
      "0000001" when "00101101001100100", -- t[23140] = 1
      "0000001" when "00101101001100101", -- t[23141] = 1
      "0000001" when "00101101001100110", -- t[23142] = 1
      "0000001" when "00101101001100111", -- t[23143] = 1
      "0000001" when "00101101001101000", -- t[23144] = 1
      "0000001" when "00101101001101001", -- t[23145] = 1
      "0000001" when "00101101001101010", -- t[23146] = 1
      "0000001" when "00101101001101011", -- t[23147] = 1
      "0000001" when "00101101001101100", -- t[23148] = 1
      "0000001" when "00101101001101101", -- t[23149] = 1
      "0000001" when "00101101001101110", -- t[23150] = 1
      "0000001" when "00101101001101111", -- t[23151] = 1
      "0000001" when "00101101001110000", -- t[23152] = 1
      "0000001" when "00101101001110001", -- t[23153] = 1
      "0000001" when "00101101001110010", -- t[23154] = 1
      "0000001" when "00101101001110011", -- t[23155] = 1
      "0000001" when "00101101001110100", -- t[23156] = 1
      "0000001" when "00101101001110101", -- t[23157] = 1
      "0000001" when "00101101001110110", -- t[23158] = 1
      "0000001" when "00101101001110111", -- t[23159] = 1
      "0000001" when "00101101001111000", -- t[23160] = 1
      "0000001" when "00101101001111001", -- t[23161] = 1
      "0000001" when "00101101001111010", -- t[23162] = 1
      "0000001" when "00101101001111011", -- t[23163] = 1
      "0000001" when "00101101001111100", -- t[23164] = 1
      "0000001" when "00101101001111101", -- t[23165] = 1
      "0000001" when "00101101001111110", -- t[23166] = 1
      "0000001" when "00101101001111111", -- t[23167] = 1
      "0000001" when "00101101010000000", -- t[23168] = 1
      "0000001" when "00101101010000001", -- t[23169] = 1
      "0000001" when "00101101010000010", -- t[23170] = 1
      "0000001" when "00101101010000011", -- t[23171] = 1
      "0000001" when "00101101010000100", -- t[23172] = 1
      "0000001" when "00101101010000101", -- t[23173] = 1
      "0000001" when "00101101010000110", -- t[23174] = 1
      "0000001" when "00101101010000111", -- t[23175] = 1
      "0000001" when "00101101010001000", -- t[23176] = 1
      "0000001" when "00101101010001001", -- t[23177] = 1
      "0000001" when "00101101010001010", -- t[23178] = 1
      "0000001" when "00101101010001011", -- t[23179] = 1
      "0000001" when "00101101010001100", -- t[23180] = 1
      "0000001" when "00101101010001101", -- t[23181] = 1
      "0000001" when "00101101010001110", -- t[23182] = 1
      "0000001" when "00101101010001111", -- t[23183] = 1
      "0000001" when "00101101010010000", -- t[23184] = 1
      "0000001" when "00101101010010001", -- t[23185] = 1
      "0000001" when "00101101010010010", -- t[23186] = 1
      "0000001" when "00101101010010011", -- t[23187] = 1
      "0000001" when "00101101010010100", -- t[23188] = 1
      "0000001" when "00101101010010101", -- t[23189] = 1
      "0000001" when "00101101010010110", -- t[23190] = 1
      "0000001" when "00101101010010111", -- t[23191] = 1
      "0000001" when "00101101010011000", -- t[23192] = 1
      "0000001" when "00101101010011001", -- t[23193] = 1
      "0000001" when "00101101010011010", -- t[23194] = 1
      "0000001" when "00101101010011011", -- t[23195] = 1
      "0000001" when "00101101010011100", -- t[23196] = 1
      "0000001" when "00101101010011101", -- t[23197] = 1
      "0000001" when "00101101010011110", -- t[23198] = 1
      "0000001" when "00101101010011111", -- t[23199] = 1
      "0000001" when "00101101010100000", -- t[23200] = 1
      "0000001" when "00101101010100001", -- t[23201] = 1
      "0000001" when "00101101010100010", -- t[23202] = 1
      "0000001" when "00101101010100011", -- t[23203] = 1
      "0000001" when "00101101010100100", -- t[23204] = 1
      "0000001" when "00101101010100101", -- t[23205] = 1
      "0000001" when "00101101010100110", -- t[23206] = 1
      "0000001" when "00101101010100111", -- t[23207] = 1
      "0000001" when "00101101010101000", -- t[23208] = 1
      "0000001" when "00101101010101001", -- t[23209] = 1
      "0000001" when "00101101010101010", -- t[23210] = 1
      "0000001" when "00101101010101011", -- t[23211] = 1
      "0000001" when "00101101010101100", -- t[23212] = 1
      "0000001" when "00101101010101101", -- t[23213] = 1
      "0000001" when "00101101010101110", -- t[23214] = 1
      "0000001" when "00101101010101111", -- t[23215] = 1
      "0000001" when "00101101010110000", -- t[23216] = 1
      "0000001" when "00101101010110001", -- t[23217] = 1
      "0000001" when "00101101010110010", -- t[23218] = 1
      "0000001" when "00101101010110011", -- t[23219] = 1
      "0000001" when "00101101010110100", -- t[23220] = 1
      "0000001" when "00101101010110101", -- t[23221] = 1
      "0000001" when "00101101010110110", -- t[23222] = 1
      "0000001" when "00101101010110111", -- t[23223] = 1
      "0000001" when "00101101010111000", -- t[23224] = 1
      "0000001" when "00101101010111001", -- t[23225] = 1
      "0000001" when "00101101010111010", -- t[23226] = 1
      "0000001" when "00101101010111011", -- t[23227] = 1
      "0000001" when "00101101010111100", -- t[23228] = 1
      "0000001" when "00101101010111101", -- t[23229] = 1
      "0000001" when "00101101010111110", -- t[23230] = 1
      "0000001" when "00101101010111111", -- t[23231] = 1
      "0000001" when "00101101011000000", -- t[23232] = 1
      "0000001" when "00101101011000001", -- t[23233] = 1
      "0000001" when "00101101011000010", -- t[23234] = 1
      "0000001" when "00101101011000011", -- t[23235] = 1
      "0000001" when "00101101011000100", -- t[23236] = 1
      "0000001" when "00101101011000101", -- t[23237] = 1
      "0000001" when "00101101011000110", -- t[23238] = 1
      "0000001" when "00101101011000111", -- t[23239] = 1
      "0000001" when "00101101011001000", -- t[23240] = 1
      "0000001" when "00101101011001001", -- t[23241] = 1
      "0000001" when "00101101011001010", -- t[23242] = 1
      "0000001" when "00101101011001011", -- t[23243] = 1
      "0000001" when "00101101011001100", -- t[23244] = 1
      "0000001" when "00101101011001101", -- t[23245] = 1
      "0000001" when "00101101011001110", -- t[23246] = 1
      "0000001" when "00101101011001111", -- t[23247] = 1
      "0000001" when "00101101011010000", -- t[23248] = 1
      "0000001" when "00101101011010001", -- t[23249] = 1
      "0000001" when "00101101011010010", -- t[23250] = 1
      "0000001" when "00101101011010011", -- t[23251] = 1
      "0000001" when "00101101011010100", -- t[23252] = 1
      "0000001" when "00101101011010101", -- t[23253] = 1
      "0000001" when "00101101011010110", -- t[23254] = 1
      "0000001" when "00101101011010111", -- t[23255] = 1
      "0000001" when "00101101011011000", -- t[23256] = 1
      "0000001" when "00101101011011001", -- t[23257] = 1
      "0000001" when "00101101011011010", -- t[23258] = 1
      "0000001" when "00101101011011011", -- t[23259] = 1
      "0000001" when "00101101011011100", -- t[23260] = 1
      "0000001" when "00101101011011101", -- t[23261] = 1
      "0000001" when "00101101011011110", -- t[23262] = 1
      "0000001" when "00101101011011111", -- t[23263] = 1
      "0000001" when "00101101011100000", -- t[23264] = 1
      "0000001" when "00101101011100001", -- t[23265] = 1
      "0000001" when "00101101011100010", -- t[23266] = 1
      "0000001" when "00101101011100011", -- t[23267] = 1
      "0000001" when "00101101011100100", -- t[23268] = 1
      "0000001" when "00101101011100101", -- t[23269] = 1
      "0000001" when "00101101011100110", -- t[23270] = 1
      "0000001" when "00101101011100111", -- t[23271] = 1
      "0000001" when "00101101011101000", -- t[23272] = 1
      "0000001" when "00101101011101001", -- t[23273] = 1
      "0000001" when "00101101011101010", -- t[23274] = 1
      "0000001" when "00101101011101011", -- t[23275] = 1
      "0000001" when "00101101011101100", -- t[23276] = 1
      "0000001" when "00101101011101101", -- t[23277] = 1
      "0000001" when "00101101011101110", -- t[23278] = 1
      "0000001" when "00101101011101111", -- t[23279] = 1
      "0000001" when "00101101011110000", -- t[23280] = 1
      "0000001" when "00101101011110001", -- t[23281] = 1
      "0000001" when "00101101011110010", -- t[23282] = 1
      "0000001" when "00101101011110011", -- t[23283] = 1
      "0000001" when "00101101011110100", -- t[23284] = 1
      "0000001" when "00101101011110101", -- t[23285] = 1
      "0000001" when "00101101011110110", -- t[23286] = 1
      "0000001" when "00101101011110111", -- t[23287] = 1
      "0000001" when "00101101011111000", -- t[23288] = 1
      "0000001" when "00101101011111001", -- t[23289] = 1
      "0000001" when "00101101011111010", -- t[23290] = 1
      "0000001" when "00101101011111011", -- t[23291] = 1
      "0000001" when "00101101011111100", -- t[23292] = 1
      "0000001" when "00101101011111101", -- t[23293] = 1
      "0000001" when "00101101011111110", -- t[23294] = 1
      "0000001" when "00101101011111111", -- t[23295] = 1
      "0000001" when "00101101100000000", -- t[23296] = 1
      "0000001" when "00101101100000001", -- t[23297] = 1
      "0000001" when "00101101100000010", -- t[23298] = 1
      "0000001" when "00101101100000011", -- t[23299] = 1
      "0000001" when "00101101100000100", -- t[23300] = 1
      "0000001" when "00101101100000101", -- t[23301] = 1
      "0000001" when "00101101100000110", -- t[23302] = 1
      "0000001" when "00101101100000111", -- t[23303] = 1
      "0000001" when "00101101100001000", -- t[23304] = 1
      "0000001" when "00101101100001001", -- t[23305] = 1
      "0000001" when "00101101100001010", -- t[23306] = 1
      "0000001" when "00101101100001011", -- t[23307] = 1
      "0000001" when "00101101100001100", -- t[23308] = 1
      "0000001" when "00101101100001101", -- t[23309] = 1
      "0000001" when "00101101100001110", -- t[23310] = 1
      "0000001" when "00101101100001111", -- t[23311] = 1
      "0000001" when "00101101100010000", -- t[23312] = 1
      "0000001" when "00101101100010001", -- t[23313] = 1
      "0000001" when "00101101100010010", -- t[23314] = 1
      "0000001" when "00101101100010011", -- t[23315] = 1
      "0000001" when "00101101100010100", -- t[23316] = 1
      "0000001" when "00101101100010101", -- t[23317] = 1
      "0000001" when "00101101100010110", -- t[23318] = 1
      "0000001" when "00101101100010111", -- t[23319] = 1
      "0000001" when "00101101100011000", -- t[23320] = 1
      "0000001" when "00101101100011001", -- t[23321] = 1
      "0000001" when "00101101100011010", -- t[23322] = 1
      "0000001" when "00101101100011011", -- t[23323] = 1
      "0000001" when "00101101100011100", -- t[23324] = 1
      "0000001" when "00101101100011101", -- t[23325] = 1
      "0000001" when "00101101100011110", -- t[23326] = 1
      "0000001" when "00101101100011111", -- t[23327] = 1
      "0000001" when "00101101100100000", -- t[23328] = 1
      "0000001" when "00101101100100001", -- t[23329] = 1
      "0000001" when "00101101100100010", -- t[23330] = 1
      "0000001" when "00101101100100011", -- t[23331] = 1
      "0000001" when "00101101100100100", -- t[23332] = 1
      "0000001" when "00101101100100101", -- t[23333] = 1
      "0000001" when "00101101100100110", -- t[23334] = 1
      "0000001" when "00101101100100111", -- t[23335] = 1
      "0000001" when "00101101100101000", -- t[23336] = 1
      "0000001" when "00101101100101001", -- t[23337] = 1
      "0000001" when "00101101100101010", -- t[23338] = 1
      "0000001" when "00101101100101011", -- t[23339] = 1
      "0000001" when "00101101100101100", -- t[23340] = 1
      "0000001" when "00101101100101101", -- t[23341] = 1
      "0000001" when "00101101100101110", -- t[23342] = 1
      "0000001" when "00101101100101111", -- t[23343] = 1
      "0000001" when "00101101100110000", -- t[23344] = 1
      "0000001" when "00101101100110001", -- t[23345] = 1
      "0000001" when "00101101100110010", -- t[23346] = 1
      "0000001" when "00101101100110011", -- t[23347] = 1
      "0000001" when "00101101100110100", -- t[23348] = 1
      "0000001" when "00101101100110101", -- t[23349] = 1
      "0000001" when "00101101100110110", -- t[23350] = 1
      "0000001" when "00101101100110111", -- t[23351] = 1
      "0000001" when "00101101100111000", -- t[23352] = 1
      "0000001" when "00101101100111001", -- t[23353] = 1
      "0000001" when "00101101100111010", -- t[23354] = 1
      "0000001" when "00101101100111011", -- t[23355] = 1
      "0000001" when "00101101100111100", -- t[23356] = 1
      "0000001" when "00101101100111101", -- t[23357] = 1
      "0000001" when "00101101100111110", -- t[23358] = 1
      "0000001" when "00101101100111111", -- t[23359] = 1
      "0000001" when "00101101101000000", -- t[23360] = 1
      "0000001" when "00101101101000001", -- t[23361] = 1
      "0000001" when "00101101101000010", -- t[23362] = 1
      "0000001" when "00101101101000011", -- t[23363] = 1
      "0000001" when "00101101101000100", -- t[23364] = 1
      "0000001" when "00101101101000101", -- t[23365] = 1
      "0000001" when "00101101101000110", -- t[23366] = 1
      "0000001" when "00101101101000111", -- t[23367] = 1
      "0000001" when "00101101101001000", -- t[23368] = 1
      "0000001" when "00101101101001001", -- t[23369] = 1
      "0000001" when "00101101101001010", -- t[23370] = 1
      "0000001" when "00101101101001011", -- t[23371] = 1
      "0000001" when "00101101101001100", -- t[23372] = 1
      "0000001" when "00101101101001101", -- t[23373] = 1
      "0000001" when "00101101101001110", -- t[23374] = 1
      "0000001" when "00101101101001111", -- t[23375] = 1
      "0000001" when "00101101101010000", -- t[23376] = 1
      "0000001" when "00101101101010001", -- t[23377] = 1
      "0000001" when "00101101101010010", -- t[23378] = 1
      "0000001" when "00101101101010011", -- t[23379] = 1
      "0000001" when "00101101101010100", -- t[23380] = 1
      "0000001" when "00101101101010101", -- t[23381] = 1
      "0000001" when "00101101101010110", -- t[23382] = 1
      "0000001" when "00101101101010111", -- t[23383] = 1
      "0000001" when "00101101101011000", -- t[23384] = 1
      "0000001" when "00101101101011001", -- t[23385] = 1
      "0000001" when "00101101101011010", -- t[23386] = 1
      "0000001" when "00101101101011011", -- t[23387] = 1
      "0000001" when "00101101101011100", -- t[23388] = 1
      "0000001" when "00101101101011101", -- t[23389] = 1
      "0000001" when "00101101101011110", -- t[23390] = 1
      "0000001" when "00101101101011111", -- t[23391] = 1
      "0000001" when "00101101101100000", -- t[23392] = 1
      "0000001" when "00101101101100001", -- t[23393] = 1
      "0000001" when "00101101101100010", -- t[23394] = 1
      "0000001" when "00101101101100011", -- t[23395] = 1
      "0000001" when "00101101101100100", -- t[23396] = 1
      "0000001" when "00101101101100101", -- t[23397] = 1
      "0000001" when "00101101101100110", -- t[23398] = 1
      "0000001" when "00101101101100111", -- t[23399] = 1
      "0000001" when "00101101101101000", -- t[23400] = 1
      "0000001" when "00101101101101001", -- t[23401] = 1
      "0000001" when "00101101101101010", -- t[23402] = 1
      "0000001" when "00101101101101011", -- t[23403] = 1
      "0000001" when "00101101101101100", -- t[23404] = 1
      "0000001" when "00101101101101101", -- t[23405] = 1
      "0000001" when "00101101101101110", -- t[23406] = 1
      "0000001" when "00101101101101111", -- t[23407] = 1
      "0000001" when "00101101101110000", -- t[23408] = 1
      "0000001" when "00101101101110001", -- t[23409] = 1
      "0000001" when "00101101101110010", -- t[23410] = 1
      "0000001" when "00101101101110011", -- t[23411] = 1
      "0000001" when "00101101101110100", -- t[23412] = 1
      "0000001" when "00101101101110101", -- t[23413] = 1
      "0000001" when "00101101101110110", -- t[23414] = 1
      "0000001" when "00101101101110111", -- t[23415] = 1
      "0000001" when "00101101101111000", -- t[23416] = 1
      "0000001" when "00101101101111001", -- t[23417] = 1
      "0000001" when "00101101101111010", -- t[23418] = 1
      "0000001" when "00101101101111011", -- t[23419] = 1
      "0000001" when "00101101101111100", -- t[23420] = 1
      "0000001" when "00101101101111101", -- t[23421] = 1
      "0000001" when "00101101101111110", -- t[23422] = 1
      "0000001" when "00101101101111111", -- t[23423] = 1
      "0000001" when "00101101110000000", -- t[23424] = 1
      "0000001" when "00101101110000001", -- t[23425] = 1
      "0000001" when "00101101110000010", -- t[23426] = 1
      "0000001" when "00101101110000011", -- t[23427] = 1
      "0000001" when "00101101110000100", -- t[23428] = 1
      "0000001" when "00101101110000101", -- t[23429] = 1
      "0000001" when "00101101110000110", -- t[23430] = 1
      "0000001" when "00101101110000111", -- t[23431] = 1
      "0000001" when "00101101110001000", -- t[23432] = 1
      "0000001" when "00101101110001001", -- t[23433] = 1
      "0000001" when "00101101110001010", -- t[23434] = 1
      "0000001" when "00101101110001011", -- t[23435] = 1
      "0000001" when "00101101110001100", -- t[23436] = 1
      "0000001" when "00101101110001101", -- t[23437] = 1
      "0000001" when "00101101110001110", -- t[23438] = 1
      "0000001" when "00101101110001111", -- t[23439] = 1
      "0000001" when "00101101110010000", -- t[23440] = 1
      "0000001" when "00101101110010001", -- t[23441] = 1
      "0000001" when "00101101110010010", -- t[23442] = 1
      "0000001" when "00101101110010011", -- t[23443] = 1
      "0000001" when "00101101110010100", -- t[23444] = 1
      "0000001" when "00101101110010101", -- t[23445] = 1
      "0000001" when "00101101110010110", -- t[23446] = 1
      "0000001" when "00101101110010111", -- t[23447] = 1
      "0000001" when "00101101110011000", -- t[23448] = 1
      "0000001" when "00101101110011001", -- t[23449] = 1
      "0000001" when "00101101110011010", -- t[23450] = 1
      "0000001" when "00101101110011011", -- t[23451] = 1
      "0000001" when "00101101110011100", -- t[23452] = 1
      "0000001" when "00101101110011101", -- t[23453] = 1
      "0000001" when "00101101110011110", -- t[23454] = 1
      "0000001" when "00101101110011111", -- t[23455] = 1
      "0000001" when "00101101110100000", -- t[23456] = 1
      "0000001" when "00101101110100001", -- t[23457] = 1
      "0000001" when "00101101110100010", -- t[23458] = 1
      "0000001" when "00101101110100011", -- t[23459] = 1
      "0000001" when "00101101110100100", -- t[23460] = 1
      "0000001" when "00101101110100101", -- t[23461] = 1
      "0000001" when "00101101110100110", -- t[23462] = 1
      "0000001" when "00101101110100111", -- t[23463] = 1
      "0000001" when "00101101110101000", -- t[23464] = 1
      "0000001" when "00101101110101001", -- t[23465] = 1
      "0000001" when "00101101110101010", -- t[23466] = 1
      "0000001" when "00101101110101011", -- t[23467] = 1
      "0000001" when "00101101110101100", -- t[23468] = 1
      "0000001" when "00101101110101101", -- t[23469] = 1
      "0000001" when "00101101110101110", -- t[23470] = 1
      "0000001" when "00101101110101111", -- t[23471] = 1
      "0000001" when "00101101110110000", -- t[23472] = 1
      "0000001" when "00101101110110001", -- t[23473] = 1
      "0000001" when "00101101110110010", -- t[23474] = 1
      "0000001" when "00101101110110011", -- t[23475] = 1
      "0000001" when "00101101110110100", -- t[23476] = 1
      "0000001" when "00101101110110101", -- t[23477] = 1
      "0000001" when "00101101110110110", -- t[23478] = 1
      "0000001" when "00101101110110111", -- t[23479] = 1
      "0000001" when "00101101110111000", -- t[23480] = 1
      "0000001" when "00101101110111001", -- t[23481] = 1
      "0000001" when "00101101110111010", -- t[23482] = 1
      "0000001" when "00101101110111011", -- t[23483] = 1
      "0000001" when "00101101110111100", -- t[23484] = 1
      "0000001" when "00101101110111101", -- t[23485] = 1
      "0000001" when "00101101110111110", -- t[23486] = 1
      "0000001" when "00101101110111111", -- t[23487] = 1
      "0000001" when "00101101111000000", -- t[23488] = 1
      "0000001" when "00101101111000001", -- t[23489] = 1
      "0000001" when "00101101111000010", -- t[23490] = 1
      "0000001" when "00101101111000011", -- t[23491] = 1
      "0000001" when "00101101111000100", -- t[23492] = 1
      "0000001" when "00101101111000101", -- t[23493] = 1
      "0000001" when "00101101111000110", -- t[23494] = 1
      "0000001" when "00101101111000111", -- t[23495] = 1
      "0000001" when "00101101111001000", -- t[23496] = 1
      "0000001" when "00101101111001001", -- t[23497] = 1
      "0000001" when "00101101111001010", -- t[23498] = 1
      "0000001" when "00101101111001011", -- t[23499] = 1
      "0000001" when "00101101111001100", -- t[23500] = 1
      "0000001" when "00101101111001101", -- t[23501] = 1
      "0000001" when "00101101111001110", -- t[23502] = 1
      "0000001" when "00101101111001111", -- t[23503] = 1
      "0000001" when "00101101111010000", -- t[23504] = 1
      "0000001" when "00101101111010001", -- t[23505] = 1
      "0000001" when "00101101111010010", -- t[23506] = 1
      "0000001" when "00101101111010011", -- t[23507] = 1
      "0000001" when "00101101111010100", -- t[23508] = 1
      "0000001" when "00101101111010101", -- t[23509] = 1
      "0000001" when "00101101111010110", -- t[23510] = 1
      "0000001" when "00101101111010111", -- t[23511] = 1
      "0000001" when "00101101111011000", -- t[23512] = 1
      "0000001" when "00101101111011001", -- t[23513] = 1
      "0000001" when "00101101111011010", -- t[23514] = 1
      "0000001" when "00101101111011011", -- t[23515] = 1
      "0000001" when "00101101111011100", -- t[23516] = 1
      "0000001" when "00101101111011101", -- t[23517] = 1
      "0000001" when "00101101111011110", -- t[23518] = 1
      "0000001" when "00101101111011111", -- t[23519] = 1
      "0000001" when "00101101111100000", -- t[23520] = 1
      "0000001" when "00101101111100001", -- t[23521] = 1
      "0000001" when "00101101111100010", -- t[23522] = 1
      "0000001" when "00101101111100011", -- t[23523] = 1
      "0000001" when "00101101111100100", -- t[23524] = 1
      "0000001" when "00101101111100101", -- t[23525] = 1
      "0000001" when "00101101111100110", -- t[23526] = 1
      "0000001" when "00101101111100111", -- t[23527] = 1
      "0000001" when "00101101111101000", -- t[23528] = 1
      "0000001" when "00101101111101001", -- t[23529] = 1
      "0000001" when "00101101111101010", -- t[23530] = 1
      "0000001" when "00101101111101011", -- t[23531] = 1
      "0000001" when "00101101111101100", -- t[23532] = 1
      "0000001" when "00101101111101101", -- t[23533] = 1
      "0000001" when "00101101111101110", -- t[23534] = 1
      "0000001" when "00101101111101111", -- t[23535] = 1
      "0000001" when "00101101111110000", -- t[23536] = 1
      "0000001" when "00101101111110001", -- t[23537] = 1
      "0000001" when "00101101111110010", -- t[23538] = 1
      "0000001" when "00101101111110011", -- t[23539] = 1
      "0000001" when "00101101111110100", -- t[23540] = 1
      "0000001" when "00101101111110101", -- t[23541] = 1
      "0000001" when "00101101111110110", -- t[23542] = 1
      "0000001" when "00101101111110111", -- t[23543] = 1
      "0000001" when "00101101111111000", -- t[23544] = 1
      "0000001" when "00101101111111001", -- t[23545] = 1
      "0000001" when "00101101111111010", -- t[23546] = 1
      "0000001" when "00101101111111011", -- t[23547] = 1
      "0000001" when "00101101111111100", -- t[23548] = 1
      "0000001" when "00101101111111101", -- t[23549] = 1
      "0000001" when "00101101111111110", -- t[23550] = 1
      "0000001" when "00101101111111111", -- t[23551] = 1
      "0000001" when "00101110000000000", -- t[23552] = 1
      "0000001" when "00101110000000001", -- t[23553] = 1
      "0000001" when "00101110000000010", -- t[23554] = 1
      "0000001" when "00101110000000011", -- t[23555] = 1
      "0000001" when "00101110000000100", -- t[23556] = 1
      "0000001" when "00101110000000101", -- t[23557] = 1
      "0000001" when "00101110000000110", -- t[23558] = 1
      "0000001" when "00101110000000111", -- t[23559] = 1
      "0000001" when "00101110000001000", -- t[23560] = 1
      "0000001" when "00101110000001001", -- t[23561] = 1
      "0000001" when "00101110000001010", -- t[23562] = 1
      "0000001" when "00101110000001011", -- t[23563] = 1
      "0000001" when "00101110000001100", -- t[23564] = 1
      "0000001" when "00101110000001101", -- t[23565] = 1
      "0000001" when "00101110000001110", -- t[23566] = 1
      "0000001" when "00101110000001111", -- t[23567] = 1
      "0000001" when "00101110000010000", -- t[23568] = 1
      "0000001" when "00101110000010001", -- t[23569] = 1
      "0000001" when "00101110000010010", -- t[23570] = 1
      "0000001" when "00101110000010011", -- t[23571] = 1
      "0000001" when "00101110000010100", -- t[23572] = 1
      "0000001" when "00101110000010101", -- t[23573] = 1
      "0000001" when "00101110000010110", -- t[23574] = 1
      "0000001" when "00101110000010111", -- t[23575] = 1
      "0000001" when "00101110000011000", -- t[23576] = 1
      "0000001" when "00101110000011001", -- t[23577] = 1
      "0000001" when "00101110000011010", -- t[23578] = 1
      "0000001" when "00101110000011011", -- t[23579] = 1
      "0000001" when "00101110000011100", -- t[23580] = 1
      "0000001" when "00101110000011101", -- t[23581] = 1
      "0000001" when "00101110000011110", -- t[23582] = 1
      "0000001" when "00101110000011111", -- t[23583] = 1
      "0000001" when "00101110000100000", -- t[23584] = 1
      "0000001" when "00101110000100001", -- t[23585] = 1
      "0000001" when "00101110000100010", -- t[23586] = 1
      "0000001" when "00101110000100011", -- t[23587] = 1
      "0000001" when "00101110000100100", -- t[23588] = 1
      "0000001" when "00101110000100101", -- t[23589] = 1
      "0000001" when "00101110000100110", -- t[23590] = 1
      "0000001" when "00101110000100111", -- t[23591] = 1
      "0000001" when "00101110000101000", -- t[23592] = 1
      "0000001" when "00101110000101001", -- t[23593] = 1
      "0000001" when "00101110000101010", -- t[23594] = 1
      "0000001" when "00101110000101011", -- t[23595] = 1
      "0000001" when "00101110000101100", -- t[23596] = 1
      "0000001" when "00101110000101101", -- t[23597] = 1
      "0000001" when "00101110000101110", -- t[23598] = 1
      "0000001" when "00101110000101111", -- t[23599] = 1
      "0000001" when "00101110000110000", -- t[23600] = 1
      "0000001" when "00101110000110001", -- t[23601] = 1
      "0000001" when "00101110000110010", -- t[23602] = 1
      "0000001" when "00101110000110011", -- t[23603] = 1
      "0000001" when "00101110000110100", -- t[23604] = 1
      "0000001" when "00101110000110101", -- t[23605] = 1
      "0000001" when "00101110000110110", -- t[23606] = 1
      "0000001" when "00101110000110111", -- t[23607] = 1
      "0000001" when "00101110000111000", -- t[23608] = 1
      "0000001" when "00101110000111001", -- t[23609] = 1
      "0000001" when "00101110000111010", -- t[23610] = 1
      "0000001" when "00101110000111011", -- t[23611] = 1
      "0000001" when "00101110000111100", -- t[23612] = 1
      "0000001" when "00101110000111101", -- t[23613] = 1
      "0000001" when "00101110000111110", -- t[23614] = 1
      "0000001" when "00101110000111111", -- t[23615] = 1
      "0000001" when "00101110001000000", -- t[23616] = 1
      "0000001" when "00101110001000001", -- t[23617] = 1
      "0000001" when "00101110001000010", -- t[23618] = 1
      "0000001" when "00101110001000011", -- t[23619] = 1
      "0000001" when "00101110001000100", -- t[23620] = 1
      "0000001" when "00101110001000101", -- t[23621] = 1
      "0000001" when "00101110001000110", -- t[23622] = 1
      "0000001" when "00101110001000111", -- t[23623] = 1
      "0000001" when "00101110001001000", -- t[23624] = 1
      "0000001" when "00101110001001001", -- t[23625] = 1
      "0000001" when "00101110001001010", -- t[23626] = 1
      "0000001" when "00101110001001011", -- t[23627] = 1
      "0000001" when "00101110001001100", -- t[23628] = 1
      "0000001" when "00101110001001101", -- t[23629] = 1
      "0000001" when "00101110001001110", -- t[23630] = 1
      "0000001" when "00101110001001111", -- t[23631] = 1
      "0000001" when "00101110001010000", -- t[23632] = 1
      "0000001" when "00101110001010001", -- t[23633] = 1
      "0000001" when "00101110001010010", -- t[23634] = 1
      "0000001" when "00101110001010011", -- t[23635] = 1
      "0000001" when "00101110001010100", -- t[23636] = 1
      "0000001" when "00101110001010101", -- t[23637] = 1
      "0000001" when "00101110001010110", -- t[23638] = 1
      "0000001" when "00101110001010111", -- t[23639] = 1
      "0000001" when "00101110001011000", -- t[23640] = 1
      "0000001" when "00101110001011001", -- t[23641] = 1
      "0000001" when "00101110001011010", -- t[23642] = 1
      "0000001" when "00101110001011011", -- t[23643] = 1
      "0000001" when "00101110001011100", -- t[23644] = 1
      "0000001" when "00101110001011101", -- t[23645] = 1
      "0000001" when "00101110001011110", -- t[23646] = 1
      "0000001" when "00101110001011111", -- t[23647] = 1
      "0000001" when "00101110001100000", -- t[23648] = 1
      "0000001" when "00101110001100001", -- t[23649] = 1
      "0000001" when "00101110001100010", -- t[23650] = 1
      "0000001" when "00101110001100011", -- t[23651] = 1
      "0000001" when "00101110001100100", -- t[23652] = 1
      "0000001" when "00101110001100101", -- t[23653] = 1
      "0000001" when "00101110001100110", -- t[23654] = 1
      "0000001" when "00101110001100111", -- t[23655] = 1
      "0000001" when "00101110001101000", -- t[23656] = 1
      "0000001" when "00101110001101001", -- t[23657] = 1
      "0000001" when "00101110001101010", -- t[23658] = 1
      "0000001" when "00101110001101011", -- t[23659] = 1
      "0000001" when "00101110001101100", -- t[23660] = 1
      "0000001" when "00101110001101101", -- t[23661] = 1
      "0000001" when "00101110001101110", -- t[23662] = 1
      "0000001" when "00101110001101111", -- t[23663] = 1
      "0000001" when "00101110001110000", -- t[23664] = 1
      "0000001" when "00101110001110001", -- t[23665] = 1
      "0000001" when "00101110001110010", -- t[23666] = 1
      "0000001" when "00101110001110011", -- t[23667] = 1
      "0000001" when "00101110001110100", -- t[23668] = 1
      "0000001" when "00101110001110101", -- t[23669] = 1
      "0000001" when "00101110001110110", -- t[23670] = 1
      "0000001" when "00101110001110111", -- t[23671] = 1
      "0000001" when "00101110001111000", -- t[23672] = 1
      "0000001" when "00101110001111001", -- t[23673] = 1
      "0000001" when "00101110001111010", -- t[23674] = 1
      "0000001" when "00101110001111011", -- t[23675] = 1
      "0000001" when "00101110001111100", -- t[23676] = 1
      "0000001" when "00101110001111101", -- t[23677] = 1
      "0000001" when "00101110001111110", -- t[23678] = 1
      "0000001" when "00101110001111111", -- t[23679] = 1
      "0000001" when "00101110010000000", -- t[23680] = 1
      "0000001" when "00101110010000001", -- t[23681] = 1
      "0000001" when "00101110010000010", -- t[23682] = 1
      "0000001" when "00101110010000011", -- t[23683] = 1
      "0000001" when "00101110010000100", -- t[23684] = 1
      "0000001" when "00101110010000101", -- t[23685] = 1
      "0000001" when "00101110010000110", -- t[23686] = 1
      "0000001" when "00101110010000111", -- t[23687] = 1
      "0000001" when "00101110010001000", -- t[23688] = 1
      "0000001" when "00101110010001001", -- t[23689] = 1
      "0000001" when "00101110010001010", -- t[23690] = 1
      "0000001" when "00101110010001011", -- t[23691] = 1
      "0000001" when "00101110010001100", -- t[23692] = 1
      "0000001" when "00101110010001101", -- t[23693] = 1
      "0000001" when "00101110010001110", -- t[23694] = 1
      "0000001" when "00101110010001111", -- t[23695] = 1
      "0000001" when "00101110010010000", -- t[23696] = 1
      "0000001" when "00101110010010001", -- t[23697] = 1
      "0000001" when "00101110010010010", -- t[23698] = 1
      "0000001" when "00101110010010011", -- t[23699] = 1
      "0000001" when "00101110010010100", -- t[23700] = 1
      "0000001" when "00101110010010101", -- t[23701] = 1
      "0000001" when "00101110010010110", -- t[23702] = 1
      "0000001" when "00101110010010111", -- t[23703] = 1
      "0000001" when "00101110010011000", -- t[23704] = 1
      "0000001" when "00101110010011001", -- t[23705] = 1
      "0000001" when "00101110010011010", -- t[23706] = 1
      "0000001" when "00101110010011011", -- t[23707] = 1
      "0000001" when "00101110010011100", -- t[23708] = 1
      "0000001" when "00101110010011101", -- t[23709] = 1
      "0000001" when "00101110010011110", -- t[23710] = 1
      "0000001" when "00101110010011111", -- t[23711] = 1
      "0000001" when "00101110010100000", -- t[23712] = 1
      "0000001" when "00101110010100001", -- t[23713] = 1
      "0000001" when "00101110010100010", -- t[23714] = 1
      "0000001" when "00101110010100011", -- t[23715] = 1
      "0000001" when "00101110010100100", -- t[23716] = 1
      "0000001" when "00101110010100101", -- t[23717] = 1
      "0000001" when "00101110010100110", -- t[23718] = 1
      "0000001" when "00101110010100111", -- t[23719] = 1
      "0000001" when "00101110010101000", -- t[23720] = 1
      "0000001" when "00101110010101001", -- t[23721] = 1
      "0000001" when "00101110010101010", -- t[23722] = 1
      "0000001" when "00101110010101011", -- t[23723] = 1
      "0000001" when "00101110010101100", -- t[23724] = 1
      "0000001" when "00101110010101101", -- t[23725] = 1
      "0000001" when "00101110010101110", -- t[23726] = 1
      "0000001" when "00101110010101111", -- t[23727] = 1
      "0000001" when "00101110010110000", -- t[23728] = 1
      "0000001" when "00101110010110001", -- t[23729] = 1
      "0000001" when "00101110010110010", -- t[23730] = 1
      "0000001" when "00101110010110011", -- t[23731] = 1
      "0000001" when "00101110010110100", -- t[23732] = 1
      "0000001" when "00101110010110101", -- t[23733] = 1
      "0000001" when "00101110010110110", -- t[23734] = 1
      "0000001" when "00101110010110111", -- t[23735] = 1
      "0000001" when "00101110010111000", -- t[23736] = 1
      "0000001" when "00101110010111001", -- t[23737] = 1
      "0000001" when "00101110010111010", -- t[23738] = 1
      "0000001" when "00101110010111011", -- t[23739] = 1
      "0000001" when "00101110010111100", -- t[23740] = 1
      "0000001" when "00101110010111101", -- t[23741] = 1
      "0000001" when "00101110010111110", -- t[23742] = 1
      "0000001" when "00101110010111111", -- t[23743] = 1
      "0000001" when "00101110011000000", -- t[23744] = 1
      "0000001" when "00101110011000001", -- t[23745] = 1
      "0000001" when "00101110011000010", -- t[23746] = 1
      "0000001" when "00101110011000011", -- t[23747] = 1
      "0000001" when "00101110011000100", -- t[23748] = 1
      "0000001" when "00101110011000101", -- t[23749] = 1
      "0000001" when "00101110011000110", -- t[23750] = 1
      "0000001" when "00101110011000111", -- t[23751] = 1
      "0000001" when "00101110011001000", -- t[23752] = 1
      "0000001" when "00101110011001001", -- t[23753] = 1
      "0000001" when "00101110011001010", -- t[23754] = 1
      "0000001" when "00101110011001011", -- t[23755] = 1
      "0000001" when "00101110011001100", -- t[23756] = 1
      "0000001" when "00101110011001101", -- t[23757] = 1
      "0000001" when "00101110011001110", -- t[23758] = 1
      "0000001" when "00101110011001111", -- t[23759] = 1
      "0000001" when "00101110011010000", -- t[23760] = 1
      "0000001" when "00101110011010001", -- t[23761] = 1
      "0000001" when "00101110011010010", -- t[23762] = 1
      "0000001" when "00101110011010011", -- t[23763] = 1
      "0000001" when "00101110011010100", -- t[23764] = 1
      "0000001" when "00101110011010101", -- t[23765] = 1
      "0000001" when "00101110011010110", -- t[23766] = 1
      "0000001" when "00101110011010111", -- t[23767] = 1
      "0000001" when "00101110011011000", -- t[23768] = 1
      "0000001" when "00101110011011001", -- t[23769] = 1
      "0000001" when "00101110011011010", -- t[23770] = 1
      "0000001" when "00101110011011011", -- t[23771] = 1
      "0000001" when "00101110011011100", -- t[23772] = 1
      "0000001" when "00101110011011101", -- t[23773] = 1
      "0000001" when "00101110011011110", -- t[23774] = 1
      "0000001" when "00101110011011111", -- t[23775] = 1
      "0000001" when "00101110011100000", -- t[23776] = 1
      "0000001" when "00101110011100001", -- t[23777] = 1
      "0000001" when "00101110011100010", -- t[23778] = 1
      "0000001" when "00101110011100011", -- t[23779] = 1
      "0000001" when "00101110011100100", -- t[23780] = 1
      "0000001" when "00101110011100101", -- t[23781] = 1
      "0000001" when "00101110011100110", -- t[23782] = 1
      "0000001" when "00101110011100111", -- t[23783] = 1
      "0000001" when "00101110011101000", -- t[23784] = 1
      "0000001" when "00101110011101001", -- t[23785] = 1
      "0000001" when "00101110011101010", -- t[23786] = 1
      "0000001" when "00101110011101011", -- t[23787] = 1
      "0000001" when "00101110011101100", -- t[23788] = 1
      "0000001" when "00101110011101101", -- t[23789] = 1
      "0000001" when "00101110011101110", -- t[23790] = 1
      "0000001" when "00101110011101111", -- t[23791] = 1
      "0000001" when "00101110011110000", -- t[23792] = 1
      "0000001" when "00101110011110001", -- t[23793] = 1
      "0000001" when "00101110011110010", -- t[23794] = 1
      "0000001" when "00101110011110011", -- t[23795] = 1
      "0000001" when "00101110011110100", -- t[23796] = 1
      "0000001" when "00101110011110101", -- t[23797] = 1
      "0000001" when "00101110011110110", -- t[23798] = 1
      "0000001" when "00101110011110111", -- t[23799] = 1
      "0000001" when "00101110011111000", -- t[23800] = 1
      "0000001" when "00101110011111001", -- t[23801] = 1
      "0000001" when "00101110011111010", -- t[23802] = 1
      "0000001" when "00101110011111011", -- t[23803] = 1
      "0000001" when "00101110011111100", -- t[23804] = 1
      "0000001" when "00101110011111101", -- t[23805] = 1
      "0000001" when "00101110011111110", -- t[23806] = 1
      "0000001" when "00101110011111111", -- t[23807] = 1
      "0000001" when "00101110100000000", -- t[23808] = 1
      "0000001" when "00101110100000001", -- t[23809] = 1
      "0000001" when "00101110100000010", -- t[23810] = 1
      "0000001" when "00101110100000011", -- t[23811] = 1
      "0000001" when "00101110100000100", -- t[23812] = 1
      "0000001" when "00101110100000101", -- t[23813] = 1
      "0000001" when "00101110100000110", -- t[23814] = 1
      "0000001" when "00101110100000111", -- t[23815] = 1
      "0000001" when "00101110100001000", -- t[23816] = 1
      "0000001" when "00101110100001001", -- t[23817] = 1
      "0000001" when "00101110100001010", -- t[23818] = 1
      "0000001" when "00101110100001011", -- t[23819] = 1
      "0000001" when "00101110100001100", -- t[23820] = 1
      "0000001" when "00101110100001101", -- t[23821] = 1
      "0000001" when "00101110100001110", -- t[23822] = 1
      "0000001" when "00101110100001111", -- t[23823] = 1
      "0000001" when "00101110100010000", -- t[23824] = 1
      "0000001" when "00101110100010001", -- t[23825] = 1
      "0000001" when "00101110100010010", -- t[23826] = 1
      "0000001" when "00101110100010011", -- t[23827] = 1
      "0000001" when "00101110100010100", -- t[23828] = 1
      "0000001" when "00101110100010101", -- t[23829] = 1
      "0000001" when "00101110100010110", -- t[23830] = 1
      "0000001" when "00101110100010111", -- t[23831] = 1
      "0000001" when "00101110100011000", -- t[23832] = 1
      "0000001" when "00101110100011001", -- t[23833] = 1
      "0000001" when "00101110100011010", -- t[23834] = 1
      "0000001" when "00101110100011011", -- t[23835] = 1
      "0000001" when "00101110100011100", -- t[23836] = 1
      "0000001" when "00101110100011101", -- t[23837] = 1
      "0000001" when "00101110100011110", -- t[23838] = 1
      "0000001" when "00101110100011111", -- t[23839] = 1
      "0000001" when "00101110100100000", -- t[23840] = 1
      "0000001" when "00101110100100001", -- t[23841] = 1
      "0000001" when "00101110100100010", -- t[23842] = 1
      "0000001" when "00101110100100011", -- t[23843] = 1
      "0000001" when "00101110100100100", -- t[23844] = 1
      "0000001" when "00101110100100101", -- t[23845] = 1
      "0000001" when "00101110100100110", -- t[23846] = 1
      "0000001" when "00101110100100111", -- t[23847] = 1
      "0000001" when "00101110100101000", -- t[23848] = 1
      "0000001" when "00101110100101001", -- t[23849] = 1
      "0000001" when "00101110100101010", -- t[23850] = 1
      "0000001" when "00101110100101011", -- t[23851] = 1
      "0000001" when "00101110100101100", -- t[23852] = 1
      "0000001" when "00101110100101101", -- t[23853] = 1
      "0000001" when "00101110100101110", -- t[23854] = 1
      "0000001" when "00101110100101111", -- t[23855] = 1
      "0000001" when "00101110100110000", -- t[23856] = 1
      "0000001" when "00101110100110001", -- t[23857] = 1
      "0000001" when "00101110100110010", -- t[23858] = 1
      "0000001" when "00101110100110011", -- t[23859] = 1
      "0000001" when "00101110100110100", -- t[23860] = 1
      "0000001" when "00101110100110101", -- t[23861] = 1
      "0000001" when "00101110100110110", -- t[23862] = 1
      "0000001" when "00101110100110111", -- t[23863] = 1
      "0000001" when "00101110100111000", -- t[23864] = 1
      "0000001" when "00101110100111001", -- t[23865] = 1
      "0000001" when "00101110100111010", -- t[23866] = 1
      "0000001" when "00101110100111011", -- t[23867] = 1
      "0000001" when "00101110100111100", -- t[23868] = 1
      "0000001" when "00101110100111101", -- t[23869] = 1
      "0000001" when "00101110100111110", -- t[23870] = 1
      "0000001" when "00101110100111111", -- t[23871] = 1
      "0000001" when "00101110101000000", -- t[23872] = 1
      "0000001" when "00101110101000001", -- t[23873] = 1
      "0000001" when "00101110101000010", -- t[23874] = 1
      "0000001" when "00101110101000011", -- t[23875] = 1
      "0000001" when "00101110101000100", -- t[23876] = 1
      "0000001" when "00101110101000101", -- t[23877] = 1
      "0000001" when "00101110101000110", -- t[23878] = 1
      "0000001" when "00101110101000111", -- t[23879] = 1
      "0000001" when "00101110101001000", -- t[23880] = 1
      "0000001" when "00101110101001001", -- t[23881] = 1
      "0000001" when "00101110101001010", -- t[23882] = 1
      "0000001" when "00101110101001011", -- t[23883] = 1
      "0000001" when "00101110101001100", -- t[23884] = 1
      "0000001" when "00101110101001101", -- t[23885] = 1
      "0000001" when "00101110101001110", -- t[23886] = 1
      "0000001" when "00101110101001111", -- t[23887] = 1
      "0000001" when "00101110101010000", -- t[23888] = 1
      "0000001" when "00101110101010001", -- t[23889] = 1
      "0000001" when "00101110101010010", -- t[23890] = 1
      "0000001" when "00101110101010011", -- t[23891] = 1
      "0000001" when "00101110101010100", -- t[23892] = 1
      "0000001" when "00101110101010101", -- t[23893] = 1
      "0000001" when "00101110101010110", -- t[23894] = 1
      "0000001" when "00101110101010111", -- t[23895] = 1
      "0000001" when "00101110101011000", -- t[23896] = 1
      "0000001" when "00101110101011001", -- t[23897] = 1
      "0000001" when "00101110101011010", -- t[23898] = 1
      "0000001" when "00101110101011011", -- t[23899] = 1
      "0000001" when "00101110101011100", -- t[23900] = 1
      "0000001" when "00101110101011101", -- t[23901] = 1
      "0000001" when "00101110101011110", -- t[23902] = 1
      "0000001" when "00101110101011111", -- t[23903] = 1
      "0000001" when "00101110101100000", -- t[23904] = 1
      "0000001" when "00101110101100001", -- t[23905] = 1
      "0000001" when "00101110101100010", -- t[23906] = 1
      "0000001" when "00101110101100011", -- t[23907] = 1
      "0000001" when "00101110101100100", -- t[23908] = 1
      "0000001" when "00101110101100101", -- t[23909] = 1
      "0000001" when "00101110101100110", -- t[23910] = 1
      "0000001" when "00101110101100111", -- t[23911] = 1
      "0000001" when "00101110101101000", -- t[23912] = 1
      "0000001" when "00101110101101001", -- t[23913] = 1
      "0000001" when "00101110101101010", -- t[23914] = 1
      "0000001" when "00101110101101011", -- t[23915] = 1
      "0000001" when "00101110101101100", -- t[23916] = 1
      "0000001" when "00101110101101101", -- t[23917] = 1
      "0000001" when "00101110101101110", -- t[23918] = 1
      "0000001" when "00101110101101111", -- t[23919] = 1
      "0000001" when "00101110101110000", -- t[23920] = 1
      "0000001" when "00101110101110001", -- t[23921] = 1
      "0000001" when "00101110101110010", -- t[23922] = 1
      "0000001" when "00101110101110011", -- t[23923] = 1
      "0000001" when "00101110101110100", -- t[23924] = 1
      "0000001" when "00101110101110101", -- t[23925] = 1
      "0000001" when "00101110101110110", -- t[23926] = 1
      "0000001" when "00101110101110111", -- t[23927] = 1
      "0000001" when "00101110101111000", -- t[23928] = 1
      "0000001" when "00101110101111001", -- t[23929] = 1
      "0000001" when "00101110101111010", -- t[23930] = 1
      "0000001" when "00101110101111011", -- t[23931] = 1
      "0000001" when "00101110101111100", -- t[23932] = 1
      "0000001" when "00101110101111101", -- t[23933] = 1
      "0000001" when "00101110101111110", -- t[23934] = 1
      "0000001" when "00101110101111111", -- t[23935] = 1
      "0000001" when "00101110110000000", -- t[23936] = 1
      "0000001" when "00101110110000001", -- t[23937] = 1
      "0000001" when "00101110110000010", -- t[23938] = 1
      "0000001" when "00101110110000011", -- t[23939] = 1
      "0000001" when "00101110110000100", -- t[23940] = 1
      "0000001" when "00101110110000101", -- t[23941] = 1
      "0000001" when "00101110110000110", -- t[23942] = 1
      "0000001" when "00101110110000111", -- t[23943] = 1
      "0000001" when "00101110110001000", -- t[23944] = 1
      "0000001" when "00101110110001001", -- t[23945] = 1
      "0000001" when "00101110110001010", -- t[23946] = 1
      "0000001" when "00101110110001011", -- t[23947] = 1
      "0000001" when "00101110110001100", -- t[23948] = 1
      "0000001" when "00101110110001101", -- t[23949] = 1
      "0000001" when "00101110110001110", -- t[23950] = 1
      "0000001" when "00101110110001111", -- t[23951] = 1
      "0000001" when "00101110110010000", -- t[23952] = 1
      "0000001" when "00101110110010001", -- t[23953] = 1
      "0000001" when "00101110110010010", -- t[23954] = 1
      "0000001" when "00101110110010011", -- t[23955] = 1
      "0000001" when "00101110110010100", -- t[23956] = 1
      "0000001" when "00101110110010101", -- t[23957] = 1
      "0000001" when "00101110110010110", -- t[23958] = 1
      "0000001" when "00101110110010111", -- t[23959] = 1
      "0000001" when "00101110110011000", -- t[23960] = 1
      "0000001" when "00101110110011001", -- t[23961] = 1
      "0000001" when "00101110110011010", -- t[23962] = 1
      "0000001" when "00101110110011011", -- t[23963] = 1
      "0000001" when "00101110110011100", -- t[23964] = 1
      "0000001" when "00101110110011101", -- t[23965] = 1
      "0000001" when "00101110110011110", -- t[23966] = 1
      "0000001" when "00101110110011111", -- t[23967] = 1
      "0000001" when "00101110110100000", -- t[23968] = 1
      "0000001" when "00101110110100001", -- t[23969] = 1
      "0000001" when "00101110110100010", -- t[23970] = 1
      "0000001" when "00101110110100011", -- t[23971] = 1
      "0000001" when "00101110110100100", -- t[23972] = 1
      "0000001" when "00101110110100101", -- t[23973] = 1
      "0000001" when "00101110110100110", -- t[23974] = 1
      "0000001" when "00101110110100111", -- t[23975] = 1
      "0000001" when "00101110110101000", -- t[23976] = 1
      "0000001" when "00101110110101001", -- t[23977] = 1
      "0000001" when "00101110110101010", -- t[23978] = 1
      "0000001" when "00101110110101011", -- t[23979] = 1
      "0000001" when "00101110110101100", -- t[23980] = 1
      "0000001" when "00101110110101101", -- t[23981] = 1
      "0000001" when "00101110110101110", -- t[23982] = 1
      "0000001" when "00101110110101111", -- t[23983] = 1
      "0000001" when "00101110110110000", -- t[23984] = 1
      "0000001" when "00101110110110001", -- t[23985] = 1
      "0000001" when "00101110110110010", -- t[23986] = 1
      "0000001" when "00101110110110011", -- t[23987] = 1
      "0000001" when "00101110110110100", -- t[23988] = 1
      "0000001" when "00101110110110101", -- t[23989] = 1
      "0000001" when "00101110110110110", -- t[23990] = 1
      "0000001" when "00101110110110111", -- t[23991] = 1
      "0000001" when "00101110110111000", -- t[23992] = 1
      "0000001" when "00101110110111001", -- t[23993] = 1
      "0000001" when "00101110110111010", -- t[23994] = 1
      "0000001" when "00101110110111011", -- t[23995] = 1
      "0000001" when "00101110110111100", -- t[23996] = 1
      "0000001" when "00101110110111101", -- t[23997] = 1
      "0000001" when "00101110110111110", -- t[23998] = 1
      "0000001" when "00101110110111111", -- t[23999] = 1
      "0000001" when "00101110111000000", -- t[24000] = 1
      "0000001" when "00101110111000001", -- t[24001] = 1
      "0000001" when "00101110111000010", -- t[24002] = 1
      "0000001" when "00101110111000011", -- t[24003] = 1
      "0000001" when "00101110111000100", -- t[24004] = 1
      "0000001" when "00101110111000101", -- t[24005] = 1
      "0000001" when "00101110111000110", -- t[24006] = 1
      "0000001" when "00101110111000111", -- t[24007] = 1
      "0000001" when "00101110111001000", -- t[24008] = 1
      "0000001" when "00101110111001001", -- t[24009] = 1
      "0000001" when "00101110111001010", -- t[24010] = 1
      "0000001" when "00101110111001011", -- t[24011] = 1
      "0000001" when "00101110111001100", -- t[24012] = 1
      "0000001" when "00101110111001101", -- t[24013] = 1
      "0000001" when "00101110111001110", -- t[24014] = 1
      "0000001" when "00101110111001111", -- t[24015] = 1
      "0000001" when "00101110111010000", -- t[24016] = 1
      "0000001" when "00101110111010001", -- t[24017] = 1
      "0000001" when "00101110111010010", -- t[24018] = 1
      "0000001" when "00101110111010011", -- t[24019] = 1
      "0000001" when "00101110111010100", -- t[24020] = 1
      "0000001" when "00101110111010101", -- t[24021] = 1
      "0000001" when "00101110111010110", -- t[24022] = 1
      "0000001" when "00101110111010111", -- t[24023] = 1
      "0000001" when "00101110111011000", -- t[24024] = 1
      "0000001" when "00101110111011001", -- t[24025] = 1
      "0000001" when "00101110111011010", -- t[24026] = 1
      "0000001" when "00101110111011011", -- t[24027] = 1
      "0000001" when "00101110111011100", -- t[24028] = 1
      "0000001" when "00101110111011101", -- t[24029] = 1
      "0000001" when "00101110111011110", -- t[24030] = 1
      "0000001" when "00101110111011111", -- t[24031] = 1
      "0000001" when "00101110111100000", -- t[24032] = 1
      "0000001" when "00101110111100001", -- t[24033] = 1
      "0000001" when "00101110111100010", -- t[24034] = 1
      "0000001" when "00101110111100011", -- t[24035] = 1
      "0000001" when "00101110111100100", -- t[24036] = 1
      "0000001" when "00101110111100101", -- t[24037] = 1
      "0000001" when "00101110111100110", -- t[24038] = 1
      "0000001" when "00101110111100111", -- t[24039] = 1
      "0000001" when "00101110111101000", -- t[24040] = 1
      "0000001" when "00101110111101001", -- t[24041] = 1
      "0000001" when "00101110111101010", -- t[24042] = 1
      "0000001" when "00101110111101011", -- t[24043] = 1
      "0000001" when "00101110111101100", -- t[24044] = 1
      "0000001" when "00101110111101101", -- t[24045] = 1
      "0000001" when "00101110111101110", -- t[24046] = 1
      "0000001" when "00101110111101111", -- t[24047] = 1
      "0000001" when "00101110111110000", -- t[24048] = 1
      "0000001" when "00101110111110001", -- t[24049] = 1
      "0000001" when "00101110111110010", -- t[24050] = 1
      "0000001" when "00101110111110011", -- t[24051] = 1
      "0000001" when "00101110111110100", -- t[24052] = 1
      "0000001" when "00101110111110101", -- t[24053] = 1
      "0000001" when "00101110111110110", -- t[24054] = 1
      "0000001" when "00101110111110111", -- t[24055] = 1
      "0000001" when "00101110111111000", -- t[24056] = 1
      "0000001" when "00101110111111001", -- t[24057] = 1
      "0000001" when "00101110111111010", -- t[24058] = 1
      "0000001" when "00101110111111011", -- t[24059] = 1
      "0000001" when "00101110111111100", -- t[24060] = 1
      "0000001" when "00101110111111101", -- t[24061] = 1
      "0000001" when "00101110111111110", -- t[24062] = 1
      "0000001" when "00101110111111111", -- t[24063] = 1
      "0000001" when "00101111000000000", -- t[24064] = 1
      "0000001" when "00101111000000001", -- t[24065] = 1
      "0000001" when "00101111000000010", -- t[24066] = 1
      "0000001" when "00101111000000011", -- t[24067] = 1
      "0000001" when "00101111000000100", -- t[24068] = 1
      "0000001" when "00101111000000101", -- t[24069] = 1
      "0000001" when "00101111000000110", -- t[24070] = 1
      "0000001" when "00101111000000111", -- t[24071] = 1
      "0000001" when "00101111000001000", -- t[24072] = 1
      "0000001" when "00101111000001001", -- t[24073] = 1
      "0000001" when "00101111000001010", -- t[24074] = 1
      "0000001" when "00101111000001011", -- t[24075] = 1
      "0000001" when "00101111000001100", -- t[24076] = 1
      "0000001" when "00101111000001101", -- t[24077] = 1
      "0000001" when "00101111000001110", -- t[24078] = 1
      "0000001" when "00101111000001111", -- t[24079] = 1
      "0000001" when "00101111000010000", -- t[24080] = 1
      "0000001" when "00101111000010001", -- t[24081] = 1
      "0000001" when "00101111000010010", -- t[24082] = 1
      "0000001" when "00101111000010011", -- t[24083] = 1
      "0000001" when "00101111000010100", -- t[24084] = 1
      "0000001" when "00101111000010101", -- t[24085] = 1
      "0000001" when "00101111000010110", -- t[24086] = 1
      "0000001" when "00101111000010111", -- t[24087] = 1
      "0000001" when "00101111000011000", -- t[24088] = 1
      "0000001" when "00101111000011001", -- t[24089] = 1
      "0000001" when "00101111000011010", -- t[24090] = 1
      "0000001" when "00101111000011011", -- t[24091] = 1
      "0000001" when "00101111000011100", -- t[24092] = 1
      "0000001" when "00101111000011101", -- t[24093] = 1
      "0000001" when "00101111000011110", -- t[24094] = 1
      "0000001" when "00101111000011111", -- t[24095] = 1
      "0000001" when "00101111000100000", -- t[24096] = 1
      "0000001" when "00101111000100001", -- t[24097] = 1
      "0000001" when "00101111000100010", -- t[24098] = 1
      "0000001" when "00101111000100011", -- t[24099] = 1
      "0000001" when "00101111000100100", -- t[24100] = 1
      "0000001" when "00101111000100101", -- t[24101] = 1
      "0000001" when "00101111000100110", -- t[24102] = 1
      "0000001" when "00101111000100111", -- t[24103] = 1
      "0000001" when "00101111000101000", -- t[24104] = 1
      "0000001" when "00101111000101001", -- t[24105] = 1
      "0000001" when "00101111000101010", -- t[24106] = 1
      "0000001" when "00101111000101011", -- t[24107] = 1
      "0000001" when "00101111000101100", -- t[24108] = 1
      "0000001" when "00101111000101101", -- t[24109] = 1
      "0000001" when "00101111000101110", -- t[24110] = 1
      "0000001" when "00101111000101111", -- t[24111] = 1
      "0000001" when "00101111000110000", -- t[24112] = 1
      "0000001" when "00101111000110001", -- t[24113] = 1
      "0000001" when "00101111000110010", -- t[24114] = 1
      "0000001" when "00101111000110011", -- t[24115] = 1
      "0000001" when "00101111000110100", -- t[24116] = 1
      "0000001" when "00101111000110101", -- t[24117] = 1
      "0000001" when "00101111000110110", -- t[24118] = 1
      "0000001" when "00101111000110111", -- t[24119] = 1
      "0000001" when "00101111000111000", -- t[24120] = 1
      "0000001" when "00101111000111001", -- t[24121] = 1
      "0000001" when "00101111000111010", -- t[24122] = 1
      "0000001" when "00101111000111011", -- t[24123] = 1
      "0000001" when "00101111000111100", -- t[24124] = 1
      "0000001" when "00101111000111101", -- t[24125] = 1
      "0000001" when "00101111000111110", -- t[24126] = 1
      "0000001" when "00101111000111111", -- t[24127] = 1
      "0000001" when "00101111001000000", -- t[24128] = 1
      "0000001" when "00101111001000001", -- t[24129] = 1
      "0000001" when "00101111001000010", -- t[24130] = 1
      "0000001" when "00101111001000011", -- t[24131] = 1
      "0000001" when "00101111001000100", -- t[24132] = 1
      "0000001" when "00101111001000101", -- t[24133] = 1
      "0000001" when "00101111001000110", -- t[24134] = 1
      "0000001" when "00101111001000111", -- t[24135] = 1
      "0000001" when "00101111001001000", -- t[24136] = 1
      "0000001" when "00101111001001001", -- t[24137] = 1
      "0000001" when "00101111001001010", -- t[24138] = 1
      "0000001" when "00101111001001011", -- t[24139] = 1
      "0000001" when "00101111001001100", -- t[24140] = 1
      "0000001" when "00101111001001101", -- t[24141] = 1
      "0000001" when "00101111001001110", -- t[24142] = 1
      "0000001" when "00101111001001111", -- t[24143] = 1
      "0000001" when "00101111001010000", -- t[24144] = 1
      "0000001" when "00101111001010001", -- t[24145] = 1
      "0000001" when "00101111001010010", -- t[24146] = 1
      "0000001" when "00101111001010011", -- t[24147] = 1
      "0000001" when "00101111001010100", -- t[24148] = 1
      "0000001" when "00101111001010101", -- t[24149] = 1
      "0000001" when "00101111001010110", -- t[24150] = 1
      "0000001" when "00101111001010111", -- t[24151] = 1
      "0000001" when "00101111001011000", -- t[24152] = 1
      "0000001" when "00101111001011001", -- t[24153] = 1
      "0000001" when "00101111001011010", -- t[24154] = 1
      "0000001" when "00101111001011011", -- t[24155] = 1
      "0000001" when "00101111001011100", -- t[24156] = 1
      "0000001" when "00101111001011101", -- t[24157] = 1
      "0000001" when "00101111001011110", -- t[24158] = 1
      "0000001" when "00101111001011111", -- t[24159] = 1
      "0000001" when "00101111001100000", -- t[24160] = 1
      "0000001" when "00101111001100001", -- t[24161] = 1
      "0000001" when "00101111001100010", -- t[24162] = 1
      "0000001" when "00101111001100011", -- t[24163] = 1
      "0000001" when "00101111001100100", -- t[24164] = 1
      "0000001" when "00101111001100101", -- t[24165] = 1
      "0000001" when "00101111001100110", -- t[24166] = 1
      "0000001" when "00101111001100111", -- t[24167] = 1
      "0000001" when "00101111001101000", -- t[24168] = 1
      "0000001" when "00101111001101001", -- t[24169] = 1
      "0000001" when "00101111001101010", -- t[24170] = 1
      "0000001" when "00101111001101011", -- t[24171] = 1
      "0000001" when "00101111001101100", -- t[24172] = 1
      "0000001" when "00101111001101101", -- t[24173] = 1
      "0000001" when "00101111001101110", -- t[24174] = 1
      "0000001" when "00101111001101111", -- t[24175] = 1
      "0000001" when "00101111001110000", -- t[24176] = 1
      "0000001" when "00101111001110001", -- t[24177] = 1
      "0000001" when "00101111001110010", -- t[24178] = 1
      "0000001" when "00101111001110011", -- t[24179] = 1
      "0000001" when "00101111001110100", -- t[24180] = 1
      "0000001" when "00101111001110101", -- t[24181] = 1
      "0000001" when "00101111001110110", -- t[24182] = 1
      "0000001" when "00101111001110111", -- t[24183] = 1
      "0000001" when "00101111001111000", -- t[24184] = 1
      "0000001" when "00101111001111001", -- t[24185] = 1
      "0000001" when "00101111001111010", -- t[24186] = 1
      "0000001" when "00101111001111011", -- t[24187] = 1
      "0000001" when "00101111001111100", -- t[24188] = 1
      "0000001" when "00101111001111101", -- t[24189] = 1
      "0000001" when "00101111001111110", -- t[24190] = 1
      "0000001" when "00101111001111111", -- t[24191] = 1
      "0000001" when "00101111010000000", -- t[24192] = 1
      "0000001" when "00101111010000001", -- t[24193] = 1
      "0000001" when "00101111010000010", -- t[24194] = 1
      "0000001" when "00101111010000011", -- t[24195] = 1
      "0000001" when "00101111010000100", -- t[24196] = 1
      "0000001" when "00101111010000101", -- t[24197] = 1
      "0000001" when "00101111010000110", -- t[24198] = 1
      "0000001" when "00101111010000111", -- t[24199] = 1
      "0000001" when "00101111010001000", -- t[24200] = 1
      "0000001" when "00101111010001001", -- t[24201] = 1
      "0000001" when "00101111010001010", -- t[24202] = 1
      "0000001" when "00101111010001011", -- t[24203] = 1
      "0000001" when "00101111010001100", -- t[24204] = 1
      "0000001" when "00101111010001101", -- t[24205] = 1
      "0000001" when "00101111010001110", -- t[24206] = 1
      "0000001" when "00101111010001111", -- t[24207] = 1
      "0000001" when "00101111010010000", -- t[24208] = 1
      "0000001" when "00101111010010001", -- t[24209] = 1
      "0000001" when "00101111010010010", -- t[24210] = 1
      "0000001" when "00101111010010011", -- t[24211] = 1
      "0000001" when "00101111010010100", -- t[24212] = 1
      "0000001" when "00101111010010101", -- t[24213] = 1
      "0000001" when "00101111010010110", -- t[24214] = 1
      "0000001" when "00101111010010111", -- t[24215] = 1
      "0000001" when "00101111010011000", -- t[24216] = 1
      "0000001" when "00101111010011001", -- t[24217] = 1
      "0000001" when "00101111010011010", -- t[24218] = 1
      "0000001" when "00101111010011011", -- t[24219] = 1
      "0000001" when "00101111010011100", -- t[24220] = 1
      "0000001" when "00101111010011101", -- t[24221] = 1
      "0000001" when "00101111010011110", -- t[24222] = 1
      "0000001" when "00101111010011111", -- t[24223] = 1
      "0000001" when "00101111010100000", -- t[24224] = 1
      "0000001" when "00101111010100001", -- t[24225] = 1
      "0000001" when "00101111010100010", -- t[24226] = 1
      "0000001" when "00101111010100011", -- t[24227] = 1
      "0000001" when "00101111010100100", -- t[24228] = 1
      "0000001" when "00101111010100101", -- t[24229] = 1
      "0000001" when "00101111010100110", -- t[24230] = 1
      "0000001" when "00101111010100111", -- t[24231] = 1
      "0000001" when "00101111010101000", -- t[24232] = 1
      "0000001" when "00101111010101001", -- t[24233] = 1
      "0000001" when "00101111010101010", -- t[24234] = 1
      "0000001" when "00101111010101011", -- t[24235] = 1
      "0000001" when "00101111010101100", -- t[24236] = 1
      "0000001" when "00101111010101101", -- t[24237] = 1
      "0000001" when "00101111010101110", -- t[24238] = 1
      "0000001" when "00101111010101111", -- t[24239] = 1
      "0000001" when "00101111010110000", -- t[24240] = 1
      "0000001" when "00101111010110001", -- t[24241] = 1
      "0000001" when "00101111010110010", -- t[24242] = 1
      "0000001" when "00101111010110011", -- t[24243] = 1
      "0000001" when "00101111010110100", -- t[24244] = 1
      "0000001" when "00101111010110101", -- t[24245] = 1
      "0000001" when "00101111010110110", -- t[24246] = 1
      "0000001" when "00101111010110111", -- t[24247] = 1
      "0000001" when "00101111010111000", -- t[24248] = 1
      "0000001" when "00101111010111001", -- t[24249] = 1
      "0000001" when "00101111010111010", -- t[24250] = 1
      "0000001" when "00101111010111011", -- t[24251] = 1
      "0000001" when "00101111010111100", -- t[24252] = 1
      "0000001" when "00101111010111101", -- t[24253] = 1
      "0000001" when "00101111010111110", -- t[24254] = 1
      "0000001" when "00101111010111111", -- t[24255] = 1
      "0000001" when "00101111011000000", -- t[24256] = 1
      "0000001" when "00101111011000001", -- t[24257] = 1
      "0000001" when "00101111011000010", -- t[24258] = 1
      "0000001" when "00101111011000011", -- t[24259] = 1
      "0000001" when "00101111011000100", -- t[24260] = 1
      "0000001" when "00101111011000101", -- t[24261] = 1
      "0000001" when "00101111011000110", -- t[24262] = 1
      "0000001" when "00101111011000111", -- t[24263] = 1
      "0000001" when "00101111011001000", -- t[24264] = 1
      "0000001" when "00101111011001001", -- t[24265] = 1
      "0000001" when "00101111011001010", -- t[24266] = 1
      "0000001" when "00101111011001011", -- t[24267] = 1
      "0000001" when "00101111011001100", -- t[24268] = 1
      "0000001" when "00101111011001101", -- t[24269] = 1
      "0000001" when "00101111011001110", -- t[24270] = 1
      "0000001" when "00101111011001111", -- t[24271] = 1
      "0000001" when "00101111011010000", -- t[24272] = 1
      "0000001" when "00101111011010001", -- t[24273] = 1
      "0000001" when "00101111011010010", -- t[24274] = 1
      "0000001" when "00101111011010011", -- t[24275] = 1
      "0000001" when "00101111011010100", -- t[24276] = 1
      "0000001" when "00101111011010101", -- t[24277] = 1
      "0000001" when "00101111011010110", -- t[24278] = 1
      "0000001" when "00101111011010111", -- t[24279] = 1
      "0000001" when "00101111011011000", -- t[24280] = 1
      "0000001" when "00101111011011001", -- t[24281] = 1
      "0000001" when "00101111011011010", -- t[24282] = 1
      "0000001" when "00101111011011011", -- t[24283] = 1
      "0000001" when "00101111011011100", -- t[24284] = 1
      "0000001" when "00101111011011101", -- t[24285] = 1
      "0000001" when "00101111011011110", -- t[24286] = 1
      "0000001" when "00101111011011111", -- t[24287] = 1
      "0000001" when "00101111011100000", -- t[24288] = 1
      "0000001" when "00101111011100001", -- t[24289] = 1
      "0000001" when "00101111011100010", -- t[24290] = 1
      "0000001" when "00101111011100011", -- t[24291] = 1
      "0000001" when "00101111011100100", -- t[24292] = 1
      "0000001" when "00101111011100101", -- t[24293] = 1
      "0000001" when "00101111011100110", -- t[24294] = 1
      "0000001" when "00101111011100111", -- t[24295] = 1
      "0000001" when "00101111011101000", -- t[24296] = 1
      "0000001" when "00101111011101001", -- t[24297] = 1
      "0000001" when "00101111011101010", -- t[24298] = 1
      "0000001" when "00101111011101011", -- t[24299] = 1
      "0000001" when "00101111011101100", -- t[24300] = 1
      "0000001" when "00101111011101101", -- t[24301] = 1
      "0000001" when "00101111011101110", -- t[24302] = 1
      "0000001" when "00101111011101111", -- t[24303] = 1
      "0000001" when "00101111011110000", -- t[24304] = 1
      "0000001" when "00101111011110001", -- t[24305] = 1
      "0000001" when "00101111011110010", -- t[24306] = 1
      "0000001" when "00101111011110011", -- t[24307] = 1
      "0000001" when "00101111011110100", -- t[24308] = 1
      "0000001" when "00101111011110101", -- t[24309] = 1
      "0000001" when "00101111011110110", -- t[24310] = 1
      "0000001" when "00101111011110111", -- t[24311] = 1
      "0000001" when "00101111011111000", -- t[24312] = 1
      "0000001" when "00101111011111001", -- t[24313] = 1
      "0000001" when "00101111011111010", -- t[24314] = 1
      "0000001" when "00101111011111011", -- t[24315] = 1
      "0000001" when "00101111011111100", -- t[24316] = 1
      "0000001" when "00101111011111101", -- t[24317] = 1
      "0000001" when "00101111011111110", -- t[24318] = 1
      "0000001" when "00101111011111111", -- t[24319] = 1
      "0000001" when "00101111100000000", -- t[24320] = 1
      "0000001" when "00101111100000001", -- t[24321] = 1
      "0000001" when "00101111100000010", -- t[24322] = 1
      "0000001" when "00101111100000011", -- t[24323] = 1
      "0000001" when "00101111100000100", -- t[24324] = 1
      "0000001" when "00101111100000101", -- t[24325] = 1
      "0000001" when "00101111100000110", -- t[24326] = 1
      "0000001" when "00101111100000111", -- t[24327] = 1
      "0000001" when "00101111100001000", -- t[24328] = 1
      "0000001" when "00101111100001001", -- t[24329] = 1
      "0000001" when "00101111100001010", -- t[24330] = 1
      "0000001" when "00101111100001011", -- t[24331] = 1
      "0000001" when "00101111100001100", -- t[24332] = 1
      "0000001" when "00101111100001101", -- t[24333] = 1
      "0000001" when "00101111100001110", -- t[24334] = 1
      "0000001" when "00101111100001111", -- t[24335] = 1
      "0000001" when "00101111100010000", -- t[24336] = 1
      "0000001" when "00101111100010001", -- t[24337] = 1
      "0000001" when "00101111100010010", -- t[24338] = 1
      "0000001" when "00101111100010011", -- t[24339] = 1
      "0000001" when "00101111100010100", -- t[24340] = 1
      "0000001" when "00101111100010101", -- t[24341] = 1
      "0000001" when "00101111100010110", -- t[24342] = 1
      "0000001" when "00101111100010111", -- t[24343] = 1
      "0000001" when "00101111100011000", -- t[24344] = 1
      "0000001" when "00101111100011001", -- t[24345] = 1
      "0000001" when "00101111100011010", -- t[24346] = 1
      "0000001" when "00101111100011011", -- t[24347] = 1
      "0000001" when "00101111100011100", -- t[24348] = 1
      "0000001" when "00101111100011101", -- t[24349] = 1
      "0000001" when "00101111100011110", -- t[24350] = 1
      "0000001" when "00101111100011111", -- t[24351] = 1
      "0000001" when "00101111100100000", -- t[24352] = 1
      "0000001" when "00101111100100001", -- t[24353] = 1
      "0000001" when "00101111100100010", -- t[24354] = 1
      "0000001" when "00101111100100011", -- t[24355] = 1
      "0000001" when "00101111100100100", -- t[24356] = 1
      "0000001" when "00101111100100101", -- t[24357] = 1
      "0000001" when "00101111100100110", -- t[24358] = 1
      "0000001" when "00101111100100111", -- t[24359] = 1
      "0000001" when "00101111100101000", -- t[24360] = 1
      "0000001" when "00101111100101001", -- t[24361] = 1
      "0000001" when "00101111100101010", -- t[24362] = 1
      "0000001" when "00101111100101011", -- t[24363] = 1
      "0000001" when "00101111100101100", -- t[24364] = 1
      "0000001" when "00101111100101101", -- t[24365] = 1
      "0000001" when "00101111100101110", -- t[24366] = 1
      "0000001" when "00101111100101111", -- t[24367] = 1
      "0000001" when "00101111100110000", -- t[24368] = 1
      "0000001" when "00101111100110001", -- t[24369] = 1
      "0000001" when "00101111100110010", -- t[24370] = 1
      "0000001" when "00101111100110011", -- t[24371] = 1
      "0000001" when "00101111100110100", -- t[24372] = 1
      "0000001" when "00101111100110101", -- t[24373] = 1
      "0000001" when "00101111100110110", -- t[24374] = 1
      "0000001" when "00101111100110111", -- t[24375] = 1
      "0000001" when "00101111100111000", -- t[24376] = 1
      "0000001" when "00101111100111001", -- t[24377] = 1
      "0000001" when "00101111100111010", -- t[24378] = 1
      "0000001" when "00101111100111011", -- t[24379] = 1
      "0000001" when "00101111100111100", -- t[24380] = 1
      "0000001" when "00101111100111101", -- t[24381] = 1
      "0000001" when "00101111100111110", -- t[24382] = 1
      "0000001" when "00101111100111111", -- t[24383] = 1
      "0000001" when "00101111101000000", -- t[24384] = 1
      "0000001" when "00101111101000001", -- t[24385] = 1
      "0000001" when "00101111101000010", -- t[24386] = 1
      "0000001" when "00101111101000011", -- t[24387] = 1
      "0000001" when "00101111101000100", -- t[24388] = 1
      "0000001" when "00101111101000101", -- t[24389] = 1
      "0000001" when "00101111101000110", -- t[24390] = 1
      "0000001" when "00101111101000111", -- t[24391] = 1
      "0000001" when "00101111101001000", -- t[24392] = 1
      "0000001" when "00101111101001001", -- t[24393] = 1
      "0000001" when "00101111101001010", -- t[24394] = 1
      "0000001" when "00101111101001011", -- t[24395] = 1
      "0000001" when "00101111101001100", -- t[24396] = 1
      "0000001" when "00101111101001101", -- t[24397] = 1
      "0000001" when "00101111101001110", -- t[24398] = 1
      "0000001" when "00101111101001111", -- t[24399] = 1
      "0000001" when "00101111101010000", -- t[24400] = 1
      "0000001" when "00101111101010001", -- t[24401] = 1
      "0000001" when "00101111101010010", -- t[24402] = 1
      "0000001" when "00101111101010011", -- t[24403] = 1
      "0000001" when "00101111101010100", -- t[24404] = 1
      "0000001" when "00101111101010101", -- t[24405] = 1
      "0000001" when "00101111101010110", -- t[24406] = 1
      "0000001" when "00101111101010111", -- t[24407] = 1
      "0000001" when "00101111101011000", -- t[24408] = 1
      "0000001" when "00101111101011001", -- t[24409] = 1
      "0000001" when "00101111101011010", -- t[24410] = 1
      "0000001" when "00101111101011011", -- t[24411] = 1
      "0000001" when "00101111101011100", -- t[24412] = 1
      "0000001" when "00101111101011101", -- t[24413] = 1
      "0000001" when "00101111101011110", -- t[24414] = 1
      "0000001" when "00101111101011111", -- t[24415] = 1
      "0000001" when "00101111101100000", -- t[24416] = 1
      "0000001" when "00101111101100001", -- t[24417] = 1
      "0000001" when "00101111101100010", -- t[24418] = 1
      "0000001" when "00101111101100011", -- t[24419] = 1
      "0000001" when "00101111101100100", -- t[24420] = 1
      "0000001" when "00101111101100101", -- t[24421] = 1
      "0000001" when "00101111101100110", -- t[24422] = 1
      "0000001" when "00101111101100111", -- t[24423] = 1
      "0000001" when "00101111101101000", -- t[24424] = 1
      "0000001" when "00101111101101001", -- t[24425] = 1
      "0000001" when "00101111101101010", -- t[24426] = 1
      "0000001" when "00101111101101011", -- t[24427] = 1
      "0000001" when "00101111101101100", -- t[24428] = 1
      "0000001" when "00101111101101101", -- t[24429] = 1
      "0000001" when "00101111101101110", -- t[24430] = 1
      "0000001" when "00101111101101111", -- t[24431] = 1
      "0000001" when "00101111101110000", -- t[24432] = 1
      "0000001" when "00101111101110001", -- t[24433] = 1
      "0000001" when "00101111101110010", -- t[24434] = 1
      "0000001" when "00101111101110011", -- t[24435] = 1
      "0000001" when "00101111101110100", -- t[24436] = 1
      "0000001" when "00101111101110101", -- t[24437] = 1
      "0000001" when "00101111101110110", -- t[24438] = 1
      "0000001" when "00101111101110111", -- t[24439] = 1
      "0000001" when "00101111101111000", -- t[24440] = 1
      "0000001" when "00101111101111001", -- t[24441] = 1
      "0000001" when "00101111101111010", -- t[24442] = 1
      "0000001" when "00101111101111011", -- t[24443] = 1
      "0000001" when "00101111101111100", -- t[24444] = 1
      "0000001" when "00101111101111101", -- t[24445] = 1
      "0000001" when "00101111101111110", -- t[24446] = 1
      "0000001" when "00101111101111111", -- t[24447] = 1
      "0000001" when "00101111110000000", -- t[24448] = 1
      "0000001" when "00101111110000001", -- t[24449] = 1
      "0000001" when "00101111110000010", -- t[24450] = 1
      "0000001" when "00101111110000011", -- t[24451] = 1
      "0000001" when "00101111110000100", -- t[24452] = 1
      "0000001" when "00101111110000101", -- t[24453] = 1
      "0000001" when "00101111110000110", -- t[24454] = 1
      "0000001" when "00101111110000111", -- t[24455] = 1
      "0000001" when "00101111110001000", -- t[24456] = 1
      "0000001" when "00101111110001001", -- t[24457] = 1
      "0000001" when "00101111110001010", -- t[24458] = 1
      "0000001" when "00101111110001011", -- t[24459] = 1
      "0000001" when "00101111110001100", -- t[24460] = 1
      "0000001" when "00101111110001101", -- t[24461] = 1
      "0000001" when "00101111110001110", -- t[24462] = 1
      "0000001" when "00101111110001111", -- t[24463] = 1
      "0000001" when "00101111110010000", -- t[24464] = 1
      "0000001" when "00101111110010001", -- t[24465] = 1
      "0000001" when "00101111110010010", -- t[24466] = 1
      "0000001" when "00101111110010011", -- t[24467] = 1
      "0000001" when "00101111110010100", -- t[24468] = 1
      "0000001" when "00101111110010101", -- t[24469] = 1
      "0000001" when "00101111110010110", -- t[24470] = 1
      "0000001" when "00101111110010111", -- t[24471] = 1
      "0000001" when "00101111110011000", -- t[24472] = 1
      "0000001" when "00101111110011001", -- t[24473] = 1
      "0000001" when "00101111110011010", -- t[24474] = 1
      "0000001" when "00101111110011011", -- t[24475] = 1
      "0000001" when "00101111110011100", -- t[24476] = 1
      "0000001" when "00101111110011101", -- t[24477] = 1
      "0000001" when "00101111110011110", -- t[24478] = 1
      "0000001" when "00101111110011111", -- t[24479] = 1
      "0000001" when "00101111110100000", -- t[24480] = 1
      "0000001" when "00101111110100001", -- t[24481] = 1
      "0000001" when "00101111110100010", -- t[24482] = 1
      "0000001" when "00101111110100011", -- t[24483] = 1
      "0000001" when "00101111110100100", -- t[24484] = 1
      "0000001" when "00101111110100101", -- t[24485] = 1
      "0000001" when "00101111110100110", -- t[24486] = 1
      "0000001" when "00101111110100111", -- t[24487] = 1
      "0000001" when "00101111110101000", -- t[24488] = 1
      "0000001" when "00101111110101001", -- t[24489] = 1
      "0000001" when "00101111110101010", -- t[24490] = 1
      "0000001" when "00101111110101011", -- t[24491] = 1
      "0000001" when "00101111110101100", -- t[24492] = 1
      "0000001" when "00101111110101101", -- t[24493] = 1
      "0000001" when "00101111110101110", -- t[24494] = 1
      "0000001" when "00101111110101111", -- t[24495] = 1
      "0000001" when "00101111110110000", -- t[24496] = 1
      "0000001" when "00101111110110001", -- t[24497] = 1
      "0000001" when "00101111110110010", -- t[24498] = 1
      "0000001" when "00101111110110011", -- t[24499] = 1
      "0000001" when "00101111110110100", -- t[24500] = 1
      "0000001" when "00101111110110101", -- t[24501] = 1
      "0000001" when "00101111110110110", -- t[24502] = 1
      "0000001" when "00101111110110111", -- t[24503] = 1
      "0000001" when "00101111110111000", -- t[24504] = 1
      "0000001" when "00101111110111001", -- t[24505] = 1
      "0000001" when "00101111110111010", -- t[24506] = 1
      "0000001" when "00101111110111011", -- t[24507] = 1
      "0000001" when "00101111110111100", -- t[24508] = 1
      "0000001" when "00101111110111101", -- t[24509] = 1
      "0000001" when "00101111110111110", -- t[24510] = 1
      "0000001" when "00101111110111111", -- t[24511] = 1
      "0000001" when "00101111111000000", -- t[24512] = 1
      "0000001" when "00101111111000001", -- t[24513] = 1
      "0000001" when "00101111111000010", -- t[24514] = 1
      "0000001" when "00101111111000011", -- t[24515] = 1
      "0000001" when "00101111111000100", -- t[24516] = 1
      "0000001" when "00101111111000101", -- t[24517] = 1
      "0000001" when "00101111111000110", -- t[24518] = 1
      "0000001" when "00101111111000111", -- t[24519] = 1
      "0000001" when "00101111111001000", -- t[24520] = 1
      "0000001" when "00101111111001001", -- t[24521] = 1
      "0000001" when "00101111111001010", -- t[24522] = 1
      "0000001" when "00101111111001011", -- t[24523] = 1
      "0000001" when "00101111111001100", -- t[24524] = 1
      "0000001" when "00101111111001101", -- t[24525] = 1
      "0000001" when "00101111111001110", -- t[24526] = 1
      "0000001" when "00101111111001111", -- t[24527] = 1
      "0000001" when "00101111111010000", -- t[24528] = 1
      "0000001" when "00101111111010001", -- t[24529] = 1
      "0000001" when "00101111111010010", -- t[24530] = 1
      "0000001" when "00101111111010011", -- t[24531] = 1
      "0000001" when "00101111111010100", -- t[24532] = 1
      "0000001" when "00101111111010101", -- t[24533] = 1
      "0000001" when "00101111111010110", -- t[24534] = 1
      "0000001" when "00101111111010111", -- t[24535] = 1
      "0000001" when "00101111111011000", -- t[24536] = 1
      "0000001" when "00101111111011001", -- t[24537] = 1
      "0000001" when "00101111111011010", -- t[24538] = 1
      "0000001" when "00101111111011011", -- t[24539] = 1
      "0000001" when "00101111111011100", -- t[24540] = 1
      "0000001" when "00101111111011101", -- t[24541] = 1
      "0000001" when "00101111111011110", -- t[24542] = 1
      "0000001" when "00101111111011111", -- t[24543] = 1
      "0000001" when "00101111111100000", -- t[24544] = 1
      "0000001" when "00101111111100001", -- t[24545] = 1
      "0000001" when "00101111111100010", -- t[24546] = 1
      "0000001" when "00101111111100011", -- t[24547] = 1
      "0000001" when "00101111111100100", -- t[24548] = 1
      "0000001" when "00101111111100101", -- t[24549] = 1
      "0000001" when "00101111111100110", -- t[24550] = 1
      "0000001" when "00101111111100111", -- t[24551] = 1
      "0000001" when "00101111111101000", -- t[24552] = 1
      "0000001" when "00101111111101001", -- t[24553] = 1
      "0000001" when "00101111111101010", -- t[24554] = 1
      "0000001" when "00101111111101011", -- t[24555] = 1
      "0000001" when "00101111111101100", -- t[24556] = 1
      "0000001" when "00101111111101101", -- t[24557] = 1
      "0000001" when "00101111111101110", -- t[24558] = 1
      "0000001" when "00101111111101111", -- t[24559] = 1
      "0000001" when "00101111111110000", -- t[24560] = 1
      "0000001" when "00101111111110001", -- t[24561] = 1
      "0000001" when "00101111111110010", -- t[24562] = 1
      "0000001" when "00101111111110011", -- t[24563] = 1
      "0000001" when "00101111111110100", -- t[24564] = 1
      "0000001" when "00101111111110101", -- t[24565] = 1
      "0000001" when "00101111111110110", -- t[24566] = 1
      "0000001" when "00101111111110111", -- t[24567] = 1
      "0000001" when "00101111111111000", -- t[24568] = 1
      "0000001" when "00101111111111001", -- t[24569] = 1
      "0000001" when "00101111111111010", -- t[24570] = 1
      "0000001" when "00101111111111011", -- t[24571] = 1
      "0000001" when "00101111111111100", -- t[24572] = 1
      "0000001" when "00101111111111101", -- t[24573] = 1
      "0000001" when "00101111111111110", -- t[24574] = 1
      "0000001" when "00101111111111111", -- t[24575] = 1
      "0000001" when "00110000000000000", -- t[24576] = 1
      "0000001" when "00110000000000001", -- t[24577] = 1
      "0000001" when "00110000000000010", -- t[24578] = 1
      "0000001" when "00110000000000011", -- t[24579] = 1
      "0000001" when "00110000000000100", -- t[24580] = 1
      "0000001" when "00110000000000101", -- t[24581] = 1
      "0000001" when "00110000000000110", -- t[24582] = 1
      "0000001" when "00110000000000111", -- t[24583] = 1
      "0000001" when "00110000000001000", -- t[24584] = 1
      "0000001" when "00110000000001001", -- t[24585] = 1
      "0000001" when "00110000000001010", -- t[24586] = 1
      "0000001" when "00110000000001011", -- t[24587] = 1
      "0000001" when "00110000000001100", -- t[24588] = 1
      "0000001" when "00110000000001101", -- t[24589] = 1
      "0000001" when "00110000000001110", -- t[24590] = 1
      "0000001" when "00110000000001111", -- t[24591] = 1
      "0000001" when "00110000000010000", -- t[24592] = 1
      "0000001" when "00110000000010001", -- t[24593] = 1
      "0000001" when "00110000000010010", -- t[24594] = 1
      "0000001" when "00110000000010011", -- t[24595] = 1
      "0000001" when "00110000000010100", -- t[24596] = 1
      "0000001" when "00110000000010101", -- t[24597] = 1
      "0000001" when "00110000000010110", -- t[24598] = 1
      "0000001" when "00110000000010111", -- t[24599] = 1
      "0000001" when "00110000000011000", -- t[24600] = 1
      "0000001" when "00110000000011001", -- t[24601] = 1
      "0000001" when "00110000000011010", -- t[24602] = 1
      "0000001" when "00110000000011011", -- t[24603] = 1
      "0000001" when "00110000000011100", -- t[24604] = 1
      "0000001" when "00110000000011101", -- t[24605] = 1
      "0000001" when "00110000000011110", -- t[24606] = 1
      "0000001" when "00110000000011111", -- t[24607] = 1
      "0000001" when "00110000000100000", -- t[24608] = 1
      "0000001" when "00110000000100001", -- t[24609] = 1
      "0000001" when "00110000000100010", -- t[24610] = 1
      "0000001" when "00110000000100011", -- t[24611] = 1
      "0000001" when "00110000000100100", -- t[24612] = 1
      "0000001" when "00110000000100101", -- t[24613] = 1
      "0000001" when "00110000000100110", -- t[24614] = 1
      "0000001" when "00110000000100111", -- t[24615] = 1
      "0000001" when "00110000000101000", -- t[24616] = 1
      "0000001" when "00110000000101001", -- t[24617] = 1
      "0000001" when "00110000000101010", -- t[24618] = 1
      "0000001" when "00110000000101011", -- t[24619] = 1
      "0000001" when "00110000000101100", -- t[24620] = 1
      "0000001" when "00110000000101101", -- t[24621] = 1
      "0000001" when "00110000000101110", -- t[24622] = 1
      "0000001" when "00110000000101111", -- t[24623] = 1
      "0000001" when "00110000000110000", -- t[24624] = 1
      "0000001" when "00110000000110001", -- t[24625] = 1
      "0000001" when "00110000000110010", -- t[24626] = 1
      "0000001" when "00110000000110011", -- t[24627] = 1
      "0000001" when "00110000000110100", -- t[24628] = 1
      "0000001" when "00110000000110101", -- t[24629] = 1
      "0000001" when "00110000000110110", -- t[24630] = 1
      "0000001" when "00110000000110111", -- t[24631] = 1
      "0000001" when "00110000000111000", -- t[24632] = 1
      "0000001" when "00110000000111001", -- t[24633] = 1
      "0000001" when "00110000000111010", -- t[24634] = 1
      "0000001" when "00110000000111011", -- t[24635] = 1
      "0000001" when "00110000000111100", -- t[24636] = 1
      "0000001" when "00110000000111101", -- t[24637] = 1
      "0000001" when "00110000000111110", -- t[24638] = 1
      "0000001" when "00110000000111111", -- t[24639] = 1
      "0000001" when "00110000001000000", -- t[24640] = 1
      "0000001" when "00110000001000001", -- t[24641] = 1
      "0000001" when "00110000001000010", -- t[24642] = 1
      "0000001" when "00110000001000011", -- t[24643] = 1
      "0000001" when "00110000001000100", -- t[24644] = 1
      "0000001" when "00110000001000101", -- t[24645] = 1
      "0000001" when "00110000001000110", -- t[24646] = 1
      "0000001" when "00110000001000111", -- t[24647] = 1
      "0000001" when "00110000001001000", -- t[24648] = 1
      "0000001" when "00110000001001001", -- t[24649] = 1
      "0000001" when "00110000001001010", -- t[24650] = 1
      "0000001" when "00110000001001011", -- t[24651] = 1
      "0000001" when "00110000001001100", -- t[24652] = 1
      "0000001" when "00110000001001101", -- t[24653] = 1
      "0000001" when "00110000001001110", -- t[24654] = 1
      "0000001" when "00110000001001111", -- t[24655] = 1
      "0000001" when "00110000001010000", -- t[24656] = 1
      "0000001" when "00110000001010001", -- t[24657] = 1
      "0000001" when "00110000001010010", -- t[24658] = 1
      "0000001" when "00110000001010011", -- t[24659] = 1
      "0000001" when "00110000001010100", -- t[24660] = 1
      "0000001" when "00110000001010101", -- t[24661] = 1
      "0000001" when "00110000001010110", -- t[24662] = 1
      "0000001" when "00110000001010111", -- t[24663] = 1
      "0000001" when "00110000001011000", -- t[24664] = 1
      "0000001" when "00110000001011001", -- t[24665] = 1
      "0000001" when "00110000001011010", -- t[24666] = 1
      "0000001" when "00110000001011011", -- t[24667] = 1
      "0000001" when "00110000001011100", -- t[24668] = 1
      "0000001" when "00110000001011101", -- t[24669] = 1
      "0000001" when "00110000001011110", -- t[24670] = 1
      "0000001" when "00110000001011111", -- t[24671] = 1
      "0000001" when "00110000001100000", -- t[24672] = 1
      "0000001" when "00110000001100001", -- t[24673] = 1
      "0000001" when "00110000001100010", -- t[24674] = 1
      "0000001" when "00110000001100011", -- t[24675] = 1
      "0000001" when "00110000001100100", -- t[24676] = 1
      "0000001" when "00110000001100101", -- t[24677] = 1
      "0000001" when "00110000001100110", -- t[24678] = 1
      "0000001" when "00110000001100111", -- t[24679] = 1
      "0000001" when "00110000001101000", -- t[24680] = 1
      "0000001" when "00110000001101001", -- t[24681] = 1
      "0000001" when "00110000001101010", -- t[24682] = 1
      "0000001" when "00110000001101011", -- t[24683] = 1
      "0000001" when "00110000001101100", -- t[24684] = 1
      "0000001" when "00110000001101101", -- t[24685] = 1
      "0000001" when "00110000001101110", -- t[24686] = 1
      "0000001" when "00110000001101111", -- t[24687] = 1
      "0000001" when "00110000001110000", -- t[24688] = 1
      "0000001" when "00110000001110001", -- t[24689] = 1
      "0000001" when "00110000001110010", -- t[24690] = 1
      "0000001" when "00110000001110011", -- t[24691] = 1
      "0000001" when "00110000001110100", -- t[24692] = 1
      "0000001" when "00110000001110101", -- t[24693] = 1
      "0000001" when "00110000001110110", -- t[24694] = 1
      "0000001" when "00110000001110111", -- t[24695] = 1
      "0000001" when "00110000001111000", -- t[24696] = 1
      "0000001" when "00110000001111001", -- t[24697] = 1
      "0000001" when "00110000001111010", -- t[24698] = 1
      "0000001" when "00110000001111011", -- t[24699] = 1
      "0000001" when "00110000001111100", -- t[24700] = 1
      "0000001" when "00110000001111101", -- t[24701] = 1
      "0000001" when "00110000001111110", -- t[24702] = 1
      "0000001" when "00110000001111111", -- t[24703] = 1
      "0000001" when "00110000010000000", -- t[24704] = 1
      "0000001" when "00110000010000001", -- t[24705] = 1
      "0000001" when "00110000010000010", -- t[24706] = 1
      "0000001" when "00110000010000011", -- t[24707] = 1
      "0000001" when "00110000010000100", -- t[24708] = 1
      "0000001" when "00110000010000101", -- t[24709] = 1
      "0000001" when "00110000010000110", -- t[24710] = 1
      "0000001" when "00110000010000111", -- t[24711] = 1
      "0000001" when "00110000010001000", -- t[24712] = 1
      "0000001" when "00110000010001001", -- t[24713] = 1
      "0000001" when "00110000010001010", -- t[24714] = 1
      "0000001" when "00110000010001011", -- t[24715] = 1
      "0000001" when "00110000010001100", -- t[24716] = 1
      "0000001" when "00110000010001101", -- t[24717] = 1
      "0000001" when "00110000010001110", -- t[24718] = 1
      "0000001" when "00110000010001111", -- t[24719] = 1
      "0000001" when "00110000010010000", -- t[24720] = 1
      "0000001" when "00110000010010001", -- t[24721] = 1
      "0000001" when "00110000010010010", -- t[24722] = 1
      "0000001" when "00110000010010011", -- t[24723] = 1
      "0000001" when "00110000010010100", -- t[24724] = 1
      "0000001" when "00110000010010101", -- t[24725] = 1
      "0000001" when "00110000010010110", -- t[24726] = 1
      "0000001" when "00110000010010111", -- t[24727] = 1
      "0000001" when "00110000010011000", -- t[24728] = 1
      "0000001" when "00110000010011001", -- t[24729] = 1
      "0000001" when "00110000010011010", -- t[24730] = 1
      "0000001" when "00110000010011011", -- t[24731] = 1
      "0000001" when "00110000010011100", -- t[24732] = 1
      "0000001" when "00110000010011101", -- t[24733] = 1
      "0000001" when "00110000010011110", -- t[24734] = 1
      "0000001" when "00110000010011111", -- t[24735] = 1
      "0000001" when "00110000010100000", -- t[24736] = 1
      "0000001" when "00110000010100001", -- t[24737] = 1
      "0000001" when "00110000010100010", -- t[24738] = 1
      "0000001" when "00110000010100011", -- t[24739] = 1
      "0000001" when "00110000010100100", -- t[24740] = 1
      "0000001" when "00110000010100101", -- t[24741] = 1
      "0000001" when "00110000010100110", -- t[24742] = 1
      "0000001" when "00110000010100111", -- t[24743] = 1
      "0000001" when "00110000010101000", -- t[24744] = 1
      "0000001" when "00110000010101001", -- t[24745] = 1
      "0000001" when "00110000010101010", -- t[24746] = 1
      "0000001" when "00110000010101011", -- t[24747] = 1
      "0000001" when "00110000010101100", -- t[24748] = 1
      "0000001" when "00110000010101101", -- t[24749] = 1
      "0000001" when "00110000010101110", -- t[24750] = 1
      "0000001" when "00110000010101111", -- t[24751] = 1
      "0000001" when "00110000010110000", -- t[24752] = 1
      "0000001" when "00110000010110001", -- t[24753] = 1
      "0000001" when "00110000010110010", -- t[24754] = 1
      "0000001" when "00110000010110011", -- t[24755] = 1
      "0000001" when "00110000010110100", -- t[24756] = 1
      "0000001" when "00110000010110101", -- t[24757] = 1
      "0000001" when "00110000010110110", -- t[24758] = 1
      "0000001" when "00110000010110111", -- t[24759] = 1
      "0000001" when "00110000010111000", -- t[24760] = 1
      "0000001" when "00110000010111001", -- t[24761] = 1
      "0000001" when "00110000010111010", -- t[24762] = 1
      "0000001" when "00110000010111011", -- t[24763] = 1
      "0000001" when "00110000010111100", -- t[24764] = 1
      "0000001" when "00110000010111101", -- t[24765] = 1
      "0000001" when "00110000010111110", -- t[24766] = 1
      "0000001" when "00110000010111111", -- t[24767] = 1
      "0000001" when "00110000011000000", -- t[24768] = 1
      "0000001" when "00110000011000001", -- t[24769] = 1
      "0000001" when "00110000011000010", -- t[24770] = 1
      "0000001" when "00110000011000011", -- t[24771] = 1
      "0000001" when "00110000011000100", -- t[24772] = 1
      "0000001" when "00110000011000101", -- t[24773] = 1
      "0000001" when "00110000011000110", -- t[24774] = 1
      "0000001" when "00110000011000111", -- t[24775] = 1
      "0000001" when "00110000011001000", -- t[24776] = 1
      "0000001" when "00110000011001001", -- t[24777] = 1
      "0000001" when "00110000011001010", -- t[24778] = 1
      "0000001" when "00110000011001011", -- t[24779] = 1
      "0000001" when "00110000011001100", -- t[24780] = 1
      "0000001" when "00110000011001101", -- t[24781] = 1
      "0000001" when "00110000011001110", -- t[24782] = 1
      "0000001" when "00110000011001111", -- t[24783] = 1
      "0000001" when "00110000011010000", -- t[24784] = 1
      "0000001" when "00110000011010001", -- t[24785] = 1
      "0000001" when "00110000011010010", -- t[24786] = 1
      "0000001" when "00110000011010011", -- t[24787] = 1
      "0000001" when "00110000011010100", -- t[24788] = 1
      "0000001" when "00110000011010101", -- t[24789] = 1
      "0000001" when "00110000011010110", -- t[24790] = 1
      "0000001" when "00110000011010111", -- t[24791] = 1
      "0000001" when "00110000011011000", -- t[24792] = 1
      "0000001" when "00110000011011001", -- t[24793] = 1
      "0000001" when "00110000011011010", -- t[24794] = 1
      "0000001" when "00110000011011011", -- t[24795] = 1
      "0000001" when "00110000011011100", -- t[24796] = 1
      "0000001" when "00110000011011101", -- t[24797] = 1
      "0000001" when "00110000011011110", -- t[24798] = 1
      "0000001" when "00110000011011111", -- t[24799] = 1
      "0000001" when "00110000011100000", -- t[24800] = 1
      "0000001" when "00110000011100001", -- t[24801] = 1
      "0000001" when "00110000011100010", -- t[24802] = 1
      "0000001" when "00110000011100011", -- t[24803] = 1
      "0000001" when "00110000011100100", -- t[24804] = 1
      "0000001" when "00110000011100101", -- t[24805] = 1
      "0000001" when "00110000011100110", -- t[24806] = 1
      "0000001" when "00110000011100111", -- t[24807] = 1
      "0000001" when "00110000011101000", -- t[24808] = 1
      "0000001" when "00110000011101001", -- t[24809] = 1
      "0000001" when "00110000011101010", -- t[24810] = 1
      "0000001" when "00110000011101011", -- t[24811] = 1
      "0000001" when "00110000011101100", -- t[24812] = 1
      "0000001" when "00110000011101101", -- t[24813] = 1
      "0000001" when "00110000011101110", -- t[24814] = 1
      "0000001" when "00110000011101111", -- t[24815] = 1
      "0000001" when "00110000011110000", -- t[24816] = 1
      "0000001" when "00110000011110001", -- t[24817] = 1
      "0000001" when "00110000011110010", -- t[24818] = 1
      "0000001" when "00110000011110011", -- t[24819] = 1
      "0000001" when "00110000011110100", -- t[24820] = 1
      "0000001" when "00110000011110101", -- t[24821] = 1
      "0000001" when "00110000011110110", -- t[24822] = 1
      "0000001" when "00110000011110111", -- t[24823] = 1
      "0000001" when "00110000011111000", -- t[24824] = 1
      "0000001" when "00110000011111001", -- t[24825] = 1
      "0000001" when "00110000011111010", -- t[24826] = 1
      "0000001" when "00110000011111011", -- t[24827] = 1
      "0000001" when "00110000011111100", -- t[24828] = 1
      "0000001" when "00110000011111101", -- t[24829] = 1
      "0000001" when "00110000011111110", -- t[24830] = 1
      "0000001" when "00110000011111111", -- t[24831] = 1
      "0000001" when "00110000100000000", -- t[24832] = 1
      "0000001" when "00110000100000001", -- t[24833] = 1
      "0000001" when "00110000100000010", -- t[24834] = 1
      "0000001" when "00110000100000011", -- t[24835] = 1
      "0000001" when "00110000100000100", -- t[24836] = 1
      "0000001" when "00110000100000101", -- t[24837] = 1
      "0000001" when "00110000100000110", -- t[24838] = 1
      "0000001" when "00110000100000111", -- t[24839] = 1
      "0000001" when "00110000100001000", -- t[24840] = 1
      "0000001" when "00110000100001001", -- t[24841] = 1
      "0000001" when "00110000100001010", -- t[24842] = 1
      "0000001" when "00110000100001011", -- t[24843] = 1
      "0000001" when "00110000100001100", -- t[24844] = 1
      "0000001" when "00110000100001101", -- t[24845] = 1
      "0000001" when "00110000100001110", -- t[24846] = 1
      "0000001" when "00110000100001111", -- t[24847] = 1
      "0000001" when "00110000100010000", -- t[24848] = 1
      "0000001" when "00110000100010001", -- t[24849] = 1
      "0000001" when "00110000100010010", -- t[24850] = 1
      "0000001" when "00110000100010011", -- t[24851] = 1
      "0000001" when "00110000100010100", -- t[24852] = 1
      "0000001" when "00110000100010101", -- t[24853] = 1
      "0000001" when "00110000100010110", -- t[24854] = 1
      "0000001" when "00110000100010111", -- t[24855] = 1
      "0000001" when "00110000100011000", -- t[24856] = 1
      "0000001" when "00110000100011001", -- t[24857] = 1
      "0000001" when "00110000100011010", -- t[24858] = 1
      "0000001" when "00110000100011011", -- t[24859] = 1
      "0000001" when "00110000100011100", -- t[24860] = 1
      "0000001" when "00110000100011101", -- t[24861] = 1
      "0000001" when "00110000100011110", -- t[24862] = 1
      "0000001" when "00110000100011111", -- t[24863] = 1
      "0000001" when "00110000100100000", -- t[24864] = 1
      "0000001" when "00110000100100001", -- t[24865] = 1
      "0000001" when "00110000100100010", -- t[24866] = 1
      "0000001" when "00110000100100011", -- t[24867] = 1
      "0000001" when "00110000100100100", -- t[24868] = 1
      "0000001" when "00110000100100101", -- t[24869] = 1
      "0000001" when "00110000100100110", -- t[24870] = 1
      "0000001" when "00110000100100111", -- t[24871] = 1
      "0000001" when "00110000100101000", -- t[24872] = 1
      "0000001" when "00110000100101001", -- t[24873] = 1
      "0000001" when "00110000100101010", -- t[24874] = 1
      "0000001" when "00110000100101011", -- t[24875] = 1
      "0000001" when "00110000100101100", -- t[24876] = 1
      "0000001" when "00110000100101101", -- t[24877] = 1
      "0000001" when "00110000100101110", -- t[24878] = 1
      "0000001" when "00110000100101111", -- t[24879] = 1
      "0000001" when "00110000100110000", -- t[24880] = 1
      "0000001" when "00110000100110001", -- t[24881] = 1
      "0000001" when "00110000100110010", -- t[24882] = 1
      "0000001" when "00110000100110011", -- t[24883] = 1
      "0000001" when "00110000100110100", -- t[24884] = 1
      "0000001" when "00110000100110101", -- t[24885] = 1
      "0000001" when "00110000100110110", -- t[24886] = 1
      "0000001" when "00110000100110111", -- t[24887] = 1
      "0000001" when "00110000100111000", -- t[24888] = 1
      "0000001" when "00110000100111001", -- t[24889] = 1
      "0000001" when "00110000100111010", -- t[24890] = 1
      "0000001" when "00110000100111011", -- t[24891] = 1
      "0000001" when "00110000100111100", -- t[24892] = 1
      "0000001" when "00110000100111101", -- t[24893] = 1
      "0000001" when "00110000100111110", -- t[24894] = 1
      "0000001" when "00110000100111111", -- t[24895] = 1
      "0000001" when "00110000101000000", -- t[24896] = 1
      "0000001" when "00110000101000001", -- t[24897] = 1
      "0000001" when "00110000101000010", -- t[24898] = 1
      "0000001" when "00110000101000011", -- t[24899] = 1
      "0000001" when "00110000101000100", -- t[24900] = 1
      "0000001" when "00110000101000101", -- t[24901] = 1
      "0000001" when "00110000101000110", -- t[24902] = 1
      "0000001" when "00110000101000111", -- t[24903] = 1
      "0000001" when "00110000101001000", -- t[24904] = 1
      "0000001" when "00110000101001001", -- t[24905] = 1
      "0000001" when "00110000101001010", -- t[24906] = 1
      "0000001" when "00110000101001011", -- t[24907] = 1
      "0000001" when "00110000101001100", -- t[24908] = 1
      "0000001" when "00110000101001101", -- t[24909] = 1
      "0000001" when "00110000101001110", -- t[24910] = 1
      "0000001" when "00110000101001111", -- t[24911] = 1
      "0000001" when "00110000101010000", -- t[24912] = 1
      "0000001" when "00110000101010001", -- t[24913] = 1
      "0000001" when "00110000101010010", -- t[24914] = 1
      "0000001" when "00110000101010011", -- t[24915] = 1
      "0000001" when "00110000101010100", -- t[24916] = 1
      "0000001" when "00110000101010101", -- t[24917] = 1
      "0000001" when "00110000101010110", -- t[24918] = 1
      "0000001" when "00110000101010111", -- t[24919] = 1
      "0000001" when "00110000101011000", -- t[24920] = 1
      "0000001" when "00110000101011001", -- t[24921] = 1
      "0000001" when "00110000101011010", -- t[24922] = 1
      "0000001" when "00110000101011011", -- t[24923] = 1
      "0000001" when "00110000101011100", -- t[24924] = 1
      "0000001" when "00110000101011101", -- t[24925] = 1
      "0000001" when "00110000101011110", -- t[24926] = 1
      "0000001" when "00110000101011111", -- t[24927] = 1
      "0000001" when "00110000101100000", -- t[24928] = 1
      "0000001" when "00110000101100001", -- t[24929] = 1
      "0000001" when "00110000101100010", -- t[24930] = 1
      "0000001" when "00110000101100011", -- t[24931] = 1
      "0000001" when "00110000101100100", -- t[24932] = 1
      "0000001" when "00110000101100101", -- t[24933] = 1
      "0000001" when "00110000101100110", -- t[24934] = 1
      "0000001" when "00110000101100111", -- t[24935] = 1
      "0000001" when "00110000101101000", -- t[24936] = 1
      "0000001" when "00110000101101001", -- t[24937] = 1
      "0000001" when "00110000101101010", -- t[24938] = 1
      "0000001" when "00110000101101011", -- t[24939] = 1
      "0000001" when "00110000101101100", -- t[24940] = 1
      "0000001" when "00110000101101101", -- t[24941] = 1
      "0000001" when "00110000101101110", -- t[24942] = 1
      "0000001" when "00110000101101111", -- t[24943] = 1
      "0000001" when "00110000101110000", -- t[24944] = 1
      "0000001" when "00110000101110001", -- t[24945] = 1
      "0000001" when "00110000101110010", -- t[24946] = 1
      "0000001" when "00110000101110011", -- t[24947] = 1
      "0000001" when "00110000101110100", -- t[24948] = 1
      "0000001" when "00110000101110101", -- t[24949] = 1
      "0000001" when "00110000101110110", -- t[24950] = 1
      "0000001" when "00110000101110111", -- t[24951] = 1
      "0000001" when "00110000101111000", -- t[24952] = 1
      "0000001" when "00110000101111001", -- t[24953] = 1
      "0000001" when "00110000101111010", -- t[24954] = 1
      "0000001" when "00110000101111011", -- t[24955] = 1
      "0000001" when "00110000101111100", -- t[24956] = 1
      "0000001" when "00110000101111101", -- t[24957] = 1
      "0000001" when "00110000101111110", -- t[24958] = 1
      "0000001" when "00110000101111111", -- t[24959] = 1
      "0000001" when "00110000110000000", -- t[24960] = 1
      "0000001" when "00110000110000001", -- t[24961] = 1
      "0000001" when "00110000110000010", -- t[24962] = 1
      "0000001" when "00110000110000011", -- t[24963] = 1
      "0000001" when "00110000110000100", -- t[24964] = 1
      "0000001" when "00110000110000101", -- t[24965] = 1
      "0000001" when "00110000110000110", -- t[24966] = 1
      "0000001" when "00110000110000111", -- t[24967] = 1
      "0000001" when "00110000110001000", -- t[24968] = 1
      "0000001" when "00110000110001001", -- t[24969] = 1
      "0000001" when "00110000110001010", -- t[24970] = 1
      "0000001" when "00110000110001011", -- t[24971] = 1
      "0000001" when "00110000110001100", -- t[24972] = 1
      "0000001" when "00110000110001101", -- t[24973] = 1
      "0000001" when "00110000110001110", -- t[24974] = 1
      "0000001" when "00110000110001111", -- t[24975] = 1
      "0000001" when "00110000110010000", -- t[24976] = 1
      "0000001" when "00110000110010001", -- t[24977] = 1
      "0000001" when "00110000110010010", -- t[24978] = 1
      "0000001" when "00110000110010011", -- t[24979] = 1
      "0000001" when "00110000110010100", -- t[24980] = 1
      "0000001" when "00110000110010101", -- t[24981] = 1
      "0000001" when "00110000110010110", -- t[24982] = 1
      "0000001" when "00110000110010111", -- t[24983] = 1
      "0000001" when "00110000110011000", -- t[24984] = 1
      "0000001" when "00110000110011001", -- t[24985] = 1
      "0000001" when "00110000110011010", -- t[24986] = 1
      "0000001" when "00110000110011011", -- t[24987] = 1
      "0000001" when "00110000110011100", -- t[24988] = 1
      "0000001" when "00110000110011101", -- t[24989] = 1
      "0000001" when "00110000110011110", -- t[24990] = 1
      "0000001" when "00110000110011111", -- t[24991] = 1
      "0000001" when "00110000110100000", -- t[24992] = 1
      "0000001" when "00110000110100001", -- t[24993] = 1
      "0000001" when "00110000110100010", -- t[24994] = 1
      "0000001" when "00110000110100011", -- t[24995] = 1
      "0000001" when "00110000110100100", -- t[24996] = 1
      "0000001" when "00110000110100101", -- t[24997] = 1
      "0000001" when "00110000110100110", -- t[24998] = 1
      "0000001" when "00110000110100111", -- t[24999] = 1
      "0000001" when "00110000110101000", -- t[25000] = 1
      "0000001" when "00110000110101001", -- t[25001] = 1
      "0000001" when "00110000110101010", -- t[25002] = 1
      "0000001" when "00110000110101011", -- t[25003] = 1
      "0000001" when "00110000110101100", -- t[25004] = 1
      "0000001" when "00110000110101101", -- t[25005] = 1
      "0000001" when "00110000110101110", -- t[25006] = 1
      "0000001" when "00110000110101111", -- t[25007] = 1
      "0000001" when "00110000110110000", -- t[25008] = 1
      "0000001" when "00110000110110001", -- t[25009] = 1
      "0000001" when "00110000110110010", -- t[25010] = 1
      "0000001" when "00110000110110011", -- t[25011] = 1
      "0000001" when "00110000110110100", -- t[25012] = 1
      "0000001" when "00110000110110101", -- t[25013] = 1
      "0000001" when "00110000110110110", -- t[25014] = 1
      "0000001" when "00110000110110111", -- t[25015] = 1
      "0000001" when "00110000110111000", -- t[25016] = 1
      "0000001" when "00110000110111001", -- t[25017] = 1
      "0000001" when "00110000110111010", -- t[25018] = 1
      "0000001" when "00110000110111011", -- t[25019] = 1
      "0000001" when "00110000110111100", -- t[25020] = 1
      "0000001" when "00110000110111101", -- t[25021] = 1
      "0000001" when "00110000110111110", -- t[25022] = 1
      "0000001" when "00110000110111111", -- t[25023] = 1
      "0000001" when "00110000111000000", -- t[25024] = 1
      "0000001" when "00110000111000001", -- t[25025] = 1
      "0000001" when "00110000111000010", -- t[25026] = 1
      "0000001" when "00110000111000011", -- t[25027] = 1
      "0000001" when "00110000111000100", -- t[25028] = 1
      "0000001" when "00110000111000101", -- t[25029] = 1
      "0000001" when "00110000111000110", -- t[25030] = 1
      "0000001" when "00110000111000111", -- t[25031] = 1
      "0000001" when "00110000111001000", -- t[25032] = 1
      "0000001" when "00110000111001001", -- t[25033] = 1
      "0000001" when "00110000111001010", -- t[25034] = 1
      "0000001" when "00110000111001011", -- t[25035] = 1
      "0000010" when "00110000111001100", -- t[25036] = 2
      "0000010" when "00110000111001101", -- t[25037] = 2
      "0000010" when "00110000111001110", -- t[25038] = 2
      "0000010" when "00110000111001111", -- t[25039] = 2
      "0000010" when "00110000111010000", -- t[25040] = 2
      "0000010" when "00110000111010001", -- t[25041] = 2
      "0000010" when "00110000111010010", -- t[25042] = 2
      "0000010" when "00110000111010011", -- t[25043] = 2
      "0000010" when "00110000111010100", -- t[25044] = 2
      "0000010" when "00110000111010101", -- t[25045] = 2
      "0000010" when "00110000111010110", -- t[25046] = 2
      "0000010" when "00110000111010111", -- t[25047] = 2
      "0000010" when "00110000111011000", -- t[25048] = 2
      "0000010" when "00110000111011001", -- t[25049] = 2
      "0000010" when "00110000111011010", -- t[25050] = 2
      "0000010" when "00110000111011011", -- t[25051] = 2
      "0000010" when "00110000111011100", -- t[25052] = 2
      "0000010" when "00110000111011101", -- t[25053] = 2
      "0000010" when "00110000111011110", -- t[25054] = 2
      "0000010" when "00110000111011111", -- t[25055] = 2
      "0000010" when "00110000111100000", -- t[25056] = 2
      "0000010" when "00110000111100001", -- t[25057] = 2
      "0000010" when "00110000111100010", -- t[25058] = 2
      "0000010" when "00110000111100011", -- t[25059] = 2
      "0000010" when "00110000111100100", -- t[25060] = 2
      "0000010" when "00110000111100101", -- t[25061] = 2
      "0000010" when "00110000111100110", -- t[25062] = 2
      "0000010" when "00110000111100111", -- t[25063] = 2
      "0000010" when "00110000111101000", -- t[25064] = 2
      "0000010" when "00110000111101001", -- t[25065] = 2
      "0000010" when "00110000111101010", -- t[25066] = 2
      "0000010" when "00110000111101011", -- t[25067] = 2
      "0000010" when "00110000111101100", -- t[25068] = 2
      "0000010" when "00110000111101101", -- t[25069] = 2
      "0000010" when "00110000111101110", -- t[25070] = 2
      "0000010" when "00110000111101111", -- t[25071] = 2
      "0000010" when "00110000111110000", -- t[25072] = 2
      "0000010" when "00110000111110001", -- t[25073] = 2
      "0000010" when "00110000111110010", -- t[25074] = 2
      "0000010" when "00110000111110011", -- t[25075] = 2
      "0000010" when "00110000111110100", -- t[25076] = 2
      "0000010" when "00110000111110101", -- t[25077] = 2
      "0000010" when "00110000111110110", -- t[25078] = 2
      "0000010" when "00110000111110111", -- t[25079] = 2
      "0000010" when "00110000111111000", -- t[25080] = 2
      "0000010" when "00110000111111001", -- t[25081] = 2
      "0000010" when "00110000111111010", -- t[25082] = 2
      "0000010" when "00110000111111011", -- t[25083] = 2
      "0000010" when "00110000111111100", -- t[25084] = 2
      "0000010" when "00110000111111101", -- t[25085] = 2
      "0000010" when "00110000111111110", -- t[25086] = 2
      "0000010" when "00110000111111111", -- t[25087] = 2
      "0000010" when "00110001000000000", -- t[25088] = 2
      "0000010" when "00110001000000001", -- t[25089] = 2
      "0000010" when "00110001000000010", -- t[25090] = 2
      "0000010" when "00110001000000011", -- t[25091] = 2
      "0000010" when "00110001000000100", -- t[25092] = 2
      "0000010" when "00110001000000101", -- t[25093] = 2
      "0000010" when "00110001000000110", -- t[25094] = 2
      "0000010" when "00110001000000111", -- t[25095] = 2
      "0000010" when "00110001000001000", -- t[25096] = 2
      "0000010" when "00110001000001001", -- t[25097] = 2
      "0000010" when "00110001000001010", -- t[25098] = 2
      "0000010" when "00110001000001011", -- t[25099] = 2
      "0000010" when "00110001000001100", -- t[25100] = 2
      "0000010" when "00110001000001101", -- t[25101] = 2
      "0000010" when "00110001000001110", -- t[25102] = 2
      "0000010" when "00110001000001111", -- t[25103] = 2
      "0000010" when "00110001000010000", -- t[25104] = 2
      "0000010" when "00110001000010001", -- t[25105] = 2
      "0000010" when "00110001000010010", -- t[25106] = 2
      "0000010" when "00110001000010011", -- t[25107] = 2
      "0000010" when "00110001000010100", -- t[25108] = 2
      "0000010" when "00110001000010101", -- t[25109] = 2
      "0000010" when "00110001000010110", -- t[25110] = 2
      "0000010" when "00110001000010111", -- t[25111] = 2
      "0000010" when "00110001000011000", -- t[25112] = 2
      "0000010" when "00110001000011001", -- t[25113] = 2
      "0000010" when "00110001000011010", -- t[25114] = 2
      "0000010" when "00110001000011011", -- t[25115] = 2
      "0000010" when "00110001000011100", -- t[25116] = 2
      "0000010" when "00110001000011101", -- t[25117] = 2
      "0000010" when "00110001000011110", -- t[25118] = 2
      "0000010" when "00110001000011111", -- t[25119] = 2
      "0000010" when "00110001000100000", -- t[25120] = 2
      "0000010" when "00110001000100001", -- t[25121] = 2
      "0000010" when "00110001000100010", -- t[25122] = 2
      "0000010" when "00110001000100011", -- t[25123] = 2
      "0000010" when "00110001000100100", -- t[25124] = 2
      "0000010" when "00110001000100101", -- t[25125] = 2
      "0000010" when "00110001000100110", -- t[25126] = 2
      "0000010" when "00110001000100111", -- t[25127] = 2
      "0000010" when "00110001000101000", -- t[25128] = 2
      "0000010" when "00110001000101001", -- t[25129] = 2
      "0000010" when "00110001000101010", -- t[25130] = 2
      "0000010" when "00110001000101011", -- t[25131] = 2
      "0000010" when "00110001000101100", -- t[25132] = 2
      "0000010" when "00110001000101101", -- t[25133] = 2
      "0000010" when "00110001000101110", -- t[25134] = 2
      "0000010" when "00110001000101111", -- t[25135] = 2
      "0000010" when "00110001000110000", -- t[25136] = 2
      "0000010" when "00110001000110001", -- t[25137] = 2
      "0000010" when "00110001000110010", -- t[25138] = 2
      "0000010" when "00110001000110011", -- t[25139] = 2
      "0000010" when "00110001000110100", -- t[25140] = 2
      "0000010" when "00110001000110101", -- t[25141] = 2
      "0000010" when "00110001000110110", -- t[25142] = 2
      "0000010" when "00110001000110111", -- t[25143] = 2
      "0000010" when "00110001000111000", -- t[25144] = 2
      "0000010" when "00110001000111001", -- t[25145] = 2
      "0000010" when "00110001000111010", -- t[25146] = 2
      "0000010" when "00110001000111011", -- t[25147] = 2
      "0000010" when "00110001000111100", -- t[25148] = 2
      "0000010" when "00110001000111101", -- t[25149] = 2
      "0000010" when "00110001000111110", -- t[25150] = 2
      "0000010" when "00110001000111111", -- t[25151] = 2
      "0000010" when "00110001001000000", -- t[25152] = 2
      "0000010" when "00110001001000001", -- t[25153] = 2
      "0000010" when "00110001001000010", -- t[25154] = 2
      "0000010" when "00110001001000011", -- t[25155] = 2
      "0000010" when "00110001001000100", -- t[25156] = 2
      "0000010" when "00110001001000101", -- t[25157] = 2
      "0000010" when "00110001001000110", -- t[25158] = 2
      "0000010" when "00110001001000111", -- t[25159] = 2
      "0000010" when "00110001001001000", -- t[25160] = 2
      "0000010" when "00110001001001001", -- t[25161] = 2
      "0000010" when "00110001001001010", -- t[25162] = 2
      "0000010" when "00110001001001011", -- t[25163] = 2
      "0000010" when "00110001001001100", -- t[25164] = 2
      "0000010" when "00110001001001101", -- t[25165] = 2
      "0000010" when "00110001001001110", -- t[25166] = 2
      "0000010" when "00110001001001111", -- t[25167] = 2
      "0000010" when "00110001001010000", -- t[25168] = 2
      "0000010" when "00110001001010001", -- t[25169] = 2
      "0000010" when "00110001001010010", -- t[25170] = 2
      "0000010" when "00110001001010011", -- t[25171] = 2
      "0000010" when "00110001001010100", -- t[25172] = 2
      "0000010" when "00110001001010101", -- t[25173] = 2
      "0000010" when "00110001001010110", -- t[25174] = 2
      "0000010" when "00110001001010111", -- t[25175] = 2
      "0000010" when "00110001001011000", -- t[25176] = 2
      "0000010" when "00110001001011001", -- t[25177] = 2
      "0000010" when "00110001001011010", -- t[25178] = 2
      "0000010" when "00110001001011011", -- t[25179] = 2
      "0000010" when "00110001001011100", -- t[25180] = 2
      "0000010" when "00110001001011101", -- t[25181] = 2
      "0000010" when "00110001001011110", -- t[25182] = 2
      "0000010" when "00110001001011111", -- t[25183] = 2
      "0000010" when "00110001001100000", -- t[25184] = 2
      "0000010" when "00110001001100001", -- t[25185] = 2
      "0000010" when "00110001001100010", -- t[25186] = 2
      "0000010" when "00110001001100011", -- t[25187] = 2
      "0000010" when "00110001001100100", -- t[25188] = 2
      "0000010" when "00110001001100101", -- t[25189] = 2
      "0000010" when "00110001001100110", -- t[25190] = 2
      "0000010" when "00110001001100111", -- t[25191] = 2
      "0000010" when "00110001001101000", -- t[25192] = 2
      "0000010" when "00110001001101001", -- t[25193] = 2
      "0000010" when "00110001001101010", -- t[25194] = 2
      "0000010" when "00110001001101011", -- t[25195] = 2
      "0000010" when "00110001001101100", -- t[25196] = 2
      "0000010" when "00110001001101101", -- t[25197] = 2
      "0000010" when "00110001001101110", -- t[25198] = 2
      "0000010" when "00110001001101111", -- t[25199] = 2
      "0000010" when "00110001001110000", -- t[25200] = 2
      "0000010" when "00110001001110001", -- t[25201] = 2
      "0000010" when "00110001001110010", -- t[25202] = 2
      "0000010" when "00110001001110011", -- t[25203] = 2
      "0000010" when "00110001001110100", -- t[25204] = 2
      "0000010" when "00110001001110101", -- t[25205] = 2
      "0000010" when "00110001001110110", -- t[25206] = 2
      "0000010" when "00110001001110111", -- t[25207] = 2
      "0000010" when "00110001001111000", -- t[25208] = 2
      "0000010" when "00110001001111001", -- t[25209] = 2
      "0000010" when "00110001001111010", -- t[25210] = 2
      "0000010" when "00110001001111011", -- t[25211] = 2
      "0000010" when "00110001001111100", -- t[25212] = 2
      "0000010" when "00110001001111101", -- t[25213] = 2
      "0000010" when "00110001001111110", -- t[25214] = 2
      "0000010" when "00110001001111111", -- t[25215] = 2
      "0000010" when "00110001010000000", -- t[25216] = 2
      "0000010" when "00110001010000001", -- t[25217] = 2
      "0000010" when "00110001010000010", -- t[25218] = 2
      "0000010" when "00110001010000011", -- t[25219] = 2
      "0000010" when "00110001010000100", -- t[25220] = 2
      "0000010" when "00110001010000101", -- t[25221] = 2
      "0000010" when "00110001010000110", -- t[25222] = 2
      "0000010" when "00110001010000111", -- t[25223] = 2
      "0000010" when "00110001010001000", -- t[25224] = 2
      "0000010" when "00110001010001001", -- t[25225] = 2
      "0000010" when "00110001010001010", -- t[25226] = 2
      "0000010" when "00110001010001011", -- t[25227] = 2
      "0000010" when "00110001010001100", -- t[25228] = 2
      "0000010" when "00110001010001101", -- t[25229] = 2
      "0000010" when "00110001010001110", -- t[25230] = 2
      "0000010" when "00110001010001111", -- t[25231] = 2
      "0000010" when "00110001010010000", -- t[25232] = 2
      "0000010" when "00110001010010001", -- t[25233] = 2
      "0000010" when "00110001010010010", -- t[25234] = 2
      "0000010" when "00110001010010011", -- t[25235] = 2
      "0000010" when "00110001010010100", -- t[25236] = 2
      "0000010" when "00110001010010101", -- t[25237] = 2
      "0000010" when "00110001010010110", -- t[25238] = 2
      "0000010" when "00110001010010111", -- t[25239] = 2
      "0000010" when "00110001010011000", -- t[25240] = 2
      "0000010" when "00110001010011001", -- t[25241] = 2
      "0000010" when "00110001010011010", -- t[25242] = 2
      "0000010" when "00110001010011011", -- t[25243] = 2
      "0000010" when "00110001010011100", -- t[25244] = 2
      "0000010" when "00110001010011101", -- t[25245] = 2
      "0000010" when "00110001010011110", -- t[25246] = 2
      "0000010" when "00110001010011111", -- t[25247] = 2
      "0000010" when "00110001010100000", -- t[25248] = 2
      "0000010" when "00110001010100001", -- t[25249] = 2
      "0000010" when "00110001010100010", -- t[25250] = 2
      "0000010" when "00110001010100011", -- t[25251] = 2
      "0000010" when "00110001010100100", -- t[25252] = 2
      "0000010" when "00110001010100101", -- t[25253] = 2
      "0000010" when "00110001010100110", -- t[25254] = 2
      "0000010" when "00110001010100111", -- t[25255] = 2
      "0000010" when "00110001010101000", -- t[25256] = 2
      "0000010" when "00110001010101001", -- t[25257] = 2
      "0000010" when "00110001010101010", -- t[25258] = 2
      "0000010" when "00110001010101011", -- t[25259] = 2
      "0000010" when "00110001010101100", -- t[25260] = 2
      "0000010" when "00110001010101101", -- t[25261] = 2
      "0000010" when "00110001010101110", -- t[25262] = 2
      "0000010" when "00110001010101111", -- t[25263] = 2
      "0000010" when "00110001010110000", -- t[25264] = 2
      "0000010" when "00110001010110001", -- t[25265] = 2
      "0000010" when "00110001010110010", -- t[25266] = 2
      "0000010" when "00110001010110011", -- t[25267] = 2
      "0000010" when "00110001010110100", -- t[25268] = 2
      "0000010" when "00110001010110101", -- t[25269] = 2
      "0000010" when "00110001010110110", -- t[25270] = 2
      "0000010" when "00110001010110111", -- t[25271] = 2
      "0000010" when "00110001010111000", -- t[25272] = 2
      "0000010" when "00110001010111001", -- t[25273] = 2
      "0000010" when "00110001010111010", -- t[25274] = 2
      "0000010" when "00110001010111011", -- t[25275] = 2
      "0000010" when "00110001010111100", -- t[25276] = 2
      "0000010" when "00110001010111101", -- t[25277] = 2
      "0000010" when "00110001010111110", -- t[25278] = 2
      "0000010" when "00110001010111111", -- t[25279] = 2
      "0000010" when "00110001011000000", -- t[25280] = 2
      "0000010" when "00110001011000001", -- t[25281] = 2
      "0000010" when "00110001011000010", -- t[25282] = 2
      "0000010" when "00110001011000011", -- t[25283] = 2
      "0000010" when "00110001011000100", -- t[25284] = 2
      "0000010" when "00110001011000101", -- t[25285] = 2
      "0000010" when "00110001011000110", -- t[25286] = 2
      "0000010" when "00110001011000111", -- t[25287] = 2
      "0000010" when "00110001011001000", -- t[25288] = 2
      "0000010" when "00110001011001001", -- t[25289] = 2
      "0000010" when "00110001011001010", -- t[25290] = 2
      "0000010" when "00110001011001011", -- t[25291] = 2
      "0000010" when "00110001011001100", -- t[25292] = 2
      "0000010" when "00110001011001101", -- t[25293] = 2
      "0000010" when "00110001011001110", -- t[25294] = 2
      "0000010" when "00110001011001111", -- t[25295] = 2
      "0000010" when "00110001011010000", -- t[25296] = 2
      "0000010" when "00110001011010001", -- t[25297] = 2
      "0000010" when "00110001011010010", -- t[25298] = 2
      "0000010" when "00110001011010011", -- t[25299] = 2
      "0000010" when "00110001011010100", -- t[25300] = 2
      "0000010" when "00110001011010101", -- t[25301] = 2
      "0000010" when "00110001011010110", -- t[25302] = 2
      "0000010" when "00110001011010111", -- t[25303] = 2
      "0000010" when "00110001011011000", -- t[25304] = 2
      "0000010" when "00110001011011001", -- t[25305] = 2
      "0000010" when "00110001011011010", -- t[25306] = 2
      "0000010" when "00110001011011011", -- t[25307] = 2
      "0000010" when "00110001011011100", -- t[25308] = 2
      "0000010" when "00110001011011101", -- t[25309] = 2
      "0000010" when "00110001011011110", -- t[25310] = 2
      "0000010" when "00110001011011111", -- t[25311] = 2
      "0000010" when "00110001011100000", -- t[25312] = 2
      "0000010" when "00110001011100001", -- t[25313] = 2
      "0000010" when "00110001011100010", -- t[25314] = 2
      "0000010" when "00110001011100011", -- t[25315] = 2
      "0000010" when "00110001011100100", -- t[25316] = 2
      "0000010" when "00110001011100101", -- t[25317] = 2
      "0000010" when "00110001011100110", -- t[25318] = 2
      "0000010" when "00110001011100111", -- t[25319] = 2
      "0000010" when "00110001011101000", -- t[25320] = 2
      "0000010" when "00110001011101001", -- t[25321] = 2
      "0000010" when "00110001011101010", -- t[25322] = 2
      "0000010" when "00110001011101011", -- t[25323] = 2
      "0000010" when "00110001011101100", -- t[25324] = 2
      "0000010" when "00110001011101101", -- t[25325] = 2
      "0000010" when "00110001011101110", -- t[25326] = 2
      "0000010" when "00110001011101111", -- t[25327] = 2
      "0000010" when "00110001011110000", -- t[25328] = 2
      "0000010" when "00110001011110001", -- t[25329] = 2
      "0000010" when "00110001011110010", -- t[25330] = 2
      "0000010" when "00110001011110011", -- t[25331] = 2
      "0000010" when "00110001011110100", -- t[25332] = 2
      "0000010" when "00110001011110101", -- t[25333] = 2
      "0000010" when "00110001011110110", -- t[25334] = 2
      "0000010" when "00110001011110111", -- t[25335] = 2
      "0000010" when "00110001011111000", -- t[25336] = 2
      "0000010" when "00110001011111001", -- t[25337] = 2
      "0000010" when "00110001011111010", -- t[25338] = 2
      "0000010" when "00110001011111011", -- t[25339] = 2
      "0000010" when "00110001011111100", -- t[25340] = 2
      "0000010" when "00110001011111101", -- t[25341] = 2
      "0000010" when "00110001011111110", -- t[25342] = 2
      "0000010" when "00110001011111111", -- t[25343] = 2
      "0000010" when "00110001100000000", -- t[25344] = 2
      "0000010" when "00110001100000001", -- t[25345] = 2
      "0000010" when "00110001100000010", -- t[25346] = 2
      "0000010" when "00110001100000011", -- t[25347] = 2
      "0000010" when "00110001100000100", -- t[25348] = 2
      "0000010" when "00110001100000101", -- t[25349] = 2
      "0000010" when "00110001100000110", -- t[25350] = 2
      "0000010" when "00110001100000111", -- t[25351] = 2
      "0000010" when "00110001100001000", -- t[25352] = 2
      "0000010" when "00110001100001001", -- t[25353] = 2
      "0000010" when "00110001100001010", -- t[25354] = 2
      "0000010" when "00110001100001011", -- t[25355] = 2
      "0000010" when "00110001100001100", -- t[25356] = 2
      "0000010" when "00110001100001101", -- t[25357] = 2
      "0000010" when "00110001100001110", -- t[25358] = 2
      "0000010" when "00110001100001111", -- t[25359] = 2
      "0000010" when "00110001100010000", -- t[25360] = 2
      "0000010" when "00110001100010001", -- t[25361] = 2
      "0000010" when "00110001100010010", -- t[25362] = 2
      "0000010" when "00110001100010011", -- t[25363] = 2
      "0000010" when "00110001100010100", -- t[25364] = 2
      "0000010" when "00110001100010101", -- t[25365] = 2
      "0000010" when "00110001100010110", -- t[25366] = 2
      "0000010" when "00110001100010111", -- t[25367] = 2
      "0000010" when "00110001100011000", -- t[25368] = 2
      "0000010" when "00110001100011001", -- t[25369] = 2
      "0000010" when "00110001100011010", -- t[25370] = 2
      "0000010" when "00110001100011011", -- t[25371] = 2
      "0000010" when "00110001100011100", -- t[25372] = 2
      "0000010" when "00110001100011101", -- t[25373] = 2
      "0000010" when "00110001100011110", -- t[25374] = 2
      "0000010" when "00110001100011111", -- t[25375] = 2
      "0000010" when "00110001100100000", -- t[25376] = 2
      "0000010" when "00110001100100001", -- t[25377] = 2
      "0000010" when "00110001100100010", -- t[25378] = 2
      "0000010" when "00110001100100011", -- t[25379] = 2
      "0000010" when "00110001100100100", -- t[25380] = 2
      "0000010" when "00110001100100101", -- t[25381] = 2
      "0000010" when "00110001100100110", -- t[25382] = 2
      "0000010" when "00110001100100111", -- t[25383] = 2
      "0000010" when "00110001100101000", -- t[25384] = 2
      "0000010" when "00110001100101001", -- t[25385] = 2
      "0000010" when "00110001100101010", -- t[25386] = 2
      "0000010" when "00110001100101011", -- t[25387] = 2
      "0000010" when "00110001100101100", -- t[25388] = 2
      "0000010" when "00110001100101101", -- t[25389] = 2
      "0000010" when "00110001100101110", -- t[25390] = 2
      "0000010" when "00110001100101111", -- t[25391] = 2
      "0000010" when "00110001100110000", -- t[25392] = 2
      "0000010" when "00110001100110001", -- t[25393] = 2
      "0000010" when "00110001100110010", -- t[25394] = 2
      "0000010" when "00110001100110011", -- t[25395] = 2
      "0000010" when "00110001100110100", -- t[25396] = 2
      "0000010" when "00110001100110101", -- t[25397] = 2
      "0000010" when "00110001100110110", -- t[25398] = 2
      "0000010" when "00110001100110111", -- t[25399] = 2
      "0000010" when "00110001100111000", -- t[25400] = 2
      "0000010" when "00110001100111001", -- t[25401] = 2
      "0000010" when "00110001100111010", -- t[25402] = 2
      "0000010" when "00110001100111011", -- t[25403] = 2
      "0000010" when "00110001100111100", -- t[25404] = 2
      "0000010" when "00110001100111101", -- t[25405] = 2
      "0000010" when "00110001100111110", -- t[25406] = 2
      "0000010" when "00110001100111111", -- t[25407] = 2
      "0000010" when "00110001101000000", -- t[25408] = 2
      "0000010" when "00110001101000001", -- t[25409] = 2
      "0000010" when "00110001101000010", -- t[25410] = 2
      "0000010" when "00110001101000011", -- t[25411] = 2
      "0000010" when "00110001101000100", -- t[25412] = 2
      "0000010" when "00110001101000101", -- t[25413] = 2
      "0000010" when "00110001101000110", -- t[25414] = 2
      "0000010" when "00110001101000111", -- t[25415] = 2
      "0000010" when "00110001101001000", -- t[25416] = 2
      "0000010" when "00110001101001001", -- t[25417] = 2
      "0000010" when "00110001101001010", -- t[25418] = 2
      "0000010" when "00110001101001011", -- t[25419] = 2
      "0000010" when "00110001101001100", -- t[25420] = 2
      "0000010" when "00110001101001101", -- t[25421] = 2
      "0000010" when "00110001101001110", -- t[25422] = 2
      "0000010" when "00110001101001111", -- t[25423] = 2
      "0000010" when "00110001101010000", -- t[25424] = 2
      "0000010" when "00110001101010001", -- t[25425] = 2
      "0000010" when "00110001101010010", -- t[25426] = 2
      "0000010" when "00110001101010011", -- t[25427] = 2
      "0000010" when "00110001101010100", -- t[25428] = 2
      "0000010" when "00110001101010101", -- t[25429] = 2
      "0000010" when "00110001101010110", -- t[25430] = 2
      "0000010" when "00110001101010111", -- t[25431] = 2
      "0000010" when "00110001101011000", -- t[25432] = 2
      "0000010" when "00110001101011001", -- t[25433] = 2
      "0000010" when "00110001101011010", -- t[25434] = 2
      "0000010" when "00110001101011011", -- t[25435] = 2
      "0000010" when "00110001101011100", -- t[25436] = 2
      "0000010" when "00110001101011101", -- t[25437] = 2
      "0000010" when "00110001101011110", -- t[25438] = 2
      "0000010" when "00110001101011111", -- t[25439] = 2
      "0000010" when "00110001101100000", -- t[25440] = 2
      "0000010" when "00110001101100001", -- t[25441] = 2
      "0000010" when "00110001101100010", -- t[25442] = 2
      "0000010" when "00110001101100011", -- t[25443] = 2
      "0000010" when "00110001101100100", -- t[25444] = 2
      "0000010" when "00110001101100101", -- t[25445] = 2
      "0000010" when "00110001101100110", -- t[25446] = 2
      "0000010" when "00110001101100111", -- t[25447] = 2
      "0000010" when "00110001101101000", -- t[25448] = 2
      "0000010" when "00110001101101001", -- t[25449] = 2
      "0000010" when "00110001101101010", -- t[25450] = 2
      "0000010" when "00110001101101011", -- t[25451] = 2
      "0000010" when "00110001101101100", -- t[25452] = 2
      "0000010" when "00110001101101101", -- t[25453] = 2
      "0000010" when "00110001101101110", -- t[25454] = 2
      "0000010" when "00110001101101111", -- t[25455] = 2
      "0000010" when "00110001101110000", -- t[25456] = 2
      "0000010" when "00110001101110001", -- t[25457] = 2
      "0000010" when "00110001101110010", -- t[25458] = 2
      "0000010" when "00110001101110011", -- t[25459] = 2
      "0000010" when "00110001101110100", -- t[25460] = 2
      "0000010" when "00110001101110101", -- t[25461] = 2
      "0000010" when "00110001101110110", -- t[25462] = 2
      "0000010" when "00110001101110111", -- t[25463] = 2
      "0000010" when "00110001101111000", -- t[25464] = 2
      "0000010" when "00110001101111001", -- t[25465] = 2
      "0000010" when "00110001101111010", -- t[25466] = 2
      "0000010" when "00110001101111011", -- t[25467] = 2
      "0000010" when "00110001101111100", -- t[25468] = 2
      "0000010" when "00110001101111101", -- t[25469] = 2
      "0000010" when "00110001101111110", -- t[25470] = 2
      "0000010" when "00110001101111111", -- t[25471] = 2
      "0000010" when "00110001110000000", -- t[25472] = 2
      "0000010" when "00110001110000001", -- t[25473] = 2
      "0000010" when "00110001110000010", -- t[25474] = 2
      "0000010" when "00110001110000011", -- t[25475] = 2
      "0000010" when "00110001110000100", -- t[25476] = 2
      "0000010" when "00110001110000101", -- t[25477] = 2
      "0000010" when "00110001110000110", -- t[25478] = 2
      "0000010" when "00110001110000111", -- t[25479] = 2
      "0000010" when "00110001110001000", -- t[25480] = 2
      "0000010" when "00110001110001001", -- t[25481] = 2
      "0000010" when "00110001110001010", -- t[25482] = 2
      "0000010" when "00110001110001011", -- t[25483] = 2
      "0000010" when "00110001110001100", -- t[25484] = 2
      "0000010" when "00110001110001101", -- t[25485] = 2
      "0000010" when "00110001110001110", -- t[25486] = 2
      "0000010" when "00110001110001111", -- t[25487] = 2
      "0000010" when "00110001110010000", -- t[25488] = 2
      "0000010" when "00110001110010001", -- t[25489] = 2
      "0000010" when "00110001110010010", -- t[25490] = 2
      "0000010" when "00110001110010011", -- t[25491] = 2
      "0000010" when "00110001110010100", -- t[25492] = 2
      "0000010" when "00110001110010101", -- t[25493] = 2
      "0000010" when "00110001110010110", -- t[25494] = 2
      "0000010" when "00110001110010111", -- t[25495] = 2
      "0000010" when "00110001110011000", -- t[25496] = 2
      "0000010" when "00110001110011001", -- t[25497] = 2
      "0000010" when "00110001110011010", -- t[25498] = 2
      "0000010" when "00110001110011011", -- t[25499] = 2
      "0000010" when "00110001110011100", -- t[25500] = 2
      "0000010" when "00110001110011101", -- t[25501] = 2
      "0000010" when "00110001110011110", -- t[25502] = 2
      "0000010" when "00110001110011111", -- t[25503] = 2
      "0000010" when "00110001110100000", -- t[25504] = 2
      "0000010" when "00110001110100001", -- t[25505] = 2
      "0000010" when "00110001110100010", -- t[25506] = 2
      "0000010" when "00110001110100011", -- t[25507] = 2
      "0000010" when "00110001110100100", -- t[25508] = 2
      "0000010" when "00110001110100101", -- t[25509] = 2
      "0000010" when "00110001110100110", -- t[25510] = 2
      "0000010" when "00110001110100111", -- t[25511] = 2
      "0000010" when "00110001110101000", -- t[25512] = 2
      "0000010" when "00110001110101001", -- t[25513] = 2
      "0000010" when "00110001110101010", -- t[25514] = 2
      "0000010" when "00110001110101011", -- t[25515] = 2
      "0000010" when "00110001110101100", -- t[25516] = 2
      "0000010" when "00110001110101101", -- t[25517] = 2
      "0000010" when "00110001110101110", -- t[25518] = 2
      "0000010" when "00110001110101111", -- t[25519] = 2
      "0000010" when "00110001110110000", -- t[25520] = 2
      "0000010" when "00110001110110001", -- t[25521] = 2
      "0000010" when "00110001110110010", -- t[25522] = 2
      "0000010" when "00110001110110011", -- t[25523] = 2
      "0000010" when "00110001110110100", -- t[25524] = 2
      "0000010" when "00110001110110101", -- t[25525] = 2
      "0000010" when "00110001110110110", -- t[25526] = 2
      "0000010" when "00110001110110111", -- t[25527] = 2
      "0000010" when "00110001110111000", -- t[25528] = 2
      "0000010" when "00110001110111001", -- t[25529] = 2
      "0000010" when "00110001110111010", -- t[25530] = 2
      "0000010" when "00110001110111011", -- t[25531] = 2
      "0000010" when "00110001110111100", -- t[25532] = 2
      "0000010" when "00110001110111101", -- t[25533] = 2
      "0000010" when "00110001110111110", -- t[25534] = 2
      "0000010" when "00110001110111111", -- t[25535] = 2
      "0000010" when "00110001111000000", -- t[25536] = 2
      "0000010" when "00110001111000001", -- t[25537] = 2
      "0000010" when "00110001111000010", -- t[25538] = 2
      "0000010" when "00110001111000011", -- t[25539] = 2
      "0000010" when "00110001111000100", -- t[25540] = 2
      "0000010" when "00110001111000101", -- t[25541] = 2
      "0000010" when "00110001111000110", -- t[25542] = 2
      "0000010" when "00110001111000111", -- t[25543] = 2
      "0000010" when "00110001111001000", -- t[25544] = 2
      "0000010" when "00110001111001001", -- t[25545] = 2
      "0000010" when "00110001111001010", -- t[25546] = 2
      "0000010" when "00110001111001011", -- t[25547] = 2
      "0000010" when "00110001111001100", -- t[25548] = 2
      "0000010" when "00110001111001101", -- t[25549] = 2
      "0000010" when "00110001111001110", -- t[25550] = 2
      "0000010" when "00110001111001111", -- t[25551] = 2
      "0000010" when "00110001111010000", -- t[25552] = 2
      "0000010" when "00110001111010001", -- t[25553] = 2
      "0000010" when "00110001111010010", -- t[25554] = 2
      "0000010" when "00110001111010011", -- t[25555] = 2
      "0000010" when "00110001111010100", -- t[25556] = 2
      "0000010" when "00110001111010101", -- t[25557] = 2
      "0000010" when "00110001111010110", -- t[25558] = 2
      "0000010" when "00110001111010111", -- t[25559] = 2
      "0000010" when "00110001111011000", -- t[25560] = 2
      "0000010" when "00110001111011001", -- t[25561] = 2
      "0000010" when "00110001111011010", -- t[25562] = 2
      "0000010" when "00110001111011011", -- t[25563] = 2
      "0000010" when "00110001111011100", -- t[25564] = 2
      "0000010" when "00110001111011101", -- t[25565] = 2
      "0000010" when "00110001111011110", -- t[25566] = 2
      "0000010" when "00110001111011111", -- t[25567] = 2
      "0000010" when "00110001111100000", -- t[25568] = 2
      "0000010" when "00110001111100001", -- t[25569] = 2
      "0000010" when "00110001111100010", -- t[25570] = 2
      "0000010" when "00110001111100011", -- t[25571] = 2
      "0000010" when "00110001111100100", -- t[25572] = 2
      "0000010" when "00110001111100101", -- t[25573] = 2
      "0000010" when "00110001111100110", -- t[25574] = 2
      "0000010" when "00110001111100111", -- t[25575] = 2
      "0000010" when "00110001111101000", -- t[25576] = 2
      "0000010" when "00110001111101001", -- t[25577] = 2
      "0000010" when "00110001111101010", -- t[25578] = 2
      "0000010" when "00110001111101011", -- t[25579] = 2
      "0000010" when "00110001111101100", -- t[25580] = 2
      "0000010" when "00110001111101101", -- t[25581] = 2
      "0000010" when "00110001111101110", -- t[25582] = 2
      "0000010" when "00110001111101111", -- t[25583] = 2
      "0000010" when "00110001111110000", -- t[25584] = 2
      "0000010" when "00110001111110001", -- t[25585] = 2
      "0000010" when "00110001111110010", -- t[25586] = 2
      "0000010" when "00110001111110011", -- t[25587] = 2
      "0000010" when "00110001111110100", -- t[25588] = 2
      "0000010" when "00110001111110101", -- t[25589] = 2
      "0000010" when "00110001111110110", -- t[25590] = 2
      "0000010" when "00110001111110111", -- t[25591] = 2
      "0000010" when "00110001111111000", -- t[25592] = 2
      "0000010" when "00110001111111001", -- t[25593] = 2
      "0000010" when "00110001111111010", -- t[25594] = 2
      "0000010" when "00110001111111011", -- t[25595] = 2
      "0000010" when "00110001111111100", -- t[25596] = 2
      "0000010" when "00110001111111101", -- t[25597] = 2
      "0000010" when "00110001111111110", -- t[25598] = 2
      "0000010" when "00110001111111111", -- t[25599] = 2
      "0000010" when "00110010000000000", -- t[25600] = 2
      "0000010" when "00110010000000001", -- t[25601] = 2
      "0000010" when "00110010000000010", -- t[25602] = 2
      "0000010" when "00110010000000011", -- t[25603] = 2
      "0000010" when "00110010000000100", -- t[25604] = 2
      "0000010" when "00110010000000101", -- t[25605] = 2
      "0000010" when "00110010000000110", -- t[25606] = 2
      "0000010" when "00110010000000111", -- t[25607] = 2
      "0000010" when "00110010000001000", -- t[25608] = 2
      "0000010" when "00110010000001001", -- t[25609] = 2
      "0000010" when "00110010000001010", -- t[25610] = 2
      "0000010" when "00110010000001011", -- t[25611] = 2
      "0000010" when "00110010000001100", -- t[25612] = 2
      "0000010" when "00110010000001101", -- t[25613] = 2
      "0000010" when "00110010000001110", -- t[25614] = 2
      "0000010" when "00110010000001111", -- t[25615] = 2
      "0000010" when "00110010000010000", -- t[25616] = 2
      "0000010" when "00110010000010001", -- t[25617] = 2
      "0000010" when "00110010000010010", -- t[25618] = 2
      "0000010" when "00110010000010011", -- t[25619] = 2
      "0000010" when "00110010000010100", -- t[25620] = 2
      "0000010" when "00110010000010101", -- t[25621] = 2
      "0000010" when "00110010000010110", -- t[25622] = 2
      "0000010" when "00110010000010111", -- t[25623] = 2
      "0000010" when "00110010000011000", -- t[25624] = 2
      "0000010" when "00110010000011001", -- t[25625] = 2
      "0000010" when "00110010000011010", -- t[25626] = 2
      "0000010" when "00110010000011011", -- t[25627] = 2
      "0000010" when "00110010000011100", -- t[25628] = 2
      "0000010" when "00110010000011101", -- t[25629] = 2
      "0000010" when "00110010000011110", -- t[25630] = 2
      "0000010" when "00110010000011111", -- t[25631] = 2
      "0000010" when "00110010000100000", -- t[25632] = 2
      "0000010" when "00110010000100001", -- t[25633] = 2
      "0000010" when "00110010000100010", -- t[25634] = 2
      "0000010" when "00110010000100011", -- t[25635] = 2
      "0000010" when "00110010000100100", -- t[25636] = 2
      "0000010" when "00110010000100101", -- t[25637] = 2
      "0000010" when "00110010000100110", -- t[25638] = 2
      "0000010" when "00110010000100111", -- t[25639] = 2
      "0000010" when "00110010000101000", -- t[25640] = 2
      "0000010" when "00110010000101001", -- t[25641] = 2
      "0000010" when "00110010000101010", -- t[25642] = 2
      "0000010" when "00110010000101011", -- t[25643] = 2
      "0000010" when "00110010000101100", -- t[25644] = 2
      "0000010" when "00110010000101101", -- t[25645] = 2
      "0000010" when "00110010000101110", -- t[25646] = 2
      "0000010" when "00110010000101111", -- t[25647] = 2
      "0000010" when "00110010000110000", -- t[25648] = 2
      "0000010" when "00110010000110001", -- t[25649] = 2
      "0000010" when "00110010000110010", -- t[25650] = 2
      "0000010" when "00110010000110011", -- t[25651] = 2
      "0000010" when "00110010000110100", -- t[25652] = 2
      "0000010" when "00110010000110101", -- t[25653] = 2
      "0000010" when "00110010000110110", -- t[25654] = 2
      "0000010" when "00110010000110111", -- t[25655] = 2
      "0000010" when "00110010000111000", -- t[25656] = 2
      "0000010" when "00110010000111001", -- t[25657] = 2
      "0000010" when "00110010000111010", -- t[25658] = 2
      "0000010" when "00110010000111011", -- t[25659] = 2
      "0000010" when "00110010000111100", -- t[25660] = 2
      "0000010" when "00110010000111101", -- t[25661] = 2
      "0000010" when "00110010000111110", -- t[25662] = 2
      "0000010" when "00110010000111111", -- t[25663] = 2
      "0000010" when "00110010001000000", -- t[25664] = 2
      "0000010" when "00110010001000001", -- t[25665] = 2
      "0000010" when "00110010001000010", -- t[25666] = 2
      "0000010" when "00110010001000011", -- t[25667] = 2
      "0000010" when "00110010001000100", -- t[25668] = 2
      "0000010" when "00110010001000101", -- t[25669] = 2
      "0000010" when "00110010001000110", -- t[25670] = 2
      "0000010" when "00110010001000111", -- t[25671] = 2
      "0000010" when "00110010001001000", -- t[25672] = 2
      "0000010" when "00110010001001001", -- t[25673] = 2
      "0000010" when "00110010001001010", -- t[25674] = 2
      "0000010" when "00110010001001011", -- t[25675] = 2
      "0000010" when "00110010001001100", -- t[25676] = 2
      "0000010" when "00110010001001101", -- t[25677] = 2
      "0000010" when "00110010001001110", -- t[25678] = 2
      "0000010" when "00110010001001111", -- t[25679] = 2
      "0000010" when "00110010001010000", -- t[25680] = 2
      "0000010" when "00110010001010001", -- t[25681] = 2
      "0000010" when "00110010001010010", -- t[25682] = 2
      "0000010" when "00110010001010011", -- t[25683] = 2
      "0000010" when "00110010001010100", -- t[25684] = 2
      "0000010" when "00110010001010101", -- t[25685] = 2
      "0000010" when "00110010001010110", -- t[25686] = 2
      "0000010" when "00110010001010111", -- t[25687] = 2
      "0000010" when "00110010001011000", -- t[25688] = 2
      "0000010" when "00110010001011001", -- t[25689] = 2
      "0000010" when "00110010001011010", -- t[25690] = 2
      "0000010" when "00110010001011011", -- t[25691] = 2
      "0000010" when "00110010001011100", -- t[25692] = 2
      "0000010" when "00110010001011101", -- t[25693] = 2
      "0000010" when "00110010001011110", -- t[25694] = 2
      "0000010" when "00110010001011111", -- t[25695] = 2
      "0000010" when "00110010001100000", -- t[25696] = 2
      "0000010" when "00110010001100001", -- t[25697] = 2
      "0000010" when "00110010001100010", -- t[25698] = 2
      "0000010" when "00110010001100011", -- t[25699] = 2
      "0000010" when "00110010001100100", -- t[25700] = 2
      "0000010" when "00110010001100101", -- t[25701] = 2
      "0000010" when "00110010001100110", -- t[25702] = 2
      "0000010" when "00110010001100111", -- t[25703] = 2
      "0000010" when "00110010001101000", -- t[25704] = 2
      "0000010" when "00110010001101001", -- t[25705] = 2
      "0000010" when "00110010001101010", -- t[25706] = 2
      "0000010" when "00110010001101011", -- t[25707] = 2
      "0000010" when "00110010001101100", -- t[25708] = 2
      "0000010" when "00110010001101101", -- t[25709] = 2
      "0000010" when "00110010001101110", -- t[25710] = 2
      "0000010" when "00110010001101111", -- t[25711] = 2
      "0000010" when "00110010001110000", -- t[25712] = 2
      "0000010" when "00110010001110001", -- t[25713] = 2
      "0000010" when "00110010001110010", -- t[25714] = 2
      "0000010" when "00110010001110011", -- t[25715] = 2
      "0000010" when "00110010001110100", -- t[25716] = 2
      "0000010" when "00110010001110101", -- t[25717] = 2
      "0000010" when "00110010001110110", -- t[25718] = 2
      "0000010" when "00110010001110111", -- t[25719] = 2
      "0000010" when "00110010001111000", -- t[25720] = 2
      "0000010" when "00110010001111001", -- t[25721] = 2
      "0000010" when "00110010001111010", -- t[25722] = 2
      "0000010" when "00110010001111011", -- t[25723] = 2
      "0000010" when "00110010001111100", -- t[25724] = 2
      "0000010" when "00110010001111101", -- t[25725] = 2
      "0000010" when "00110010001111110", -- t[25726] = 2
      "0000010" when "00110010001111111", -- t[25727] = 2
      "0000010" when "00110010010000000", -- t[25728] = 2
      "0000010" when "00110010010000001", -- t[25729] = 2
      "0000010" when "00110010010000010", -- t[25730] = 2
      "0000010" when "00110010010000011", -- t[25731] = 2
      "0000010" when "00110010010000100", -- t[25732] = 2
      "0000010" when "00110010010000101", -- t[25733] = 2
      "0000010" when "00110010010000110", -- t[25734] = 2
      "0000010" when "00110010010000111", -- t[25735] = 2
      "0000010" when "00110010010001000", -- t[25736] = 2
      "0000010" when "00110010010001001", -- t[25737] = 2
      "0000010" when "00110010010001010", -- t[25738] = 2
      "0000010" when "00110010010001011", -- t[25739] = 2
      "0000010" when "00110010010001100", -- t[25740] = 2
      "0000010" when "00110010010001101", -- t[25741] = 2
      "0000010" when "00110010010001110", -- t[25742] = 2
      "0000010" when "00110010010001111", -- t[25743] = 2
      "0000010" when "00110010010010000", -- t[25744] = 2
      "0000010" when "00110010010010001", -- t[25745] = 2
      "0000010" when "00110010010010010", -- t[25746] = 2
      "0000010" when "00110010010010011", -- t[25747] = 2
      "0000010" when "00110010010010100", -- t[25748] = 2
      "0000010" when "00110010010010101", -- t[25749] = 2
      "0000010" when "00110010010010110", -- t[25750] = 2
      "0000010" when "00110010010010111", -- t[25751] = 2
      "0000010" when "00110010010011000", -- t[25752] = 2
      "0000010" when "00110010010011001", -- t[25753] = 2
      "0000010" when "00110010010011010", -- t[25754] = 2
      "0000010" when "00110010010011011", -- t[25755] = 2
      "0000010" when "00110010010011100", -- t[25756] = 2
      "0000010" when "00110010010011101", -- t[25757] = 2
      "0000010" when "00110010010011110", -- t[25758] = 2
      "0000010" when "00110010010011111", -- t[25759] = 2
      "0000010" when "00110010010100000", -- t[25760] = 2
      "0000010" when "00110010010100001", -- t[25761] = 2
      "0000010" when "00110010010100010", -- t[25762] = 2
      "0000010" when "00110010010100011", -- t[25763] = 2
      "0000010" when "00110010010100100", -- t[25764] = 2
      "0000010" when "00110010010100101", -- t[25765] = 2
      "0000010" when "00110010010100110", -- t[25766] = 2
      "0000010" when "00110010010100111", -- t[25767] = 2
      "0000010" when "00110010010101000", -- t[25768] = 2
      "0000010" when "00110010010101001", -- t[25769] = 2
      "0000010" when "00110010010101010", -- t[25770] = 2
      "0000010" when "00110010010101011", -- t[25771] = 2
      "0000010" when "00110010010101100", -- t[25772] = 2
      "0000010" when "00110010010101101", -- t[25773] = 2
      "0000010" when "00110010010101110", -- t[25774] = 2
      "0000010" when "00110010010101111", -- t[25775] = 2
      "0000010" when "00110010010110000", -- t[25776] = 2
      "0000010" when "00110010010110001", -- t[25777] = 2
      "0000010" when "00110010010110010", -- t[25778] = 2
      "0000010" when "00110010010110011", -- t[25779] = 2
      "0000010" when "00110010010110100", -- t[25780] = 2
      "0000010" when "00110010010110101", -- t[25781] = 2
      "0000010" when "00110010010110110", -- t[25782] = 2
      "0000010" when "00110010010110111", -- t[25783] = 2
      "0000010" when "00110010010111000", -- t[25784] = 2
      "0000010" when "00110010010111001", -- t[25785] = 2
      "0000010" when "00110010010111010", -- t[25786] = 2
      "0000010" when "00110010010111011", -- t[25787] = 2
      "0000010" when "00110010010111100", -- t[25788] = 2
      "0000010" when "00110010010111101", -- t[25789] = 2
      "0000010" when "00110010010111110", -- t[25790] = 2
      "0000010" when "00110010010111111", -- t[25791] = 2
      "0000010" when "00110010011000000", -- t[25792] = 2
      "0000010" when "00110010011000001", -- t[25793] = 2
      "0000010" when "00110010011000010", -- t[25794] = 2
      "0000010" when "00110010011000011", -- t[25795] = 2
      "0000010" when "00110010011000100", -- t[25796] = 2
      "0000010" when "00110010011000101", -- t[25797] = 2
      "0000010" when "00110010011000110", -- t[25798] = 2
      "0000010" when "00110010011000111", -- t[25799] = 2
      "0000010" when "00110010011001000", -- t[25800] = 2
      "0000010" when "00110010011001001", -- t[25801] = 2
      "0000010" when "00110010011001010", -- t[25802] = 2
      "0000010" when "00110010011001011", -- t[25803] = 2
      "0000010" when "00110010011001100", -- t[25804] = 2
      "0000010" when "00110010011001101", -- t[25805] = 2
      "0000010" when "00110010011001110", -- t[25806] = 2
      "0000010" when "00110010011001111", -- t[25807] = 2
      "0000010" when "00110010011010000", -- t[25808] = 2
      "0000010" when "00110010011010001", -- t[25809] = 2
      "0000010" when "00110010011010010", -- t[25810] = 2
      "0000010" when "00110010011010011", -- t[25811] = 2
      "0000010" when "00110010011010100", -- t[25812] = 2
      "0000010" when "00110010011010101", -- t[25813] = 2
      "0000010" when "00110010011010110", -- t[25814] = 2
      "0000010" when "00110010011010111", -- t[25815] = 2
      "0000010" when "00110010011011000", -- t[25816] = 2
      "0000010" when "00110010011011001", -- t[25817] = 2
      "0000010" when "00110010011011010", -- t[25818] = 2
      "0000010" when "00110010011011011", -- t[25819] = 2
      "0000010" when "00110010011011100", -- t[25820] = 2
      "0000010" when "00110010011011101", -- t[25821] = 2
      "0000010" when "00110010011011110", -- t[25822] = 2
      "0000010" when "00110010011011111", -- t[25823] = 2
      "0000010" when "00110010011100000", -- t[25824] = 2
      "0000010" when "00110010011100001", -- t[25825] = 2
      "0000010" when "00110010011100010", -- t[25826] = 2
      "0000010" when "00110010011100011", -- t[25827] = 2
      "0000010" when "00110010011100100", -- t[25828] = 2
      "0000010" when "00110010011100101", -- t[25829] = 2
      "0000010" when "00110010011100110", -- t[25830] = 2
      "0000010" when "00110010011100111", -- t[25831] = 2
      "0000010" when "00110010011101000", -- t[25832] = 2
      "0000010" when "00110010011101001", -- t[25833] = 2
      "0000010" when "00110010011101010", -- t[25834] = 2
      "0000010" when "00110010011101011", -- t[25835] = 2
      "0000010" when "00110010011101100", -- t[25836] = 2
      "0000010" when "00110010011101101", -- t[25837] = 2
      "0000010" when "00110010011101110", -- t[25838] = 2
      "0000010" when "00110010011101111", -- t[25839] = 2
      "0000010" when "00110010011110000", -- t[25840] = 2
      "0000010" when "00110010011110001", -- t[25841] = 2
      "0000010" when "00110010011110010", -- t[25842] = 2
      "0000010" when "00110010011110011", -- t[25843] = 2
      "0000010" when "00110010011110100", -- t[25844] = 2
      "0000010" when "00110010011110101", -- t[25845] = 2
      "0000010" when "00110010011110110", -- t[25846] = 2
      "0000010" when "00110010011110111", -- t[25847] = 2
      "0000010" when "00110010011111000", -- t[25848] = 2
      "0000010" when "00110010011111001", -- t[25849] = 2
      "0000010" when "00110010011111010", -- t[25850] = 2
      "0000010" when "00110010011111011", -- t[25851] = 2
      "0000010" when "00110010011111100", -- t[25852] = 2
      "0000010" when "00110010011111101", -- t[25853] = 2
      "0000010" when "00110010011111110", -- t[25854] = 2
      "0000010" when "00110010011111111", -- t[25855] = 2
      "0000010" when "00110010100000000", -- t[25856] = 2
      "0000010" when "00110010100000001", -- t[25857] = 2
      "0000010" when "00110010100000010", -- t[25858] = 2
      "0000010" when "00110010100000011", -- t[25859] = 2
      "0000010" when "00110010100000100", -- t[25860] = 2
      "0000010" when "00110010100000101", -- t[25861] = 2
      "0000010" when "00110010100000110", -- t[25862] = 2
      "0000010" when "00110010100000111", -- t[25863] = 2
      "0000010" when "00110010100001000", -- t[25864] = 2
      "0000010" when "00110010100001001", -- t[25865] = 2
      "0000010" when "00110010100001010", -- t[25866] = 2
      "0000010" when "00110010100001011", -- t[25867] = 2
      "0000010" when "00110010100001100", -- t[25868] = 2
      "0000010" when "00110010100001101", -- t[25869] = 2
      "0000010" when "00110010100001110", -- t[25870] = 2
      "0000010" when "00110010100001111", -- t[25871] = 2
      "0000010" when "00110010100010000", -- t[25872] = 2
      "0000010" when "00110010100010001", -- t[25873] = 2
      "0000010" when "00110010100010010", -- t[25874] = 2
      "0000010" when "00110010100010011", -- t[25875] = 2
      "0000010" when "00110010100010100", -- t[25876] = 2
      "0000010" when "00110010100010101", -- t[25877] = 2
      "0000010" when "00110010100010110", -- t[25878] = 2
      "0000010" when "00110010100010111", -- t[25879] = 2
      "0000010" when "00110010100011000", -- t[25880] = 2
      "0000010" when "00110010100011001", -- t[25881] = 2
      "0000010" when "00110010100011010", -- t[25882] = 2
      "0000010" when "00110010100011011", -- t[25883] = 2
      "0000010" when "00110010100011100", -- t[25884] = 2
      "0000010" when "00110010100011101", -- t[25885] = 2
      "0000010" when "00110010100011110", -- t[25886] = 2
      "0000010" when "00110010100011111", -- t[25887] = 2
      "0000010" when "00110010100100000", -- t[25888] = 2
      "0000010" when "00110010100100001", -- t[25889] = 2
      "0000010" when "00110010100100010", -- t[25890] = 2
      "0000010" when "00110010100100011", -- t[25891] = 2
      "0000010" when "00110010100100100", -- t[25892] = 2
      "0000010" when "00110010100100101", -- t[25893] = 2
      "0000010" when "00110010100100110", -- t[25894] = 2
      "0000010" when "00110010100100111", -- t[25895] = 2
      "0000010" when "00110010100101000", -- t[25896] = 2
      "0000010" when "00110010100101001", -- t[25897] = 2
      "0000010" when "00110010100101010", -- t[25898] = 2
      "0000010" when "00110010100101011", -- t[25899] = 2
      "0000010" when "00110010100101100", -- t[25900] = 2
      "0000010" when "00110010100101101", -- t[25901] = 2
      "0000010" when "00110010100101110", -- t[25902] = 2
      "0000010" when "00110010100101111", -- t[25903] = 2
      "0000010" when "00110010100110000", -- t[25904] = 2
      "0000010" when "00110010100110001", -- t[25905] = 2
      "0000010" when "00110010100110010", -- t[25906] = 2
      "0000010" when "00110010100110011", -- t[25907] = 2
      "0000010" when "00110010100110100", -- t[25908] = 2
      "0000010" when "00110010100110101", -- t[25909] = 2
      "0000010" when "00110010100110110", -- t[25910] = 2
      "0000010" when "00110010100110111", -- t[25911] = 2
      "0000010" when "00110010100111000", -- t[25912] = 2
      "0000010" when "00110010100111001", -- t[25913] = 2
      "0000010" when "00110010100111010", -- t[25914] = 2
      "0000010" when "00110010100111011", -- t[25915] = 2
      "0000010" when "00110010100111100", -- t[25916] = 2
      "0000010" when "00110010100111101", -- t[25917] = 2
      "0000010" when "00110010100111110", -- t[25918] = 2
      "0000010" when "00110010100111111", -- t[25919] = 2
      "0000010" when "00110010101000000", -- t[25920] = 2
      "0000010" when "00110010101000001", -- t[25921] = 2
      "0000010" when "00110010101000010", -- t[25922] = 2
      "0000010" when "00110010101000011", -- t[25923] = 2
      "0000010" when "00110010101000100", -- t[25924] = 2
      "0000010" when "00110010101000101", -- t[25925] = 2
      "0000010" when "00110010101000110", -- t[25926] = 2
      "0000010" when "00110010101000111", -- t[25927] = 2
      "0000010" when "00110010101001000", -- t[25928] = 2
      "0000010" when "00110010101001001", -- t[25929] = 2
      "0000010" when "00110010101001010", -- t[25930] = 2
      "0000010" when "00110010101001011", -- t[25931] = 2
      "0000010" when "00110010101001100", -- t[25932] = 2
      "0000010" when "00110010101001101", -- t[25933] = 2
      "0000010" when "00110010101001110", -- t[25934] = 2
      "0000010" when "00110010101001111", -- t[25935] = 2
      "0000010" when "00110010101010000", -- t[25936] = 2
      "0000010" when "00110010101010001", -- t[25937] = 2
      "0000010" when "00110010101010010", -- t[25938] = 2
      "0000010" when "00110010101010011", -- t[25939] = 2
      "0000010" when "00110010101010100", -- t[25940] = 2
      "0000010" when "00110010101010101", -- t[25941] = 2
      "0000010" when "00110010101010110", -- t[25942] = 2
      "0000010" when "00110010101010111", -- t[25943] = 2
      "0000010" when "00110010101011000", -- t[25944] = 2
      "0000010" when "00110010101011001", -- t[25945] = 2
      "0000010" when "00110010101011010", -- t[25946] = 2
      "0000010" when "00110010101011011", -- t[25947] = 2
      "0000010" when "00110010101011100", -- t[25948] = 2
      "0000010" when "00110010101011101", -- t[25949] = 2
      "0000010" when "00110010101011110", -- t[25950] = 2
      "0000010" when "00110010101011111", -- t[25951] = 2
      "0000010" when "00110010101100000", -- t[25952] = 2
      "0000010" when "00110010101100001", -- t[25953] = 2
      "0000010" when "00110010101100010", -- t[25954] = 2
      "0000010" when "00110010101100011", -- t[25955] = 2
      "0000010" when "00110010101100100", -- t[25956] = 2
      "0000010" when "00110010101100101", -- t[25957] = 2
      "0000010" when "00110010101100110", -- t[25958] = 2
      "0000010" when "00110010101100111", -- t[25959] = 2
      "0000010" when "00110010101101000", -- t[25960] = 2
      "0000010" when "00110010101101001", -- t[25961] = 2
      "0000010" when "00110010101101010", -- t[25962] = 2
      "0000010" when "00110010101101011", -- t[25963] = 2
      "0000010" when "00110010101101100", -- t[25964] = 2
      "0000010" when "00110010101101101", -- t[25965] = 2
      "0000010" when "00110010101101110", -- t[25966] = 2
      "0000010" when "00110010101101111", -- t[25967] = 2
      "0000010" when "00110010101110000", -- t[25968] = 2
      "0000010" when "00110010101110001", -- t[25969] = 2
      "0000010" when "00110010101110010", -- t[25970] = 2
      "0000010" when "00110010101110011", -- t[25971] = 2
      "0000010" when "00110010101110100", -- t[25972] = 2
      "0000010" when "00110010101110101", -- t[25973] = 2
      "0000010" when "00110010101110110", -- t[25974] = 2
      "0000010" when "00110010101110111", -- t[25975] = 2
      "0000010" when "00110010101111000", -- t[25976] = 2
      "0000010" when "00110010101111001", -- t[25977] = 2
      "0000010" when "00110010101111010", -- t[25978] = 2
      "0000010" when "00110010101111011", -- t[25979] = 2
      "0000010" when "00110010101111100", -- t[25980] = 2
      "0000010" when "00110010101111101", -- t[25981] = 2
      "0000010" when "00110010101111110", -- t[25982] = 2
      "0000010" when "00110010101111111", -- t[25983] = 2
      "0000010" when "00110010110000000", -- t[25984] = 2
      "0000010" when "00110010110000001", -- t[25985] = 2
      "0000010" when "00110010110000010", -- t[25986] = 2
      "0000010" when "00110010110000011", -- t[25987] = 2
      "0000010" when "00110010110000100", -- t[25988] = 2
      "0000010" when "00110010110000101", -- t[25989] = 2
      "0000010" when "00110010110000110", -- t[25990] = 2
      "0000010" when "00110010110000111", -- t[25991] = 2
      "0000010" when "00110010110001000", -- t[25992] = 2
      "0000010" when "00110010110001001", -- t[25993] = 2
      "0000010" when "00110010110001010", -- t[25994] = 2
      "0000010" when "00110010110001011", -- t[25995] = 2
      "0000010" when "00110010110001100", -- t[25996] = 2
      "0000010" when "00110010110001101", -- t[25997] = 2
      "0000010" when "00110010110001110", -- t[25998] = 2
      "0000010" when "00110010110001111", -- t[25999] = 2
      "0000010" when "00110010110010000", -- t[26000] = 2
      "0000010" when "00110010110010001", -- t[26001] = 2
      "0000010" when "00110010110010010", -- t[26002] = 2
      "0000010" when "00110010110010011", -- t[26003] = 2
      "0000010" when "00110010110010100", -- t[26004] = 2
      "0000010" when "00110010110010101", -- t[26005] = 2
      "0000010" when "00110010110010110", -- t[26006] = 2
      "0000010" when "00110010110010111", -- t[26007] = 2
      "0000010" when "00110010110011000", -- t[26008] = 2
      "0000010" when "00110010110011001", -- t[26009] = 2
      "0000010" when "00110010110011010", -- t[26010] = 2
      "0000010" when "00110010110011011", -- t[26011] = 2
      "0000010" when "00110010110011100", -- t[26012] = 2
      "0000010" when "00110010110011101", -- t[26013] = 2
      "0000010" when "00110010110011110", -- t[26014] = 2
      "0000010" when "00110010110011111", -- t[26015] = 2
      "0000010" when "00110010110100000", -- t[26016] = 2
      "0000010" when "00110010110100001", -- t[26017] = 2
      "0000010" when "00110010110100010", -- t[26018] = 2
      "0000010" when "00110010110100011", -- t[26019] = 2
      "0000010" when "00110010110100100", -- t[26020] = 2
      "0000010" when "00110010110100101", -- t[26021] = 2
      "0000010" when "00110010110100110", -- t[26022] = 2
      "0000010" when "00110010110100111", -- t[26023] = 2
      "0000010" when "00110010110101000", -- t[26024] = 2
      "0000010" when "00110010110101001", -- t[26025] = 2
      "0000010" when "00110010110101010", -- t[26026] = 2
      "0000010" when "00110010110101011", -- t[26027] = 2
      "0000010" when "00110010110101100", -- t[26028] = 2
      "0000010" when "00110010110101101", -- t[26029] = 2
      "0000010" when "00110010110101110", -- t[26030] = 2
      "0000010" when "00110010110101111", -- t[26031] = 2
      "0000010" when "00110010110110000", -- t[26032] = 2
      "0000010" when "00110010110110001", -- t[26033] = 2
      "0000010" when "00110010110110010", -- t[26034] = 2
      "0000010" when "00110010110110011", -- t[26035] = 2
      "0000010" when "00110010110110100", -- t[26036] = 2
      "0000010" when "00110010110110101", -- t[26037] = 2
      "0000010" when "00110010110110110", -- t[26038] = 2
      "0000010" when "00110010110110111", -- t[26039] = 2
      "0000010" when "00110010110111000", -- t[26040] = 2
      "0000010" when "00110010110111001", -- t[26041] = 2
      "0000010" when "00110010110111010", -- t[26042] = 2
      "0000010" when "00110010110111011", -- t[26043] = 2
      "0000010" when "00110010110111100", -- t[26044] = 2
      "0000010" when "00110010110111101", -- t[26045] = 2
      "0000010" when "00110010110111110", -- t[26046] = 2
      "0000010" when "00110010110111111", -- t[26047] = 2
      "0000010" when "00110010111000000", -- t[26048] = 2
      "0000010" when "00110010111000001", -- t[26049] = 2
      "0000010" when "00110010111000010", -- t[26050] = 2
      "0000010" when "00110010111000011", -- t[26051] = 2
      "0000010" when "00110010111000100", -- t[26052] = 2
      "0000010" when "00110010111000101", -- t[26053] = 2
      "0000010" when "00110010111000110", -- t[26054] = 2
      "0000010" when "00110010111000111", -- t[26055] = 2
      "0000010" when "00110010111001000", -- t[26056] = 2
      "0000010" when "00110010111001001", -- t[26057] = 2
      "0000010" when "00110010111001010", -- t[26058] = 2
      "0000010" when "00110010111001011", -- t[26059] = 2
      "0000010" when "00110010111001100", -- t[26060] = 2
      "0000010" when "00110010111001101", -- t[26061] = 2
      "0000010" when "00110010111001110", -- t[26062] = 2
      "0000010" when "00110010111001111", -- t[26063] = 2
      "0000010" when "00110010111010000", -- t[26064] = 2
      "0000010" when "00110010111010001", -- t[26065] = 2
      "0000010" when "00110010111010010", -- t[26066] = 2
      "0000010" when "00110010111010011", -- t[26067] = 2
      "0000010" when "00110010111010100", -- t[26068] = 2
      "0000010" when "00110010111010101", -- t[26069] = 2
      "0000010" when "00110010111010110", -- t[26070] = 2
      "0000010" when "00110010111010111", -- t[26071] = 2
      "0000010" when "00110010111011000", -- t[26072] = 2
      "0000010" when "00110010111011001", -- t[26073] = 2
      "0000010" when "00110010111011010", -- t[26074] = 2
      "0000010" when "00110010111011011", -- t[26075] = 2
      "0000010" when "00110010111011100", -- t[26076] = 2
      "0000010" when "00110010111011101", -- t[26077] = 2
      "0000010" when "00110010111011110", -- t[26078] = 2
      "0000010" when "00110010111011111", -- t[26079] = 2
      "0000010" when "00110010111100000", -- t[26080] = 2
      "0000010" when "00110010111100001", -- t[26081] = 2
      "0000010" when "00110010111100010", -- t[26082] = 2
      "0000010" when "00110010111100011", -- t[26083] = 2
      "0000010" when "00110010111100100", -- t[26084] = 2
      "0000010" when "00110010111100101", -- t[26085] = 2
      "0000010" when "00110010111100110", -- t[26086] = 2
      "0000010" when "00110010111100111", -- t[26087] = 2
      "0000010" when "00110010111101000", -- t[26088] = 2
      "0000010" when "00110010111101001", -- t[26089] = 2
      "0000010" when "00110010111101010", -- t[26090] = 2
      "0000010" when "00110010111101011", -- t[26091] = 2
      "0000010" when "00110010111101100", -- t[26092] = 2
      "0000010" when "00110010111101101", -- t[26093] = 2
      "0000010" when "00110010111101110", -- t[26094] = 2
      "0000010" when "00110010111101111", -- t[26095] = 2
      "0000010" when "00110010111110000", -- t[26096] = 2
      "0000010" when "00110010111110001", -- t[26097] = 2
      "0000010" when "00110010111110010", -- t[26098] = 2
      "0000010" when "00110010111110011", -- t[26099] = 2
      "0000010" when "00110010111110100", -- t[26100] = 2
      "0000010" when "00110010111110101", -- t[26101] = 2
      "0000010" when "00110010111110110", -- t[26102] = 2
      "0000010" when "00110010111110111", -- t[26103] = 2
      "0000010" when "00110010111111000", -- t[26104] = 2
      "0000010" when "00110010111111001", -- t[26105] = 2
      "0000010" when "00110010111111010", -- t[26106] = 2
      "0000010" when "00110010111111011", -- t[26107] = 2
      "0000010" when "00110010111111100", -- t[26108] = 2
      "0000010" when "00110010111111101", -- t[26109] = 2
      "0000010" when "00110010111111110", -- t[26110] = 2
      "0000010" when "00110010111111111", -- t[26111] = 2
      "0000010" when "00110011000000000", -- t[26112] = 2
      "0000010" when "00110011000000001", -- t[26113] = 2
      "0000010" when "00110011000000010", -- t[26114] = 2
      "0000010" when "00110011000000011", -- t[26115] = 2
      "0000010" when "00110011000000100", -- t[26116] = 2
      "0000010" when "00110011000000101", -- t[26117] = 2
      "0000010" when "00110011000000110", -- t[26118] = 2
      "0000010" when "00110011000000111", -- t[26119] = 2
      "0000010" when "00110011000001000", -- t[26120] = 2
      "0000010" when "00110011000001001", -- t[26121] = 2
      "0000010" when "00110011000001010", -- t[26122] = 2
      "0000010" when "00110011000001011", -- t[26123] = 2
      "0000010" when "00110011000001100", -- t[26124] = 2
      "0000010" when "00110011000001101", -- t[26125] = 2
      "0000010" when "00110011000001110", -- t[26126] = 2
      "0000010" when "00110011000001111", -- t[26127] = 2
      "0000010" when "00110011000010000", -- t[26128] = 2
      "0000010" when "00110011000010001", -- t[26129] = 2
      "0000010" when "00110011000010010", -- t[26130] = 2
      "0000010" when "00110011000010011", -- t[26131] = 2
      "0000010" when "00110011000010100", -- t[26132] = 2
      "0000010" when "00110011000010101", -- t[26133] = 2
      "0000010" when "00110011000010110", -- t[26134] = 2
      "0000010" when "00110011000010111", -- t[26135] = 2
      "0000010" when "00110011000011000", -- t[26136] = 2
      "0000010" when "00110011000011001", -- t[26137] = 2
      "0000010" when "00110011000011010", -- t[26138] = 2
      "0000010" when "00110011000011011", -- t[26139] = 2
      "0000010" when "00110011000011100", -- t[26140] = 2
      "0000010" when "00110011000011101", -- t[26141] = 2
      "0000010" when "00110011000011110", -- t[26142] = 2
      "0000010" when "00110011000011111", -- t[26143] = 2
      "0000010" when "00110011000100000", -- t[26144] = 2
      "0000010" when "00110011000100001", -- t[26145] = 2
      "0000010" when "00110011000100010", -- t[26146] = 2
      "0000010" when "00110011000100011", -- t[26147] = 2
      "0000010" when "00110011000100100", -- t[26148] = 2
      "0000010" when "00110011000100101", -- t[26149] = 2
      "0000010" when "00110011000100110", -- t[26150] = 2
      "0000010" when "00110011000100111", -- t[26151] = 2
      "0000010" when "00110011000101000", -- t[26152] = 2
      "0000010" when "00110011000101001", -- t[26153] = 2
      "0000010" when "00110011000101010", -- t[26154] = 2
      "0000010" when "00110011000101011", -- t[26155] = 2
      "0000010" when "00110011000101100", -- t[26156] = 2
      "0000010" when "00110011000101101", -- t[26157] = 2
      "0000010" when "00110011000101110", -- t[26158] = 2
      "0000010" when "00110011000101111", -- t[26159] = 2
      "0000010" when "00110011000110000", -- t[26160] = 2
      "0000010" when "00110011000110001", -- t[26161] = 2
      "0000010" when "00110011000110010", -- t[26162] = 2
      "0000010" when "00110011000110011", -- t[26163] = 2
      "0000010" when "00110011000110100", -- t[26164] = 2
      "0000010" when "00110011000110101", -- t[26165] = 2
      "0000010" when "00110011000110110", -- t[26166] = 2
      "0000010" when "00110011000110111", -- t[26167] = 2
      "0000010" when "00110011000111000", -- t[26168] = 2
      "0000010" when "00110011000111001", -- t[26169] = 2
      "0000010" when "00110011000111010", -- t[26170] = 2
      "0000010" when "00110011000111011", -- t[26171] = 2
      "0000010" when "00110011000111100", -- t[26172] = 2
      "0000010" when "00110011000111101", -- t[26173] = 2
      "0000010" when "00110011000111110", -- t[26174] = 2
      "0000010" when "00110011000111111", -- t[26175] = 2
      "0000010" when "00110011001000000", -- t[26176] = 2
      "0000010" when "00110011001000001", -- t[26177] = 2
      "0000010" when "00110011001000010", -- t[26178] = 2
      "0000010" when "00110011001000011", -- t[26179] = 2
      "0000010" when "00110011001000100", -- t[26180] = 2
      "0000010" when "00110011001000101", -- t[26181] = 2
      "0000010" when "00110011001000110", -- t[26182] = 2
      "0000010" when "00110011001000111", -- t[26183] = 2
      "0000010" when "00110011001001000", -- t[26184] = 2
      "0000010" when "00110011001001001", -- t[26185] = 2
      "0000010" when "00110011001001010", -- t[26186] = 2
      "0000010" when "00110011001001011", -- t[26187] = 2
      "0000010" when "00110011001001100", -- t[26188] = 2
      "0000010" when "00110011001001101", -- t[26189] = 2
      "0000010" when "00110011001001110", -- t[26190] = 2
      "0000010" when "00110011001001111", -- t[26191] = 2
      "0000010" when "00110011001010000", -- t[26192] = 2
      "0000010" when "00110011001010001", -- t[26193] = 2
      "0000010" when "00110011001010010", -- t[26194] = 2
      "0000010" when "00110011001010011", -- t[26195] = 2
      "0000010" when "00110011001010100", -- t[26196] = 2
      "0000010" when "00110011001010101", -- t[26197] = 2
      "0000010" when "00110011001010110", -- t[26198] = 2
      "0000010" when "00110011001010111", -- t[26199] = 2
      "0000010" when "00110011001011000", -- t[26200] = 2
      "0000010" when "00110011001011001", -- t[26201] = 2
      "0000010" when "00110011001011010", -- t[26202] = 2
      "0000010" when "00110011001011011", -- t[26203] = 2
      "0000010" when "00110011001011100", -- t[26204] = 2
      "0000010" when "00110011001011101", -- t[26205] = 2
      "0000010" when "00110011001011110", -- t[26206] = 2
      "0000010" when "00110011001011111", -- t[26207] = 2
      "0000010" when "00110011001100000", -- t[26208] = 2
      "0000010" when "00110011001100001", -- t[26209] = 2
      "0000010" when "00110011001100010", -- t[26210] = 2
      "0000010" when "00110011001100011", -- t[26211] = 2
      "0000010" when "00110011001100100", -- t[26212] = 2
      "0000010" when "00110011001100101", -- t[26213] = 2
      "0000010" when "00110011001100110", -- t[26214] = 2
      "0000010" when "00110011001100111", -- t[26215] = 2
      "0000010" when "00110011001101000", -- t[26216] = 2
      "0000010" when "00110011001101001", -- t[26217] = 2
      "0000010" when "00110011001101010", -- t[26218] = 2
      "0000010" when "00110011001101011", -- t[26219] = 2
      "0000010" when "00110011001101100", -- t[26220] = 2
      "0000010" when "00110011001101101", -- t[26221] = 2
      "0000010" when "00110011001101110", -- t[26222] = 2
      "0000010" when "00110011001101111", -- t[26223] = 2
      "0000010" when "00110011001110000", -- t[26224] = 2
      "0000010" when "00110011001110001", -- t[26225] = 2
      "0000010" when "00110011001110010", -- t[26226] = 2
      "0000010" when "00110011001110011", -- t[26227] = 2
      "0000010" when "00110011001110100", -- t[26228] = 2
      "0000010" when "00110011001110101", -- t[26229] = 2
      "0000010" when "00110011001110110", -- t[26230] = 2
      "0000010" when "00110011001110111", -- t[26231] = 2
      "0000010" when "00110011001111000", -- t[26232] = 2
      "0000010" when "00110011001111001", -- t[26233] = 2
      "0000010" when "00110011001111010", -- t[26234] = 2
      "0000010" when "00110011001111011", -- t[26235] = 2
      "0000010" when "00110011001111100", -- t[26236] = 2
      "0000010" when "00110011001111101", -- t[26237] = 2
      "0000010" when "00110011001111110", -- t[26238] = 2
      "0000010" when "00110011001111111", -- t[26239] = 2
      "0000010" when "00110011010000000", -- t[26240] = 2
      "0000010" when "00110011010000001", -- t[26241] = 2
      "0000010" when "00110011010000010", -- t[26242] = 2
      "0000010" when "00110011010000011", -- t[26243] = 2
      "0000010" when "00110011010000100", -- t[26244] = 2
      "0000010" when "00110011010000101", -- t[26245] = 2
      "0000010" when "00110011010000110", -- t[26246] = 2
      "0000010" when "00110011010000111", -- t[26247] = 2
      "0000010" when "00110011010001000", -- t[26248] = 2
      "0000010" when "00110011010001001", -- t[26249] = 2
      "0000010" when "00110011010001010", -- t[26250] = 2
      "0000010" when "00110011010001011", -- t[26251] = 2
      "0000010" when "00110011010001100", -- t[26252] = 2
      "0000010" when "00110011010001101", -- t[26253] = 2
      "0000010" when "00110011010001110", -- t[26254] = 2
      "0000010" when "00110011010001111", -- t[26255] = 2
      "0000010" when "00110011010010000", -- t[26256] = 2
      "0000010" when "00110011010010001", -- t[26257] = 2
      "0000010" when "00110011010010010", -- t[26258] = 2
      "0000010" when "00110011010010011", -- t[26259] = 2
      "0000010" when "00110011010010100", -- t[26260] = 2
      "0000010" when "00110011010010101", -- t[26261] = 2
      "0000010" when "00110011010010110", -- t[26262] = 2
      "0000010" when "00110011010010111", -- t[26263] = 2
      "0000010" when "00110011010011000", -- t[26264] = 2
      "0000010" when "00110011010011001", -- t[26265] = 2
      "0000010" when "00110011010011010", -- t[26266] = 2
      "0000010" when "00110011010011011", -- t[26267] = 2
      "0000010" when "00110011010011100", -- t[26268] = 2
      "0000010" when "00110011010011101", -- t[26269] = 2
      "0000010" when "00110011010011110", -- t[26270] = 2
      "0000010" when "00110011010011111", -- t[26271] = 2
      "0000010" when "00110011010100000", -- t[26272] = 2
      "0000010" when "00110011010100001", -- t[26273] = 2
      "0000010" when "00110011010100010", -- t[26274] = 2
      "0000010" when "00110011010100011", -- t[26275] = 2
      "0000010" when "00110011010100100", -- t[26276] = 2
      "0000010" when "00110011010100101", -- t[26277] = 2
      "0000010" when "00110011010100110", -- t[26278] = 2
      "0000010" when "00110011010100111", -- t[26279] = 2
      "0000010" when "00110011010101000", -- t[26280] = 2
      "0000010" when "00110011010101001", -- t[26281] = 2
      "0000010" when "00110011010101010", -- t[26282] = 2
      "0000010" when "00110011010101011", -- t[26283] = 2
      "0000010" when "00110011010101100", -- t[26284] = 2
      "0000010" when "00110011010101101", -- t[26285] = 2
      "0000010" when "00110011010101110", -- t[26286] = 2
      "0000010" when "00110011010101111", -- t[26287] = 2
      "0000010" when "00110011010110000", -- t[26288] = 2
      "0000010" when "00110011010110001", -- t[26289] = 2
      "0000010" when "00110011010110010", -- t[26290] = 2
      "0000010" when "00110011010110011", -- t[26291] = 2
      "0000010" when "00110011010110100", -- t[26292] = 2
      "0000010" when "00110011010110101", -- t[26293] = 2
      "0000010" when "00110011010110110", -- t[26294] = 2
      "0000010" when "00110011010110111", -- t[26295] = 2
      "0000010" when "00110011010111000", -- t[26296] = 2
      "0000010" when "00110011010111001", -- t[26297] = 2
      "0000010" when "00110011010111010", -- t[26298] = 2
      "0000010" when "00110011010111011", -- t[26299] = 2
      "0000010" when "00110011010111100", -- t[26300] = 2
      "0000010" when "00110011010111101", -- t[26301] = 2
      "0000010" when "00110011010111110", -- t[26302] = 2
      "0000010" when "00110011010111111", -- t[26303] = 2
      "0000010" when "00110011011000000", -- t[26304] = 2
      "0000010" when "00110011011000001", -- t[26305] = 2
      "0000010" when "00110011011000010", -- t[26306] = 2
      "0000010" when "00110011011000011", -- t[26307] = 2
      "0000010" when "00110011011000100", -- t[26308] = 2
      "0000010" when "00110011011000101", -- t[26309] = 2
      "0000010" when "00110011011000110", -- t[26310] = 2
      "0000010" when "00110011011000111", -- t[26311] = 2
      "0000010" when "00110011011001000", -- t[26312] = 2
      "0000010" when "00110011011001001", -- t[26313] = 2
      "0000010" when "00110011011001010", -- t[26314] = 2
      "0000010" when "00110011011001011", -- t[26315] = 2
      "0000010" when "00110011011001100", -- t[26316] = 2
      "0000010" when "00110011011001101", -- t[26317] = 2
      "0000010" when "00110011011001110", -- t[26318] = 2
      "0000010" when "00110011011001111", -- t[26319] = 2
      "0000010" when "00110011011010000", -- t[26320] = 2
      "0000010" when "00110011011010001", -- t[26321] = 2
      "0000010" when "00110011011010010", -- t[26322] = 2
      "0000010" when "00110011011010011", -- t[26323] = 2
      "0000010" when "00110011011010100", -- t[26324] = 2
      "0000010" when "00110011011010101", -- t[26325] = 2
      "0000010" when "00110011011010110", -- t[26326] = 2
      "0000010" when "00110011011010111", -- t[26327] = 2
      "0000010" when "00110011011011000", -- t[26328] = 2
      "0000010" when "00110011011011001", -- t[26329] = 2
      "0000010" when "00110011011011010", -- t[26330] = 2
      "0000010" when "00110011011011011", -- t[26331] = 2
      "0000010" when "00110011011011100", -- t[26332] = 2
      "0000010" when "00110011011011101", -- t[26333] = 2
      "0000010" when "00110011011011110", -- t[26334] = 2
      "0000010" when "00110011011011111", -- t[26335] = 2
      "0000010" when "00110011011100000", -- t[26336] = 2
      "0000010" when "00110011011100001", -- t[26337] = 2
      "0000010" when "00110011011100010", -- t[26338] = 2
      "0000010" when "00110011011100011", -- t[26339] = 2
      "0000010" when "00110011011100100", -- t[26340] = 2
      "0000010" when "00110011011100101", -- t[26341] = 2
      "0000010" when "00110011011100110", -- t[26342] = 2
      "0000010" when "00110011011100111", -- t[26343] = 2
      "0000010" when "00110011011101000", -- t[26344] = 2
      "0000010" when "00110011011101001", -- t[26345] = 2
      "0000010" when "00110011011101010", -- t[26346] = 2
      "0000010" when "00110011011101011", -- t[26347] = 2
      "0000010" when "00110011011101100", -- t[26348] = 2
      "0000010" when "00110011011101101", -- t[26349] = 2
      "0000010" when "00110011011101110", -- t[26350] = 2
      "0000010" when "00110011011101111", -- t[26351] = 2
      "0000010" when "00110011011110000", -- t[26352] = 2
      "0000010" when "00110011011110001", -- t[26353] = 2
      "0000010" when "00110011011110010", -- t[26354] = 2
      "0000010" when "00110011011110011", -- t[26355] = 2
      "0000010" when "00110011011110100", -- t[26356] = 2
      "0000010" when "00110011011110101", -- t[26357] = 2
      "0000010" when "00110011011110110", -- t[26358] = 2
      "0000010" when "00110011011110111", -- t[26359] = 2
      "0000010" when "00110011011111000", -- t[26360] = 2
      "0000010" when "00110011011111001", -- t[26361] = 2
      "0000010" when "00110011011111010", -- t[26362] = 2
      "0000010" when "00110011011111011", -- t[26363] = 2
      "0000010" when "00110011011111100", -- t[26364] = 2
      "0000010" when "00110011011111101", -- t[26365] = 2
      "0000010" when "00110011011111110", -- t[26366] = 2
      "0000010" when "00110011011111111", -- t[26367] = 2
      "0000010" when "00110011100000000", -- t[26368] = 2
      "0000010" when "00110011100000001", -- t[26369] = 2
      "0000010" when "00110011100000010", -- t[26370] = 2
      "0000010" when "00110011100000011", -- t[26371] = 2
      "0000010" when "00110011100000100", -- t[26372] = 2
      "0000010" when "00110011100000101", -- t[26373] = 2
      "0000010" when "00110011100000110", -- t[26374] = 2
      "0000010" when "00110011100000111", -- t[26375] = 2
      "0000010" when "00110011100001000", -- t[26376] = 2
      "0000010" when "00110011100001001", -- t[26377] = 2
      "0000010" when "00110011100001010", -- t[26378] = 2
      "0000010" when "00110011100001011", -- t[26379] = 2
      "0000010" when "00110011100001100", -- t[26380] = 2
      "0000010" when "00110011100001101", -- t[26381] = 2
      "0000010" when "00110011100001110", -- t[26382] = 2
      "0000010" when "00110011100001111", -- t[26383] = 2
      "0000010" when "00110011100010000", -- t[26384] = 2
      "0000010" when "00110011100010001", -- t[26385] = 2
      "0000010" when "00110011100010010", -- t[26386] = 2
      "0000010" when "00110011100010011", -- t[26387] = 2
      "0000010" when "00110011100010100", -- t[26388] = 2
      "0000010" when "00110011100010101", -- t[26389] = 2
      "0000010" when "00110011100010110", -- t[26390] = 2
      "0000010" when "00110011100010111", -- t[26391] = 2
      "0000010" when "00110011100011000", -- t[26392] = 2
      "0000010" when "00110011100011001", -- t[26393] = 2
      "0000010" when "00110011100011010", -- t[26394] = 2
      "0000010" when "00110011100011011", -- t[26395] = 2
      "0000010" when "00110011100011100", -- t[26396] = 2
      "0000010" when "00110011100011101", -- t[26397] = 2
      "0000010" when "00110011100011110", -- t[26398] = 2
      "0000010" when "00110011100011111", -- t[26399] = 2
      "0000010" when "00110011100100000", -- t[26400] = 2
      "0000010" when "00110011100100001", -- t[26401] = 2
      "0000010" when "00110011100100010", -- t[26402] = 2
      "0000010" when "00110011100100011", -- t[26403] = 2
      "0000010" when "00110011100100100", -- t[26404] = 2
      "0000010" when "00110011100100101", -- t[26405] = 2
      "0000010" when "00110011100100110", -- t[26406] = 2
      "0000010" when "00110011100100111", -- t[26407] = 2
      "0000010" when "00110011100101000", -- t[26408] = 2
      "0000010" when "00110011100101001", -- t[26409] = 2
      "0000010" when "00110011100101010", -- t[26410] = 2
      "0000010" when "00110011100101011", -- t[26411] = 2
      "0000010" when "00110011100101100", -- t[26412] = 2
      "0000010" when "00110011100101101", -- t[26413] = 2
      "0000010" when "00110011100101110", -- t[26414] = 2
      "0000010" when "00110011100101111", -- t[26415] = 2
      "0000010" when "00110011100110000", -- t[26416] = 2
      "0000010" when "00110011100110001", -- t[26417] = 2
      "0000010" when "00110011100110010", -- t[26418] = 2
      "0000010" when "00110011100110011", -- t[26419] = 2
      "0000010" when "00110011100110100", -- t[26420] = 2
      "0000010" when "00110011100110101", -- t[26421] = 2
      "0000010" when "00110011100110110", -- t[26422] = 2
      "0000010" when "00110011100110111", -- t[26423] = 2
      "0000010" when "00110011100111000", -- t[26424] = 2
      "0000010" when "00110011100111001", -- t[26425] = 2
      "0000010" when "00110011100111010", -- t[26426] = 2
      "0000010" when "00110011100111011", -- t[26427] = 2
      "0000010" when "00110011100111100", -- t[26428] = 2
      "0000010" when "00110011100111101", -- t[26429] = 2
      "0000010" when "00110011100111110", -- t[26430] = 2
      "0000010" when "00110011100111111", -- t[26431] = 2
      "0000010" when "00110011101000000", -- t[26432] = 2
      "0000010" when "00110011101000001", -- t[26433] = 2
      "0000010" when "00110011101000010", -- t[26434] = 2
      "0000010" when "00110011101000011", -- t[26435] = 2
      "0000010" when "00110011101000100", -- t[26436] = 2
      "0000010" when "00110011101000101", -- t[26437] = 2
      "0000010" when "00110011101000110", -- t[26438] = 2
      "0000010" when "00110011101000111", -- t[26439] = 2
      "0000010" when "00110011101001000", -- t[26440] = 2
      "0000010" when "00110011101001001", -- t[26441] = 2
      "0000010" when "00110011101001010", -- t[26442] = 2
      "0000010" when "00110011101001011", -- t[26443] = 2
      "0000010" when "00110011101001100", -- t[26444] = 2
      "0000010" when "00110011101001101", -- t[26445] = 2
      "0000010" when "00110011101001110", -- t[26446] = 2
      "0000010" when "00110011101001111", -- t[26447] = 2
      "0000010" when "00110011101010000", -- t[26448] = 2
      "0000010" when "00110011101010001", -- t[26449] = 2
      "0000010" when "00110011101010010", -- t[26450] = 2
      "0000010" when "00110011101010011", -- t[26451] = 2
      "0000010" when "00110011101010100", -- t[26452] = 2
      "0000010" when "00110011101010101", -- t[26453] = 2
      "0000010" when "00110011101010110", -- t[26454] = 2
      "0000010" when "00110011101010111", -- t[26455] = 2
      "0000010" when "00110011101011000", -- t[26456] = 2
      "0000010" when "00110011101011001", -- t[26457] = 2
      "0000010" when "00110011101011010", -- t[26458] = 2
      "0000010" when "00110011101011011", -- t[26459] = 2
      "0000010" when "00110011101011100", -- t[26460] = 2
      "0000010" when "00110011101011101", -- t[26461] = 2
      "0000010" when "00110011101011110", -- t[26462] = 2
      "0000010" when "00110011101011111", -- t[26463] = 2
      "0000010" when "00110011101100000", -- t[26464] = 2
      "0000010" when "00110011101100001", -- t[26465] = 2
      "0000010" when "00110011101100010", -- t[26466] = 2
      "0000010" when "00110011101100011", -- t[26467] = 2
      "0000010" when "00110011101100100", -- t[26468] = 2
      "0000010" when "00110011101100101", -- t[26469] = 2
      "0000010" when "00110011101100110", -- t[26470] = 2
      "0000010" when "00110011101100111", -- t[26471] = 2
      "0000010" when "00110011101101000", -- t[26472] = 2
      "0000010" when "00110011101101001", -- t[26473] = 2
      "0000010" when "00110011101101010", -- t[26474] = 2
      "0000010" when "00110011101101011", -- t[26475] = 2
      "0000010" when "00110011101101100", -- t[26476] = 2
      "0000010" when "00110011101101101", -- t[26477] = 2
      "0000010" when "00110011101101110", -- t[26478] = 2
      "0000010" when "00110011101101111", -- t[26479] = 2
      "0000010" when "00110011101110000", -- t[26480] = 2
      "0000010" when "00110011101110001", -- t[26481] = 2
      "0000010" when "00110011101110010", -- t[26482] = 2
      "0000010" when "00110011101110011", -- t[26483] = 2
      "0000010" when "00110011101110100", -- t[26484] = 2
      "0000010" when "00110011101110101", -- t[26485] = 2
      "0000010" when "00110011101110110", -- t[26486] = 2
      "0000010" when "00110011101110111", -- t[26487] = 2
      "0000010" when "00110011101111000", -- t[26488] = 2
      "0000010" when "00110011101111001", -- t[26489] = 2
      "0000010" when "00110011101111010", -- t[26490] = 2
      "0000010" when "00110011101111011", -- t[26491] = 2
      "0000010" when "00110011101111100", -- t[26492] = 2
      "0000010" when "00110011101111101", -- t[26493] = 2
      "0000010" when "00110011101111110", -- t[26494] = 2
      "0000010" when "00110011101111111", -- t[26495] = 2
      "0000010" when "00110011110000000", -- t[26496] = 2
      "0000010" when "00110011110000001", -- t[26497] = 2
      "0000010" when "00110011110000010", -- t[26498] = 2
      "0000010" when "00110011110000011", -- t[26499] = 2
      "0000010" when "00110011110000100", -- t[26500] = 2
      "0000010" when "00110011110000101", -- t[26501] = 2
      "0000010" when "00110011110000110", -- t[26502] = 2
      "0000010" when "00110011110000111", -- t[26503] = 2
      "0000010" when "00110011110001000", -- t[26504] = 2
      "0000010" when "00110011110001001", -- t[26505] = 2
      "0000010" when "00110011110001010", -- t[26506] = 2
      "0000010" when "00110011110001011", -- t[26507] = 2
      "0000010" when "00110011110001100", -- t[26508] = 2
      "0000010" when "00110011110001101", -- t[26509] = 2
      "0000010" when "00110011110001110", -- t[26510] = 2
      "0000010" when "00110011110001111", -- t[26511] = 2
      "0000010" when "00110011110010000", -- t[26512] = 2
      "0000010" when "00110011110010001", -- t[26513] = 2
      "0000010" when "00110011110010010", -- t[26514] = 2
      "0000010" when "00110011110010011", -- t[26515] = 2
      "0000010" when "00110011110010100", -- t[26516] = 2
      "0000010" when "00110011110010101", -- t[26517] = 2
      "0000010" when "00110011110010110", -- t[26518] = 2
      "0000010" when "00110011110010111", -- t[26519] = 2
      "0000010" when "00110011110011000", -- t[26520] = 2
      "0000010" when "00110011110011001", -- t[26521] = 2
      "0000010" when "00110011110011010", -- t[26522] = 2
      "0000010" when "00110011110011011", -- t[26523] = 2
      "0000010" when "00110011110011100", -- t[26524] = 2
      "0000010" when "00110011110011101", -- t[26525] = 2
      "0000010" when "00110011110011110", -- t[26526] = 2
      "0000010" when "00110011110011111", -- t[26527] = 2
      "0000010" when "00110011110100000", -- t[26528] = 2
      "0000010" when "00110011110100001", -- t[26529] = 2
      "0000010" when "00110011110100010", -- t[26530] = 2
      "0000010" when "00110011110100011", -- t[26531] = 2
      "0000010" when "00110011110100100", -- t[26532] = 2
      "0000010" when "00110011110100101", -- t[26533] = 2
      "0000010" when "00110011110100110", -- t[26534] = 2
      "0000010" when "00110011110100111", -- t[26535] = 2
      "0000010" when "00110011110101000", -- t[26536] = 2
      "0000010" when "00110011110101001", -- t[26537] = 2
      "0000010" when "00110011110101010", -- t[26538] = 2
      "0000010" when "00110011110101011", -- t[26539] = 2
      "0000010" when "00110011110101100", -- t[26540] = 2
      "0000010" when "00110011110101101", -- t[26541] = 2
      "0000010" when "00110011110101110", -- t[26542] = 2
      "0000010" when "00110011110101111", -- t[26543] = 2
      "0000010" when "00110011110110000", -- t[26544] = 2
      "0000010" when "00110011110110001", -- t[26545] = 2
      "0000010" when "00110011110110010", -- t[26546] = 2
      "0000010" when "00110011110110011", -- t[26547] = 2
      "0000010" when "00110011110110100", -- t[26548] = 2
      "0000010" when "00110011110110101", -- t[26549] = 2
      "0000010" when "00110011110110110", -- t[26550] = 2
      "0000010" when "00110011110110111", -- t[26551] = 2
      "0000010" when "00110011110111000", -- t[26552] = 2
      "0000010" when "00110011110111001", -- t[26553] = 2
      "0000010" when "00110011110111010", -- t[26554] = 2
      "0000010" when "00110011110111011", -- t[26555] = 2
      "0000010" when "00110011110111100", -- t[26556] = 2
      "0000010" when "00110011110111101", -- t[26557] = 2
      "0000010" when "00110011110111110", -- t[26558] = 2
      "0000010" when "00110011110111111", -- t[26559] = 2
      "0000010" when "00110011111000000", -- t[26560] = 2
      "0000010" when "00110011111000001", -- t[26561] = 2
      "0000010" when "00110011111000010", -- t[26562] = 2
      "0000010" when "00110011111000011", -- t[26563] = 2
      "0000010" when "00110011111000100", -- t[26564] = 2
      "0000010" when "00110011111000101", -- t[26565] = 2
      "0000010" when "00110011111000110", -- t[26566] = 2
      "0000010" when "00110011111000111", -- t[26567] = 2
      "0000010" when "00110011111001000", -- t[26568] = 2
      "0000010" when "00110011111001001", -- t[26569] = 2
      "0000010" when "00110011111001010", -- t[26570] = 2
      "0000010" when "00110011111001011", -- t[26571] = 2
      "0000010" when "00110011111001100", -- t[26572] = 2
      "0000010" when "00110011111001101", -- t[26573] = 2
      "0000010" when "00110011111001110", -- t[26574] = 2
      "0000010" when "00110011111001111", -- t[26575] = 2
      "0000010" when "00110011111010000", -- t[26576] = 2
      "0000010" when "00110011111010001", -- t[26577] = 2
      "0000010" when "00110011111010010", -- t[26578] = 2
      "0000010" when "00110011111010011", -- t[26579] = 2
      "0000010" when "00110011111010100", -- t[26580] = 2
      "0000010" when "00110011111010101", -- t[26581] = 2
      "0000010" when "00110011111010110", -- t[26582] = 2
      "0000010" when "00110011111010111", -- t[26583] = 2
      "0000010" when "00110011111011000", -- t[26584] = 2
      "0000010" when "00110011111011001", -- t[26585] = 2
      "0000010" when "00110011111011010", -- t[26586] = 2
      "0000010" when "00110011111011011", -- t[26587] = 2
      "0000010" when "00110011111011100", -- t[26588] = 2
      "0000010" when "00110011111011101", -- t[26589] = 2
      "0000010" when "00110011111011110", -- t[26590] = 2
      "0000010" when "00110011111011111", -- t[26591] = 2
      "0000010" when "00110011111100000", -- t[26592] = 2
      "0000010" when "00110011111100001", -- t[26593] = 2
      "0000010" when "00110011111100010", -- t[26594] = 2
      "0000010" when "00110011111100011", -- t[26595] = 2
      "0000010" when "00110011111100100", -- t[26596] = 2
      "0000010" when "00110011111100101", -- t[26597] = 2
      "0000010" when "00110011111100110", -- t[26598] = 2
      "0000010" when "00110011111100111", -- t[26599] = 2
      "0000010" when "00110011111101000", -- t[26600] = 2
      "0000010" when "00110011111101001", -- t[26601] = 2
      "0000010" when "00110011111101010", -- t[26602] = 2
      "0000010" when "00110011111101011", -- t[26603] = 2
      "0000010" when "00110011111101100", -- t[26604] = 2
      "0000010" when "00110011111101101", -- t[26605] = 2
      "0000010" when "00110011111101110", -- t[26606] = 2
      "0000010" when "00110011111101111", -- t[26607] = 2
      "0000010" when "00110011111110000", -- t[26608] = 2
      "0000010" when "00110011111110001", -- t[26609] = 2
      "0000010" when "00110011111110010", -- t[26610] = 2
      "0000010" when "00110011111110011", -- t[26611] = 2
      "0000010" when "00110011111110100", -- t[26612] = 2
      "0000010" when "00110011111110101", -- t[26613] = 2
      "0000010" when "00110011111110110", -- t[26614] = 2
      "0000010" when "00110011111110111", -- t[26615] = 2
      "0000010" when "00110011111111000", -- t[26616] = 2
      "0000010" when "00110011111111001", -- t[26617] = 2
      "0000010" when "00110011111111010", -- t[26618] = 2
      "0000010" when "00110011111111011", -- t[26619] = 2
      "0000010" when "00110011111111100", -- t[26620] = 2
      "0000010" when "00110011111111101", -- t[26621] = 2
      "0000010" when "00110011111111110", -- t[26622] = 2
      "0000010" when "00110011111111111", -- t[26623] = 2
      "0000010" when "00110100000000000", -- t[26624] = 2
      "0000010" when "00110100000000001", -- t[26625] = 2
      "0000010" when "00110100000000010", -- t[26626] = 2
      "0000010" when "00110100000000011", -- t[26627] = 2
      "0000010" when "00110100000000100", -- t[26628] = 2
      "0000010" when "00110100000000101", -- t[26629] = 2
      "0000010" when "00110100000000110", -- t[26630] = 2
      "0000010" when "00110100000000111", -- t[26631] = 2
      "0000010" when "00110100000001000", -- t[26632] = 2
      "0000010" when "00110100000001001", -- t[26633] = 2
      "0000010" when "00110100000001010", -- t[26634] = 2
      "0000010" when "00110100000001011", -- t[26635] = 2
      "0000010" when "00110100000001100", -- t[26636] = 2
      "0000010" when "00110100000001101", -- t[26637] = 2
      "0000010" when "00110100000001110", -- t[26638] = 2
      "0000010" when "00110100000001111", -- t[26639] = 2
      "0000010" when "00110100000010000", -- t[26640] = 2
      "0000010" when "00110100000010001", -- t[26641] = 2
      "0000010" when "00110100000010010", -- t[26642] = 2
      "0000010" when "00110100000010011", -- t[26643] = 2
      "0000010" when "00110100000010100", -- t[26644] = 2
      "0000010" when "00110100000010101", -- t[26645] = 2
      "0000010" when "00110100000010110", -- t[26646] = 2
      "0000010" when "00110100000010111", -- t[26647] = 2
      "0000010" when "00110100000011000", -- t[26648] = 2
      "0000010" when "00110100000011001", -- t[26649] = 2
      "0000010" when "00110100000011010", -- t[26650] = 2
      "0000010" when "00110100000011011", -- t[26651] = 2
      "0000010" when "00110100000011100", -- t[26652] = 2
      "0000010" when "00110100000011101", -- t[26653] = 2
      "0000010" when "00110100000011110", -- t[26654] = 2
      "0000010" when "00110100000011111", -- t[26655] = 2
      "0000010" when "00110100000100000", -- t[26656] = 2
      "0000010" when "00110100000100001", -- t[26657] = 2
      "0000010" when "00110100000100010", -- t[26658] = 2
      "0000010" when "00110100000100011", -- t[26659] = 2
      "0000010" when "00110100000100100", -- t[26660] = 2
      "0000010" when "00110100000100101", -- t[26661] = 2
      "0000010" when "00110100000100110", -- t[26662] = 2
      "0000010" when "00110100000100111", -- t[26663] = 2
      "0000010" when "00110100000101000", -- t[26664] = 2
      "0000010" when "00110100000101001", -- t[26665] = 2
      "0000010" when "00110100000101010", -- t[26666] = 2
      "0000010" when "00110100000101011", -- t[26667] = 2
      "0000010" when "00110100000101100", -- t[26668] = 2
      "0000010" when "00110100000101101", -- t[26669] = 2
      "0000010" when "00110100000101110", -- t[26670] = 2
      "0000010" when "00110100000101111", -- t[26671] = 2
      "0000010" when "00110100000110000", -- t[26672] = 2
      "0000010" when "00110100000110001", -- t[26673] = 2
      "0000010" when "00110100000110010", -- t[26674] = 2
      "0000010" when "00110100000110011", -- t[26675] = 2
      "0000010" when "00110100000110100", -- t[26676] = 2
      "0000010" when "00110100000110101", -- t[26677] = 2
      "0000010" when "00110100000110110", -- t[26678] = 2
      "0000010" when "00110100000110111", -- t[26679] = 2
      "0000010" when "00110100000111000", -- t[26680] = 2
      "0000010" when "00110100000111001", -- t[26681] = 2
      "0000010" when "00110100000111010", -- t[26682] = 2
      "0000010" when "00110100000111011", -- t[26683] = 2
      "0000010" when "00110100000111100", -- t[26684] = 2
      "0000010" when "00110100000111101", -- t[26685] = 2
      "0000010" when "00110100000111110", -- t[26686] = 2
      "0000010" when "00110100000111111", -- t[26687] = 2
      "0000010" when "00110100001000000", -- t[26688] = 2
      "0000010" when "00110100001000001", -- t[26689] = 2
      "0000010" when "00110100001000010", -- t[26690] = 2
      "0000010" when "00110100001000011", -- t[26691] = 2
      "0000010" when "00110100001000100", -- t[26692] = 2
      "0000010" when "00110100001000101", -- t[26693] = 2
      "0000010" when "00110100001000110", -- t[26694] = 2
      "0000010" when "00110100001000111", -- t[26695] = 2
      "0000010" when "00110100001001000", -- t[26696] = 2
      "0000010" when "00110100001001001", -- t[26697] = 2
      "0000010" when "00110100001001010", -- t[26698] = 2
      "0000010" when "00110100001001011", -- t[26699] = 2
      "0000010" when "00110100001001100", -- t[26700] = 2
      "0000010" when "00110100001001101", -- t[26701] = 2
      "0000010" when "00110100001001110", -- t[26702] = 2
      "0000010" when "00110100001001111", -- t[26703] = 2
      "0000010" when "00110100001010000", -- t[26704] = 2
      "0000010" when "00110100001010001", -- t[26705] = 2
      "0000010" when "00110100001010010", -- t[26706] = 2
      "0000010" when "00110100001010011", -- t[26707] = 2
      "0000010" when "00110100001010100", -- t[26708] = 2
      "0000010" when "00110100001010101", -- t[26709] = 2
      "0000010" when "00110100001010110", -- t[26710] = 2
      "0000010" when "00110100001010111", -- t[26711] = 2
      "0000010" when "00110100001011000", -- t[26712] = 2
      "0000010" when "00110100001011001", -- t[26713] = 2
      "0000010" when "00110100001011010", -- t[26714] = 2
      "0000010" when "00110100001011011", -- t[26715] = 2
      "0000010" when "00110100001011100", -- t[26716] = 2
      "0000010" when "00110100001011101", -- t[26717] = 2
      "0000010" when "00110100001011110", -- t[26718] = 2
      "0000010" when "00110100001011111", -- t[26719] = 2
      "0000010" when "00110100001100000", -- t[26720] = 2
      "0000010" when "00110100001100001", -- t[26721] = 2
      "0000010" when "00110100001100010", -- t[26722] = 2
      "0000010" when "00110100001100011", -- t[26723] = 2
      "0000010" when "00110100001100100", -- t[26724] = 2
      "0000010" when "00110100001100101", -- t[26725] = 2
      "0000010" when "00110100001100110", -- t[26726] = 2
      "0000010" when "00110100001100111", -- t[26727] = 2
      "0000010" when "00110100001101000", -- t[26728] = 2
      "0000010" when "00110100001101001", -- t[26729] = 2
      "0000010" when "00110100001101010", -- t[26730] = 2
      "0000010" when "00110100001101011", -- t[26731] = 2
      "0000010" when "00110100001101100", -- t[26732] = 2
      "0000010" when "00110100001101101", -- t[26733] = 2
      "0000010" when "00110100001101110", -- t[26734] = 2
      "0000010" when "00110100001101111", -- t[26735] = 2
      "0000010" when "00110100001110000", -- t[26736] = 2
      "0000010" when "00110100001110001", -- t[26737] = 2
      "0000010" when "00110100001110010", -- t[26738] = 2
      "0000010" when "00110100001110011", -- t[26739] = 2
      "0000010" when "00110100001110100", -- t[26740] = 2
      "0000010" when "00110100001110101", -- t[26741] = 2
      "0000010" when "00110100001110110", -- t[26742] = 2
      "0000010" when "00110100001110111", -- t[26743] = 2
      "0000010" when "00110100001111000", -- t[26744] = 2
      "0000010" when "00110100001111001", -- t[26745] = 2
      "0000010" when "00110100001111010", -- t[26746] = 2
      "0000010" when "00110100001111011", -- t[26747] = 2
      "0000010" when "00110100001111100", -- t[26748] = 2
      "0000010" when "00110100001111101", -- t[26749] = 2
      "0000010" when "00110100001111110", -- t[26750] = 2
      "0000010" when "00110100001111111", -- t[26751] = 2
      "0000010" when "00110100010000000", -- t[26752] = 2
      "0000010" when "00110100010000001", -- t[26753] = 2
      "0000010" when "00110100010000010", -- t[26754] = 2
      "0000010" when "00110100010000011", -- t[26755] = 2
      "0000010" when "00110100010000100", -- t[26756] = 2
      "0000010" when "00110100010000101", -- t[26757] = 2
      "0000010" when "00110100010000110", -- t[26758] = 2
      "0000010" when "00110100010000111", -- t[26759] = 2
      "0000010" when "00110100010001000", -- t[26760] = 2
      "0000010" when "00110100010001001", -- t[26761] = 2
      "0000010" when "00110100010001010", -- t[26762] = 2
      "0000010" when "00110100010001011", -- t[26763] = 2
      "0000010" when "00110100010001100", -- t[26764] = 2
      "0000010" when "00110100010001101", -- t[26765] = 2
      "0000010" when "00110100010001110", -- t[26766] = 2
      "0000010" when "00110100010001111", -- t[26767] = 2
      "0000010" when "00110100010010000", -- t[26768] = 2
      "0000010" when "00110100010010001", -- t[26769] = 2
      "0000010" when "00110100010010010", -- t[26770] = 2
      "0000010" when "00110100010010011", -- t[26771] = 2
      "0000010" when "00110100010010100", -- t[26772] = 2
      "0000010" when "00110100010010101", -- t[26773] = 2
      "0000010" when "00110100010010110", -- t[26774] = 2
      "0000010" when "00110100010010111", -- t[26775] = 2
      "0000010" when "00110100010011000", -- t[26776] = 2
      "0000010" when "00110100010011001", -- t[26777] = 2
      "0000010" when "00110100010011010", -- t[26778] = 2
      "0000010" when "00110100010011011", -- t[26779] = 2
      "0000010" when "00110100010011100", -- t[26780] = 2
      "0000010" when "00110100010011101", -- t[26781] = 2
      "0000010" when "00110100010011110", -- t[26782] = 2
      "0000010" when "00110100010011111", -- t[26783] = 2
      "0000010" when "00110100010100000", -- t[26784] = 2
      "0000010" when "00110100010100001", -- t[26785] = 2
      "0000010" when "00110100010100010", -- t[26786] = 2
      "0000010" when "00110100010100011", -- t[26787] = 2
      "0000010" when "00110100010100100", -- t[26788] = 2
      "0000010" when "00110100010100101", -- t[26789] = 2
      "0000010" when "00110100010100110", -- t[26790] = 2
      "0000010" when "00110100010100111", -- t[26791] = 2
      "0000010" when "00110100010101000", -- t[26792] = 2
      "0000010" when "00110100010101001", -- t[26793] = 2
      "0000010" when "00110100010101010", -- t[26794] = 2
      "0000010" when "00110100010101011", -- t[26795] = 2
      "0000010" when "00110100010101100", -- t[26796] = 2
      "0000010" when "00110100010101101", -- t[26797] = 2
      "0000010" when "00110100010101110", -- t[26798] = 2
      "0000010" when "00110100010101111", -- t[26799] = 2
      "0000010" when "00110100010110000", -- t[26800] = 2
      "0000010" when "00110100010110001", -- t[26801] = 2
      "0000010" when "00110100010110010", -- t[26802] = 2
      "0000010" when "00110100010110011", -- t[26803] = 2
      "0000010" when "00110100010110100", -- t[26804] = 2
      "0000010" when "00110100010110101", -- t[26805] = 2
      "0000010" when "00110100010110110", -- t[26806] = 2
      "0000010" when "00110100010110111", -- t[26807] = 2
      "0000010" when "00110100010111000", -- t[26808] = 2
      "0000010" when "00110100010111001", -- t[26809] = 2
      "0000010" when "00110100010111010", -- t[26810] = 2
      "0000010" when "00110100010111011", -- t[26811] = 2
      "0000010" when "00110100010111100", -- t[26812] = 2
      "0000010" when "00110100010111101", -- t[26813] = 2
      "0000010" when "00110100010111110", -- t[26814] = 2
      "0000010" when "00110100010111111", -- t[26815] = 2
      "0000010" when "00110100011000000", -- t[26816] = 2
      "0000010" when "00110100011000001", -- t[26817] = 2
      "0000010" when "00110100011000010", -- t[26818] = 2
      "0000010" when "00110100011000011", -- t[26819] = 2
      "0000010" when "00110100011000100", -- t[26820] = 2
      "0000010" when "00110100011000101", -- t[26821] = 2
      "0000010" when "00110100011000110", -- t[26822] = 2
      "0000010" when "00110100011000111", -- t[26823] = 2
      "0000010" when "00110100011001000", -- t[26824] = 2
      "0000010" when "00110100011001001", -- t[26825] = 2
      "0000010" when "00110100011001010", -- t[26826] = 2
      "0000010" when "00110100011001011", -- t[26827] = 2
      "0000010" when "00110100011001100", -- t[26828] = 2
      "0000010" when "00110100011001101", -- t[26829] = 2
      "0000010" when "00110100011001110", -- t[26830] = 2
      "0000010" when "00110100011001111", -- t[26831] = 2
      "0000010" when "00110100011010000", -- t[26832] = 2
      "0000010" when "00110100011010001", -- t[26833] = 2
      "0000010" when "00110100011010010", -- t[26834] = 2
      "0000010" when "00110100011010011", -- t[26835] = 2
      "0000010" when "00110100011010100", -- t[26836] = 2
      "0000010" when "00110100011010101", -- t[26837] = 2
      "0000010" when "00110100011010110", -- t[26838] = 2
      "0000010" when "00110100011010111", -- t[26839] = 2
      "0000010" when "00110100011011000", -- t[26840] = 2
      "0000010" when "00110100011011001", -- t[26841] = 2
      "0000010" when "00110100011011010", -- t[26842] = 2
      "0000010" when "00110100011011011", -- t[26843] = 2
      "0000010" when "00110100011011100", -- t[26844] = 2
      "0000010" when "00110100011011101", -- t[26845] = 2
      "0000010" when "00110100011011110", -- t[26846] = 2
      "0000010" when "00110100011011111", -- t[26847] = 2
      "0000010" when "00110100011100000", -- t[26848] = 2
      "0000010" when "00110100011100001", -- t[26849] = 2
      "0000010" when "00110100011100010", -- t[26850] = 2
      "0000010" when "00110100011100011", -- t[26851] = 2
      "0000010" when "00110100011100100", -- t[26852] = 2
      "0000010" when "00110100011100101", -- t[26853] = 2
      "0000010" when "00110100011100110", -- t[26854] = 2
      "0000010" when "00110100011100111", -- t[26855] = 2
      "0000010" when "00110100011101000", -- t[26856] = 2
      "0000010" when "00110100011101001", -- t[26857] = 2
      "0000010" when "00110100011101010", -- t[26858] = 2
      "0000010" when "00110100011101011", -- t[26859] = 2
      "0000010" when "00110100011101100", -- t[26860] = 2
      "0000010" when "00110100011101101", -- t[26861] = 2
      "0000010" when "00110100011101110", -- t[26862] = 2
      "0000010" when "00110100011101111", -- t[26863] = 2
      "0000010" when "00110100011110000", -- t[26864] = 2
      "0000010" when "00110100011110001", -- t[26865] = 2
      "0000010" when "00110100011110010", -- t[26866] = 2
      "0000010" when "00110100011110011", -- t[26867] = 2
      "0000010" when "00110100011110100", -- t[26868] = 2
      "0000010" when "00110100011110101", -- t[26869] = 2
      "0000010" when "00110100011110110", -- t[26870] = 2
      "0000010" when "00110100011110111", -- t[26871] = 2
      "0000010" when "00110100011111000", -- t[26872] = 2
      "0000010" when "00110100011111001", -- t[26873] = 2
      "0000010" when "00110100011111010", -- t[26874] = 2
      "0000010" when "00110100011111011", -- t[26875] = 2
      "0000010" when "00110100011111100", -- t[26876] = 2
      "0000010" when "00110100011111101", -- t[26877] = 2
      "0000010" when "00110100011111110", -- t[26878] = 2
      "0000010" when "00110100011111111", -- t[26879] = 2
      "0000010" when "00110100100000000", -- t[26880] = 2
      "0000010" when "00110100100000001", -- t[26881] = 2
      "0000010" when "00110100100000010", -- t[26882] = 2
      "0000010" when "00110100100000011", -- t[26883] = 2
      "0000010" when "00110100100000100", -- t[26884] = 2
      "0000010" when "00110100100000101", -- t[26885] = 2
      "0000010" when "00110100100000110", -- t[26886] = 2
      "0000010" when "00110100100000111", -- t[26887] = 2
      "0000010" when "00110100100001000", -- t[26888] = 2
      "0000010" when "00110100100001001", -- t[26889] = 2
      "0000010" when "00110100100001010", -- t[26890] = 2
      "0000010" when "00110100100001011", -- t[26891] = 2
      "0000010" when "00110100100001100", -- t[26892] = 2
      "0000010" when "00110100100001101", -- t[26893] = 2
      "0000010" when "00110100100001110", -- t[26894] = 2
      "0000010" when "00110100100001111", -- t[26895] = 2
      "0000010" when "00110100100010000", -- t[26896] = 2
      "0000010" when "00110100100010001", -- t[26897] = 2
      "0000010" when "00110100100010010", -- t[26898] = 2
      "0000010" when "00110100100010011", -- t[26899] = 2
      "0000010" when "00110100100010100", -- t[26900] = 2
      "0000010" when "00110100100010101", -- t[26901] = 2
      "0000010" when "00110100100010110", -- t[26902] = 2
      "0000010" when "00110100100010111", -- t[26903] = 2
      "0000010" when "00110100100011000", -- t[26904] = 2
      "0000010" when "00110100100011001", -- t[26905] = 2
      "0000010" when "00110100100011010", -- t[26906] = 2
      "0000010" when "00110100100011011", -- t[26907] = 2
      "0000010" when "00110100100011100", -- t[26908] = 2
      "0000010" when "00110100100011101", -- t[26909] = 2
      "0000010" when "00110100100011110", -- t[26910] = 2
      "0000010" when "00110100100011111", -- t[26911] = 2
      "0000010" when "00110100100100000", -- t[26912] = 2
      "0000010" when "00110100100100001", -- t[26913] = 2
      "0000010" when "00110100100100010", -- t[26914] = 2
      "0000010" when "00110100100100011", -- t[26915] = 2
      "0000010" when "00110100100100100", -- t[26916] = 2
      "0000010" when "00110100100100101", -- t[26917] = 2
      "0000010" when "00110100100100110", -- t[26918] = 2
      "0000010" when "00110100100100111", -- t[26919] = 2
      "0000010" when "00110100100101000", -- t[26920] = 2
      "0000010" when "00110100100101001", -- t[26921] = 2
      "0000010" when "00110100100101010", -- t[26922] = 2
      "0000010" when "00110100100101011", -- t[26923] = 2
      "0000010" when "00110100100101100", -- t[26924] = 2
      "0000010" when "00110100100101101", -- t[26925] = 2
      "0000010" when "00110100100101110", -- t[26926] = 2
      "0000010" when "00110100100101111", -- t[26927] = 2
      "0000010" when "00110100100110000", -- t[26928] = 2
      "0000010" when "00110100100110001", -- t[26929] = 2
      "0000010" when "00110100100110010", -- t[26930] = 2
      "0000010" when "00110100100110011", -- t[26931] = 2
      "0000010" when "00110100100110100", -- t[26932] = 2
      "0000010" when "00110100100110101", -- t[26933] = 2
      "0000010" when "00110100100110110", -- t[26934] = 2
      "0000010" when "00110100100110111", -- t[26935] = 2
      "0000010" when "00110100100111000", -- t[26936] = 2
      "0000010" when "00110100100111001", -- t[26937] = 2
      "0000010" when "00110100100111010", -- t[26938] = 2
      "0000010" when "00110100100111011", -- t[26939] = 2
      "0000010" when "00110100100111100", -- t[26940] = 2
      "0000010" when "00110100100111101", -- t[26941] = 2
      "0000010" when "00110100100111110", -- t[26942] = 2
      "0000010" when "00110100100111111", -- t[26943] = 2
      "0000010" when "00110100101000000", -- t[26944] = 2
      "0000010" when "00110100101000001", -- t[26945] = 2
      "0000010" when "00110100101000010", -- t[26946] = 2
      "0000010" when "00110100101000011", -- t[26947] = 2
      "0000010" when "00110100101000100", -- t[26948] = 2
      "0000010" when "00110100101000101", -- t[26949] = 2
      "0000010" when "00110100101000110", -- t[26950] = 2
      "0000010" when "00110100101000111", -- t[26951] = 2
      "0000010" when "00110100101001000", -- t[26952] = 2
      "0000010" when "00110100101001001", -- t[26953] = 2
      "0000010" when "00110100101001010", -- t[26954] = 2
      "0000010" when "00110100101001011", -- t[26955] = 2
      "0000010" when "00110100101001100", -- t[26956] = 2
      "0000010" when "00110100101001101", -- t[26957] = 2
      "0000010" when "00110100101001110", -- t[26958] = 2
      "0000010" when "00110100101001111", -- t[26959] = 2
      "0000010" when "00110100101010000", -- t[26960] = 2
      "0000010" when "00110100101010001", -- t[26961] = 2
      "0000010" when "00110100101010010", -- t[26962] = 2
      "0000010" when "00110100101010011", -- t[26963] = 2
      "0000010" when "00110100101010100", -- t[26964] = 2
      "0000010" when "00110100101010101", -- t[26965] = 2
      "0000010" when "00110100101010110", -- t[26966] = 2
      "0000010" when "00110100101010111", -- t[26967] = 2
      "0000010" when "00110100101011000", -- t[26968] = 2
      "0000010" when "00110100101011001", -- t[26969] = 2
      "0000010" when "00110100101011010", -- t[26970] = 2
      "0000010" when "00110100101011011", -- t[26971] = 2
      "0000010" when "00110100101011100", -- t[26972] = 2
      "0000010" when "00110100101011101", -- t[26973] = 2
      "0000010" when "00110100101011110", -- t[26974] = 2
      "0000010" when "00110100101011111", -- t[26975] = 2
      "0000010" when "00110100101100000", -- t[26976] = 2
      "0000010" when "00110100101100001", -- t[26977] = 2
      "0000010" when "00110100101100010", -- t[26978] = 2
      "0000010" when "00110100101100011", -- t[26979] = 2
      "0000010" when "00110100101100100", -- t[26980] = 2
      "0000010" when "00110100101100101", -- t[26981] = 2
      "0000010" when "00110100101100110", -- t[26982] = 2
      "0000010" when "00110100101100111", -- t[26983] = 2
      "0000010" when "00110100101101000", -- t[26984] = 2
      "0000010" when "00110100101101001", -- t[26985] = 2
      "0000010" when "00110100101101010", -- t[26986] = 2
      "0000010" when "00110100101101011", -- t[26987] = 2
      "0000010" when "00110100101101100", -- t[26988] = 2
      "0000010" when "00110100101101101", -- t[26989] = 2
      "0000010" when "00110100101101110", -- t[26990] = 2
      "0000010" when "00110100101101111", -- t[26991] = 2
      "0000010" when "00110100101110000", -- t[26992] = 2
      "0000010" when "00110100101110001", -- t[26993] = 2
      "0000010" when "00110100101110010", -- t[26994] = 2
      "0000010" when "00110100101110011", -- t[26995] = 2
      "0000010" when "00110100101110100", -- t[26996] = 2
      "0000010" when "00110100101110101", -- t[26997] = 2
      "0000010" when "00110100101110110", -- t[26998] = 2
      "0000010" when "00110100101110111", -- t[26999] = 2
      "0000010" when "00110100101111000", -- t[27000] = 2
      "0000010" when "00110100101111001", -- t[27001] = 2
      "0000010" when "00110100101111010", -- t[27002] = 2
      "0000010" when "00110100101111011", -- t[27003] = 2
      "0000010" when "00110100101111100", -- t[27004] = 2
      "0000010" when "00110100101111101", -- t[27005] = 2
      "0000010" when "00110100101111110", -- t[27006] = 2
      "0000010" when "00110100101111111", -- t[27007] = 2
      "0000010" when "00110100110000000", -- t[27008] = 2
      "0000010" when "00110100110000001", -- t[27009] = 2
      "0000010" when "00110100110000010", -- t[27010] = 2
      "0000010" when "00110100110000011", -- t[27011] = 2
      "0000010" when "00110100110000100", -- t[27012] = 2
      "0000010" when "00110100110000101", -- t[27013] = 2
      "0000010" when "00110100110000110", -- t[27014] = 2
      "0000010" when "00110100110000111", -- t[27015] = 2
      "0000010" when "00110100110001000", -- t[27016] = 2
      "0000010" when "00110100110001001", -- t[27017] = 2
      "0000010" when "00110100110001010", -- t[27018] = 2
      "0000010" when "00110100110001011", -- t[27019] = 2
      "0000010" when "00110100110001100", -- t[27020] = 2
      "0000010" when "00110100110001101", -- t[27021] = 2
      "0000010" when "00110100110001110", -- t[27022] = 2
      "0000010" when "00110100110001111", -- t[27023] = 2
      "0000010" when "00110100110010000", -- t[27024] = 2
      "0000010" when "00110100110010001", -- t[27025] = 2
      "0000010" when "00110100110010010", -- t[27026] = 2
      "0000010" when "00110100110010011", -- t[27027] = 2
      "0000010" when "00110100110010100", -- t[27028] = 2
      "0000010" when "00110100110010101", -- t[27029] = 2
      "0000010" when "00110100110010110", -- t[27030] = 2
      "0000010" when "00110100110010111", -- t[27031] = 2
      "0000010" when "00110100110011000", -- t[27032] = 2
      "0000010" when "00110100110011001", -- t[27033] = 2
      "0000010" when "00110100110011010", -- t[27034] = 2
      "0000010" when "00110100110011011", -- t[27035] = 2
      "0000010" when "00110100110011100", -- t[27036] = 2
      "0000010" when "00110100110011101", -- t[27037] = 2
      "0000010" when "00110100110011110", -- t[27038] = 2
      "0000010" when "00110100110011111", -- t[27039] = 2
      "0000010" when "00110100110100000", -- t[27040] = 2
      "0000010" when "00110100110100001", -- t[27041] = 2
      "0000010" when "00110100110100010", -- t[27042] = 2
      "0000010" when "00110100110100011", -- t[27043] = 2
      "0000010" when "00110100110100100", -- t[27044] = 2
      "0000010" when "00110100110100101", -- t[27045] = 2
      "0000010" when "00110100110100110", -- t[27046] = 2
      "0000010" when "00110100110100111", -- t[27047] = 2
      "0000010" when "00110100110101000", -- t[27048] = 2
      "0000010" when "00110100110101001", -- t[27049] = 2
      "0000010" when "00110100110101010", -- t[27050] = 2
      "0000010" when "00110100110101011", -- t[27051] = 2
      "0000010" when "00110100110101100", -- t[27052] = 2
      "0000010" when "00110100110101101", -- t[27053] = 2
      "0000010" when "00110100110101110", -- t[27054] = 2
      "0000010" when "00110100110101111", -- t[27055] = 2
      "0000010" when "00110100110110000", -- t[27056] = 2
      "0000010" when "00110100110110001", -- t[27057] = 2
      "0000010" when "00110100110110010", -- t[27058] = 2
      "0000010" when "00110100110110011", -- t[27059] = 2
      "0000010" when "00110100110110100", -- t[27060] = 2
      "0000010" when "00110100110110101", -- t[27061] = 2
      "0000010" when "00110100110110110", -- t[27062] = 2
      "0000010" when "00110100110110111", -- t[27063] = 2
      "0000010" when "00110100110111000", -- t[27064] = 2
      "0000010" when "00110100110111001", -- t[27065] = 2
      "0000010" when "00110100110111010", -- t[27066] = 2
      "0000010" when "00110100110111011", -- t[27067] = 2
      "0000010" when "00110100110111100", -- t[27068] = 2
      "0000010" when "00110100110111101", -- t[27069] = 2
      "0000010" when "00110100110111110", -- t[27070] = 2
      "0000010" when "00110100110111111", -- t[27071] = 2
      "0000010" when "00110100111000000", -- t[27072] = 2
      "0000010" when "00110100111000001", -- t[27073] = 2
      "0000010" when "00110100111000010", -- t[27074] = 2
      "0000010" when "00110100111000011", -- t[27075] = 2
      "0000010" when "00110100111000100", -- t[27076] = 2
      "0000010" when "00110100111000101", -- t[27077] = 2
      "0000010" when "00110100111000110", -- t[27078] = 2
      "0000010" when "00110100111000111", -- t[27079] = 2
      "0000010" when "00110100111001000", -- t[27080] = 2
      "0000010" when "00110100111001001", -- t[27081] = 2
      "0000010" when "00110100111001010", -- t[27082] = 2
      "0000010" when "00110100111001011", -- t[27083] = 2
      "0000010" when "00110100111001100", -- t[27084] = 2
      "0000010" when "00110100111001101", -- t[27085] = 2
      "0000010" when "00110100111001110", -- t[27086] = 2
      "0000010" when "00110100111001111", -- t[27087] = 2
      "0000010" when "00110100111010000", -- t[27088] = 2
      "0000010" when "00110100111010001", -- t[27089] = 2
      "0000010" when "00110100111010010", -- t[27090] = 2
      "0000010" when "00110100111010011", -- t[27091] = 2
      "0000010" when "00110100111010100", -- t[27092] = 2
      "0000010" when "00110100111010101", -- t[27093] = 2
      "0000010" when "00110100111010110", -- t[27094] = 2
      "0000010" when "00110100111010111", -- t[27095] = 2
      "0000010" when "00110100111011000", -- t[27096] = 2
      "0000010" when "00110100111011001", -- t[27097] = 2
      "0000010" when "00110100111011010", -- t[27098] = 2
      "0000010" when "00110100111011011", -- t[27099] = 2
      "0000010" when "00110100111011100", -- t[27100] = 2
      "0000010" when "00110100111011101", -- t[27101] = 2
      "0000010" when "00110100111011110", -- t[27102] = 2
      "0000010" when "00110100111011111", -- t[27103] = 2
      "0000010" when "00110100111100000", -- t[27104] = 2
      "0000010" when "00110100111100001", -- t[27105] = 2
      "0000010" when "00110100111100010", -- t[27106] = 2
      "0000010" when "00110100111100011", -- t[27107] = 2
      "0000010" when "00110100111100100", -- t[27108] = 2
      "0000010" when "00110100111100101", -- t[27109] = 2
      "0000010" when "00110100111100110", -- t[27110] = 2
      "0000010" when "00110100111100111", -- t[27111] = 2
      "0000010" when "00110100111101000", -- t[27112] = 2
      "0000010" when "00110100111101001", -- t[27113] = 2
      "0000010" when "00110100111101010", -- t[27114] = 2
      "0000010" when "00110100111101011", -- t[27115] = 2
      "0000010" when "00110100111101100", -- t[27116] = 2
      "0000010" when "00110100111101101", -- t[27117] = 2
      "0000010" when "00110100111101110", -- t[27118] = 2
      "0000010" when "00110100111101111", -- t[27119] = 2
      "0000010" when "00110100111110000", -- t[27120] = 2
      "0000010" when "00110100111110001", -- t[27121] = 2
      "0000010" when "00110100111110010", -- t[27122] = 2
      "0000010" when "00110100111110011", -- t[27123] = 2
      "0000010" when "00110100111110100", -- t[27124] = 2
      "0000010" when "00110100111110101", -- t[27125] = 2
      "0000010" when "00110100111110110", -- t[27126] = 2
      "0000010" when "00110100111110111", -- t[27127] = 2
      "0000010" when "00110100111111000", -- t[27128] = 2
      "0000010" when "00110100111111001", -- t[27129] = 2
      "0000010" when "00110100111111010", -- t[27130] = 2
      "0000010" when "00110100111111011", -- t[27131] = 2
      "0000010" when "00110100111111100", -- t[27132] = 2
      "0000010" when "00110100111111101", -- t[27133] = 2
      "0000010" when "00110100111111110", -- t[27134] = 2
      "0000010" when "00110100111111111", -- t[27135] = 2
      "0000010" when "00110101000000000", -- t[27136] = 2
      "0000010" when "00110101000000001", -- t[27137] = 2
      "0000010" when "00110101000000010", -- t[27138] = 2
      "0000010" when "00110101000000011", -- t[27139] = 2
      "0000010" when "00110101000000100", -- t[27140] = 2
      "0000010" when "00110101000000101", -- t[27141] = 2
      "0000010" when "00110101000000110", -- t[27142] = 2
      "0000010" when "00110101000000111", -- t[27143] = 2
      "0000010" when "00110101000001000", -- t[27144] = 2
      "0000010" when "00110101000001001", -- t[27145] = 2
      "0000010" when "00110101000001010", -- t[27146] = 2
      "0000010" when "00110101000001011", -- t[27147] = 2
      "0000010" when "00110101000001100", -- t[27148] = 2
      "0000010" when "00110101000001101", -- t[27149] = 2
      "0000010" when "00110101000001110", -- t[27150] = 2
      "0000010" when "00110101000001111", -- t[27151] = 2
      "0000010" when "00110101000010000", -- t[27152] = 2
      "0000010" when "00110101000010001", -- t[27153] = 2
      "0000010" when "00110101000010010", -- t[27154] = 2
      "0000010" when "00110101000010011", -- t[27155] = 2
      "0000010" when "00110101000010100", -- t[27156] = 2
      "0000010" when "00110101000010101", -- t[27157] = 2
      "0000010" when "00110101000010110", -- t[27158] = 2
      "0000010" when "00110101000010111", -- t[27159] = 2
      "0000010" when "00110101000011000", -- t[27160] = 2
      "0000010" when "00110101000011001", -- t[27161] = 2
      "0000010" when "00110101000011010", -- t[27162] = 2
      "0000010" when "00110101000011011", -- t[27163] = 2
      "0000010" when "00110101000011100", -- t[27164] = 2
      "0000010" when "00110101000011101", -- t[27165] = 2
      "0000010" when "00110101000011110", -- t[27166] = 2
      "0000010" when "00110101000011111", -- t[27167] = 2
      "0000010" when "00110101000100000", -- t[27168] = 2
      "0000010" when "00110101000100001", -- t[27169] = 2
      "0000010" when "00110101000100010", -- t[27170] = 2
      "0000010" when "00110101000100011", -- t[27171] = 2
      "0000010" when "00110101000100100", -- t[27172] = 2
      "0000010" when "00110101000100101", -- t[27173] = 2
      "0000010" when "00110101000100110", -- t[27174] = 2
      "0000010" when "00110101000100111", -- t[27175] = 2
      "0000010" when "00110101000101000", -- t[27176] = 2
      "0000010" when "00110101000101001", -- t[27177] = 2
      "0000010" when "00110101000101010", -- t[27178] = 2
      "0000010" when "00110101000101011", -- t[27179] = 2
      "0000010" when "00110101000101100", -- t[27180] = 2
      "0000010" when "00110101000101101", -- t[27181] = 2
      "0000010" when "00110101000101110", -- t[27182] = 2
      "0000010" when "00110101000101111", -- t[27183] = 2
      "0000010" when "00110101000110000", -- t[27184] = 2
      "0000010" when "00110101000110001", -- t[27185] = 2
      "0000010" when "00110101000110010", -- t[27186] = 2
      "0000010" when "00110101000110011", -- t[27187] = 2
      "0000010" when "00110101000110100", -- t[27188] = 2
      "0000010" when "00110101000110101", -- t[27189] = 2
      "0000010" when "00110101000110110", -- t[27190] = 2
      "0000010" when "00110101000110111", -- t[27191] = 2
      "0000010" when "00110101000111000", -- t[27192] = 2
      "0000010" when "00110101000111001", -- t[27193] = 2
      "0000010" when "00110101000111010", -- t[27194] = 2
      "0000010" when "00110101000111011", -- t[27195] = 2
      "0000010" when "00110101000111100", -- t[27196] = 2
      "0000010" when "00110101000111101", -- t[27197] = 2
      "0000010" when "00110101000111110", -- t[27198] = 2
      "0000010" when "00110101000111111", -- t[27199] = 2
      "0000010" when "00110101001000000", -- t[27200] = 2
      "0000010" when "00110101001000001", -- t[27201] = 2
      "0000010" when "00110101001000010", -- t[27202] = 2
      "0000010" when "00110101001000011", -- t[27203] = 2
      "0000010" when "00110101001000100", -- t[27204] = 2
      "0000010" when "00110101001000101", -- t[27205] = 2
      "0000010" when "00110101001000110", -- t[27206] = 2
      "0000010" when "00110101001000111", -- t[27207] = 2
      "0000010" when "00110101001001000", -- t[27208] = 2
      "0000010" when "00110101001001001", -- t[27209] = 2
      "0000010" when "00110101001001010", -- t[27210] = 2
      "0000010" when "00110101001001011", -- t[27211] = 2
      "0000010" when "00110101001001100", -- t[27212] = 2
      "0000010" when "00110101001001101", -- t[27213] = 2
      "0000010" when "00110101001001110", -- t[27214] = 2
      "0000010" when "00110101001001111", -- t[27215] = 2
      "0000010" when "00110101001010000", -- t[27216] = 2
      "0000010" when "00110101001010001", -- t[27217] = 2
      "0000010" when "00110101001010010", -- t[27218] = 2
      "0000010" when "00110101001010011", -- t[27219] = 2
      "0000010" when "00110101001010100", -- t[27220] = 2
      "0000010" when "00110101001010101", -- t[27221] = 2
      "0000010" when "00110101001010110", -- t[27222] = 2
      "0000010" when "00110101001010111", -- t[27223] = 2
      "0000010" when "00110101001011000", -- t[27224] = 2
      "0000010" when "00110101001011001", -- t[27225] = 2
      "0000010" when "00110101001011010", -- t[27226] = 2
      "0000010" when "00110101001011011", -- t[27227] = 2
      "0000010" when "00110101001011100", -- t[27228] = 2
      "0000010" when "00110101001011101", -- t[27229] = 2
      "0000010" when "00110101001011110", -- t[27230] = 2
      "0000010" when "00110101001011111", -- t[27231] = 2
      "0000010" when "00110101001100000", -- t[27232] = 2
      "0000010" when "00110101001100001", -- t[27233] = 2
      "0000010" when "00110101001100010", -- t[27234] = 2
      "0000010" when "00110101001100011", -- t[27235] = 2
      "0000010" when "00110101001100100", -- t[27236] = 2
      "0000010" when "00110101001100101", -- t[27237] = 2
      "0000010" when "00110101001100110", -- t[27238] = 2
      "0000010" when "00110101001100111", -- t[27239] = 2
      "0000010" when "00110101001101000", -- t[27240] = 2
      "0000010" when "00110101001101001", -- t[27241] = 2
      "0000010" when "00110101001101010", -- t[27242] = 2
      "0000010" when "00110101001101011", -- t[27243] = 2
      "0000010" when "00110101001101100", -- t[27244] = 2
      "0000010" when "00110101001101101", -- t[27245] = 2
      "0000010" when "00110101001101110", -- t[27246] = 2
      "0000010" when "00110101001101111", -- t[27247] = 2
      "0000010" when "00110101001110000", -- t[27248] = 2
      "0000010" when "00110101001110001", -- t[27249] = 2
      "0000010" when "00110101001110010", -- t[27250] = 2
      "0000010" when "00110101001110011", -- t[27251] = 2
      "0000010" when "00110101001110100", -- t[27252] = 2
      "0000010" when "00110101001110101", -- t[27253] = 2
      "0000010" when "00110101001110110", -- t[27254] = 2
      "0000010" when "00110101001110111", -- t[27255] = 2
      "0000010" when "00110101001111000", -- t[27256] = 2
      "0000010" when "00110101001111001", -- t[27257] = 2
      "0000010" when "00110101001111010", -- t[27258] = 2
      "0000010" when "00110101001111011", -- t[27259] = 2
      "0000010" when "00110101001111100", -- t[27260] = 2
      "0000010" when "00110101001111101", -- t[27261] = 2
      "0000010" when "00110101001111110", -- t[27262] = 2
      "0000010" when "00110101001111111", -- t[27263] = 2
      "0000010" when "00110101010000000", -- t[27264] = 2
      "0000010" when "00110101010000001", -- t[27265] = 2
      "0000010" when "00110101010000010", -- t[27266] = 2
      "0000010" when "00110101010000011", -- t[27267] = 2
      "0000010" when "00110101010000100", -- t[27268] = 2
      "0000010" when "00110101010000101", -- t[27269] = 2
      "0000010" when "00110101010000110", -- t[27270] = 2
      "0000010" when "00110101010000111", -- t[27271] = 2
      "0000010" when "00110101010001000", -- t[27272] = 2
      "0000010" when "00110101010001001", -- t[27273] = 2
      "0000010" when "00110101010001010", -- t[27274] = 2
      "0000010" when "00110101010001011", -- t[27275] = 2
      "0000010" when "00110101010001100", -- t[27276] = 2
      "0000010" when "00110101010001101", -- t[27277] = 2
      "0000010" when "00110101010001110", -- t[27278] = 2
      "0000010" when "00110101010001111", -- t[27279] = 2
      "0000010" when "00110101010010000", -- t[27280] = 2
      "0000010" when "00110101010010001", -- t[27281] = 2
      "0000010" when "00110101010010010", -- t[27282] = 2
      "0000010" when "00110101010010011", -- t[27283] = 2
      "0000010" when "00110101010010100", -- t[27284] = 2
      "0000010" when "00110101010010101", -- t[27285] = 2
      "0000010" when "00110101010010110", -- t[27286] = 2
      "0000010" when "00110101010010111", -- t[27287] = 2
      "0000010" when "00110101010011000", -- t[27288] = 2
      "0000010" when "00110101010011001", -- t[27289] = 2
      "0000010" when "00110101010011010", -- t[27290] = 2
      "0000010" when "00110101010011011", -- t[27291] = 2
      "0000010" when "00110101010011100", -- t[27292] = 2
      "0000010" when "00110101010011101", -- t[27293] = 2
      "0000010" when "00110101010011110", -- t[27294] = 2
      "0000010" when "00110101010011111", -- t[27295] = 2
      "0000010" when "00110101010100000", -- t[27296] = 2
      "0000010" when "00110101010100001", -- t[27297] = 2
      "0000010" when "00110101010100010", -- t[27298] = 2
      "0000010" when "00110101010100011", -- t[27299] = 2
      "0000010" when "00110101010100100", -- t[27300] = 2
      "0000010" when "00110101010100101", -- t[27301] = 2
      "0000010" when "00110101010100110", -- t[27302] = 2
      "0000010" when "00110101010100111", -- t[27303] = 2
      "0000010" when "00110101010101000", -- t[27304] = 2
      "0000010" when "00110101010101001", -- t[27305] = 2
      "0000010" when "00110101010101010", -- t[27306] = 2
      "0000010" when "00110101010101011", -- t[27307] = 2
      "0000010" when "00110101010101100", -- t[27308] = 2
      "0000010" when "00110101010101101", -- t[27309] = 2
      "0000010" when "00110101010101110", -- t[27310] = 2
      "0000010" when "00110101010101111", -- t[27311] = 2
      "0000010" when "00110101010110000", -- t[27312] = 2
      "0000010" when "00110101010110001", -- t[27313] = 2
      "0000010" when "00110101010110010", -- t[27314] = 2
      "0000010" when "00110101010110011", -- t[27315] = 2
      "0000010" when "00110101010110100", -- t[27316] = 2
      "0000010" when "00110101010110101", -- t[27317] = 2
      "0000010" when "00110101010110110", -- t[27318] = 2
      "0000010" when "00110101010110111", -- t[27319] = 2
      "0000010" when "00110101010111000", -- t[27320] = 2
      "0000010" when "00110101010111001", -- t[27321] = 2
      "0000010" when "00110101010111010", -- t[27322] = 2
      "0000010" when "00110101010111011", -- t[27323] = 2
      "0000010" when "00110101010111100", -- t[27324] = 2
      "0000010" when "00110101010111101", -- t[27325] = 2
      "0000010" when "00110101010111110", -- t[27326] = 2
      "0000010" when "00110101010111111", -- t[27327] = 2
      "0000010" when "00110101011000000", -- t[27328] = 2
      "0000010" when "00110101011000001", -- t[27329] = 2
      "0000010" when "00110101011000010", -- t[27330] = 2
      "0000010" when "00110101011000011", -- t[27331] = 2
      "0000010" when "00110101011000100", -- t[27332] = 2
      "0000010" when "00110101011000101", -- t[27333] = 2
      "0000010" when "00110101011000110", -- t[27334] = 2
      "0000010" when "00110101011000111", -- t[27335] = 2
      "0000010" when "00110101011001000", -- t[27336] = 2
      "0000010" when "00110101011001001", -- t[27337] = 2
      "0000010" when "00110101011001010", -- t[27338] = 2
      "0000010" when "00110101011001011", -- t[27339] = 2
      "0000010" when "00110101011001100", -- t[27340] = 2
      "0000010" when "00110101011001101", -- t[27341] = 2
      "0000010" when "00110101011001110", -- t[27342] = 2
      "0000010" when "00110101011001111", -- t[27343] = 2
      "0000010" when "00110101011010000", -- t[27344] = 2
      "0000010" when "00110101011010001", -- t[27345] = 2
      "0000010" when "00110101011010010", -- t[27346] = 2
      "0000010" when "00110101011010011", -- t[27347] = 2
      "0000010" when "00110101011010100", -- t[27348] = 2
      "0000010" when "00110101011010101", -- t[27349] = 2
      "0000010" when "00110101011010110", -- t[27350] = 2
      "0000010" when "00110101011010111", -- t[27351] = 2
      "0000010" when "00110101011011000", -- t[27352] = 2
      "0000010" when "00110101011011001", -- t[27353] = 2
      "0000010" when "00110101011011010", -- t[27354] = 2
      "0000010" when "00110101011011011", -- t[27355] = 2
      "0000010" when "00110101011011100", -- t[27356] = 2
      "0000010" when "00110101011011101", -- t[27357] = 2
      "0000010" when "00110101011011110", -- t[27358] = 2
      "0000010" when "00110101011011111", -- t[27359] = 2
      "0000010" when "00110101011100000", -- t[27360] = 2
      "0000010" when "00110101011100001", -- t[27361] = 2
      "0000010" when "00110101011100010", -- t[27362] = 2
      "0000010" when "00110101011100011", -- t[27363] = 2
      "0000010" when "00110101011100100", -- t[27364] = 2
      "0000010" when "00110101011100101", -- t[27365] = 2
      "0000010" when "00110101011100110", -- t[27366] = 2
      "0000010" when "00110101011100111", -- t[27367] = 2
      "0000010" when "00110101011101000", -- t[27368] = 2
      "0000010" when "00110101011101001", -- t[27369] = 2
      "0000010" when "00110101011101010", -- t[27370] = 2
      "0000010" when "00110101011101011", -- t[27371] = 2
      "0000010" when "00110101011101100", -- t[27372] = 2
      "0000010" when "00110101011101101", -- t[27373] = 2
      "0000010" when "00110101011101110", -- t[27374] = 2
      "0000010" when "00110101011101111", -- t[27375] = 2
      "0000010" when "00110101011110000", -- t[27376] = 2
      "0000010" when "00110101011110001", -- t[27377] = 2
      "0000010" when "00110101011110010", -- t[27378] = 2
      "0000010" when "00110101011110011", -- t[27379] = 2
      "0000010" when "00110101011110100", -- t[27380] = 2
      "0000010" when "00110101011110101", -- t[27381] = 2
      "0000010" when "00110101011110110", -- t[27382] = 2
      "0000010" when "00110101011110111", -- t[27383] = 2
      "0000010" when "00110101011111000", -- t[27384] = 2
      "0000010" when "00110101011111001", -- t[27385] = 2
      "0000010" when "00110101011111010", -- t[27386] = 2
      "0000010" when "00110101011111011", -- t[27387] = 2
      "0000010" when "00110101011111100", -- t[27388] = 2
      "0000010" when "00110101011111101", -- t[27389] = 2
      "0000010" when "00110101011111110", -- t[27390] = 2
      "0000010" when "00110101011111111", -- t[27391] = 2
      "0000010" when "00110101100000000", -- t[27392] = 2
      "0000010" when "00110101100000001", -- t[27393] = 2
      "0000010" when "00110101100000010", -- t[27394] = 2
      "0000010" when "00110101100000011", -- t[27395] = 2
      "0000010" when "00110101100000100", -- t[27396] = 2
      "0000010" when "00110101100000101", -- t[27397] = 2
      "0000010" when "00110101100000110", -- t[27398] = 2
      "0000010" when "00110101100000111", -- t[27399] = 2
      "0000010" when "00110101100001000", -- t[27400] = 2
      "0000010" when "00110101100001001", -- t[27401] = 2
      "0000010" when "00110101100001010", -- t[27402] = 2
      "0000010" when "00110101100001011", -- t[27403] = 2
      "0000010" when "00110101100001100", -- t[27404] = 2
      "0000010" when "00110101100001101", -- t[27405] = 2
      "0000010" when "00110101100001110", -- t[27406] = 2
      "0000010" when "00110101100001111", -- t[27407] = 2
      "0000010" when "00110101100010000", -- t[27408] = 2
      "0000010" when "00110101100010001", -- t[27409] = 2
      "0000010" when "00110101100010010", -- t[27410] = 2
      "0000010" when "00110101100010011", -- t[27411] = 2
      "0000010" when "00110101100010100", -- t[27412] = 2
      "0000010" when "00110101100010101", -- t[27413] = 2
      "0000010" when "00110101100010110", -- t[27414] = 2
      "0000010" when "00110101100010111", -- t[27415] = 2
      "0000010" when "00110101100011000", -- t[27416] = 2
      "0000010" when "00110101100011001", -- t[27417] = 2
      "0000010" when "00110101100011010", -- t[27418] = 2
      "0000010" when "00110101100011011", -- t[27419] = 2
      "0000010" when "00110101100011100", -- t[27420] = 2
      "0000010" when "00110101100011101", -- t[27421] = 2
      "0000010" when "00110101100011110", -- t[27422] = 2
      "0000010" when "00110101100011111", -- t[27423] = 2
      "0000010" when "00110101100100000", -- t[27424] = 2
      "0000010" when "00110101100100001", -- t[27425] = 2
      "0000010" when "00110101100100010", -- t[27426] = 2
      "0000010" when "00110101100100011", -- t[27427] = 2
      "0000010" when "00110101100100100", -- t[27428] = 2
      "0000010" when "00110101100100101", -- t[27429] = 2
      "0000010" when "00110101100100110", -- t[27430] = 2
      "0000010" when "00110101100100111", -- t[27431] = 2
      "0000010" when "00110101100101000", -- t[27432] = 2
      "0000010" when "00110101100101001", -- t[27433] = 2
      "0000010" when "00110101100101010", -- t[27434] = 2
      "0000010" when "00110101100101011", -- t[27435] = 2
      "0000010" when "00110101100101100", -- t[27436] = 2
      "0000010" when "00110101100101101", -- t[27437] = 2
      "0000010" when "00110101100101110", -- t[27438] = 2
      "0000010" when "00110101100101111", -- t[27439] = 2
      "0000010" when "00110101100110000", -- t[27440] = 2
      "0000010" when "00110101100110001", -- t[27441] = 2
      "0000010" when "00110101100110010", -- t[27442] = 2
      "0000010" when "00110101100110011", -- t[27443] = 2
      "0000010" when "00110101100110100", -- t[27444] = 2
      "0000010" when "00110101100110101", -- t[27445] = 2
      "0000010" when "00110101100110110", -- t[27446] = 2
      "0000010" when "00110101100110111", -- t[27447] = 2
      "0000010" when "00110101100111000", -- t[27448] = 2
      "0000010" when "00110101100111001", -- t[27449] = 2
      "0000010" when "00110101100111010", -- t[27450] = 2
      "0000010" when "00110101100111011", -- t[27451] = 2
      "0000010" when "00110101100111100", -- t[27452] = 2
      "0000010" when "00110101100111101", -- t[27453] = 2
      "0000010" when "00110101100111110", -- t[27454] = 2
      "0000010" when "00110101100111111", -- t[27455] = 2
      "0000010" when "00110101101000000", -- t[27456] = 2
      "0000010" when "00110101101000001", -- t[27457] = 2
      "0000010" when "00110101101000010", -- t[27458] = 2
      "0000010" when "00110101101000011", -- t[27459] = 2
      "0000010" when "00110101101000100", -- t[27460] = 2
      "0000010" when "00110101101000101", -- t[27461] = 2
      "0000010" when "00110101101000110", -- t[27462] = 2
      "0000010" when "00110101101000111", -- t[27463] = 2
      "0000010" when "00110101101001000", -- t[27464] = 2
      "0000010" when "00110101101001001", -- t[27465] = 2
      "0000010" when "00110101101001010", -- t[27466] = 2
      "0000010" when "00110101101001011", -- t[27467] = 2
      "0000010" when "00110101101001100", -- t[27468] = 2
      "0000010" when "00110101101001101", -- t[27469] = 2
      "0000010" when "00110101101001110", -- t[27470] = 2
      "0000010" when "00110101101001111", -- t[27471] = 2
      "0000010" when "00110101101010000", -- t[27472] = 2
      "0000010" when "00110101101010001", -- t[27473] = 2
      "0000010" when "00110101101010010", -- t[27474] = 2
      "0000010" when "00110101101010011", -- t[27475] = 2
      "0000010" when "00110101101010100", -- t[27476] = 2
      "0000010" when "00110101101010101", -- t[27477] = 2
      "0000010" when "00110101101010110", -- t[27478] = 2
      "0000010" when "00110101101010111", -- t[27479] = 2
      "0000010" when "00110101101011000", -- t[27480] = 2
      "0000010" when "00110101101011001", -- t[27481] = 2
      "0000010" when "00110101101011010", -- t[27482] = 2
      "0000010" when "00110101101011011", -- t[27483] = 2
      "0000010" when "00110101101011100", -- t[27484] = 2
      "0000010" when "00110101101011101", -- t[27485] = 2
      "0000010" when "00110101101011110", -- t[27486] = 2
      "0000010" when "00110101101011111", -- t[27487] = 2
      "0000010" when "00110101101100000", -- t[27488] = 2
      "0000010" when "00110101101100001", -- t[27489] = 2
      "0000010" when "00110101101100010", -- t[27490] = 2
      "0000010" when "00110101101100011", -- t[27491] = 2
      "0000010" when "00110101101100100", -- t[27492] = 2
      "0000010" when "00110101101100101", -- t[27493] = 2
      "0000010" when "00110101101100110", -- t[27494] = 2
      "0000010" when "00110101101100111", -- t[27495] = 2
      "0000010" when "00110101101101000", -- t[27496] = 2
      "0000010" when "00110101101101001", -- t[27497] = 2
      "0000010" when "00110101101101010", -- t[27498] = 2
      "0000010" when "00110101101101011", -- t[27499] = 2
      "0000010" when "00110101101101100", -- t[27500] = 2
      "0000010" when "00110101101101101", -- t[27501] = 2
      "0000010" when "00110101101101110", -- t[27502] = 2
      "0000010" when "00110101101101111", -- t[27503] = 2
      "0000010" when "00110101101110000", -- t[27504] = 2
      "0000010" when "00110101101110001", -- t[27505] = 2
      "0000010" when "00110101101110010", -- t[27506] = 2
      "0000010" when "00110101101110011", -- t[27507] = 2
      "0000010" when "00110101101110100", -- t[27508] = 2
      "0000010" when "00110101101110101", -- t[27509] = 2
      "0000010" when "00110101101110110", -- t[27510] = 2
      "0000010" when "00110101101110111", -- t[27511] = 2
      "0000010" when "00110101101111000", -- t[27512] = 2
      "0000010" when "00110101101111001", -- t[27513] = 2
      "0000010" when "00110101101111010", -- t[27514] = 2
      "0000010" when "00110101101111011", -- t[27515] = 2
      "0000010" when "00110101101111100", -- t[27516] = 2
      "0000010" when "00110101101111101", -- t[27517] = 2
      "0000010" when "00110101101111110", -- t[27518] = 2
      "0000010" when "00110101101111111", -- t[27519] = 2
      "0000010" when "00110101110000000", -- t[27520] = 2
      "0000010" when "00110101110000001", -- t[27521] = 2
      "0000010" when "00110101110000010", -- t[27522] = 2
      "0000010" when "00110101110000011", -- t[27523] = 2
      "0000010" when "00110101110000100", -- t[27524] = 2
      "0000010" when "00110101110000101", -- t[27525] = 2
      "0000010" when "00110101110000110", -- t[27526] = 2
      "0000010" when "00110101110000111", -- t[27527] = 2
      "0000010" when "00110101110001000", -- t[27528] = 2
      "0000010" when "00110101110001001", -- t[27529] = 2
      "0000010" when "00110101110001010", -- t[27530] = 2
      "0000010" when "00110101110001011", -- t[27531] = 2
      "0000010" when "00110101110001100", -- t[27532] = 2
      "0000010" when "00110101110001101", -- t[27533] = 2
      "0000010" when "00110101110001110", -- t[27534] = 2
      "0000010" when "00110101110001111", -- t[27535] = 2
      "0000010" when "00110101110010000", -- t[27536] = 2
      "0000010" when "00110101110010001", -- t[27537] = 2
      "0000010" when "00110101110010010", -- t[27538] = 2
      "0000010" when "00110101110010011", -- t[27539] = 2
      "0000010" when "00110101110010100", -- t[27540] = 2
      "0000010" when "00110101110010101", -- t[27541] = 2
      "0000010" when "00110101110010110", -- t[27542] = 2
      "0000010" when "00110101110010111", -- t[27543] = 2
      "0000010" when "00110101110011000", -- t[27544] = 2
      "0000010" when "00110101110011001", -- t[27545] = 2
      "0000010" when "00110101110011010", -- t[27546] = 2
      "0000010" when "00110101110011011", -- t[27547] = 2
      "0000010" when "00110101110011100", -- t[27548] = 2
      "0000010" when "00110101110011101", -- t[27549] = 2
      "0000010" when "00110101110011110", -- t[27550] = 2
      "0000010" when "00110101110011111", -- t[27551] = 2
      "0000010" when "00110101110100000", -- t[27552] = 2
      "0000010" when "00110101110100001", -- t[27553] = 2
      "0000010" when "00110101110100010", -- t[27554] = 2
      "0000010" when "00110101110100011", -- t[27555] = 2
      "0000010" when "00110101110100100", -- t[27556] = 2
      "0000010" when "00110101110100101", -- t[27557] = 2
      "0000010" when "00110101110100110", -- t[27558] = 2
      "0000010" when "00110101110100111", -- t[27559] = 2
      "0000010" when "00110101110101000", -- t[27560] = 2
      "0000010" when "00110101110101001", -- t[27561] = 2
      "0000010" when "00110101110101010", -- t[27562] = 2
      "0000010" when "00110101110101011", -- t[27563] = 2
      "0000010" when "00110101110101100", -- t[27564] = 2
      "0000010" when "00110101110101101", -- t[27565] = 2
      "0000010" when "00110101110101110", -- t[27566] = 2
      "0000010" when "00110101110101111", -- t[27567] = 2
      "0000010" when "00110101110110000", -- t[27568] = 2
      "0000010" when "00110101110110001", -- t[27569] = 2
      "0000010" when "00110101110110010", -- t[27570] = 2
      "0000010" when "00110101110110011", -- t[27571] = 2
      "0000010" when "00110101110110100", -- t[27572] = 2
      "0000010" when "00110101110110101", -- t[27573] = 2
      "0000010" when "00110101110110110", -- t[27574] = 2
      "0000010" when "00110101110110111", -- t[27575] = 2
      "0000010" when "00110101110111000", -- t[27576] = 2
      "0000010" when "00110101110111001", -- t[27577] = 2
      "0000010" when "00110101110111010", -- t[27578] = 2
      "0000010" when "00110101110111011", -- t[27579] = 2
      "0000010" when "00110101110111100", -- t[27580] = 2
      "0000010" when "00110101110111101", -- t[27581] = 2
      "0000010" when "00110101110111110", -- t[27582] = 2
      "0000010" when "00110101110111111", -- t[27583] = 2
      "0000010" when "00110101111000000", -- t[27584] = 2
      "0000010" when "00110101111000001", -- t[27585] = 2
      "0000010" when "00110101111000010", -- t[27586] = 2
      "0000010" when "00110101111000011", -- t[27587] = 2
      "0000010" when "00110101111000100", -- t[27588] = 2
      "0000010" when "00110101111000101", -- t[27589] = 2
      "0000010" when "00110101111000110", -- t[27590] = 2
      "0000010" when "00110101111000111", -- t[27591] = 2
      "0000010" when "00110101111001000", -- t[27592] = 2
      "0000010" when "00110101111001001", -- t[27593] = 2
      "0000010" when "00110101111001010", -- t[27594] = 2
      "0000010" when "00110101111001011", -- t[27595] = 2
      "0000010" when "00110101111001100", -- t[27596] = 2
      "0000010" when "00110101111001101", -- t[27597] = 2
      "0000010" when "00110101111001110", -- t[27598] = 2
      "0000010" when "00110101111001111", -- t[27599] = 2
      "0000010" when "00110101111010000", -- t[27600] = 2
      "0000010" when "00110101111010001", -- t[27601] = 2
      "0000010" when "00110101111010010", -- t[27602] = 2
      "0000010" when "00110101111010011", -- t[27603] = 2
      "0000010" when "00110101111010100", -- t[27604] = 2
      "0000010" when "00110101111010101", -- t[27605] = 2
      "0000010" when "00110101111010110", -- t[27606] = 2
      "0000010" when "00110101111010111", -- t[27607] = 2
      "0000010" when "00110101111011000", -- t[27608] = 2
      "0000010" when "00110101111011001", -- t[27609] = 2
      "0000010" when "00110101111011010", -- t[27610] = 2
      "0000010" when "00110101111011011", -- t[27611] = 2
      "0000010" when "00110101111011100", -- t[27612] = 2
      "0000010" when "00110101111011101", -- t[27613] = 2
      "0000010" when "00110101111011110", -- t[27614] = 2
      "0000010" when "00110101111011111", -- t[27615] = 2
      "0000010" when "00110101111100000", -- t[27616] = 2
      "0000010" when "00110101111100001", -- t[27617] = 2
      "0000010" when "00110101111100010", -- t[27618] = 2
      "0000010" when "00110101111100011", -- t[27619] = 2
      "0000010" when "00110101111100100", -- t[27620] = 2
      "0000010" when "00110101111100101", -- t[27621] = 2
      "0000010" when "00110101111100110", -- t[27622] = 2
      "0000010" when "00110101111100111", -- t[27623] = 2
      "0000010" when "00110101111101000", -- t[27624] = 2
      "0000010" when "00110101111101001", -- t[27625] = 2
      "0000010" when "00110101111101010", -- t[27626] = 2
      "0000010" when "00110101111101011", -- t[27627] = 2
      "0000010" when "00110101111101100", -- t[27628] = 2
      "0000010" when "00110101111101101", -- t[27629] = 2
      "0000010" when "00110101111101110", -- t[27630] = 2
      "0000010" when "00110101111101111", -- t[27631] = 2
      "0000010" when "00110101111110000", -- t[27632] = 2
      "0000010" when "00110101111110001", -- t[27633] = 2
      "0000010" when "00110101111110010", -- t[27634] = 2
      "0000010" when "00110101111110011", -- t[27635] = 2
      "0000010" when "00110101111110100", -- t[27636] = 2
      "0000010" when "00110101111110101", -- t[27637] = 2
      "0000010" when "00110101111110110", -- t[27638] = 2
      "0000010" when "00110101111110111", -- t[27639] = 2
      "0000010" when "00110101111111000", -- t[27640] = 2
      "0000010" when "00110101111111001", -- t[27641] = 2
      "0000010" when "00110101111111010", -- t[27642] = 2
      "0000010" when "00110101111111011", -- t[27643] = 2
      "0000010" when "00110101111111100", -- t[27644] = 2
      "0000010" when "00110101111111101", -- t[27645] = 2
      "0000010" when "00110101111111110", -- t[27646] = 2
      "0000010" when "00110101111111111", -- t[27647] = 2
      "0000010" when "00110110000000000", -- t[27648] = 2
      "0000010" when "00110110000000001", -- t[27649] = 2
      "0000010" when "00110110000000010", -- t[27650] = 2
      "0000010" when "00110110000000011", -- t[27651] = 2
      "0000010" when "00110110000000100", -- t[27652] = 2
      "0000010" when "00110110000000101", -- t[27653] = 2
      "0000010" when "00110110000000110", -- t[27654] = 2
      "0000010" when "00110110000000111", -- t[27655] = 2
      "0000010" when "00110110000001000", -- t[27656] = 2
      "0000010" when "00110110000001001", -- t[27657] = 2
      "0000010" when "00110110000001010", -- t[27658] = 2
      "0000010" when "00110110000001011", -- t[27659] = 2
      "0000010" when "00110110000001100", -- t[27660] = 2
      "0000010" when "00110110000001101", -- t[27661] = 2
      "0000010" when "00110110000001110", -- t[27662] = 2
      "0000010" when "00110110000001111", -- t[27663] = 2
      "0000010" when "00110110000010000", -- t[27664] = 2
      "0000010" when "00110110000010001", -- t[27665] = 2
      "0000010" when "00110110000010010", -- t[27666] = 2
      "0000010" when "00110110000010011", -- t[27667] = 2
      "0000010" when "00110110000010100", -- t[27668] = 2
      "0000010" when "00110110000010101", -- t[27669] = 2
      "0000010" when "00110110000010110", -- t[27670] = 2
      "0000010" when "00110110000010111", -- t[27671] = 2
      "0000010" when "00110110000011000", -- t[27672] = 2
      "0000010" when "00110110000011001", -- t[27673] = 2
      "0000010" when "00110110000011010", -- t[27674] = 2
      "0000010" when "00110110000011011", -- t[27675] = 2
      "0000010" when "00110110000011100", -- t[27676] = 2
      "0000010" when "00110110000011101", -- t[27677] = 2
      "0000010" when "00110110000011110", -- t[27678] = 2
      "0000010" when "00110110000011111", -- t[27679] = 2
      "0000010" when "00110110000100000", -- t[27680] = 2
      "0000010" when "00110110000100001", -- t[27681] = 2
      "0000010" when "00110110000100010", -- t[27682] = 2
      "0000010" when "00110110000100011", -- t[27683] = 2
      "0000010" when "00110110000100100", -- t[27684] = 2
      "0000010" when "00110110000100101", -- t[27685] = 2
      "0000010" when "00110110000100110", -- t[27686] = 2
      "0000010" when "00110110000100111", -- t[27687] = 2
      "0000010" when "00110110000101000", -- t[27688] = 2
      "0000010" when "00110110000101001", -- t[27689] = 2
      "0000010" when "00110110000101010", -- t[27690] = 2
      "0000010" when "00110110000101011", -- t[27691] = 2
      "0000010" when "00110110000101100", -- t[27692] = 2
      "0000010" when "00110110000101101", -- t[27693] = 2
      "0000010" when "00110110000101110", -- t[27694] = 2
      "0000010" when "00110110000101111", -- t[27695] = 2
      "0000010" when "00110110000110000", -- t[27696] = 2
      "0000010" when "00110110000110001", -- t[27697] = 2
      "0000010" when "00110110000110010", -- t[27698] = 2
      "0000010" when "00110110000110011", -- t[27699] = 2
      "0000010" when "00110110000110100", -- t[27700] = 2
      "0000010" when "00110110000110101", -- t[27701] = 2
      "0000010" when "00110110000110110", -- t[27702] = 2
      "0000010" when "00110110000110111", -- t[27703] = 2
      "0000010" when "00110110000111000", -- t[27704] = 2
      "0000010" when "00110110000111001", -- t[27705] = 2
      "0000010" when "00110110000111010", -- t[27706] = 2
      "0000010" when "00110110000111011", -- t[27707] = 2
      "0000010" when "00110110000111100", -- t[27708] = 2
      "0000010" when "00110110000111101", -- t[27709] = 2
      "0000010" when "00110110000111110", -- t[27710] = 2
      "0000010" when "00110110000111111", -- t[27711] = 2
      "0000010" when "00110110001000000", -- t[27712] = 2
      "0000010" when "00110110001000001", -- t[27713] = 2
      "0000010" when "00110110001000010", -- t[27714] = 2
      "0000010" when "00110110001000011", -- t[27715] = 2
      "0000010" when "00110110001000100", -- t[27716] = 2
      "0000010" when "00110110001000101", -- t[27717] = 2
      "0000010" when "00110110001000110", -- t[27718] = 2
      "0000010" when "00110110001000111", -- t[27719] = 2
      "0000010" when "00110110001001000", -- t[27720] = 2
      "0000010" when "00110110001001001", -- t[27721] = 2
      "0000010" when "00110110001001010", -- t[27722] = 2
      "0000010" when "00110110001001011", -- t[27723] = 2
      "0000010" when "00110110001001100", -- t[27724] = 2
      "0000010" when "00110110001001101", -- t[27725] = 2
      "0000010" when "00110110001001110", -- t[27726] = 2
      "0000010" when "00110110001001111", -- t[27727] = 2
      "0000010" when "00110110001010000", -- t[27728] = 2
      "0000010" when "00110110001010001", -- t[27729] = 2
      "0000010" when "00110110001010010", -- t[27730] = 2
      "0000010" when "00110110001010011", -- t[27731] = 2
      "0000010" when "00110110001010100", -- t[27732] = 2
      "0000010" when "00110110001010101", -- t[27733] = 2
      "0000010" when "00110110001010110", -- t[27734] = 2
      "0000010" when "00110110001010111", -- t[27735] = 2
      "0000010" when "00110110001011000", -- t[27736] = 2
      "0000010" when "00110110001011001", -- t[27737] = 2
      "0000010" when "00110110001011010", -- t[27738] = 2
      "0000010" when "00110110001011011", -- t[27739] = 2
      "0000010" when "00110110001011100", -- t[27740] = 2
      "0000010" when "00110110001011101", -- t[27741] = 2
      "0000010" when "00110110001011110", -- t[27742] = 2
      "0000010" when "00110110001011111", -- t[27743] = 2
      "0000010" when "00110110001100000", -- t[27744] = 2
      "0000010" when "00110110001100001", -- t[27745] = 2
      "0000010" when "00110110001100010", -- t[27746] = 2
      "0000010" when "00110110001100011", -- t[27747] = 2
      "0000010" when "00110110001100100", -- t[27748] = 2
      "0000010" when "00110110001100101", -- t[27749] = 2
      "0000010" when "00110110001100110", -- t[27750] = 2
      "0000010" when "00110110001100111", -- t[27751] = 2
      "0000010" when "00110110001101000", -- t[27752] = 2
      "0000010" when "00110110001101001", -- t[27753] = 2
      "0000010" when "00110110001101010", -- t[27754] = 2
      "0000010" when "00110110001101011", -- t[27755] = 2
      "0000010" when "00110110001101100", -- t[27756] = 2
      "0000010" when "00110110001101101", -- t[27757] = 2
      "0000010" when "00110110001101110", -- t[27758] = 2
      "0000010" when "00110110001101111", -- t[27759] = 2
      "0000010" when "00110110001110000", -- t[27760] = 2
      "0000010" when "00110110001110001", -- t[27761] = 2
      "0000010" when "00110110001110010", -- t[27762] = 2
      "0000010" when "00110110001110011", -- t[27763] = 2
      "0000010" when "00110110001110100", -- t[27764] = 2
      "0000010" when "00110110001110101", -- t[27765] = 2
      "0000010" when "00110110001110110", -- t[27766] = 2
      "0000010" when "00110110001110111", -- t[27767] = 2
      "0000010" when "00110110001111000", -- t[27768] = 2
      "0000010" when "00110110001111001", -- t[27769] = 2
      "0000010" when "00110110001111010", -- t[27770] = 2
      "0000010" when "00110110001111011", -- t[27771] = 2
      "0000010" when "00110110001111100", -- t[27772] = 2
      "0000010" when "00110110001111101", -- t[27773] = 2
      "0000010" when "00110110001111110", -- t[27774] = 2
      "0000010" when "00110110001111111", -- t[27775] = 2
      "0000010" when "00110110010000000", -- t[27776] = 2
      "0000010" when "00110110010000001", -- t[27777] = 2
      "0000010" when "00110110010000010", -- t[27778] = 2
      "0000010" when "00110110010000011", -- t[27779] = 2
      "0000010" when "00110110010000100", -- t[27780] = 2
      "0000010" when "00110110010000101", -- t[27781] = 2
      "0000010" when "00110110010000110", -- t[27782] = 2
      "0000010" when "00110110010000111", -- t[27783] = 2
      "0000010" when "00110110010001000", -- t[27784] = 2
      "0000010" when "00110110010001001", -- t[27785] = 2
      "0000010" when "00110110010001010", -- t[27786] = 2
      "0000010" when "00110110010001011", -- t[27787] = 2
      "0000010" when "00110110010001100", -- t[27788] = 2
      "0000010" when "00110110010001101", -- t[27789] = 2
      "0000010" when "00110110010001110", -- t[27790] = 2
      "0000010" when "00110110010001111", -- t[27791] = 2
      "0000010" when "00110110010010000", -- t[27792] = 2
      "0000010" when "00110110010010001", -- t[27793] = 2
      "0000010" when "00110110010010010", -- t[27794] = 2
      "0000010" when "00110110010010011", -- t[27795] = 2
      "0000010" when "00110110010010100", -- t[27796] = 2
      "0000010" when "00110110010010101", -- t[27797] = 2
      "0000010" when "00110110010010110", -- t[27798] = 2
      "0000010" when "00110110010010111", -- t[27799] = 2
      "0000010" when "00110110010011000", -- t[27800] = 2
      "0000010" when "00110110010011001", -- t[27801] = 2
      "0000010" when "00110110010011010", -- t[27802] = 2
      "0000010" when "00110110010011011", -- t[27803] = 2
      "0000010" when "00110110010011100", -- t[27804] = 2
      "0000010" when "00110110010011101", -- t[27805] = 2
      "0000010" when "00110110010011110", -- t[27806] = 2
      "0000010" when "00110110010011111", -- t[27807] = 2
      "0000010" when "00110110010100000", -- t[27808] = 2
      "0000010" when "00110110010100001", -- t[27809] = 2
      "0000010" when "00110110010100010", -- t[27810] = 2
      "0000010" when "00110110010100011", -- t[27811] = 2
      "0000010" when "00110110010100100", -- t[27812] = 2
      "0000010" when "00110110010100101", -- t[27813] = 2
      "0000010" when "00110110010100110", -- t[27814] = 2
      "0000010" when "00110110010100111", -- t[27815] = 2
      "0000010" when "00110110010101000", -- t[27816] = 2
      "0000010" when "00110110010101001", -- t[27817] = 2
      "0000010" when "00110110010101010", -- t[27818] = 2
      "0000010" when "00110110010101011", -- t[27819] = 2
      "0000010" when "00110110010101100", -- t[27820] = 2
      "0000010" when "00110110010101101", -- t[27821] = 2
      "0000010" when "00110110010101110", -- t[27822] = 2
      "0000010" when "00110110010101111", -- t[27823] = 2
      "0000010" when "00110110010110000", -- t[27824] = 2
      "0000010" when "00110110010110001", -- t[27825] = 2
      "0000010" when "00110110010110010", -- t[27826] = 2
      "0000010" when "00110110010110011", -- t[27827] = 2
      "0000010" when "00110110010110100", -- t[27828] = 2
      "0000010" when "00110110010110101", -- t[27829] = 2
      "0000010" when "00110110010110110", -- t[27830] = 2
      "0000010" when "00110110010110111", -- t[27831] = 2
      "0000010" when "00110110010111000", -- t[27832] = 2
      "0000010" when "00110110010111001", -- t[27833] = 2
      "0000010" when "00110110010111010", -- t[27834] = 2
      "0000010" when "00110110010111011", -- t[27835] = 2
      "0000010" when "00110110010111100", -- t[27836] = 2
      "0000010" when "00110110010111101", -- t[27837] = 2
      "0000010" when "00110110010111110", -- t[27838] = 2
      "0000010" when "00110110010111111", -- t[27839] = 2
      "0000010" when "00110110011000000", -- t[27840] = 2
      "0000010" when "00110110011000001", -- t[27841] = 2
      "0000010" when "00110110011000010", -- t[27842] = 2
      "0000010" when "00110110011000011", -- t[27843] = 2
      "0000010" when "00110110011000100", -- t[27844] = 2
      "0000010" when "00110110011000101", -- t[27845] = 2
      "0000010" when "00110110011000110", -- t[27846] = 2
      "0000010" when "00110110011000111", -- t[27847] = 2
      "0000010" when "00110110011001000", -- t[27848] = 2
      "0000010" when "00110110011001001", -- t[27849] = 2
      "0000010" when "00110110011001010", -- t[27850] = 2
      "0000010" when "00110110011001011", -- t[27851] = 2
      "0000010" when "00110110011001100", -- t[27852] = 2
      "0000010" when "00110110011001101", -- t[27853] = 2
      "0000010" when "00110110011001110", -- t[27854] = 2
      "0000010" when "00110110011001111", -- t[27855] = 2
      "0000010" when "00110110011010000", -- t[27856] = 2
      "0000010" when "00110110011010001", -- t[27857] = 2
      "0000010" when "00110110011010010", -- t[27858] = 2
      "0000010" when "00110110011010011", -- t[27859] = 2
      "0000010" when "00110110011010100", -- t[27860] = 2
      "0000010" when "00110110011010101", -- t[27861] = 2
      "0000010" when "00110110011010110", -- t[27862] = 2
      "0000010" when "00110110011010111", -- t[27863] = 2
      "0000010" when "00110110011011000", -- t[27864] = 2
      "0000010" when "00110110011011001", -- t[27865] = 2
      "0000010" when "00110110011011010", -- t[27866] = 2
      "0000010" when "00110110011011011", -- t[27867] = 2
      "0000010" when "00110110011011100", -- t[27868] = 2
      "0000010" when "00110110011011101", -- t[27869] = 2
      "0000010" when "00110110011011110", -- t[27870] = 2
      "0000010" when "00110110011011111", -- t[27871] = 2
      "0000010" when "00110110011100000", -- t[27872] = 2
      "0000010" when "00110110011100001", -- t[27873] = 2
      "0000010" when "00110110011100010", -- t[27874] = 2
      "0000010" when "00110110011100011", -- t[27875] = 2
      "0000010" when "00110110011100100", -- t[27876] = 2
      "0000010" when "00110110011100101", -- t[27877] = 2
      "0000010" when "00110110011100110", -- t[27878] = 2
      "0000010" when "00110110011100111", -- t[27879] = 2
      "0000010" when "00110110011101000", -- t[27880] = 2
      "0000010" when "00110110011101001", -- t[27881] = 2
      "0000010" when "00110110011101010", -- t[27882] = 2
      "0000010" when "00110110011101011", -- t[27883] = 2
      "0000010" when "00110110011101100", -- t[27884] = 2
      "0000010" when "00110110011101101", -- t[27885] = 2
      "0000010" when "00110110011101110", -- t[27886] = 2
      "0000010" when "00110110011101111", -- t[27887] = 2
      "0000010" when "00110110011110000", -- t[27888] = 2
      "0000010" when "00110110011110001", -- t[27889] = 2
      "0000010" when "00110110011110010", -- t[27890] = 2
      "0000010" when "00110110011110011", -- t[27891] = 2
      "0000010" when "00110110011110100", -- t[27892] = 2
      "0000010" when "00110110011110101", -- t[27893] = 2
      "0000010" when "00110110011110110", -- t[27894] = 2
      "0000010" when "00110110011110111", -- t[27895] = 2
      "0000010" when "00110110011111000", -- t[27896] = 2
      "0000010" when "00110110011111001", -- t[27897] = 2
      "0000010" when "00110110011111010", -- t[27898] = 2
      "0000010" when "00110110011111011", -- t[27899] = 2
      "0000010" when "00110110011111100", -- t[27900] = 2
      "0000010" when "00110110011111101", -- t[27901] = 2
      "0000010" when "00110110011111110", -- t[27902] = 2
      "0000010" when "00110110011111111", -- t[27903] = 2
      "0000010" when "00110110100000000", -- t[27904] = 2
      "0000010" when "00110110100000001", -- t[27905] = 2
      "0000010" when "00110110100000010", -- t[27906] = 2
      "0000010" when "00110110100000011", -- t[27907] = 2
      "0000010" when "00110110100000100", -- t[27908] = 2
      "0000010" when "00110110100000101", -- t[27909] = 2
      "0000010" when "00110110100000110", -- t[27910] = 2
      "0000010" when "00110110100000111", -- t[27911] = 2
      "0000010" when "00110110100001000", -- t[27912] = 2
      "0000010" when "00110110100001001", -- t[27913] = 2
      "0000010" when "00110110100001010", -- t[27914] = 2
      "0000010" when "00110110100001011", -- t[27915] = 2
      "0000010" when "00110110100001100", -- t[27916] = 2
      "0000010" when "00110110100001101", -- t[27917] = 2
      "0000010" when "00110110100001110", -- t[27918] = 2
      "0000010" when "00110110100001111", -- t[27919] = 2
      "0000010" when "00110110100010000", -- t[27920] = 2
      "0000010" when "00110110100010001", -- t[27921] = 2
      "0000010" when "00110110100010010", -- t[27922] = 2
      "0000010" when "00110110100010011", -- t[27923] = 2
      "0000010" when "00110110100010100", -- t[27924] = 2
      "0000010" when "00110110100010101", -- t[27925] = 2
      "0000010" when "00110110100010110", -- t[27926] = 2
      "0000010" when "00110110100010111", -- t[27927] = 2
      "0000010" when "00110110100011000", -- t[27928] = 2
      "0000010" when "00110110100011001", -- t[27929] = 2
      "0000010" when "00110110100011010", -- t[27930] = 2
      "0000010" when "00110110100011011", -- t[27931] = 2
      "0000010" when "00110110100011100", -- t[27932] = 2
      "0000010" when "00110110100011101", -- t[27933] = 2
      "0000010" when "00110110100011110", -- t[27934] = 2
      "0000010" when "00110110100011111", -- t[27935] = 2
      "0000010" when "00110110100100000", -- t[27936] = 2
      "0000010" when "00110110100100001", -- t[27937] = 2
      "0000010" when "00110110100100010", -- t[27938] = 2
      "0000010" when "00110110100100011", -- t[27939] = 2
      "0000010" when "00110110100100100", -- t[27940] = 2
      "0000010" when "00110110100100101", -- t[27941] = 2
      "0000010" when "00110110100100110", -- t[27942] = 2
      "0000010" when "00110110100100111", -- t[27943] = 2
      "0000010" when "00110110100101000", -- t[27944] = 2
      "0000010" when "00110110100101001", -- t[27945] = 2
      "0000010" when "00110110100101010", -- t[27946] = 2
      "0000010" when "00110110100101011", -- t[27947] = 2
      "0000010" when "00110110100101100", -- t[27948] = 2
      "0000010" when "00110110100101101", -- t[27949] = 2
      "0000010" when "00110110100101110", -- t[27950] = 2
      "0000010" when "00110110100101111", -- t[27951] = 2
      "0000010" when "00110110100110000", -- t[27952] = 2
      "0000010" when "00110110100110001", -- t[27953] = 2
      "0000010" when "00110110100110010", -- t[27954] = 2
      "0000010" when "00110110100110011", -- t[27955] = 2
      "0000010" when "00110110100110100", -- t[27956] = 2
      "0000010" when "00110110100110101", -- t[27957] = 2
      "0000010" when "00110110100110110", -- t[27958] = 2
      "0000010" when "00110110100110111", -- t[27959] = 2
      "0000010" when "00110110100111000", -- t[27960] = 2
      "0000010" when "00110110100111001", -- t[27961] = 2
      "0000010" when "00110110100111010", -- t[27962] = 2
      "0000010" when "00110110100111011", -- t[27963] = 2
      "0000010" when "00110110100111100", -- t[27964] = 2
      "0000010" when "00110110100111101", -- t[27965] = 2
      "0000010" when "00110110100111110", -- t[27966] = 2
      "0000010" when "00110110100111111", -- t[27967] = 2
      "0000010" when "00110110101000000", -- t[27968] = 2
      "0000010" when "00110110101000001", -- t[27969] = 2
      "0000010" when "00110110101000010", -- t[27970] = 2
      "0000010" when "00110110101000011", -- t[27971] = 2
      "0000010" when "00110110101000100", -- t[27972] = 2
      "0000010" when "00110110101000101", -- t[27973] = 2
      "0000010" when "00110110101000110", -- t[27974] = 2
      "0000010" when "00110110101000111", -- t[27975] = 2
      "0000010" when "00110110101001000", -- t[27976] = 2
      "0000010" when "00110110101001001", -- t[27977] = 2
      "0000010" when "00110110101001010", -- t[27978] = 2
      "0000010" when "00110110101001011", -- t[27979] = 2
      "0000010" when "00110110101001100", -- t[27980] = 2
      "0000010" when "00110110101001101", -- t[27981] = 2
      "0000010" when "00110110101001110", -- t[27982] = 2
      "0000010" when "00110110101001111", -- t[27983] = 2
      "0000010" when "00110110101010000", -- t[27984] = 2
      "0000010" when "00110110101010001", -- t[27985] = 2
      "0000010" when "00110110101010010", -- t[27986] = 2
      "0000010" when "00110110101010011", -- t[27987] = 2
      "0000010" when "00110110101010100", -- t[27988] = 2
      "0000010" when "00110110101010101", -- t[27989] = 2
      "0000010" when "00110110101010110", -- t[27990] = 2
      "0000010" when "00110110101010111", -- t[27991] = 2
      "0000010" when "00110110101011000", -- t[27992] = 2
      "0000010" when "00110110101011001", -- t[27993] = 2
      "0000010" when "00110110101011010", -- t[27994] = 2
      "0000010" when "00110110101011011", -- t[27995] = 2
      "0000010" when "00110110101011100", -- t[27996] = 2
      "0000010" when "00110110101011101", -- t[27997] = 2
      "0000010" when "00110110101011110", -- t[27998] = 2
      "0000010" when "00110110101011111", -- t[27999] = 2
      "0000010" when "00110110101100000", -- t[28000] = 2
      "0000010" when "00110110101100001", -- t[28001] = 2
      "0000010" when "00110110101100010", -- t[28002] = 2
      "0000010" when "00110110101100011", -- t[28003] = 2
      "0000010" when "00110110101100100", -- t[28004] = 2
      "0000010" when "00110110101100101", -- t[28005] = 2
      "0000010" when "00110110101100110", -- t[28006] = 2
      "0000010" when "00110110101100111", -- t[28007] = 2
      "0000010" when "00110110101101000", -- t[28008] = 2
      "0000010" when "00110110101101001", -- t[28009] = 2
      "0000010" when "00110110101101010", -- t[28010] = 2
      "0000010" when "00110110101101011", -- t[28011] = 2
      "0000010" when "00110110101101100", -- t[28012] = 2
      "0000010" when "00110110101101101", -- t[28013] = 2
      "0000010" when "00110110101101110", -- t[28014] = 2
      "0000010" when "00110110101101111", -- t[28015] = 2
      "0000010" when "00110110101110000", -- t[28016] = 2
      "0000010" when "00110110101110001", -- t[28017] = 2
      "0000010" when "00110110101110010", -- t[28018] = 2
      "0000010" when "00110110101110011", -- t[28019] = 2
      "0000010" when "00110110101110100", -- t[28020] = 2
      "0000010" when "00110110101110101", -- t[28021] = 2
      "0000010" when "00110110101110110", -- t[28022] = 2
      "0000010" when "00110110101110111", -- t[28023] = 2
      "0000010" when "00110110101111000", -- t[28024] = 2
      "0000010" when "00110110101111001", -- t[28025] = 2
      "0000010" when "00110110101111010", -- t[28026] = 2
      "0000010" when "00110110101111011", -- t[28027] = 2
      "0000010" when "00110110101111100", -- t[28028] = 2
      "0000010" when "00110110101111101", -- t[28029] = 2
      "0000010" when "00110110101111110", -- t[28030] = 2
      "0000010" when "00110110101111111", -- t[28031] = 2
      "0000010" when "00110110110000000", -- t[28032] = 2
      "0000010" when "00110110110000001", -- t[28033] = 2
      "0000010" when "00110110110000010", -- t[28034] = 2
      "0000010" when "00110110110000011", -- t[28035] = 2
      "0000010" when "00110110110000100", -- t[28036] = 2
      "0000010" when "00110110110000101", -- t[28037] = 2
      "0000010" when "00110110110000110", -- t[28038] = 2
      "0000010" when "00110110110000111", -- t[28039] = 2
      "0000010" when "00110110110001000", -- t[28040] = 2
      "0000010" when "00110110110001001", -- t[28041] = 2
      "0000010" when "00110110110001010", -- t[28042] = 2
      "0000010" when "00110110110001011", -- t[28043] = 2
      "0000010" when "00110110110001100", -- t[28044] = 2
      "0000010" when "00110110110001101", -- t[28045] = 2
      "0000010" when "00110110110001110", -- t[28046] = 2
      "0000010" when "00110110110001111", -- t[28047] = 2
      "0000010" when "00110110110010000", -- t[28048] = 2
      "0000010" when "00110110110010001", -- t[28049] = 2
      "0000010" when "00110110110010010", -- t[28050] = 2
      "0000010" when "00110110110010011", -- t[28051] = 2
      "0000010" when "00110110110010100", -- t[28052] = 2
      "0000010" when "00110110110010101", -- t[28053] = 2
      "0000010" when "00110110110010110", -- t[28054] = 2
      "0000010" when "00110110110010111", -- t[28055] = 2
      "0000010" when "00110110110011000", -- t[28056] = 2
      "0000010" when "00110110110011001", -- t[28057] = 2
      "0000010" when "00110110110011010", -- t[28058] = 2
      "0000010" when "00110110110011011", -- t[28059] = 2
      "0000010" when "00110110110011100", -- t[28060] = 2
      "0000010" when "00110110110011101", -- t[28061] = 2
      "0000010" when "00110110110011110", -- t[28062] = 2
      "0000010" when "00110110110011111", -- t[28063] = 2
      "0000010" when "00110110110100000", -- t[28064] = 2
      "0000010" when "00110110110100001", -- t[28065] = 2
      "0000010" when "00110110110100010", -- t[28066] = 2
      "0000010" when "00110110110100011", -- t[28067] = 2
      "0000010" when "00110110110100100", -- t[28068] = 2
      "0000010" when "00110110110100101", -- t[28069] = 2
      "0000010" when "00110110110100110", -- t[28070] = 2
      "0000010" when "00110110110100111", -- t[28071] = 2
      "0000010" when "00110110110101000", -- t[28072] = 2
      "0000010" when "00110110110101001", -- t[28073] = 2
      "0000010" when "00110110110101010", -- t[28074] = 2
      "0000010" when "00110110110101011", -- t[28075] = 2
      "0000010" when "00110110110101100", -- t[28076] = 2
      "0000010" when "00110110110101101", -- t[28077] = 2
      "0000010" when "00110110110101110", -- t[28078] = 2
      "0000010" when "00110110110101111", -- t[28079] = 2
      "0000010" when "00110110110110000", -- t[28080] = 2
      "0000010" when "00110110110110001", -- t[28081] = 2
      "0000010" when "00110110110110010", -- t[28082] = 2
      "0000010" when "00110110110110011", -- t[28083] = 2
      "0000010" when "00110110110110100", -- t[28084] = 2
      "0000010" when "00110110110110101", -- t[28085] = 2
      "0000010" when "00110110110110110", -- t[28086] = 2
      "0000010" when "00110110110110111", -- t[28087] = 2
      "0000010" when "00110110110111000", -- t[28088] = 2
      "0000010" when "00110110110111001", -- t[28089] = 2
      "0000010" when "00110110110111010", -- t[28090] = 2
      "0000010" when "00110110110111011", -- t[28091] = 2
      "0000010" when "00110110110111100", -- t[28092] = 2
      "0000010" when "00110110110111101", -- t[28093] = 2
      "0000010" when "00110110110111110", -- t[28094] = 2
      "0000010" when "00110110110111111", -- t[28095] = 2
      "0000010" when "00110110111000000", -- t[28096] = 2
      "0000010" when "00110110111000001", -- t[28097] = 2
      "0000010" when "00110110111000010", -- t[28098] = 2
      "0000010" when "00110110111000011", -- t[28099] = 2
      "0000010" when "00110110111000100", -- t[28100] = 2
      "0000010" when "00110110111000101", -- t[28101] = 2
      "0000010" when "00110110111000110", -- t[28102] = 2
      "0000010" when "00110110111000111", -- t[28103] = 2
      "0000010" when "00110110111001000", -- t[28104] = 2
      "0000010" when "00110110111001001", -- t[28105] = 2
      "0000010" when "00110110111001010", -- t[28106] = 2
      "0000010" when "00110110111001011", -- t[28107] = 2
      "0000010" when "00110110111001100", -- t[28108] = 2
      "0000010" when "00110110111001101", -- t[28109] = 2
      "0000010" when "00110110111001110", -- t[28110] = 2
      "0000010" when "00110110111001111", -- t[28111] = 2
      "0000010" when "00110110111010000", -- t[28112] = 2
      "0000010" when "00110110111010001", -- t[28113] = 2
      "0000010" when "00110110111010010", -- t[28114] = 2
      "0000010" when "00110110111010011", -- t[28115] = 2
      "0000010" when "00110110111010100", -- t[28116] = 2
      "0000010" when "00110110111010101", -- t[28117] = 2
      "0000010" when "00110110111010110", -- t[28118] = 2
      "0000010" when "00110110111010111", -- t[28119] = 2
      "0000010" when "00110110111011000", -- t[28120] = 2
      "0000010" when "00110110111011001", -- t[28121] = 2
      "0000010" when "00110110111011010", -- t[28122] = 2
      "0000010" when "00110110111011011", -- t[28123] = 2
      "0000010" when "00110110111011100", -- t[28124] = 2
      "0000010" when "00110110111011101", -- t[28125] = 2
      "0000010" when "00110110111011110", -- t[28126] = 2
      "0000010" when "00110110111011111", -- t[28127] = 2
      "0000010" when "00110110111100000", -- t[28128] = 2
      "0000010" when "00110110111100001", -- t[28129] = 2
      "0000010" when "00110110111100010", -- t[28130] = 2
      "0000010" when "00110110111100011", -- t[28131] = 2
      "0000010" when "00110110111100100", -- t[28132] = 2
      "0000010" when "00110110111100101", -- t[28133] = 2
      "0000010" when "00110110111100110", -- t[28134] = 2
      "0000010" when "00110110111100111", -- t[28135] = 2
      "0000010" when "00110110111101000", -- t[28136] = 2
      "0000010" when "00110110111101001", -- t[28137] = 2
      "0000010" when "00110110111101010", -- t[28138] = 2
      "0000010" when "00110110111101011", -- t[28139] = 2
      "0000010" when "00110110111101100", -- t[28140] = 2
      "0000010" when "00110110111101101", -- t[28141] = 2
      "0000010" when "00110110111101110", -- t[28142] = 2
      "0000010" when "00110110111101111", -- t[28143] = 2
      "0000010" when "00110110111110000", -- t[28144] = 2
      "0000010" when "00110110111110001", -- t[28145] = 2
      "0000010" when "00110110111110010", -- t[28146] = 2
      "0000010" when "00110110111110011", -- t[28147] = 2
      "0000010" when "00110110111110100", -- t[28148] = 2
      "0000010" when "00110110111110101", -- t[28149] = 2
      "0000010" when "00110110111110110", -- t[28150] = 2
      "0000010" when "00110110111110111", -- t[28151] = 2
      "0000010" when "00110110111111000", -- t[28152] = 2
      "0000010" when "00110110111111001", -- t[28153] = 2
      "0000010" when "00110110111111010", -- t[28154] = 2
      "0000010" when "00110110111111011", -- t[28155] = 2
      "0000010" when "00110110111111100", -- t[28156] = 2
      "0000010" when "00110110111111101", -- t[28157] = 2
      "0000010" when "00110110111111110", -- t[28158] = 2
      "0000010" when "00110110111111111", -- t[28159] = 2
      "0000010" when "00110111000000000", -- t[28160] = 2
      "0000010" when "00110111000000001", -- t[28161] = 2
      "0000010" when "00110111000000010", -- t[28162] = 2
      "0000010" when "00110111000000011", -- t[28163] = 2
      "0000010" when "00110111000000100", -- t[28164] = 2
      "0000010" when "00110111000000101", -- t[28165] = 2
      "0000010" when "00110111000000110", -- t[28166] = 2
      "0000010" when "00110111000000111", -- t[28167] = 2
      "0000010" when "00110111000001000", -- t[28168] = 2
      "0000010" when "00110111000001001", -- t[28169] = 2
      "0000010" when "00110111000001010", -- t[28170] = 2
      "0000010" when "00110111000001011", -- t[28171] = 2
      "0000010" when "00110111000001100", -- t[28172] = 2
      "0000010" when "00110111000001101", -- t[28173] = 2
      "0000010" when "00110111000001110", -- t[28174] = 2
      "0000010" when "00110111000001111", -- t[28175] = 2
      "0000010" when "00110111000010000", -- t[28176] = 2
      "0000010" when "00110111000010001", -- t[28177] = 2
      "0000010" when "00110111000010010", -- t[28178] = 2
      "0000010" when "00110111000010011", -- t[28179] = 2
      "0000010" when "00110111000010100", -- t[28180] = 2
      "0000010" when "00110111000010101", -- t[28181] = 2
      "0000010" when "00110111000010110", -- t[28182] = 2
      "0000010" when "00110111000010111", -- t[28183] = 2
      "0000010" when "00110111000011000", -- t[28184] = 2
      "0000010" when "00110111000011001", -- t[28185] = 2
      "0000010" when "00110111000011010", -- t[28186] = 2
      "0000010" when "00110111000011011", -- t[28187] = 2
      "0000010" when "00110111000011100", -- t[28188] = 2
      "0000010" when "00110111000011101", -- t[28189] = 2
      "0000010" when "00110111000011110", -- t[28190] = 2
      "0000010" when "00110111000011111", -- t[28191] = 2
      "0000010" when "00110111000100000", -- t[28192] = 2
      "0000010" when "00110111000100001", -- t[28193] = 2
      "0000010" when "00110111000100010", -- t[28194] = 2
      "0000010" when "00110111000100011", -- t[28195] = 2
      "0000010" when "00110111000100100", -- t[28196] = 2
      "0000010" when "00110111000100101", -- t[28197] = 2
      "0000010" when "00110111000100110", -- t[28198] = 2
      "0000010" when "00110111000100111", -- t[28199] = 2
      "0000010" when "00110111000101000", -- t[28200] = 2
      "0000010" when "00110111000101001", -- t[28201] = 2
      "0000010" when "00110111000101010", -- t[28202] = 2
      "0000010" when "00110111000101011", -- t[28203] = 2
      "0000010" when "00110111000101100", -- t[28204] = 2
      "0000010" when "00110111000101101", -- t[28205] = 2
      "0000010" when "00110111000101110", -- t[28206] = 2
      "0000010" when "00110111000101111", -- t[28207] = 2
      "0000010" when "00110111000110000", -- t[28208] = 2
      "0000010" when "00110111000110001", -- t[28209] = 2
      "0000010" when "00110111000110010", -- t[28210] = 2
      "0000010" when "00110111000110011", -- t[28211] = 2
      "0000010" when "00110111000110100", -- t[28212] = 2
      "0000010" when "00110111000110101", -- t[28213] = 2
      "0000010" when "00110111000110110", -- t[28214] = 2
      "0000010" when "00110111000110111", -- t[28215] = 2
      "0000010" when "00110111000111000", -- t[28216] = 2
      "0000010" when "00110111000111001", -- t[28217] = 2
      "0000010" when "00110111000111010", -- t[28218] = 2
      "0000010" when "00110111000111011", -- t[28219] = 2
      "0000010" when "00110111000111100", -- t[28220] = 2
      "0000010" when "00110111000111101", -- t[28221] = 2
      "0000010" when "00110111000111110", -- t[28222] = 2
      "0000010" when "00110111000111111", -- t[28223] = 2
      "0000010" when "00110111001000000", -- t[28224] = 2
      "0000010" when "00110111001000001", -- t[28225] = 2
      "0000010" when "00110111001000010", -- t[28226] = 2
      "0000010" when "00110111001000011", -- t[28227] = 2
      "0000010" when "00110111001000100", -- t[28228] = 2
      "0000010" when "00110111001000101", -- t[28229] = 2
      "0000010" when "00110111001000110", -- t[28230] = 2
      "0000010" when "00110111001000111", -- t[28231] = 2
      "0000010" when "00110111001001000", -- t[28232] = 2
      "0000010" when "00110111001001001", -- t[28233] = 2
      "0000010" when "00110111001001010", -- t[28234] = 2
      "0000010" when "00110111001001011", -- t[28235] = 2
      "0000010" when "00110111001001100", -- t[28236] = 2
      "0000010" when "00110111001001101", -- t[28237] = 2
      "0000010" when "00110111001001110", -- t[28238] = 2
      "0000010" when "00110111001001111", -- t[28239] = 2
      "0000010" when "00110111001010000", -- t[28240] = 2
      "0000010" when "00110111001010001", -- t[28241] = 2
      "0000010" when "00110111001010010", -- t[28242] = 2
      "0000010" when "00110111001010011", -- t[28243] = 2
      "0000010" when "00110111001010100", -- t[28244] = 2
      "0000010" when "00110111001010101", -- t[28245] = 2
      "0000010" when "00110111001010110", -- t[28246] = 2
      "0000010" when "00110111001010111", -- t[28247] = 2
      "0000010" when "00110111001011000", -- t[28248] = 2
      "0000010" when "00110111001011001", -- t[28249] = 2
      "0000010" when "00110111001011010", -- t[28250] = 2
      "0000010" when "00110111001011011", -- t[28251] = 2
      "0000010" when "00110111001011100", -- t[28252] = 2
      "0000010" when "00110111001011101", -- t[28253] = 2
      "0000010" when "00110111001011110", -- t[28254] = 2
      "0000010" when "00110111001011111", -- t[28255] = 2
      "0000010" when "00110111001100000", -- t[28256] = 2
      "0000010" when "00110111001100001", -- t[28257] = 2
      "0000010" when "00110111001100010", -- t[28258] = 2
      "0000010" when "00110111001100011", -- t[28259] = 2
      "0000010" when "00110111001100100", -- t[28260] = 2
      "0000010" when "00110111001100101", -- t[28261] = 2
      "0000010" when "00110111001100110", -- t[28262] = 2
      "0000010" when "00110111001100111", -- t[28263] = 2
      "0000010" when "00110111001101000", -- t[28264] = 2
      "0000010" when "00110111001101001", -- t[28265] = 2
      "0000010" when "00110111001101010", -- t[28266] = 2
      "0000010" when "00110111001101011", -- t[28267] = 2
      "0000010" when "00110111001101100", -- t[28268] = 2
      "0000010" when "00110111001101101", -- t[28269] = 2
      "0000010" when "00110111001101110", -- t[28270] = 2
      "0000010" when "00110111001101111", -- t[28271] = 2
      "0000010" when "00110111001110000", -- t[28272] = 2
      "0000010" when "00110111001110001", -- t[28273] = 2
      "0000010" when "00110111001110010", -- t[28274] = 2
      "0000010" when "00110111001110011", -- t[28275] = 2
      "0000010" when "00110111001110100", -- t[28276] = 2
      "0000010" when "00110111001110101", -- t[28277] = 2
      "0000010" when "00110111001110110", -- t[28278] = 2
      "0000010" when "00110111001110111", -- t[28279] = 2
      "0000010" when "00110111001111000", -- t[28280] = 2
      "0000010" when "00110111001111001", -- t[28281] = 2
      "0000010" when "00110111001111010", -- t[28282] = 2
      "0000010" when "00110111001111011", -- t[28283] = 2
      "0000010" when "00110111001111100", -- t[28284] = 2
      "0000010" when "00110111001111101", -- t[28285] = 2
      "0000010" when "00110111001111110", -- t[28286] = 2
      "0000010" when "00110111001111111", -- t[28287] = 2
      "0000010" when "00110111010000000", -- t[28288] = 2
      "0000010" when "00110111010000001", -- t[28289] = 2
      "0000010" when "00110111010000010", -- t[28290] = 2
      "0000010" when "00110111010000011", -- t[28291] = 2
      "0000010" when "00110111010000100", -- t[28292] = 2
      "0000010" when "00110111010000101", -- t[28293] = 2
      "0000010" when "00110111010000110", -- t[28294] = 2
      "0000010" when "00110111010000111", -- t[28295] = 2
      "0000010" when "00110111010001000", -- t[28296] = 2
      "0000010" when "00110111010001001", -- t[28297] = 2
      "0000010" when "00110111010001010", -- t[28298] = 2
      "0000010" when "00110111010001011", -- t[28299] = 2
      "0000010" when "00110111010001100", -- t[28300] = 2
      "0000010" when "00110111010001101", -- t[28301] = 2
      "0000010" when "00110111010001110", -- t[28302] = 2
      "0000010" when "00110111010001111", -- t[28303] = 2
      "0000010" when "00110111010010000", -- t[28304] = 2
      "0000010" when "00110111010010001", -- t[28305] = 2
      "0000010" when "00110111010010010", -- t[28306] = 2
      "0000010" when "00110111010010011", -- t[28307] = 2
      "0000010" when "00110111010010100", -- t[28308] = 2
      "0000010" when "00110111010010101", -- t[28309] = 2
      "0000010" when "00110111010010110", -- t[28310] = 2
      "0000010" when "00110111010010111", -- t[28311] = 2
      "0000010" when "00110111010011000", -- t[28312] = 2
      "0000010" when "00110111010011001", -- t[28313] = 2
      "0000010" when "00110111010011010", -- t[28314] = 2
      "0000010" when "00110111010011011", -- t[28315] = 2
      "0000010" when "00110111010011100", -- t[28316] = 2
      "0000010" when "00110111010011101", -- t[28317] = 2
      "0000010" when "00110111010011110", -- t[28318] = 2
      "0000010" when "00110111010011111", -- t[28319] = 2
      "0000010" when "00110111010100000", -- t[28320] = 2
      "0000010" when "00110111010100001", -- t[28321] = 2
      "0000010" when "00110111010100010", -- t[28322] = 2
      "0000010" when "00110111010100011", -- t[28323] = 2
      "0000010" when "00110111010100100", -- t[28324] = 2
      "0000010" when "00110111010100101", -- t[28325] = 2
      "0000010" when "00110111010100110", -- t[28326] = 2
      "0000010" when "00110111010100111", -- t[28327] = 2
      "0000010" when "00110111010101000", -- t[28328] = 2
      "0000010" when "00110111010101001", -- t[28329] = 2
      "0000010" when "00110111010101010", -- t[28330] = 2
      "0000010" when "00110111010101011", -- t[28331] = 2
      "0000010" when "00110111010101100", -- t[28332] = 2
      "0000010" when "00110111010101101", -- t[28333] = 2
      "0000010" when "00110111010101110", -- t[28334] = 2
      "0000010" when "00110111010101111", -- t[28335] = 2
      "0000010" when "00110111010110000", -- t[28336] = 2
      "0000010" when "00110111010110001", -- t[28337] = 2
      "0000010" when "00110111010110010", -- t[28338] = 2
      "0000010" when "00110111010110011", -- t[28339] = 2
      "0000010" when "00110111010110100", -- t[28340] = 2
      "0000010" when "00110111010110101", -- t[28341] = 2
      "0000010" when "00110111010110110", -- t[28342] = 2
      "0000010" when "00110111010110111", -- t[28343] = 2
      "0000010" when "00110111010111000", -- t[28344] = 2
      "0000010" when "00110111010111001", -- t[28345] = 2
      "0000010" when "00110111010111010", -- t[28346] = 2
      "0000010" when "00110111010111011", -- t[28347] = 2
      "0000010" when "00110111010111100", -- t[28348] = 2
      "0000010" when "00110111010111101", -- t[28349] = 2
      "0000010" when "00110111010111110", -- t[28350] = 2
      "0000010" when "00110111010111111", -- t[28351] = 2
      "0000010" when "00110111011000000", -- t[28352] = 2
      "0000010" when "00110111011000001", -- t[28353] = 2
      "0000010" when "00110111011000010", -- t[28354] = 2
      "0000010" when "00110111011000011", -- t[28355] = 2
      "0000010" when "00110111011000100", -- t[28356] = 2
      "0000010" when "00110111011000101", -- t[28357] = 2
      "0000010" when "00110111011000110", -- t[28358] = 2
      "0000010" when "00110111011000111", -- t[28359] = 2
      "0000010" when "00110111011001000", -- t[28360] = 2
      "0000010" when "00110111011001001", -- t[28361] = 2
      "0000010" when "00110111011001010", -- t[28362] = 2
      "0000010" when "00110111011001011", -- t[28363] = 2
      "0000010" when "00110111011001100", -- t[28364] = 2
      "0000010" when "00110111011001101", -- t[28365] = 2
      "0000010" when "00110111011001110", -- t[28366] = 2
      "0000010" when "00110111011001111", -- t[28367] = 2
      "0000010" when "00110111011010000", -- t[28368] = 2
      "0000010" when "00110111011010001", -- t[28369] = 2
      "0000010" when "00110111011010010", -- t[28370] = 2
      "0000010" when "00110111011010011", -- t[28371] = 2
      "0000010" when "00110111011010100", -- t[28372] = 2
      "0000010" when "00110111011010101", -- t[28373] = 2
      "0000010" when "00110111011010110", -- t[28374] = 2
      "0000010" when "00110111011010111", -- t[28375] = 2
      "0000010" when "00110111011011000", -- t[28376] = 2
      "0000010" when "00110111011011001", -- t[28377] = 2
      "0000010" when "00110111011011010", -- t[28378] = 2
      "0000010" when "00110111011011011", -- t[28379] = 2
      "0000010" when "00110111011011100", -- t[28380] = 2
      "0000010" when "00110111011011101", -- t[28381] = 2
      "0000010" when "00110111011011110", -- t[28382] = 2
      "0000010" when "00110111011011111", -- t[28383] = 2
      "0000010" when "00110111011100000", -- t[28384] = 2
      "0000010" when "00110111011100001", -- t[28385] = 2
      "0000010" when "00110111011100010", -- t[28386] = 2
      "0000010" when "00110111011100011", -- t[28387] = 2
      "0000010" when "00110111011100100", -- t[28388] = 2
      "0000010" when "00110111011100101", -- t[28389] = 2
      "0000010" when "00110111011100110", -- t[28390] = 2
      "0000010" when "00110111011100111", -- t[28391] = 2
      "0000010" when "00110111011101000", -- t[28392] = 2
      "0000010" when "00110111011101001", -- t[28393] = 2
      "0000010" when "00110111011101010", -- t[28394] = 2
      "0000010" when "00110111011101011", -- t[28395] = 2
      "0000010" when "00110111011101100", -- t[28396] = 2
      "0000010" when "00110111011101101", -- t[28397] = 2
      "0000010" when "00110111011101110", -- t[28398] = 2
      "0000010" when "00110111011101111", -- t[28399] = 2
      "0000010" when "00110111011110000", -- t[28400] = 2
      "0000010" when "00110111011110001", -- t[28401] = 2
      "0000010" when "00110111011110010", -- t[28402] = 2
      "0000010" when "00110111011110011", -- t[28403] = 2
      "0000010" when "00110111011110100", -- t[28404] = 2
      "0000010" when "00110111011110101", -- t[28405] = 2
      "0000010" when "00110111011110110", -- t[28406] = 2
      "0000010" when "00110111011110111", -- t[28407] = 2
      "0000010" when "00110111011111000", -- t[28408] = 2
      "0000010" when "00110111011111001", -- t[28409] = 2
      "0000010" when "00110111011111010", -- t[28410] = 2
      "0000010" when "00110111011111011", -- t[28411] = 2
      "0000010" when "00110111011111100", -- t[28412] = 2
      "0000010" when "00110111011111101", -- t[28413] = 2
      "0000010" when "00110111011111110", -- t[28414] = 2
      "0000010" when "00110111011111111", -- t[28415] = 2
      "0000010" when "00110111100000000", -- t[28416] = 2
      "0000010" when "00110111100000001", -- t[28417] = 2
      "0000010" when "00110111100000010", -- t[28418] = 2
      "0000010" when "00110111100000011", -- t[28419] = 2
      "0000010" when "00110111100000100", -- t[28420] = 2
      "0000010" when "00110111100000101", -- t[28421] = 2
      "0000010" when "00110111100000110", -- t[28422] = 2
      "0000010" when "00110111100000111", -- t[28423] = 2
      "0000010" when "00110111100001000", -- t[28424] = 2
      "0000010" when "00110111100001001", -- t[28425] = 2
      "0000010" when "00110111100001010", -- t[28426] = 2
      "0000010" when "00110111100001011", -- t[28427] = 2
      "0000010" when "00110111100001100", -- t[28428] = 2
      "0000010" when "00110111100001101", -- t[28429] = 2
      "0000010" when "00110111100001110", -- t[28430] = 2
      "0000010" when "00110111100001111", -- t[28431] = 2
      "0000010" when "00110111100010000", -- t[28432] = 2
      "0000010" when "00110111100010001", -- t[28433] = 2
      "0000010" when "00110111100010010", -- t[28434] = 2
      "0000010" when "00110111100010011", -- t[28435] = 2
      "0000010" when "00110111100010100", -- t[28436] = 2
      "0000010" when "00110111100010101", -- t[28437] = 2
      "0000010" when "00110111100010110", -- t[28438] = 2
      "0000010" when "00110111100010111", -- t[28439] = 2
      "0000010" when "00110111100011000", -- t[28440] = 2
      "0000010" when "00110111100011001", -- t[28441] = 2
      "0000010" when "00110111100011010", -- t[28442] = 2
      "0000010" when "00110111100011011", -- t[28443] = 2
      "0000010" when "00110111100011100", -- t[28444] = 2
      "0000010" when "00110111100011101", -- t[28445] = 2
      "0000010" when "00110111100011110", -- t[28446] = 2
      "0000010" when "00110111100011111", -- t[28447] = 2
      "0000010" when "00110111100100000", -- t[28448] = 2
      "0000010" when "00110111100100001", -- t[28449] = 2
      "0000010" when "00110111100100010", -- t[28450] = 2
      "0000010" when "00110111100100011", -- t[28451] = 2
      "0000010" when "00110111100100100", -- t[28452] = 2
      "0000010" when "00110111100100101", -- t[28453] = 2
      "0000010" when "00110111100100110", -- t[28454] = 2
      "0000010" when "00110111100100111", -- t[28455] = 2
      "0000010" when "00110111100101000", -- t[28456] = 2
      "0000010" when "00110111100101001", -- t[28457] = 2
      "0000010" when "00110111100101010", -- t[28458] = 2
      "0000010" when "00110111100101011", -- t[28459] = 2
      "0000010" when "00110111100101100", -- t[28460] = 2
      "0000010" when "00110111100101101", -- t[28461] = 2
      "0000010" when "00110111100101110", -- t[28462] = 2
      "0000010" when "00110111100101111", -- t[28463] = 2
      "0000010" when "00110111100110000", -- t[28464] = 2
      "0000010" when "00110111100110001", -- t[28465] = 2
      "0000010" when "00110111100110010", -- t[28466] = 2
      "0000010" when "00110111100110011", -- t[28467] = 2
      "0000010" when "00110111100110100", -- t[28468] = 2
      "0000010" when "00110111100110101", -- t[28469] = 2
      "0000010" when "00110111100110110", -- t[28470] = 2
      "0000010" when "00110111100110111", -- t[28471] = 2
      "0000010" when "00110111100111000", -- t[28472] = 2
      "0000010" when "00110111100111001", -- t[28473] = 2
      "0000010" when "00110111100111010", -- t[28474] = 2
      "0000010" when "00110111100111011", -- t[28475] = 2
      "0000010" when "00110111100111100", -- t[28476] = 2
      "0000010" when "00110111100111101", -- t[28477] = 2
      "0000010" when "00110111100111110", -- t[28478] = 2
      "0000010" when "00110111100111111", -- t[28479] = 2
      "0000010" when "00110111101000000", -- t[28480] = 2
      "0000010" when "00110111101000001", -- t[28481] = 2
      "0000010" when "00110111101000010", -- t[28482] = 2
      "0000010" when "00110111101000011", -- t[28483] = 2
      "0000010" when "00110111101000100", -- t[28484] = 2
      "0000010" when "00110111101000101", -- t[28485] = 2
      "0000010" when "00110111101000110", -- t[28486] = 2
      "0000010" when "00110111101000111", -- t[28487] = 2
      "0000010" when "00110111101001000", -- t[28488] = 2
      "0000010" when "00110111101001001", -- t[28489] = 2
      "0000010" when "00110111101001010", -- t[28490] = 2
      "0000010" when "00110111101001011", -- t[28491] = 2
      "0000010" when "00110111101001100", -- t[28492] = 2
      "0000010" when "00110111101001101", -- t[28493] = 2
      "0000010" when "00110111101001110", -- t[28494] = 2
      "0000010" when "00110111101001111", -- t[28495] = 2
      "0000010" when "00110111101010000", -- t[28496] = 2
      "0000010" when "00110111101010001", -- t[28497] = 2
      "0000010" when "00110111101010010", -- t[28498] = 2
      "0000010" when "00110111101010011", -- t[28499] = 2
      "0000010" when "00110111101010100", -- t[28500] = 2
      "0000010" when "00110111101010101", -- t[28501] = 2
      "0000010" when "00110111101010110", -- t[28502] = 2
      "0000010" when "00110111101010111", -- t[28503] = 2
      "0000010" when "00110111101011000", -- t[28504] = 2
      "0000010" when "00110111101011001", -- t[28505] = 2
      "0000010" when "00110111101011010", -- t[28506] = 2
      "0000010" when "00110111101011011", -- t[28507] = 2
      "0000010" when "00110111101011100", -- t[28508] = 2
      "0000010" when "00110111101011101", -- t[28509] = 2
      "0000010" when "00110111101011110", -- t[28510] = 2
      "0000010" when "00110111101011111", -- t[28511] = 2
      "0000010" when "00110111101100000", -- t[28512] = 2
      "0000010" when "00110111101100001", -- t[28513] = 2
      "0000010" when "00110111101100010", -- t[28514] = 2
      "0000010" when "00110111101100011", -- t[28515] = 2
      "0000010" when "00110111101100100", -- t[28516] = 2
      "0000010" when "00110111101100101", -- t[28517] = 2
      "0000010" when "00110111101100110", -- t[28518] = 2
      "0000010" when "00110111101100111", -- t[28519] = 2
      "0000010" when "00110111101101000", -- t[28520] = 2
      "0000010" when "00110111101101001", -- t[28521] = 2
      "0000010" when "00110111101101010", -- t[28522] = 2
      "0000010" when "00110111101101011", -- t[28523] = 2
      "0000010" when "00110111101101100", -- t[28524] = 2
      "0000010" when "00110111101101101", -- t[28525] = 2
      "0000010" when "00110111101101110", -- t[28526] = 2
      "0000010" when "00110111101101111", -- t[28527] = 2
      "0000010" when "00110111101110000", -- t[28528] = 2
      "0000010" when "00110111101110001", -- t[28529] = 2
      "0000010" when "00110111101110010", -- t[28530] = 2
      "0000010" when "00110111101110011", -- t[28531] = 2
      "0000010" when "00110111101110100", -- t[28532] = 2
      "0000010" when "00110111101110101", -- t[28533] = 2
      "0000010" when "00110111101110110", -- t[28534] = 2
      "0000010" when "00110111101110111", -- t[28535] = 2
      "0000010" when "00110111101111000", -- t[28536] = 2
      "0000010" when "00110111101111001", -- t[28537] = 2
      "0000010" when "00110111101111010", -- t[28538] = 2
      "0000010" when "00110111101111011", -- t[28539] = 2
      "0000010" when "00110111101111100", -- t[28540] = 2
      "0000010" when "00110111101111101", -- t[28541] = 2
      "0000010" when "00110111101111110", -- t[28542] = 2
      "0000010" when "00110111101111111", -- t[28543] = 2
      "0000010" when "00110111110000000", -- t[28544] = 2
      "0000010" when "00110111110000001", -- t[28545] = 2
      "0000010" when "00110111110000010", -- t[28546] = 2
      "0000010" when "00110111110000011", -- t[28547] = 2
      "0000010" when "00110111110000100", -- t[28548] = 2
      "0000010" when "00110111110000101", -- t[28549] = 2
      "0000010" when "00110111110000110", -- t[28550] = 2
      "0000010" when "00110111110000111", -- t[28551] = 2
      "0000010" when "00110111110001000", -- t[28552] = 2
      "0000010" when "00110111110001001", -- t[28553] = 2
      "0000010" when "00110111110001010", -- t[28554] = 2
      "0000010" when "00110111110001011", -- t[28555] = 2
      "0000010" when "00110111110001100", -- t[28556] = 2
      "0000010" when "00110111110001101", -- t[28557] = 2
      "0000010" when "00110111110001110", -- t[28558] = 2
      "0000010" when "00110111110001111", -- t[28559] = 2
      "0000010" when "00110111110010000", -- t[28560] = 2
      "0000010" when "00110111110010001", -- t[28561] = 2
      "0000010" when "00110111110010010", -- t[28562] = 2
      "0000010" when "00110111110010011", -- t[28563] = 2
      "0000010" when "00110111110010100", -- t[28564] = 2
      "0000010" when "00110111110010101", -- t[28565] = 2
      "0000010" when "00110111110010110", -- t[28566] = 2
      "0000010" when "00110111110010111", -- t[28567] = 2
      "0000010" when "00110111110011000", -- t[28568] = 2
      "0000010" when "00110111110011001", -- t[28569] = 2
      "0000010" when "00110111110011010", -- t[28570] = 2
      "0000010" when "00110111110011011", -- t[28571] = 2
      "0000010" when "00110111110011100", -- t[28572] = 2
      "0000010" when "00110111110011101", -- t[28573] = 2
      "0000010" when "00110111110011110", -- t[28574] = 2
      "0000010" when "00110111110011111", -- t[28575] = 2
      "0000010" when "00110111110100000", -- t[28576] = 2
      "0000010" when "00110111110100001", -- t[28577] = 2
      "0000010" when "00110111110100010", -- t[28578] = 2
      "0000010" when "00110111110100011", -- t[28579] = 2
      "0000010" when "00110111110100100", -- t[28580] = 2
      "0000010" when "00110111110100101", -- t[28581] = 2
      "0000010" when "00110111110100110", -- t[28582] = 2
      "0000010" when "00110111110100111", -- t[28583] = 2
      "0000010" when "00110111110101000", -- t[28584] = 2
      "0000010" when "00110111110101001", -- t[28585] = 2
      "0000010" when "00110111110101010", -- t[28586] = 2
      "0000010" when "00110111110101011", -- t[28587] = 2
      "0000010" when "00110111110101100", -- t[28588] = 2
      "0000010" when "00110111110101101", -- t[28589] = 2
      "0000010" when "00110111110101110", -- t[28590] = 2
      "0000010" when "00110111110101111", -- t[28591] = 2
      "0000010" when "00110111110110000", -- t[28592] = 2
      "0000010" when "00110111110110001", -- t[28593] = 2
      "0000010" when "00110111110110010", -- t[28594] = 2
      "0000010" when "00110111110110011", -- t[28595] = 2
      "0000010" when "00110111110110100", -- t[28596] = 2
      "0000010" when "00110111110110101", -- t[28597] = 2
      "0000010" when "00110111110110110", -- t[28598] = 2
      "0000010" when "00110111110110111", -- t[28599] = 2
      "0000010" when "00110111110111000", -- t[28600] = 2
      "0000010" when "00110111110111001", -- t[28601] = 2
      "0000010" when "00110111110111010", -- t[28602] = 2
      "0000010" when "00110111110111011", -- t[28603] = 2
      "0000010" when "00110111110111100", -- t[28604] = 2
      "0000010" when "00110111110111101", -- t[28605] = 2
      "0000010" when "00110111110111110", -- t[28606] = 2
      "0000010" when "00110111110111111", -- t[28607] = 2
      "0000010" when "00110111111000000", -- t[28608] = 2
      "0000010" when "00110111111000001", -- t[28609] = 2
      "0000010" when "00110111111000010", -- t[28610] = 2
      "0000010" when "00110111111000011", -- t[28611] = 2
      "0000010" when "00110111111000100", -- t[28612] = 2
      "0000010" when "00110111111000101", -- t[28613] = 2
      "0000010" when "00110111111000110", -- t[28614] = 2
      "0000010" when "00110111111000111", -- t[28615] = 2
      "0000010" when "00110111111001000", -- t[28616] = 2
      "0000010" when "00110111111001001", -- t[28617] = 2
      "0000010" when "00110111111001010", -- t[28618] = 2
      "0000010" when "00110111111001011", -- t[28619] = 2
      "0000010" when "00110111111001100", -- t[28620] = 2
      "0000010" when "00110111111001101", -- t[28621] = 2
      "0000010" when "00110111111001110", -- t[28622] = 2
      "0000010" when "00110111111001111", -- t[28623] = 2
      "0000010" when "00110111111010000", -- t[28624] = 2
      "0000010" when "00110111111010001", -- t[28625] = 2
      "0000010" when "00110111111010010", -- t[28626] = 2
      "0000010" when "00110111111010011", -- t[28627] = 2
      "0000010" when "00110111111010100", -- t[28628] = 2
      "0000010" when "00110111111010101", -- t[28629] = 2
      "0000010" when "00110111111010110", -- t[28630] = 2
      "0000010" when "00110111111010111", -- t[28631] = 2
      "0000010" when "00110111111011000", -- t[28632] = 2
      "0000010" when "00110111111011001", -- t[28633] = 2
      "0000010" when "00110111111011010", -- t[28634] = 2
      "0000010" when "00110111111011011", -- t[28635] = 2
      "0000010" when "00110111111011100", -- t[28636] = 2
      "0000010" when "00110111111011101", -- t[28637] = 2
      "0000010" when "00110111111011110", -- t[28638] = 2
      "0000010" when "00110111111011111", -- t[28639] = 2
      "0000010" when "00110111111100000", -- t[28640] = 2
      "0000010" when "00110111111100001", -- t[28641] = 2
      "0000010" when "00110111111100010", -- t[28642] = 2
      "0000010" when "00110111111100011", -- t[28643] = 2
      "0000010" when "00110111111100100", -- t[28644] = 2
      "0000010" when "00110111111100101", -- t[28645] = 2
      "0000010" when "00110111111100110", -- t[28646] = 2
      "0000010" when "00110111111100111", -- t[28647] = 2
      "0000010" when "00110111111101000", -- t[28648] = 2
      "0000010" when "00110111111101001", -- t[28649] = 2
      "0000010" when "00110111111101010", -- t[28650] = 2
      "0000010" when "00110111111101011", -- t[28651] = 2
      "0000010" when "00110111111101100", -- t[28652] = 2
      "0000010" when "00110111111101101", -- t[28653] = 2
      "0000010" when "00110111111101110", -- t[28654] = 2
      "0000010" when "00110111111101111", -- t[28655] = 2
      "0000010" when "00110111111110000", -- t[28656] = 2
      "0000010" when "00110111111110001", -- t[28657] = 2
      "0000010" when "00110111111110010", -- t[28658] = 2
      "0000010" when "00110111111110011", -- t[28659] = 2
      "0000010" when "00110111111110100", -- t[28660] = 2
      "0000010" when "00110111111110101", -- t[28661] = 2
      "0000010" when "00110111111110110", -- t[28662] = 2
      "0000010" when "00110111111110111", -- t[28663] = 2
      "0000010" when "00110111111111000", -- t[28664] = 2
      "0000010" when "00110111111111001", -- t[28665] = 2
      "0000010" when "00110111111111010", -- t[28666] = 2
      "0000010" when "00110111111111011", -- t[28667] = 2
      "0000010" when "00110111111111100", -- t[28668] = 2
      "0000010" when "00110111111111101", -- t[28669] = 2
      "0000010" when "00110111111111110", -- t[28670] = 2
      "0000010" when "00110111111111111", -- t[28671] = 2
      "0000010" when "00111000000000000", -- t[28672] = 2
      "0000010" when "00111000000000001", -- t[28673] = 2
      "0000010" when "00111000000000010", -- t[28674] = 2
      "0000010" when "00111000000000011", -- t[28675] = 2
      "0000010" when "00111000000000100", -- t[28676] = 2
      "0000010" when "00111000000000101", -- t[28677] = 2
      "0000010" when "00111000000000110", -- t[28678] = 2
      "0000010" when "00111000000000111", -- t[28679] = 2
      "0000010" when "00111000000001000", -- t[28680] = 2
      "0000010" when "00111000000001001", -- t[28681] = 2
      "0000010" when "00111000000001010", -- t[28682] = 2
      "0000010" when "00111000000001011", -- t[28683] = 2
      "0000010" when "00111000000001100", -- t[28684] = 2
      "0000010" when "00111000000001101", -- t[28685] = 2
      "0000010" when "00111000000001110", -- t[28686] = 2
      "0000010" when "00111000000001111", -- t[28687] = 2
      "0000010" when "00111000000010000", -- t[28688] = 2
      "0000010" when "00111000000010001", -- t[28689] = 2
      "0000010" when "00111000000010010", -- t[28690] = 2
      "0000010" when "00111000000010011", -- t[28691] = 2
      "0000010" when "00111000000010100", -- t[28692] = 2
      "0000010" when "00111000000010101", -- t[28693] = 2
      "0000010" when "00111000000010110", -- t[28694] = 2
      "0000010" when "00111000000010111", -- t[28695] = 2
      "0000010" when "00111000000011000", -- t[28696] = 2
      "0000010" when "00111000000011001", -- t[28697] = 2
      "0000010" when "00111000000011010", -- t[28698] = 2
      "0000010" when "00111000000011011", -- t[28699] = 2
      "0000010" when "00111000000011100", -- t[28700] = 2
      "0000010" when "00111000000011101", -- t[28701] = 2
      "0000010" when "00111000000011110", -- t[28702] = 2
      "0000010" when "00111000000011111", -- t[28703] = 2
      "0000010" when "00111000000100000", -- t[28704] = 2
      "0000010" when "00111000000100001", -- t[28705] = 2
      "0000010" when "00111000000100010", -- t[28706] = 2
      "0000010" when "00111000000100011", -- t[28707] = 2
      "0000010" when "00111000000100100", -- t[28708] = 2
      "0000010" when "00111000000100101", -- t[28709] = 2
      "0000010" when "00111000000100110", -- t[28710] = 2
      "0000010" when "00111000000100111", -- t[28711] = 2
      "0000010" when "00111000000101000", -- t[28712] = 2
      "0000010" when "00111000000101001", -- t[28713] = 2
      "0000010" when "00111000000101010", -- t[28714] = 2
      "0000010" when "00111000000101011", -- t[28715] = 2
      "0000010" when "00111000000101100", -- t[28716] = 2
      "0000010" when "00111000000101101", -- t[28717] = 2
      "0000010" when "00111000000101110", -- t[28718] = 2
      "0000010" when "00111000000101111", -- t[28719] = 2
      "0000010" when "00111000000110000", -- t[28720] = 2
      "0000010" when "00111000000110001", -- t[28721] = 2
      "0000010" when "00111000000110010", -- t[28722] = 2
      "0000010" when "00111000000110011", -- t[28723] = 2
      "0000010" when "00111000000110100", -- t[28724] = 2
      "0000010" when "00111000000110101", -- t[28725] = 2
      "0000010" when "00111000000110110", -- t[28726] = 2
      "0000010" when "00111000000110111", -- t[28727] = 2
      "0000010" when "00111000000111000", -- t[28728] = 2
      "0000010" when "00111000000111001", -- t[28729] = 2
      "0000010" when "00111000000111010", -- t[28730] = 2
      "0000010" when "00111000000111011", -- t[28731] = 2
      "0000010" when "00111000000111100", -- t[28732] = 2
      "0000010" when "00111000000111101", -- t[28733] = 2
      "0000010" when "00111000000111110", -- t[28734] = 2
      "0000010" when "00111000000111111", -- t[28735] = 2
      "0000010" when "00111000001000000", -- t[28736] = 2
      "0000010" when "00111000001000001", -- t[28737] = 2
      "0000010" when "00111000001000010", -- t[28738] = 2
      "0000010" when "00111000001000011", -- t[28739] = 2
      "0000010" when "00111000001000100", -- t[28740] = 2
      "0000010" when "00111000001000101", -- t[28741] = 2
      "0000010" when "00111000001000110", -- t[28742] = 2
      "0000010" when "00111000001000111", -- t[28743] = 2
      "0000010" when "00111000001001000", -- t[28744] = 2
      "0000010" when "00111000001001001", -- t[28745] = 2
      "0000010" when "00111000001001010", -- t[28746] = 2
      "0000010" when "00111000001001011", -- t[28747] = 2
      "0000010" when "00111000001001100", -- t[28748] = 2
      "0000010" when "00111000001001101", -- t[28749] = 2
      "0000010" when "00111000001001110", -- t[28750] = 2
      "0000010" when "00111000001001111", -- t[28751] = 2
      "0000010" when "00111000001010000", -- t[28752] = 2
      "0000010" when "00111000001010001", -- t[28753] = 2
      "0000010" when "00111000001010010", -- t[28754] = 2
      "0000010" when "00111000001010011", -- t[28755] = 2
      "0000010" when "00111000001010100", -- t[28756] = 2
      "0000010" when "00111000001010101", -- t[28757] = 2
      "0000010" when "00111000001010110", -- t[28758] = 2
      "0000010" when "00111000001010111", -- t[28759] = 2
      "0000010" when "00111000001011000", -- t[28760] = 2
      "0000010" when "00111000001011001", -- t[28761] = 2
      "0000010" when "00111000001011010", -- t[28762] = 2
      "0000010" when "00111000001011011", -- t[28763] = 2
      "0000010" when "00111000001011100", -- t[28764] = 2
      "0000010" when "00111000001011101", -- t[28765] = 2
      "0000010" when "00111000001011110", -- t[28766] = 2
      "0000010" when "00111000001011111", -- t[28767] = 2
      "0000010" when "00111000001100000", -- t[28768] = 2
      "0000010" when "00111000001100001", -- t[28769] = 2
      "0000010" when "00111000001100010", -- t[28770] = 2
      "0000010" when "00111000001100011", -- t[28771] = 2
      "0000010" when "00111000001100100", -- t[28772] = 2
      "0000010" when "00111000001100101", -- t[28773] = 2
      "0000010" when "00111000001100110", -- t[28774] = 2
      "0000010" when "00111000001100111", -- t[28775] = 2
      "0000010" when "00111000001101000", -- t[28776] = 2
      "0000010" when "00111000001101001", -- t[28777] = 2
      "0000010" when "00111000001101010", -- t[28778] = 2
      "0000010" when "00111000001101011", -- t[28779] = 2
      "0000010" when "00111000001101100", -- t[28780] = 2
      "0000010" when "00111000001101101", -- t[28781] = 2
      "0000010" when "00111000001101110", -- t[28782] = 2
      "0000010" when "00111000001101111", -- t[28783] = 2
      "0000010" when "00111000001110000", -- t[28784] = 2
      "0000010" when "00111000001110001", -- t[28785] = 2
      "0000010" when "00111000001110010", -- t[28786] = 2
      "0000010" when "00111000001110011", -- t[28787] = 2
      "0000010" when "00111000001110100", -- t[28788] = 2
      "0000010" when "00111000001110101", -- t[28789] = 2
      "0000010" when "00111000001110110", -- t[28790] = 2
      "0000010" when "00111000001110111", -- t[28791] = 2
      "0000010" when "00111000001111000", -- t[28792] = 2
      "0000010" when "00111000001111001", -- t[28793] = 2
      "0000010" when "00111000001111010", -- t[28794] = 2
      "0000010" when "00111000001111011", -- t[28795] = 2
      "0000010" when "00111000001111100", -- t[28796] = 2
      "0000010" when "00111000001111101", -- t[28797] = 2
      "0000010" when "00111000001111110", -- t[28798] = 2
      "0000010" when "00111000001111111", -- t[28799] = 2
      "0000010" when "00111000010000000", -- t[28800] = 2
      "0000010" when "00111000010000001", -- t[28801] = 2
      "0000010" when "00111000010000010", -- t[28802] = 2
      "0000010" when "00111000010000011", -- t[28803] = 2
      "0000010" when "00111000010000100", -- t[28804] = 2
      "0000010" when "00111000010000101", -- t[28805] = 2
      "0000010" when "00111000010000110", -- t[28806] = 2
      "0000010" when "00111000010000111", -- t[28807] = 2
      "0000010" when "00111000010001000", -- t[28808] = 2
      "0000010" when "00111000010001001", -- t[28809] = 2
      "0000010" when "00111000010001010", -- t[28810] = 2
      "0000010" when "00111000010001011", -- t[28811] = 2
      "0000010" when "00111000010001100", -- t[28812] = 2
      "0000010" when "00111000010001101", -- t[28813] = 2
      "0000010" when "00111000010001110", -- t[28814] = 2
      "0000010" when "00111000010001111", -- t[28815] = 2
      "0000010" when "00111000010010000", -- t[28816] = 2
      "0000010" when "00111000010010001", -- t[28817] = 2
      "0000010" when "00111000010010010", -- t[28818] = 2
      "0000010" when "00111000010010011", -- t[28819] = 2
      "0000010" when "00111000010010100", -- t[28820] = 2
      "0000010" when "00111000010010101", -- t[28821] = 2
      "0000010" when "00111000010010110", -- t[28822] = 2
      "0000010" when "00111000010010111", -- t[28823] = 2
      "0000010" when "00111000010011000", -- t[28824] = 2
      "0000010" when "00111000010011001", -- t[28825] = 2
      "0000010" when "00111000010011010", -- t[28826] = 2
      "0000010" when "00111000010011011", -- t[28827] = 2
      "0000010" when "00111000010011100", -- t[28828] = 2
      "0000010" when "00111000010011101", -- t[28829] = 2
      "0000010" when "00111000010011110", -- t[28830] = 2
      "0000010" when "00111000010011111", -- t[28831] = 2
      "0000010" when "00111000010100000", -- t[28832] = 2
      "0000010" when "00111000010100001", -- t[28833] = 2
      "0000010" when "00111000010100010", -- t[28834] = 2
      "0000010" when "00111000010100011", -- t[28835] = 2
      "0000010" when "00111000010100100", -- t[28836] = 2
      "0000010" when "00111000010100101", -- t[28837] = 2
      "0000010" when "00111000010100110", -- t[28838] = 2
      "0000010" when "00111000010100111", -- t[28839] = 2
      "0000010" when "00111000010101000", -- t[28840] = 2
      "0000010" when "00111000010101001", -- t[28841] = 2
      "0000010" when "00111000010101010", -- t[28842] = 2
      "0000010" when "00111000010101011", -- t[28843] = 2
      "0000010" when "00111000010101100", -- t[28844] = 2
      "0000010" when "00111000010101101", -- t[28845] = 2
      "0000010" when "00111000010101110", -- t[28846] = 2
      "0000010" when "00111000010101111", -- t[28847] = 2
      "0000010" when "00111000010110000", -- t[28848] = 2
      "0000010" when "00111000010110001", -- t[28849] = 2
      "0000010" when "00111000010110010", -- t[28850] = 2
      "0000010" when "00111000010110011", -- t[28851] = 2
      "0000010" when "00111000010110100", -- t[28852] = 2
      "0000010" when "00111000010110101", -- t[28853] = 2
      "0000010" when "00111000010110110", -- t[28854] = 2
      "0000010" when "00111000010110111", -- t[28855] = 2
      "0000010" when "00111000010111000", -- t[28856] = 2
      "0000010" when "00111000010111001", -- t[28857] = 2
      "0000010" when "00111000010111010", -- t[28858] = 2
      "0000010" when "00111000010111011", -- t[28859] = 2
      "0000010" when "00111000010111100", -- t[28860] = 2
      "0000010" when "00111000010111101", -- t[28861] = 2
      "0000010" when "00111000010111110", -- t[28862] = 2
      "0000010" when "00111000010111111", -- t[28863] = 2
      "0000010" when "00111000011000000", -- t[28864] = 2
      "0000010" when "00111000011000001", -- t[28865] = 2
      "0000010" when "00111000011000010", -- t[28866] = 2
      "0000010" when "00111000011000011", -- t[28867] = 2
      "0000010" when "00111000011000100", -- t[28868] = 2
      "0000010" when "00111000011000101", -- t[28869] = 2
      "0000010" when "00111000011000110", -- t[28870] = 2
      "0000010" when "00111000011000111", -- t[28871] = 2
      "0000010" when "00111000011001000", -- t[28872] = 2
      "0000010" when "00111000011001001", -- t[28873] = 2
      "0000010" when "00111000011001010", -- t[28874] = 2
      "0000010" when "00111000011001011", -- t[28875] = 2
      "0000010" when "00111000011001100", -- t[28876] = 2
      "0000010" when "00111000011001101", -- t[28877] = 2
      "0000010" when "00111000011001110", -- t[28878] = 2
      "0000010" when "00111000011001111", -- t[28879] = 2
      "0000010" when "00111000011010000", -- t[28880] = 2
      "0000010" when "00111000011010001", -- t[28881] = 2
      "0000010" when "00111000011010010", -- t[28882] = 2
      "0000010" when "00111000011010011", -- t[28883] = 2
      "0000010" when "00111000011010100", -- t[28884] = 2
      "0000010" when "00111000011010101", -- t[28885] = 2
      "0000010" when "00111000011010110", -- t[28886] = 2
      "0000010" when "00111000011010111", -- t[28887] = 2
      "0000010" when "00111000011011000", -- t[28888] = 2
      "0000010" when "00111000011011001", -- t[28889] = 2
      "0000010" when "00111000011011010", -- t[28890] = 2
      "0000010" when "00111000011011011", -- t[28891] = 2
      "0000010" when "00111000011011100", -- t[28892] = 2
      "0000010" when "00111000011011101", -- t[28893] = 2
      "0000010" when "00111000011011110", -- t[28894] = 2
      "0000010" when "00111000011011111", -- t[28895] = 2
      "0000010" when "00111000011100000", -- t[28896] = 2
      "0000010" when "00111000011100001", -- t[28897] = 2
      "0000010" when "00111000011100010", -- t[28898] = 2
      "0000010" when "00111000011100011", -- t[28899] = 2
      "0000010" when "00111000011100100", -- t[28900] = 2
      "0000010" when "00111000011100101", -- t[28901] = 2
      "0000010" when "00111000011100110", -- t[28902] = 2
      "0000010" when "00111000011100111", -- t[28903] = 2
      "0000010" when "00111000011101000", -- t[28904] = 2
      "0000010" when "00111000011101001", -- t[28905] = 2
      "0000010" when "00111000011101010", -- t[28906] = 2
      "0000010" when "00111000011101011", -- t[28907] = 2
      "0000010" when "00111000011101100", -- t[28908] = 2
      "0000010" when "00111000011101101", -- t[28909] = 2
      "0000010" when "00111000011101110", -- t[28910] = 2
      "0000010" when "00111000011101111", -- t[28911] = 2
      "0000010" when "00111000011110000", -- t[28912] = 2
      "0000010" when "00111000011110001", -- t[28913] = 2
      "0000010" when "00111000011110010", -- t[28914] = 2
      "0000010" when "00111000011110011", -- t[28915] = 2
      "0000010" when "00111000011110100", -- t[28916] = 2
      "0000010" when "00111000011110101", -- t[28917] = 2
      "0000010" when "00111000011110110", -- t[28918] = 2
      "0000010" when "00111000011110111", -- t[28919] = 2
      "0000010" when "00111000011111000", -- t[28920] = 2
      "0000010" when "00111000011111001", -- t[28921] = 2
      "0000010" when "00111000011111010", -- t[28922] = 2
      "0000010" when "00111000011111011", -- t[28923] = 2
      "0000010" when "00111000011111100", -- t[28924] = 2
      "0000010" when "00111000011111101", -- t[28925] = 2
      "0000010" when "00111000011111110", -- t[28926] = 2
      "0000010" when "00111000011111111", -- t[28927] = 2
      "0000010" when "00111000100000000", -- t[28928] = 2
      "0000010" when "00111000100000001", -- t[28929] = 2
      "0000010" when "00111000100000010", -- t[28930] = 2
      "0000010" when "00111000100000011", -- t[28931] = 2
      "0000010" when "00111000100000100", -- t[28932] = 2
      "0000010" when "00111000100000101", -- t[28933] = 2
      "0000010" when "00111000100000110", -- t[28934] = 2
      "0000010" when "00111000100000111", -- t[28935] = 2
      "0000010" when "00111000100001000", -- t[28936] = 2
      "0000010" when "00111000100001001", -- t[28937] = 2
      "0000010" when "00111000100001010", -- t[28938] = 2
      "0000010" when "00111000100001011", -- t[28939] = 2
      "0000010" when "00111000100001100", -- t[28940] = 2
      "0000010" when "00111000100001101", -- t[28941] = 2
      "0000010" when "00111000100001110", -- t[28942] = 2
      "0000010" when "00111000100001111", -- t[28943] = 2
      "0000010" when "00111000100010000", -- t[28944] = 2
      "0000010" when "00111000100010001", -- t[28945] = 2
      "0000010" when "00111000100010010", -- t[28946] = 2
      "0000010" when "00111000100010011", -- t[28947] = 2
      "0000010" when "00111000100010100", -- t[28948] = 2
      "0000010" when "00111000100010101", -- t[28949] = 2
      "0000010" when "00111000100010110", -- t[28950] = 2
      "0000010" when "00111000100010111", -- t[28951] = 2
      "0000010" when "00111000100011000", -- t[28952] = 2
      "0000010" when "00111000100011001", -- t[28953] = 2
      "0000010" when "00111000100011010", -- t[28954] = 2
      "0000010" when "00111000100011011", -- t[28955] = 2
      "0000010" when "00111000100011100", -- t[28956] = 2
      "0000010" when "00111000100011101", -- t[28957] = 2
      "0000010" when "00111000100011110", -- t[28958] = 2
      "0000010" when "00111000100011111", -- t[28959] = 2
      "0000010" when "00111000100100000", -- t[28960] = 2
      "0000010" when "00111000100100001", -- t[28961] = 2
      "0000010" when "00111000100100010", -- t[28962] = 2
      "0000010" when "00111000100100011", -- t[28963] = 2
      "0000010" when "00111000100100100", -- t[28964] = 2
      "0000010" when "00111000100100101", -- t[28965] = 2
      "0000010" when "00111000100100110", -- t[28966] = 2
      "0000010" when "00111000100100111", -- t[28967] = 2
      "0000010" when "00111000100101000", -- t[28968] = 2
      "0000010" when "00111000100101001", -- t[28969] = 2
      "0000010" when "00111000100101010", -- t[28970] = 2
      "0000010" when "00111000100101011", -- t[28971] = 2
      "0000010" when "00111000100101100", -- t[28972] = 2
      "0000010" when "00111000100101101", -- t[28973] = 2
      "0000010" when "00111000100101110", -- t[28974] = 2
      "0000010" when "00111000100101111", -- t[28975] = 2
      "0000010" when "00111000100110000", -- t[28976] = 2
      "0000010" when "00111000100110001", -- t[28977] = 2
      "0000010" when "00111000100110010", -- t[28978] = 2
      "0000010" when "00111000100110011", -- t[28979] = 2
      "0000010" when "00111000100110100", -- t[28980] = 2
      "0000010" when "00111000100110101", -- t[28981] = 2
      "0000010" when "00111000100110110", -- t[28982] = 2
      "0000010" when "00111000100110111", -- t[28983] = 2
      "0000010" when "00111000100111000", -- t[28984] = 2
      "0000010" when "00111000100111001", -- t[28985] = 2
      "0000010" when "00111000100111010", -- t[28986] = 2
      "0000010" when "00111000100111011", -- t[28987] = 2
      "0000010" when "00111000100111100", -- t[28988] = 2
      "0000010" when "00111000100111101", -- t[28989] = 2
      "0000010" when "00111000100111110", -- t[28990] = 2
      "0000010" when "00111000100111111", -- t[28991] = 2
      "0000010" when "00111000101000000", -- t[28992] = 2
      "0000010" when "00111000101000001", -- t[28993] = 2
      "0000010" when "00111000101000010", -- t[28994] = 2
      "0000010" when "00111000101000011", -- t[28995] = 2
      "0000010" when "00111000101000100", -- t[28996] = 2
      "0000010" when "00111000101000101", -- t[28997] = 2
      "0000010" when "00111000101000110", -- t[28998] = 2
      "0000010" when "00111000101000111", -- t[28999] = 2
      "0000010" when "00111000101001000", -- t[29000] = 2
      "0000010" when "00111000101001001", -- t[29001] = 2
      "0000010" when "00111000101001010", -- t[29002] = 2
      "0000010" when "00111000101001011", -- t[29003] = 2
      "0000010" when "00111000101001100", -- t[29004] = 2
      "0000010" when "00111000101001101", -- t[29005] = 2
      "0000010" when "00111000101001110", -- t[29006] = 2
      "0000010" when "00111000101001111", -- t[29007] = 2
      "0000010" when "00111000101010000", -- t[29008] = 2
      "0000010" when "00111000101010001", -- t[29009] = 2
      "0000010" when "00111000101010010", -- t[29010] = 2
      "0000010" when "00111000101010011", -- t[29011] = 2
      "0000010" when "00111000101010100", -- t[29012] = 2
      "0000010" when "00111000101010101", -- t[29013] = 2
      "0000010" when "00111000101010110", -- t[29014] = 2
      "0000010" when "00111000101010111", -- t[29015] = 2
      "0000010" when "00111000101011000", -- t[29016] = 2
      "0000010" when "00111000101011001", -- t[29017] = 2
      "0000010" when "00111000101011010", -- t[29018] = 2
      "0000010" when "00111000101011011", -- t[29019] = 2
      "0000010" when "00111000101011100", -- t[29020] = 2
      "0000010" when "00111000101011101", -- t[29021] = 2
      "0000010" when "00111000101011110", -- t[29022] = 2
      "0000010" when "00111000101011111", -- t[29023] = 2
      "0000010" when "00111000101100000", -- t[29024] = 2
      "0000010" when "00111000101100001", -- t[29025] = 2
      "0000010" when "00111000101100010", -- t[29026] = 2
      "0000010" when "00111000101100011", -- t[29027] = 2
      "0000010" when "00111000101100100", -- t[29028] = 2
      "0000010" when "00111000101100101", -- t[29029] = 2
      "0000010" when "00111000101100110", -- t[29030] = 2
      "0000010" when "00111000101100111", -- t[29031] = 2
      "0000010" when "00111000101101000", -- t[29032] = 2
      "0000010" when "00111000101101001", -- t[29033] = 2
      "0000010" when "00111000101101010", -- t[29034] = 2
      "0000010" when "00111000101101011", -- t[29035] = 2
      "0000010" when "00111000101101100", -- t[29036] = 2
      "0000010" when "00111000101101101", -- t[29037] = 2
      "0000010" when "00111000101101110", -- t[29038] = 2
      "0000010" when "00111000101101111", -- t[29039] = 2
      "0000010" when "00111000101110000", -- t[29040] = 2
      "0000010" when "00111000101110001", -- t[29041] = 2
      "0000010" when "00111000101110010", -- t[29042] = 2
      "0000010" when "00111000101110011", -- t[29043] = 2
      "0000010" when "00111000101110100", -- t[29044] = 2
      "0000010" when "00111000101110101", -- t[29045] = 2
      "0000010" when "00111000101110110", -- t[29046] = 2
      "0000010" when "00111000101110111", -- t[29047] = 2
      "0000010" when "00111000101111000", -- t[29048] = 2
      "0000010" when "00111000101111001", -- t[29049] = 2
      "0000010" when "00111000101111010", -- t[29050] = 2
      "0000010" when "00111000101111011", -- t[29051] = 2
      "0000010" when "00111000101111100", -- t[29052] = 2
      "0000010" when "00111000101111101", -- t[29053] = 2
      "0000010" when "00111000101111110", -- t[29054] = 2
      "0000010" when "00111000101111111", -- t[29055] = 2
      "0000010" when "00111000110000000", -- t[29056] = 2
      "0000010" when "00111000110000001", -- t[29057] = 2
      "0000010" when "00111000110000010", -- t[29058] = 2
      "0000010" when "00111000110000011", -- t[29059] = 2
      "0000010" when "00111000110000100", -- t[29060] = 2
      "0000010" when "00111000110000101", -- t[29061] = 2
      "0000010" when "00111000110000110", -- t[29062] = 2
      "0000010" when "00111000110000111", -- t[29063] = 2
      "0000010" when "00111000110001000", -- t[29064] = 2
      "0000010" when "00111000110001001", -- t[29065] = 2
      "0000010" when "00111000110001010", -- t[29066] = 2
      "0000010" when "00111000110001011", -- t[29067] = 2
      "0000010" when "00111000110001100", -- t[29068] = 2
      "0000010" when "00111000110001101", -- t[29069] = 2
      "0000010" when "00111000110001110", -- t[29070] = 2
      "0000010" when "00111000110001111", -- t[29071] = 2
      "0000010" when "00111000110010000", -- t[29072] = 2
      "0000010" when "00111000110010001", -- t[29073] = 2
      "0000010" when "00111000110010010", -- t[29074] = 2
      "0000010" when "00111000110010011", -- t[29075] = 2
      "0000010" when "00111000110010100", -- t[29076] = 2
      "0000010" when "00111000110010101", -- t[29077] = 2
      "0000010" when "00111000110010110", -- t[29078] = 2
      "0000010" when "00111000110010111", -- t[29079] = 2
      "0000010" when "00111000110011000", -- t[29080] = 2
      "0000010" when "00111000110011001", -- t[29081] = 2
      "0000010" when "00111000110011010", -- t[29082] = 2
      "0000010" when "00111000110011011", -- t[29083] = 2
      "0000010" when "00111000110011100", -- t[29084] = 2
      "0000010" when "00111000110011101", -- t[29085] = 2
      "0000010" when "00111000110011110", -- t[29086] = 2
      "0000010" when "00111000110011111", -- t[29087] = 2
      "0000010" when "00111000110100000", -- t[29088] = 2
      "0000010" when "00111000110100001", -- t[29089] = 2
      "0000010" when "00111000110100010", -- t[29090] = 2
      "0000010" when "00111000110100011", -- t[29091] = 2
      "0000010" when "00111000110100100", -- t[29092] = 2
      "0000010" when "00111000110100101", -- t[29093] = 2
      "0000010" when "00111000110100110", -- t[29094] = 2
      "0000010" when "00111000110100111", -- t[29095] = 2
      "0000010" when "00111000110101000", -- t[29096] = 2
      "0000010" when "00111000110101001", -- t[29097] = 2
      "0000010" when "00111000110101010", -- t[29098] = 2
      "0000010" when "00111000110101011", -- t[29099] = 2
      "0000010" when "00111000110101100", -- t[29100] = 2
      "0000010" when "00111000110101101", -- t[29101] = 2
      "0000010" when "00111000110101110", -- t[29102] = 2
      "0000010" when "00111000110101111", -- t[29103] = 2
      "0000010" when "00111000110110000", -- t[29104] = 2
      "0000010" when "00111000110110001", -- t[29105] = 2
      "0000010" when "00111000110110010", -- t[29106] = 2
      "0000010" when "00111000110110011", -- t[29107] = 2
      "0000010" when "00111000110110100", -- t[29108] = 2
      "0000010" when "00111000110110101", -- t[29109] = 2
      "0000010" when "00111000110110110", -- t[29110] = 2
      "0000010" when "00111000110110111", -- t[29111] = 2
      "0000010" when "00111000110111000", -- t[29112] = 2
      "0000010" when "00111000110111001", -- t[29113] = 2
      "0000010" when "00111000110111010", -- t[29114] = 2
      "0000010" when "00111000110111011", -- t[29115] = 2
      "0000010" when "00111000110111100", -- t[29116] = 2
      "0000010" when "00111000110111101", -- t[29117] = 2
      "0000010" when "00111000110111110", -- t[29118] = 2
      "0000010" when "00111000110111111", -- t[29119] = 2
      "0000010" when "00111000111000000", -- t[29120] = 2
      "0000010" when "00111000111000001", -- t[29121] = 2
      "0000010" when "00111000111000010", -- t[29122] = 2
      "0000010" when "00111000111000011", -- t[29123] = 2
      "0000010" when "00111000111000100", -- t[29124] = 2
      "0000010" when "00111000111000101", -- t[29125] = 2
      "0000010" when "00111000111000110", -- t[29126] = 2
      "0000010" when "00111000111000111", -- t[29127] = 2
      "0000010" when "00111000111001000", -- t[29128] = 2
      "0000010" when "00111000111001001", -- t[29129] = 2
      "0000010" when "00111000111001010", -- t[29130] = 2
      "0000010" when "00111000111001011", -- t[29131] = 2
      "0000010" when "00111000111001100", -- t[29132] = 2
      "0000010" when "00111000111001101", -- t[29133] = 2
      "0000010" when "00111000111001110", -- t[29134] = 2
      "0000010" when "00111000111001111", -- t[29135] = 2
      "0000010" when "00111000111010000", -- t[29136] = 2
      "0000010" when "00111000111010001", -- t[29137] = 2
      "0000010" when "00111000111010010", -- t[29138] = 2
      "0000010" when "00111000111010011", -- t[29139] = 2
      "0000010" when "00111000111010100", -- t[29140] = 2
      "0000010" when "00111000111010101", -- t[29141] = 2
      "0000010" when "00111000111010110", -- t[29142] = 2
      "0000010" when "00111000111010111", -- t[29143] = 2
      "0000010" when "00111000111011000", -- t[29144] = 2
      "0000010" when "00111000111011001", -- t[29145] = 2
      "0000010" when "00111000111011010", -- t[29146] = 2
      "0000010" when "00111000111011011", -- t[29147] = 2
      "0000010" when "00111000111011100", -- t[29148] = 2
      "0000010" when "00111000111011101", -- t[29149] = 2
      "0000010" when "00111000111011110", -- t[29150] = 2
      "0000010" when "00111000111011111", -- t[29151] = 2
      "0000010" when "00111000111100000", -- t[29152] = 2
      "0000010" when "00111000111100001", -- t[29153] = 2
      "0000010" when "00111000111100010", -- t[29154] = 2
      "0000010" when "00111000111100011", -- t[29155] = 2
      "0000010" when "00111000111100100", -- t[29156] = 2
      "0000010" when "00111000111100101", -- t[29157] = 2
      "0000010" when "00111000111100110", -- t[29158] = 2
      "0000010" when "00111000111100111", -- t[29159] = 2
      "0000010" when "00111000111101000", -- t[29160] = 2
      "0000010" when "00111000111101001", -- t[29161] = 2
      "0000010" when "00111000111101010", -- t[29162] = 2
      "0000010" when "00111000111101011", -- t[29163] = 2
      "0000010" when "00111000111101100", -- t[29164] = 2
      "0000010" when "00111000111101101", -- t[29165] = 2
      "0000010" when "00111000111101110", -- t[29166] = 2
      "0000010" when "00111000111101111", -- t[29167] = 2
      "0000010" when "00111000111110000", -- t[29168] = 2
      "0000010" when "00111000111110001", -- t[29169] = 2
      "0000010" when "00111000111110010", -- t[29170] = 2
      "0000010" when "00111000111110011", -- t[29171] = 2
      "0000010" when "00111000111110100", -- t[29172] = 2
      "0000010" when "00111000111110101", -- t[29173] = 2
      "0000010" when "00111000111110110", -- t[29174] = 2
      "0000010" when "00111000111110111", -- t[29175] = 2
      "0000010" when "00111000111111000", -- t[29176] = 2
      "0000010" when "00111000111111001", -- t[29177] = 2
      "0000010" when "00111000111111010", -- t[29178] = 2
      "0000010" when "00111000111111011", -- t[29179] = 2
      "0000010" when "00111000111111100", -- t[29180] = 2
      "0000010" when "00111000111111101", -- t[29181] = 2
      "0000010" when "00111000111111110", -- t[29182] = 2
      "0000010" when "00111000111111111", -- t[29183] = 2
      "0000010" when "00111001000000000", -- t[29184] = 2
      "0000010" when "00111001000000001", -- t[29185] = 2
      "0000010" when "00111001000000010", -- t[29186] = 2
      "0000010" when "00111001000000011", -- t[29187] = 2
      "0000010" when "00111001000000100", -- t[29188] = 2
      "0000010" when "00111001000000101", -- t[29189] = 2
      "0000010" when "00111001000000110", -- t[29190] = 2
      "0000010" when "00111001000000111", -- t[29191] = 2
      "0000010" when "00111001000001000", -- t[29192] = 2
      "0000010" when "00111001000001001", -- t[29193] = 2
      "0000010" when "00111001000001010", -- t[29194] = 2
      "0000010" when "00111001000001011", -- t[29195] = 2
      "0000010" when "00111001000001100", -- t[29196] = 2
      "0000010" when "00111001000001101", -- t[29197] = 2
      "0000010" when "00111001000001110", -- t[29198] = 2
      "0000010" when "00111001000001111", -- t[29199] = 2
      "0000010" when "00111001000010000", -- t[29200] = 2
      "0000010" when "00111001000010001", -- t[29201] = 2
      "0000010" when "00111001000010010", -- t[29202] = 2
      "0000010" when "00111001000010011", -- t[29203] = 2
      "0000010" when "00111001000010100", -- t[29204] = 2
      "0000010" when "00111001000010101", -- t[29205] = 2
      "0000010" when "00111001000010110", -- t[29206] = 2
      "0000010" when "00111001000010111", -- t[29207] = 2
      "0000010" when "00111001000011000", -- t[29208] = 2
      "0000010" when "00111001000011001", -- t[29209] = 2
      "0000010" when "00111001000011010", -- t[29210] = 2
      "0000010" when "00111001000011011", -- t[29211] = 2
      "0000010" when "00111001000011100", -- t[29212] = 2
      "0000010" when "00111001000011101", -- t[29213] = 2
      "0000010" when "00111001000011110", -- t[29214] = 2
      "0000010" when "00111001000011111", -- t[29215] = 2
      "0000010" when "00111001000100000", -- t[29216] = 2
      "0000010" when "00111001000100001", -- t[29217] = 2
      "0000010" when "00111001000100010", -- t[29218] = 2
      "0000010" when "00111001000100011", -- t[29219] = 2
      "0000010" when "00111001000100100", -- t[29220] = 2
      "0000010" when "00111001000100101", -- t[29221] = 2
      "0000010" when "00111001000100110", -- t[29222] = 2
      "0000010" when "00111001000100111", -- t[29223] = 2
      "0000010" when "00111001000101000", -- t[29224] = 2
      "0000010" when "00111001000101001", -- t[29225] = 2
      "0000010" when "00111001000101010", -- t[29226] = 2
      "0000010" when "00111001000101011", -- t[29227] = 2
      "0000010" when "00111001000101100", -- t[29228] = 2
      "0000010" when "00111001000101101", -- t[29229] = 2
      "0000010" when "00111001000101110", -- t[29230] = 2
      "0000010" when "00111001000101111", -- t[29231] = 2
      "0000010" when "00111001000110000", -- t[29232] = 2
      "0000010" when "00111001000110001", -- t[29233] = 2
      "0000010" when "00111001000110010", -- t[29234] = 2
      "0000010" when "00111001000110011", -- t[29235] = 2
      "0000010" when "00111001000110100", -- t[29236] = 2
      "0000010" when "00111001000110101", -- t[29237] = 2
      "0000010" when "00111001000110110", -- t[29238] = 2
      "0000010" when "00111001000110111", -- t[29239] = 2
      "0000010" when "00111001000111000", -- t[29240] = 2
      "0000010" when "00111001000111001", -- t[29241] = 2
      "0000010" when "00111001000111010", -- t[29242] = 2
      "0000010" when "00111001000111011", -- t[29243] = 2
      "0000010" when "00111001000111100", -- t[29244] = 2
      "0000010" when "00111001000111101", -- t[29245] = 2
      "0000010" when "00111001000111110", -- t[29246] = 2
      "0000010" when "00111001000111111", -- t[29247] = 2
      "0000010" when "00111001001000000", -- t[29248] = 2
      "0000010" when "00111001001000001", -- t[29249] = 2
      "0000010" when "00111001001000010", -- t[29250] = 2
      "0000010" when "00111001001000011", -- t[29251] = 2
      "0000010" when "00111001001000100", -- t[29252] = 2
      "0000010" when "00111001001000101", -- t[29253] = 2
      "0000010" when "00111001001000110", -- t[29254] = 2
      "0000010" when "00111001001000111", -- t[29255] = 2
      "0000010" when "00111001001001000", -- t[29256] = 2
      "0000010" when "00111001001001001", -- t[29257] = 2
      "0000010" when "00111001001001010", -- t[29258] = 2
      "0000010" when "00111001001001011", -- t[29259] = 2
      "0000010" when "00111001001001100", -- t[29260] = 2
      "0000010" when "00111001001001101", -- t[29261] = 2
      "0000010" when "00111001001001110", -- t[29262] = 2
      "0000010" when "00111001001001111", -- t[29263] = 2
      "0000010" when "00111001001010000", -- t[29264] = 2
      "0000010" when "00111001001010001", -- t[29265] = 2
      "0000010" when "00111001001010010", -- t[29266] = 2
      "0000010" when "00111001001010011", -- t[29267] = 2
      "0000010" when "00111001001010100", -- t[29268] = 2
      "0000010" when "00111001001010101", -- t[29269] = 2
      "0000010" when "00111001001010110", -- t[29270] = 2
      "0000010" when "00111001001010111", -- t[29271] = 2
      "0000010" when "00111001001011000", -- t[29272] = 2
      "0000010" when "00111001001011001", -- t[29273] = 2
      "0000010" when "00111001001011010", -- t[29274] = 2
      "0000010" when "00111001001011011", -- t[29275] = 2
      "0000010" when "00111001001011100", -- t[29276] = 2
      "0000010" when "00111001001011101", -- t[29277] = 2
      "0000010" when "00111001001011110", -- t[29278] = 2
      "0000010" when "00111001001011111", -- t[29279] = 2
      "0000010" when "00111001001100000", -- t[29280] = 2
      "0000010" when "00111001001100001", -- t[29281] = 2
      "0000010" when "00111001001100010", -- t[29282] = 2
      "0000010" when "00111001001100011", -- t[29283] = 2
      "0000010" when "00111001001100100", -- t[29284] = 2
      "0000010" when "00111001001100101", -- t[29285] = 2
      "0000010" when "00111001001100110", -- t[29286] = 2
      "0000010" when "00111001001100111", -- t[29287] = 2
      "0000010" when "00111001001101000", -- t[29288] = 2
      "0000010" when "00111001001101001", -- t[29289] = 2
      "0000010" when "00111001001101010", -- t[29290] = 2
      "0000010" when "00111001001101011", -- t[29291] = 2
      "0000010" when "00111001001101100", -- t[29292] = 2
      "0000010" when "00111001001101101", -- t[29293] = 2
      "0000010" when "00111001001101110", -- t[29294] = 2
      "0000010" when "00111001001101111", -- t[29295] = 2
      "0000010" when "00111001001110000", -- t[29296] = 2
      "0000010" when "00111001001110001", -- t[29297] = 2
      "0000010" when "00111001001110010", -- t[29298] = 2
      "0000010" when "00111001001110011", -- t[29299] = 2
      "0000010" when "00111001001110100", -- t[29300] = 2
      "0000010" when "00111001001110101", -- t[29301] = 2
      "0000010" when "00111001001110110", -- t[29302] = 2
      "0000010" when "00111001001110111", -- t[29303] = 2
      "0000010" when "00111001001111000", -- t[29304] = 2
      "0000010" when "00111001001111001", -- t[29305] = 2
      "0000010" when "00111001001111010", -- t[29306] = 2
      "0000010" when "00111001001111011", -- t[29307] = 2
      "0000010" when "00111001001111100", -- t[29308] = 2
      "0000010" when "00111001001111101", -- t[29309] = 2
      "0000010" when "00111001001111110", -- t[29310] = 2
      "0000010" when "00111001001111111", -- t[29311] = 2
      "0000010" when "00111001010000000", -- t[29312] = 2
      "0000010" when "00111001010000001", -- t[29313] = 2
      "0000010" when "00111001010000010", -- t[29314] = 2
      "0000010" when "00111001010000011", -- t[29315] = 2
      "0000010" when "00111001010000100", -- t[29316] = 2
      "0000010" when "00111001010000101", -- t[29317] = 2
      "0000010" when "00111001010000110", -- t[29318] = 2
      "0000010" when "00111001010000111", -- t[29319] = 2
      "0000010" when "00111001010001000", -- t[29320] = 2
      "0000010" when "00111001010001001", -- t[29321] = 2
      "0000010" when "00111001010001010", -- t[29322] = 2
      "0000010" when "00111001010001011", -- t[29323] = 2
      "0000010" when "00111001010001100", -- t[29324] = 2
      "0000010" when "00111001010001101", -- t[29325] = 2
      "0000010" when "00111001010001110", -- t[29326] = 2
      "0000010" when "00111001010001111", -- t[29327] = 2
      "0000010" when "00111001010010000", -- t[29328] = 2
      "0000010" when "00111001010010001", -- t[29329] = 2
      "0000010" when "00111001010010010", -- t[29330] = 2
      "0000010" when "00111001010010011", -- t[29331] = 2
      "0000010" when "00111001010010100", -- t[29332] = 2
      "0000010" when "00111001010010101", -- t[29333] = 2
      "0000010" when "00111001010010110", -- t[29334] = 2
      "0000010" when "00111001010010111", -- t[29335] = 2
      "0000010" when "00111001010011000", -- t[29336] = 2
      "0000010" when "00111001010011001", -- t[29337] = 2
      "0000010" when "00111001010011010", -- t[29338] = 2
      "0000010" when "00111001010011011", -- t[29339] = 2
      "0000010" when "00111001010011100", -- t[29340] = 2
      "0000010" when "00111001010011101", -- t[29341] = 2
      "0000010" when "00111001010011110", -- t[29342] = 2
      "0000010" when "00111001010011111", -- t[29343] = 2
      "0000010" when "00111001010100000", -- t[29344] = 2
      "0000010" when "00111001010100001", -- t[29345] = 2
      "0000010" when "00111001010100010", -- t[29346] = 2
      "0000010" when "00111001010100011", -- t[29347] = 2
      "0000010" when "00111001010100100", -- t[29348] = 2
      "0000010" when "00111001010100101", -- t[29349] = 2
      "0000010" when "00111001010100110", -- t[29350] = 2
      "0000010" when "00111001010100111", -- t[29351] = 2
      "0000010" when "00111001010101000", -- t[29352] = 2
      "0000010" when "00111001010101001", -- t[29353] = 2
      "0000010" when "00111001010101010", -- t[29354] = 2
      "0000010" when "00111001010101011", -- t[29355] = 2
      "0000010" when "00111001010101100", -- t[29356] = 2
      "0000010" when "00111001010101101", -- t[29357] = 2
      "0000010" when "00111001010101110", -- t[29358] = 2
      "0000010" when "00111001010101111", -- t[29359] = 2
      "0000010" when "00111001010110000", -- t[29360] = 2
      "0000010" when "00111001010110001", -- t[29361] = 2
      "0000010" when "00111001010110010", -- t[29362] = 2
      "0000010" when "00111001010110011", -- t[29363] = 2
      "0000010" when "00111001010110100", -- t[29364] = 2
      "0000010" when "00111001010110101", -- t[29365] = 2
      "0000010" when "00111001010110110", -- t[29366] = 2
      "0000010" when "00111001010110111", -- t[29367] = 2
      "0000010" when "00111001010111000", -- t[29368] = 2
      "0000010" when "00111001010111001", -- t[29369] = 2
      "0000010" when "00111001010111010", -- t[29370] = 2
      "0000010" when "00111001010111011", -- t[29371] = 2
      "0000010" when "00111001010111100", -- t[29372] = 2
      "0000010" when "00111001010111101", -- t[29373] = 2
      "0000010" when "00111001010111110", -- t[29374] = 2
      "0000010" when "00111001010111111", -- t[29375] = 2
      "0000010" when "00111001011000000", -- t[29376] = 2
      "0000010" when "00111001011000001", -- t[29377] = 2
      "0000010" when "00111001011000010", -- t[29378] = 2
      "0000010" when "00111001011000011", -- t[29379] = 2
      "0000010" when "00111001011000100", -- t[29380] = 2
      "0000010" when "00111001011000101", -- t[29381] = 2
      "0000010" when "00111001011000110", -- t[29382] = 2
      "0000010" when "00111001011000111", -- t[29383] = 2
      "0000010" when "00111001011001000", -- t[29384] = 2
      "0000010" when "00111001011001001", -- t[29385] = 2
      "0000010" when "00111001011001010", -- t[29386] = 2
      "0000010" when "00111001011001011", -- t[29387] = 2
      "0000010" when "00111001011001100", -- t[29388] = 2
      "0000010" when "00111001011001101", -- t[29389] = 2
      "0000010" when "00111001011001110", -- t[29390] = 2
      "0000010" when "00111001011001111", -- t[29391] = 2
      "0000010" when "00111001011010000", -- t[29392] = 2
      "0000010" when "00111001011010001", -- t[29393] = 2
      "0000010" when "00111001011010010", -- t[29394] = 2
      "0000010" when "00111001011010011", -- t[29395] = 2
      "0000010" when "00111001011010100", -- t[29396] = 2
      "0000010" when "00111001011010101", -- t[29397] = 2
      "0000010" when "00111001011010110", -- t[29398] = 2
      "0000010" when "00111001011010111", -- t[29399] = 2
      "0000010" when "00111001011011000", -- t[29400] = 2
      "0000010" when "00111001011011001", -- t[29401] = 2
      "0000010" when "00111001011011010", -- t[29402] = 2
      "0000010" when "00111001011011011", -- t[29403] = 2
      "0000010" when "00111001011011100", -- t[29404] = 2
      "0000010" when "00111001011011101", -- t[29405] = 2
      "0000010" when "00111001011011110", -- t[29406] = 2
      "0000010" when "00111001011011111", -- t[29407] = 2
      "0000010" when "00111001011100000", -- t[29408] = 2
      "0000010" when "00111001011100001", -- t[29409] = 2
      "0000010" when "00111001011100010", -- t[29410] = 2
      "0000010" when "00111001011100011", -- t[29411] = 2
      "0000010" when "00111001011100100", -- t[29412] = 2
      "0000010" when "00111001011100101", -- t[29413] = 2
      "0000010" when "00111001011100110", -- t[29414] = 2
      "0000010" when "00111001011100111", -- t[29415] = 2
      "0000010" when "00111001011101000", -- t[29416] = 2
      "0000010" when "00111001011101001", -- t[29417] = 2
      "0000010" when "00111001011101010", -- t[29418] = 2
      "0000010" when "00111001011101011", -- t[29419] = 2
      "0000010" when "00111001011101100", -- t[29420] = 2
      "0000010" when "00111001011101101", -- t[29421] = 2
      "0000010" when "00111001011101110", -- t[29422] = 2
      "0000010" when "00111001011101111", -- t[29423] = 2
      "0000010" when "00111001011110000", -- t[29424] = 2
      "0000010" when "00111001011110001", -- t[29425] = 2
      "0000010" when "00111001011110010", -- t[29426] = 2
      "0000010" when "00111001011110011", -- t[29427] = 2
      "0000010" when "00111001011110100", -- t[29428] = 2
      "0000010" when "00111001011110101", -- t[29429] = 2
      "0000010" when "00111001011110110", -- t[29430] = 2
      "0000010" when "00111001011110111", -- t[29431] = 2
      "0000010" when "00111001011111000", -- t[29432] = 2
      "0000010" when "00111001011111001", -- t[29433] = 2
      "0000010" when "00111001011111010", -- t[29434] = 2
      "0000010" when "00111001011111011", -- t[29435] = 2
      "0000010" when "00111001011111100", -- t[29436] = 2
      "0000010" when "00111001011111101", -- t[29437] = 2
      "0000010" when "00111001011111110", -- t[29438] = 2
      "0000010" when "00111001011111111", -- t[29439] = 2
      "0000010" when "00111001100000000", -- t[29440] = 2
      "0000010" when "00111001100000001", -- t[29441] = 2
      "0000010" when "00111001100000010", -- t[29442] = 2
      "0000010" when "00111001100000011", -- t[29443] = 2
      "0000010" when "00111001100000100", -- t[29444] = 2
      "0000010" when "00111001100000101", -- t[29445] = 2
      "0000010" when "00111001100000110", -- t[29446] = 2
      "0000010" when "00111001100000111", -- t[29447] = 2
      "0000010" when "00111001100001000", -- t[29448] = 2
      "0000010" when "00111001100001001", -- t[29449] = 2
      "0000010" when "00111001100001010", -- t[29450] = 2
      "0000010" when "00111001100001011", -- t[29451] = 2
      "0000010" when "00111001100001100", -- t[29452] = 2
      "0000010" when "00111001100001101", -- t[29453] = 2
      "0000010" when "00111001100001110", -- t[29454] = 2
      "0000010" when "00111001100001111", -- t[29455] = 2
      "0000010" when "00111001100010000", -- t[29456] = 2
      "0000010" when "00111001100010001", -- t[29457] = 2
      "0000010" when "00111001100010010", -- t[29458] = 2
      "0000010" when "00111001100010011", -- t[29459] = 2
      "0000010" when "00111001100010100", -- t[29460] = 2
      "0000010" when "00111001100010101", -- t[29461] = 2
      "0000010" when "00111001100010110", -- t[29462] = 2
      "0000010" when "00111001100010111", -- t[29463] = 2
      "0000010" when "00111001100011000", -- t[29464] = 2
      "0000010" when "00111001100011001", -- t[29465] = 2
      "0000010" when "00111001100011010", -- t[29466] = 2
      "0000010" when "00111001100011011", -- t[29467] = 2
      "0000010" when "00111001100011100", -- t[29468] = 2
      "0000010" when "00111001100011101", -- t[29469] = 2
      "0000010" when "00111001100011110", -- t[29470] = 2
      "0000010" when "00111001100011111", -- t[29471] = 2
      "0000010" when "00111001100100000", -- t[29472] = 2
      "0000010" when "00111001100100001", -- t[29473] = 2
      "0000010" when "00111001100100010", -- t[29474] = 2
      "0000010" when "00111001100100011", -- t[29475] = 2
      "0000010" when "00111001100100100", -- t[29476] = 2
      "0000010" when "00111001100100101", -- t[29477] = 2
      "0000010" when "00111001100100110", -- t[29478] = 2
      "0000010" when "00111001100100111", -- t[29479] = 2
      "0000010" when "00111001100101000", -- t[29480] = 2
      "0000010" when "00111001100101001", -- t[29481] = 2
      "0000010" when "00111001100101010", -- t[29482] = 2
      "0000010" when "00111001100101011", -- t[29483] = 2
      "0000010" when "00111001100101100", -- t[29484] = 2
      "0000010" when "00111001100101101", -- t[29485] = 2
      "0000010" when "00111001100101110", -- t[29486] = 2
      "0000010" when "00111001100101111", -- t[29487] = 2
      "0000010" when "00111001100110000", -- t[29488] = 2
      "0000010" when "00111001100110001", -- t[29489] = 2
      "0000010" when "00111001100110010", -- t[29490] = 2
      "0000010" when "00111001100110011", -- t[29491] = 2
      "0000010" when "00111001100110100", -- t[29492] = 2
      "0000010" when "00111001100110101", -- t[29493] = 2
      "0000010" when "00111001100110110", -- t[29494] = 2
      "0000010" when "00111001100110111", -- t[29495] = 2
      "0000010" when "00111001100111000", -- t[29496] = 2
      "0000010" when "00111001100111001", -- t[29497] = 2
      "0000010" when "00111001100111010", -- t[29498] = 2
      "0000010" when "00111001100111011", -- t[29499] = 2
      "0000010" when "00111001100111100", -- t[29500] = 2
      "0000010" when "00111001100111101", -- t[29501] = 2
      "0000010" when "00111001100111110", -- t[29502] = 2
      "0000010" when "00111001100111111", -- t[29503] = 2
      "0000010" when "00111001101000000", -- t[29504] = 2
      "0000010" when "00111001101000001", -- t[29505] = 2
      "0000010" when "00111001101000010", -- t[29506] = 2
      "0000010" when "00111001101000011", -- t[29507] = 2
      "0000010" when "00111001101000100", -- t[29508] = 2
      "0000010" when "00111001101000101", -- t[29509] = 2
      "0000010" when "00111001101000110", -- t[29510] = 2
      "0000010" when "00111001101000111", -- t[29511] = 2
      "0000010" when "00111001101001000", -- t[29512] = 2
      "0000010" when "00111001101001001", -- t[29513] = 2
      "0000010" when "00111001101001010", -- t[29514] = 2
      "0000010" when "00111001101001011", -- t[29515] = 2
      "0000010" when "00111001101001100", -- t[29516] = 2
      "0000010" when "00111001101001101", -- t[29517] = 2
      "0000010" when "00111001101001110", -- t[29518] = 2
      "0000010" when "00111001101001111", -- t[29519] = 2
      "0000010" when "00111001101010000", -- t[29520] = 2
      "0000010" when "00111001101010001", -- t[29521] = 2
      "0000010" when "00111001101010010", -- t[29522] = 2
      "0000010" when "00111001101010011", -- t[29523] = 2
      "0000010" when "00111001101010100", -- t[29524] = 2
      "0000010" when "00111001101010101", -- t[29525] = 2
      "0000010" when "00111001101010110", -- t[29526] = 2
      "0000010" when "00111001101010111", -- t[29527] = 2
      "0000010" when "00111001101011000", -- t[29528] = 2
      "0000010" when "00111001101011001", -- t[29529] = 2
      "0000010" when "00111001101011010", -- t[29530] = 2
      "0000010" when "00111001101011011", -- t[29531] = 2
      "0000010" when "00111001101011100", -- t[29532] = 2
      "0000010" when "00111001101011101", -- t[29533] = 2
      "0000010" when "00111001101011110", -- t[29534] = 2
      "0000010" when "00111001101011111", -- t[29535] = 2
      "0000010" when "00111001101100000", -- t[29536] = 2
      "0000010" when "00111001101100001", -- t[29537] = 2
      "0000010" when "00111001101100010", -- t[29538] = 2
      "0000010" when "00111001101100011", -- t[29539] = 2
      "0000010" when "00111001101100100", -- t[29540] = 2
      "0000010" when "00111001101100101", -- t[29541] = 2
      "0000010" when "00111001101100110", -- t[29542] = 2
      "0000010" when "00111001101100111", -- t[29543] = 2
      "0000010" when "00111001101101000", -- t[29544] = 2
      "0000010" when "00111001101101001", -- t[29545] = 2
      "0000010" when "00111001101101010", -- t[29546] = 2
      "0000010" when "00111001101101011", -- t[29547] = 2
      "0000010" when "00111001101101100", -- t[29548] = 2
      "0000010" when "00111001101101101", -- t[29549] = 2
      "0000010" when "00111001101101110", -- t[29550] = 2
      "0000010" when "00111001101101111", -- t[29551] = 2
      "0000010" when "00111001101110000", -- t[29552] = 2
      "0000010" when "00111001101110001", -- t[29553] = 2
      "0000010" when "00111001101110010", -- t[29554] = 2
      "0000010" when "00111001101110011", -- t[29555] = 2
      "0000010" when "00111001101110100", -- t[29556] = 2
      "0000010" when "00111001101110101", -- t[29557] = 2
      "0000010" when "00111001101110110", -- t[29558] = 2
      "0000010" when "00111001101110111", -- t[29559] = 2
      "0000010" when "00111001101111000", -- t[29560] = 2
      "0000010" when "00111001101111001", -- t[29561] = 2
      "0000010" when "00111001101111010", -- t[29562] = 2
      "0000010" when "00111001101111011", -- t[29563] = 2
      "0000010" when "00111001101111100", -- t[29564] = 2
      "0000010" when "00111001101111101", -- t[29565] = 2
      "0000010" when "00111001101111110", -- t[29566] = 2
      "0000010" when "00111001101111111", -- t[29567] = 2
      "0000010" when "00111001110000000", -- t[29568] = 2
      "0000010" when "00111001110000001", -- t[29569] = 2
      "0000010" when "00111001110000010", -- t[29570] = 2
      "0000010" when "00111001110000011", -- t[29571] = 2
      "0000010" when "00111001110000100", -- t[29572] = 2
      "0000010" when "00111001110000101", -- t[29573] = 2
      "0000010" when "00111001110000110", -- t[29574] = 2
      "0000010" when "00111001110000111", -- t[29575] = 2
      "0000010" when "00111001110001000", -- t[29576] = 2
      "0000010" when "00111001110001001", -- t[29577] = 2
      "0000010" when "00111001110001010", -- t[29578] = 2
      "0000010" when "00111001110001011", -- t[29579] = 2
      "0000010" when "00111001110001100", -- t[29580] = 2
      "0000010" when "00111001110001101", -- t[29581] = 2
      "0000010" when "00111001110001110", -- t[29582] = 2
      "0000010" when "00111001110001111", -- t[29583] = 2
      "0000010" when "00111001110010000", -- t[29584] = 2
      "0000010" when "00111001110010001", -- t[29585] = 2
      "0000010" when "00111001110010010", -- t[29586] = 2
      "0000010" when "00111001110010011", -- t[29587] = 2
      "0000010" when "00111001110010100", -- t[29588] = 2
      "0000010" when "00111001110010101", -- t[29589] = 2
      "0000010" when "00111001110010110", -- t[29590] = 2
      "0000010" when "00111001110010111", -- t[29591] = 2
      "0000010" when "00111001110011000", -- t[29592] = 2
      "0000010" when "00111001110011001", -- t[29593] = 2
      "0000010" when "00111001110011010", -- t[29594] = 2
      "0000010" when "00111001110011011", -- t[29595] = 2
      "0000010" when "00111001110011100", -- t[29596] = 2
      "0000010" when "00111001110011101", -- t[29597] = 2
      "0000010" when "00111001110011110", -- t[29598] = 2
      "0000010" when "00111001110011111", -- t[29599] = 2
      "0000010" when "00111001110100000", -- t[29600] = 2
      "0000010" when "00111001110100001", -- t[29601] = 2
      "0000010" when "00111001110100010", -- t[29602] = 2
      "0000010" when "00111001110100011", -- t[29603] = 2
      "0000010" when "00111001110100100", -- t[29604] = 2
      "0000010" when "00111001110100101", -- t[29605] = 2
      "0000010" when "00111001110100110", -- t[29606] = 2
      "0000010" when "00111001110100111", -- t[29607] = 2
      "0000010" when "00111001110101000", -- t[29608] = 2
      "0000010" when "00111001110101001", -- t[29609] = 2
      "0000010" when "00111001110101010", -- t[29610] = 2
      "0000010" when "00111001110101011", -- t[29611] = 2
      "0000010" when "00111001110101100", -- t[29612] = 2
      "0000010" when "00111001110101101", -- t[29613] = 2
      "0000010" when "00111001110101110", -- t[29614] = 2
      "0000010" when "00111001110101111", -- t[29615] = 2
      "0000010" when "00111001110110000", -- t[29616] = 2
      "0000010" when "00111001110110001", -- t[29617] = 2
      "0000010" when "00111001110110010", -- t[29618] = 2
      "0000010" when "00111001110110011", -- t[29619] = 2
      "0000010" when "00111001110110100", -- t[29620] = 2
      "0000010" when "00111001110110101", -- t[29621] = 2
      "0000010" when "00111001110110110", -- t[29622] = 2
      "0000010" when "00111001110110111", -- t[29623] = 2
      "0000010" when "00111001110111000", -- t[29624] = 2
      "0000010" when "00111001110111001", -- t[29625] = 2
      "0000010" when "00111001110111010", -- t[29626] = 2
      "0000010" when "00111001110111011", -- t[29627] = 2
      "0000010" when "00111001110111100", -- t[29628] = 2
      "0000010" when "00111001110111101", -- t[29629] = 2
      "0000010" when "00111001110111110", -- t[29630] = 2
      "0000010" when "00111001110111111", -- t[29631] = 2
      "0000010" when "00111001111000000", -- t[29632] = 2
      "0000010" when "00111001111000001", -- t[29633] = 2
      "0000010" when "00111001111000010", -- t[29634] = 2
      "0000010" when "00111001111000011", -- t[29635] = 2
      "0000010" when "00111001111000100", -- t[29636] = 2
      "0000010" when "00111001111000101", -- t[29637] = 2
      "0000010" when "00111001111000110", -- t[29638] = 2
      "0000010" when "00111001111000111", -- t[29639] = 2
      "0000010" when "00111001111001000", -- t[29640] = 2
      "0000010" when "00111001111001001", -- t[29641] = 2
      "0000010" when "00111001111001010", -- t[29642] = 2
      "0000010" when "00111001111001011", -- t[29643] = 2
      "0000010" when "00111001111001100", -- t[29644] = 2
      "0000010" when "00111001111001101", -- t[29645] = 2
      "0000010" when "00111001111001110", -- t[29646] = 2
      "0000010" when "00111001111001111", -- t[29647] = 2
      "0000010" when "00111001111010000", -- t[29648] = 2
      "0000010" when "00111001111010001", -- t[29649] = 2
      "0000010" when "00111001111010010", -- t[29650] = 2
      "0000010" when "00111001111010011", -- t[29651] = 2
      "0000010" when "00111001111010100", -- t[29652] = 2
      "0000010" when "00111001111010101", -- t[29653] = 2
      "0000010" when "00111001111010110", -- t[29654] = 2
      "0000010" when "00111001111010111", -- t[29655] = 2
      "0000010" when "00111001111011000", -- t[29656] = 2
      "0000010" when "00111001111011001", -- t[29657] = 2
      "0000010" when "00111001111011010", -- t[29658] = 2
      "0000010" when "00111001111011011", -- t[29659] = 2
      "0000010" when "00111001111011100", -- t[29660] = 2
      "0000010" when "00111001111011101", -- t[29661] = 2
      "0000010" when "00111001111011110", -- t[29662] = 2
      "0000010" when "00111001111011111", -- t[29663] = 2
      "0000010" when "00111001111100000", -- t[29664] = 2
      "0000010" when "00111001111100001", -- t[29665] = 2
      "0000010" when "00111001111100010", -- t[29666] = 2
      "0000010" when "00111001111100011", -- t[29667] = 2
      "0000010" when "00111001111100100", -- t[29668] = 2
      "0000010" when "00111001111100101", -- t[29669] = 2
      "0000010" when "00111001111100110", -- t[29670] = 2
      "0000010" when "00111001111100111", -- t[29671] = 2
      "0000010" when "00111001111101000", -- t[29672] = 2
      "0000010" when "00111001111101001", -- t[29673] = 2
      "0000010" when "00111001111101010", -- t[29674] = 2
      "0000010" when "00111001111101011", -- t[29675] = 2
      "0000010" when "00111001111101100", -- t[29676] = 2
      "0000010" when "00111001111101101", -- t[29677] = 2
      "0000010" when "00111001111101110", -- t[29678] = 2
      "0000010" when "00111001111101111", -- t[29679] = 2
      "0000010" when "00111001111110000", -- t[29680] = 2
      "0000010" when "00111001111110001", -- t[29681] = 2
      "0000010" when "00111001111110010", -- t[29682] = 2
      "0000010" when "00111001111110011", -- t[29683] = 2
      "0000010" when "00111001111110100", -- t[29684] = 2
      "0000010" when "00111001111110101", -- t[29685] = 2
      "0000010" when "00111001111110110", -- t[29686] = 2
      "0000010" when "00111001111110111", -- t[29687] = 2
      "0000010" when "00111001111111000", -- t[29688] = 2
      "0000010" when "00111001111111001", -- t[29689] = 2
      "0000010" when "00111001111111010", -- t[29690] = 2
      "0000010" when "00111001111111011", -- t[29691] = 2
      "0000010" when "00111001111111100", -- t[29692] = 2
      "0000010" when "00111001111111101", -- t[29693] = 2
      "0000010" when "00111001111111110", -- t[29694] = 2
      "0000010" when "00111001111111111", -- t[29695] = 2
      "0000010" when "00111010000000000", -- t[29696] = 2
      "0000010" when "00111010000000001", -- t[29697] = 2
      "0000010" when "00111010000000010", -- t[29698] = 2
      "0000010" when "00111010000000011", -- t[29699] = 2
      "0000010" when "00111010000000100", -- t[29700] = 2
      "0000010" when "00111010000000101", -- t[29701] = 2
      "0000010" when "00111010000000110", -- t[29702] = 2
      "0000010" when "00111010000000111", -- t[29703] = 2
      "0000010" when "00111010000001000", -- t[29704] = 2
      "0000010" when "00111010000001001", -- t[29705] = 2
      "0000010" when "00111010000001010", -- t[29706] = 2
      "0000010" when "00111010000001011", -- t[29707] = 2
      "0000010" when "00111010000001100", -- t[29708] = 2
      "0000010" when "00111010000001101", -- t[29709] = 2
      "0000010" when "00111010000001110", -- t[29710] = 2
      "0000010" when "00111010000001111", -- t[29711] = 2
      "0000010" when "00111010000010000", -- t[29712] = 2
      "0000010" when "00111010000010001", -- t[29713] = 2
      "0000010" when "00111010000010010", -- t[29714] = 2
      "0000010" when "00111010000010011", -- t[29715] = 2
      "0000010" when "00111010000010100", -- t[29716] = 2
      "0000010" when "00111010000010101", -- t[29717] = 2
      "0000010" when "00111010000010110", -- t[29718] = 2
      "0000010" when "00111010000010111", -- t[29719] = 2
      "0000010" when "00111010000011000", -- t[29720] = 2
      "0000010" when "00111010000011001", -- t[29721] = 2
      "0000010" when "00111010000011010", -- t[29722] = 2
      "0000010" when "00111010000011011", -- t[29723] = 2
      "0000010" when "00111010000011100", -- t[29724] = 2
      "0000010" when "00111010000011101", -- t[29725] = 2
      "0000010" when "00111010000011110", -- t[29726] = 2
      "0000010" when "00111010000011111", -- t[29727] = 2
      "0000010" when "00111010000100000", -- t[29728] = 2
      "0000010" when "00111010000100001", -- t[29729] = 2
      "0000010" when "00111010000100010", -- t[29730] = 2
      "0000010" when "00111010000100011", -- t[29731] = 2
      "0000010" when "00111010000100100", -- t[29732] = 2
      "0000010" when "00111010000100101", -- t[29733] = 2
      "0000010" when "00111010000100110", -- t[29734] = 2
      "0000010" when "00111010000100111", -- t[29735] = 2
      "0000010" when "00111010000101000", -- t[29736] = 2
      "0000010" when "00111010000101001", -- t[29737] = 2
      "0000010" when "00111010000101010", -- t[29738] = 2
      "0000010" when "00111010000101011", -- t[29739] = 2
      "0000010" when "00111010000101100", -- t[29740] = 2
      "0000010" when "00111010000101101", -- t[29741] = 2
      "0000010" when "00111010000101110", -- t[29742] = 2
      "0000010" when "00111010000101111", -- t[29743] = 2
      "0000010" when "00111010000110000", -- t[29744] = 2
      "0000010" when "00111010000110001", -- t[29745] = 2
      "0000010" when "00111010000110010", -- t[29746] = 2
      "0000010" when "00111010000110011", -- t[29747] = 2
      "0000010" when "00111010000110100", -- t[29748] = 2
      "0000010" when "00111010000110101", -- t[29749] = 2
      "0000010" when "00111010000110110", -- t[29750] = 2
      "0000010" when "00111010000110111", -- t[29751] = 2
      "0000010" when "00111010000111000", -- t[29752] = 2
      "0000010" when "00111010000111001", -- t[29753] = 2
      "0000010" when "00111010000111010", -- t[29754] = 2
      "0000010" when "00111010000111011", -- t[29755] = 2
      "0000010" when "00111010000111100", -- t[29756] = 2
      "0000010" when "00111010000111101", -- t[29757] = 2
      "0000010" when "00111010000111110", -- t[29758] = 2
      "0000010" when "00111010000111111", -- t[29759] = 2
      "0000010" when "00111010001000000", -- t[29760] = 2
      "0000010" when "00111010001000001", -- t[29761] = 2
      "0000010" when "00111010001000010", -- t[29762] = 2
      "0000010" when "00111010001000011", -- t[29763] = 2
      "0000010" when "00111010001000100", -- t[29764] = 2
      "0000010" when "00111010001000101", -- t[29765] = 2
      "0000010" when "00111010001000110", -- t[29766] = 2
      "0000010" when "00111010001000111", -- t[29767] = 2
      "0000010" when "00111010001001000", -- t[29768] = 2
      "0000010" when "00111010001001001", -- t[29769] = 2
      "0000010" when "00111010001001010", -- t[29770] = 2
      "0000010" when "00111010001001011", -- t[29771] = 2
      "0000010" when "00111010001001100", -- t[29772] = 2
      "0000010" when "00111010001001101", -- t[29773] = 2
      "0000010" when "00111010001001110", -- t[29774] = 2
      "0000010" when "00111010001001111", -- t[29775] = 2
      "0000010" when "00111010001010000", -- t[29776] = 2
      "0000010" when "00111010001010001", -- t[29777] = 2
      "0000010" when "00111010001010010", -- t[29778] = 2
      "0000010" when "00111010001010011", -- t[29779] = 2
      "0000010" when "00111010001010100", -- t[29780] = 2
      "0000010" when "00111010001010101", -- t[29781] = 2
      "0000010" when "00111010001010110", -- t[29782] = 2
      "0000010" when "00111010001010111", -- t[29783] = 2
      "0000010" when "00111010001011000", -- t[29784] = 2
      "0000010" when "00111010001011001", -- t[29785] = 2
      "0000010" when "00111010001011010", -- t[29786] = 2
      "0000010" when "00111010001011011", -- t[29787] = 2
      "0000010" when "00111010001011100", -- t[29788] = 2
      "0000010" when "00111010001011101", -- t[29789] = 2
      "0000010" when "00111010001011110", -- t[29790] = 2
      "0000010" when "00111010001011111", -- t[29791] = 2
      "0000010" when "00111010001100000", -- t[29792] = 2
      "0000010" when "00111010001100001", -- t[29793] = 2
      "0000010" when "00111010001100010", -- t[29794] = 2
      "0000010" when "00111010001100011", -- t[29795] = 2
      "0000010" when "00111010001100100", -- t[29796] = 2
      "0000010" when "00111010001100101", -- t[29797] = 2
      "0000010" when "00111010001100110", -- t[29798] = 2
      "0000010" when "00111010001100111", -- t[29799] = 2
      "0000010" when "00111010001101000", -- t[29800] = 2
      "0000010" when "00111010001101001", -- t[29801] = 2
      "0000010" when "00111010001101010", -- t[29802] = 2
      "0000010" when "00111010001101011", -- t[29803] = 2
      "0000010" when "00111010001101100", -- t[29804] = 2
      "0000010" when "00111010001101101", -- t[29805] = 2
      "0000010" when "00111010001101110", -- t[29806] = 2
      "0000010" when "00111010001101111", -- t[29807] = 2
      "0000010" when "00111010001110000", -- t[29808] = 2
      "0000010" when "00111010001110001", -- t[29809] = 2
      "0000010" when "00111010001110010", -- t[29810] = 2
      "0000010" when "00111010001110011", -- t[29811] = 2
      "0000010" when "00111010001110100", -- t[29812] = 2
      "0000010" when "00111010001110101", -- t[29813] = 2
      "0000010" when "00111010001110110", -- t[29814] = 2
      "0000010" when "00111010001110111", -- t[29815] = 2
      "0000010" when "00111010001111000", -- t[29816] = 2
      "0000010" when "00111010001111001", -- t[29817] = 2
      "0000010" when "00111010001111010", -- t[29818] = 2
      "0000010" when "00111010001111011", -- t[29819] = 2
      "0000010" when "00111010001111100", -- t[29820] = 2
      "0000010" when "00111010001111101", -- t[29821] = 2
      "0000010" when "00111010001111110", -- t[29822] = 2
      "0000010" when "00111010001111111", -- t[29823] = 2
      "0000010" when "00111010010000000", -- t[29824] = 2
      "0000010" when "00111010010000001", -- t[29825] = 2
      "0000010" when "00111010010000010", -- t[29826] = 2
      "0000010" when "00111010010000011", -- t[29827] = 2
      "0000010" when "00111010010000100", -- t[29828] = 2
      "0000010" when "00111010010000101", -- t[29829] = 2
      "0000010" when "00111010010000110", -- t[29830] = 2
      "0000010" when "00111010010000111", -- t[29831] = 2
      "0000010" when "00111010010001000", -- t[29832] = 2
      "0000010" when "00111010010001001", -- t[29833] = 2
      "0000010" when "00111010010001010", -- t[29834] = 2
      "0000010" when "00111010010001011", -- t[29835] = 2
      "0000010" when "00111010010001100", -- t[29836] = 2
      "0000010" when "00111010010001101", -- t[29837] = 2
      "0000010" when "00111010010001110", -- t[29838] = 2
      "0000010" when "00111010010001111", -- t[29839] = 2
      "0000010" when "00111010010010000", -- t[29840] = 2
      "0000010" when "00111010010010001", -- t[29841] = 2
      "0000010" when "00111010010010010", -- t[29842] = 2
      "0000010" when "00111010010010011", -- t[29843] = 2
      "0000010" when "00111010010010100", -- t[29844] = 2
      "0000010" when "00111010010010101", -- t[29845] = 2
      "0000010" when "00111010010010110", -- t[29846] = 2
      "0000010" when "00111010010010111", -- t[29847] = 2
      "0000010" when "00111010010011000", -- t[29848] = 2
      "0000010" when "00111010010011001", -- t[29849] = 2
      "0000010" when "00111010010011010", -- t[29850] = 2
      "0000010" when "00111010010011011", -- t[29851] = 2
      "0000010" when "00111010010011100", -- t[29852] = 2
      "0000010" when "00111010010011101", -- t[29853] = 2
      "0000010" when "00111010010011110", -- t[29854] = 2
      "0000010" when "00111010010011111", -- t[29855] = 2
      "0000010" when "00111010010100000", -- t[29856] = 2
      "0000010" when "00111010010100001", -- t[29857] = 2
      "0000010" when "00111010010100010", -- t[29858] = 2
      "0000010" when "00111010010100011", -- t[29859] = 2
      "0000010" when "00111010010100100", -- t[29860] = 2
      "0000010" when "00111010010100101", -- t[29861] = 2
      "0000010" when "00111010010100110", -- t[29862] = 2
      "0000010" when "00111010010100111", -- t[29863] = 2
      "0000010" when "00111010010101000", -- t[29864] = 2
      "0000010" when "00111010010101001", -- t[29865] = 2
      "0000010" when "00111010010101010", -- t[29866] = 2
      "0000010" when "00111010010101011", -- t[29867] = 2
      "0000010" when "00111010010101100", -- t[29868] = 2
      "0000010" when "00111010010101101", -- t[29869] = 2
      "0000010" when "00111010010101110", -- t[29870] = 2
      "0000010" when "00111010010101111", -- t[29871] = 2
      "0000010" when "00111010010110000", -- t[29872] = 2
      "0000010" when "00111010010110001", -- t[29873] = 2
      "0000010" when "00111010010110010", -- t[29874] = 2
      "0000010" when "00111010010110011", -- t[29875] = 2
      "0000010" when "00111010010110100", -- t[29876] = 2
      "0000010" when "00111010010110101", -- t[29877] = 2
      "0000010" when "00111010010110110", -- t[29878] = 2
      "0000010" when "00111010010110111", -- t[29879] = 2
      "0000010" when "00111010010111000", -- t[29880] = 2
      "0000010" when "00111010010111001", -- t[29881] = 2
      "0000010" when "00111010010111010", -- t[29882] = 2
      "0000010" when "00111010010111011", -- t[29883] = 2
      "0000010" when "00111010010111100", -- t[29884] = 2
      "0000010" when "00111010010111101", -- t[29885] = 2
      "0000010" when "00111010010111110", -- t[29886] = 2
      "0000010" when "00111010010111111", -- t[29887] = 2
      "0000010" when "00111010011000000", -- t[29888] = 2
      "0000010" when "00111010011000001", -- t[29889] = 2
      "0000010" when "00111010011000010", -- t[29890] = 2
      "0000010" when "00111010011000011", -- t[29891] = 2
      "0000010" when "00111010011000100", -- t[29892] = 2
      "0000010" when "00111010011000101", -- t[29893] = 2
      "0000010" when "00111010011000110", -- t[29894] = 2
      "0000010" when "00111010011000111", -- t[29895] = 2
      "0000010" when "00111010011001000", -- t[29896] = 2
      "0000010" when "00111010011001001", -- t[29897] = 2
      "0000010" when "00111010011001010", -- t[29898] = 2
      "0000010" when "00111010011001011", -- t[29899] = 2
      "0000010" when "00111010011001100", -- t[29900] = 2
      "0000010" when "00111010011001101", -- t[29901] = 2
      "0000010" when "00111010011001110", -- t[29902] = 2
      "0000010" when "00111010011001111", -- t[29903] = 2
      "0000010" when "00111010011010000", -- t[29904] = 2
      "0000010" when "00111010011010001", -- t[29905] = 2
      "0000010" when "00111010011010010", -- t[29906] = 2
      "0000010" when "00111010011010011", -- t[29907] = 2
      "0000010" when "00111010011010100", -- t[29908] = 2
      "0000010" when "00111010011010101", -- t[29909] = 2
      "0000010" when "00111010011010110", -- t[29910] = 2
      "0000010" when "00111010011010111", -- t[29911] = 2
      "0000010" when "00111010011011000", -- t[29912] = 2
      "0000010" when "00111010011011001", -- t[29913] = 2
      "0000010" when "00111010011011010", -- t[29914] = 2
      "0000010" when "00111010011011011", -- t[29915] = 2
      "0000010" when "00111010011011100", -- t[29916] = 2
      "0000010" when "00111010011011101", -- t[29917] = 2
      "0000010" when "00111010011011110", -- t[29918] = 2
      "0000010" when "00111010011011111", -- t[29919] = 2
      "0000010" when "00111010011100000", -- t[29920] = 2
      "0000010" when "00111010011100001", -- t[29921] = 2
      "0000010" when "00111010011100010", -- t[29922] = 2
      "0000010" when "00111010011100011", -- t[29923] = 2
      "0000010" when "00111010011100100", -- t[29924] = 2
      "0000010" when "00111010011100101", -- t[29925] = 2
      "0000010" when "00111010011100110", -- t[29926] = 2
      "0000010" when "00111010011100111", -- t[29927] = 2
      "0000010" when "00111010011101000", -- t[29928] = 2
      "0000010" when "00111010011101001", -- t[29929] = 2
      "0000010" when "00111010011101010", -- t[29930] = 2
      "0000010" when "00111010011101011", -- t[29931] = 2
      "0000010" when "00111010011101100", -- t[29932] = 2
      "0000010" when "00111010011101101", -- t[29933] = 2
      "0000010" when "00111010011101110", -- t[29934] = 2
      "0000010" when "00111010011101111", -- t[29935] = 2
      "0000010" when "00111010011110000", -- t[29936] = 2
      "0000010" when "00111010011110001", -- t[29937] = 2
      "0000010" when "00111010011110010", -- t[29938] = 2
      "0000010" when "00111010011110011", -- t[29939] = 2
      "0000010" when "00111010011110100", -- t[29940] = 2
      "0000010" when "00111010011110101", -- t[29941] = 2
      "0000010" when "00111010011110110", -- t[29942] = 2
      "0000010" when "00111010011110111", -- t[29943] = 2
      "0000010" when "00111010011111000", -- t[29944] = 2
      "0000010" when "00111010011111001", -- t[29945] = 2
      "0000010" when "00111010011111010", -- t[29946] = 2
      "0000010" when "00111010011111011", -- t[29947] = 2
      "0000010" when "00111010011111100", -- t[29948] = 2
      "0000010" when "00111010011111101", -- t[29949] = 2
      "0000010" when "00111010011111110", -- t[29950] = 2
      "0000010" when "00111010011111111", -- t[29951] = 2
      "0000010" when "00111010100000000", -- t[29952] = 2
      "0000010" when "00111010100000001", -- t[29953] = 2
      "0000010" when "00111010100000010", -- t[29954] = 2
      "0000010" when "00111010100000011", -- t[29955] = 2
      "0000010" when "00111010100000100", -- t[29956] = 2
      "0000010" when "00111010100000101", -- t[29957] = 2
      "0000010" when "00111010100000110", -- t[29958] = 2
      "0000010" when "00111010100000111", -- t[29959] = 2
      "0000010" when "00111010100001000", -- t[29960] = 2
      "0000010" when "00111010100001001", -- t[29961] = 2
      "0000010" when "00111010100001010", -- t[29962] = 2
      "0000010" when "00111010100001011", -- t[29963] = 2
      "0000010" when "00111010100001100", -- t[29964] = 2
      "0000010" when "00111010100001101", -- t[29965] = 2
      "0000010" when "00111010100001110", -- t[29966] = 2
      "0000010" when "00111010100001111", -- t[29967] = 2
      "0000010" when "00111010100010000", -- t[29968] = 2
      "0000010" when "00111010100010001", -- t[29969] = 2
      "0000010" when "00111010100010010", -- t[29970] = 2
      "0000010" when "00111010100010011", -- t[29971] = 2
      "0000010" when "00111010100010100", -- t[29972] = 2
      "0000010" when "00111010100010101", -- t[29973] = 2
      "0000010" when "00111010100010110", -- t[29974] = 2
      "0000010" when "00111010100010111", -- t[29975] = 2
      "0000010" when "00111010100011000", -- t[29976] = 2
      "0000010" when "00111010100011001", -- t[29977] = 2
      "0000010" when "00111010100011010", -- t[29978] = 2
      "0000010" when "00111010100011011", -- t[29979] = 2
      "0000010" when "00111010100011100", -- t[29980] = 2
      "0000010" when "00111010100011101", -- t[29981] = 2
      "0000010" when "00111010100011110", -- t[29982] = 2
      "0000010" when "00111010100011111", -- t[29983] = 2
      "0000010" when "00111010100100000", -- t[29984] = 2
      "0000010" when "00111010100100001", -- t[29985] = 2
      "0000010" when "00111010100100010", -- t[29986] = 2
      "0000010" when "00111010100100011", -- t[29987] = 2
      "0000010" when "00111010100100100", -- t[29988] = 2
      "0000010" when "00111010100100101", -- t[29989] = 2
      "0000010" when "00111010100100110", -- t[29990] = 2
      "0000010" when "00111010100100111", -- t[29991] = 2
      "0000010" when "00111010100101000", -- t[29992] = 2
      "0000010" when "00111010100101001", -- t[29993] = 2
      "0000010" when "00111010100101010", -- t[29994] = 2
      "0000010" when "00111010100101011", -- t[29995] = 2
      "0000010" when "00111010100101100", -- t[29996] = 2
      "0000010" when "00111010100101101", -- t[29997] = 2
      "0000010" when "00111010100101110", -- t[29998] = 2
      "0000010" when "00111010100101111", -- t[29999] = 2
      "0000010" when "00111010100110000", -- t[30000] = 2
      "0000010" when "00111010100110001", -- t[30001] = 2
      "0000010" when "00111010100110010", -- t[30002] = 2
      "0000010" when "00111010100110011", -- t[30003] = 2
      "0000010" when "00111010100110100", -- t[30004] = 2
      "0000010" when "00111010100110101", -- t[30005] = 2
      "0000010" when "00111010100110110", -- t[30006] = 2
      "0000010" when "00111010100110111", -- t[30007] = 2
      "0000010" when "00111010100111000", -- t[30008] = 2
      "0000010" when "00111010100111001", -- t[30009] = 2
      "0000010" when "00111010100111010", -- t[30010] = 2
      "0000010" when "00111010100111011", -- t[30011] = 2
      "0000010" when "00111010100111100", -- t[30012] = 2
      "0000010" when "00111010100111101", -- t[30013] = 2
      "0000010" when "00111010100111110", -- t[30014] = 2
      "0000010" when "00111010100111111", -- t[30015] = 2
      "0000010" when "00111010101000000", -- t[30016] = 2
      "0000010" when "00111010101000001", -- t[30017] = 2
      "0000010" when "00111010101000010", -- t[30018] = 2
      "0000010" when "00111010101000011", -- t[30019] = 2
      "0000010" when "00111010101000100", -- t[30020] = 2
      "0000010" when "00111010101000101", -- t[30021] = 2
      "0000010" when "00111010101000110", -- t[30022] = 2
      "0000010" when "00111010101000111", -- t[30023] = 2
      "0000010" when "00111010101001000", -- t[30024] = 2
      "0000010" when "00111010101001001", -- t[30025] = 2
      "0000010" when "00111010101001010", -- t[30026] = 2
      "0000010" when "00111010101001011", -- t[30027] = 2
      "0000010" when "00111010101001100", -- t[30028] = 2
      "0000010" when "00111010101001101", -- t[30029] = 2
      "0000010" when "00111010101001110", -- t[30030] = 2
      "0000010" when "00111010101001111", -- t[30031] = 2
      "0000010" when "00111010101010000", -- t[30032] = 2
      "0000010" when "00111010101010001", -- t[30033] = 2
      "0000010" when "00111010101010010", -- t[30034] = 2
      "0000010" when "00111010101010011", -- t[30035] = 2
      "0000010" when "00111010101010100", -- t[30036] = 2
      "0000010" when "00111010101010101", -- t[30037] = 2
      "0000010" when "00111010101010110", -- t[30038] = 2
      "0000010" when "00111010101010111", -- t[30039] = 2
      "0000010" when "00111010101011000", -- t[30040] = 2
      "0000010" when "00111010101011001", -- t[30041] = 2
      "0000010" when "00111010101011010", -- t[30042] = 2
      "0000010" when "00111010101011011", -- t[30043] = 2
      "0000010" when "00111010101011100", -- t[30044] = 2
      "0000010" when "00111010101011101", -- t[30045] = 2
      "0000010" when "00111010101011110", -- t[30046] = 2
      "0000010" when "00111010101011111", -- t[30047] = 2
      "0000010" when "00111010101100000", -- t[30048] = 2
      "0000010" when "00111010101100001", -- t[30049] = 2
      "0000010" when "00111010101100010", -- t[30050] = 2
      "0000010" when "00111010101100011", -- t[30051] = 2
      "0000010" when "00111010101100100", -- t[30052] = 2
      "0000010" when "00111010101100101", -- t[30053] = 2
      "0000010" when "00111010101100110", -- t[30054] = 2
      "0000010" when "00111010101100111", -- t[30055] = 2
      "0000010" when "00111010101101000", -- t[30056] = 2
      "0000010" when "00111010101101001", -- t[30057] = 2
      "0000010" when "00111010101101010", -- t[30058] = 2
      "0000010" when "00111010101101011", -- t[30059] = 2
      "0000010" when "00111010101101100", -- t[30060] = 2
      "0000010" when "00111010101101101", -- t[30061] = 2
      "0000010" when "00111010101101110", -- t[30062] = 2
      "0000010" when "00111010101101111", -- t[30063] = 2
      "0000010" when "00111010101110000", -- t[30064] = 2
      "0000010" when "00111010101110001", -- t[30065] = 2
      "0000010" when "00111010101110010", -- t[30066] = 2
      "0000010" when "00111010101110011", -- t[30067] = 2
      "0000010" when "00111010101110100", -- t[30068] = 2
      "0000010" when "00111010101110101", -- t[30069] = 2
      "0000010" when "00111010101110110", -- t[30070] = 2
      "0000010" when "00111010101110111", -- t[30071] = 2
      "0000010" when "00111010101111000", -- t[30072] = 2
      "0000010" when "00111010101111001", -- t[30073] = 2
      "0000010" when "00111010101111010", -- t[30074] = 2
      "0000010" when "00111010101111011", -- t[30075] = 2
      "0000010" when "00111010101111100", -- t[30076] = 2
      "0000010" when "00111010101111101", -- t[30077] = 2
      "0000010" when "00111010101111110", -- t[30078] = 2
      "0000010" when "00111010101111111", -- t[30079] = 2
      "0000010" when "00111010110000000", -- t[30080] = 2
      "0000010" when "00111010110000001", -- t[30081] = 2
      "0000010" when "00111010110000010", -- t[30082] = 2
      "0000010" when "00111010110000011", -- t[30083] = 2
      "0000010" when "00111010110000100", -- t[30084] = 2
      "0000010" when "00111010110000101", -- t[30085] = 2
      "0000010" when "00111010110000110", -- t[30086] = 2
      "0000010" when "00111010110000111", -- t[30087] = 2
      "0000010" when "00111010110001000", -- t[30088] = 2
      "0000010" when "00111010110001001", -- t[30089] = 2
      "0000010" when "00111010110001010", -- t[30090] = 2
      "0000010" when "00111010110001011", -- t[30091] = 2
      "0000010" when "00111010110001100", -- t[30092] = 2
      "0000010" when "00111010110001101", -- t[30093] = 2
      "0000010" when "00111010110001110", -- t[30094] = 2
      "0000010" when "00111010110001111", -- t[30095] = 2
      "0000010" when "00111010110010000", -- t[30096] = 2
      "0000010" when "00111010110010001", -- t[30097] = 2
      "0000010" when "00111010110010010", -- t[30098] = 2
      "0000010" when "00111010110010011", -- t[30099] = 2
      "0000010" when "00111010110010100", -- t[30100] = 2
      "0000010" when "00111010110010101", -- t[30101] = 2
      "0000010" when "00111010110010110", -- t[30102] = 2
      "0000010" when "00111010110010111", -- t[30103] = 2
      "0000010" when "00111010110011000", -- t[30104] = 2
      "0000010" when "00111010110011001", -- t[30105] = 2
      "0000010" when "00111010110011010", -- t[30106] = 2
      "0000010" when "00111010110011011", -- t[30107] = 2
      "0000010" when "00111010110011100", -- t[30108] = 2
      "0000010" when "00111010110011101", -- t[30109] = 2
      "0000010" when "00111010110011110", -- t[30110] = 2
      "0000010" when "00111010110011111", -- t[30111] = 2
      "0000010" when "00111010110100000", -- t[30112] = 2
      "0000010" when "00111010110100001", -- t[30113] = 2
      "0000010" when "00111010110100010", -- t[30114] = 2
      "0000010" when "00111010110100011", -- t[30115] = 2
      "0000010" when "00111010110100100", -- t[30116] = 2
      "0000010" when "00111010110100101", -- t[30117] = 2
      "0000010" when "00111010110100110", -- t[30118] = 2
      "0000010" when "00111010110100111", -- t[30119] = 2
      "0000010" when "00111010110101000", -- t[30120] = 2
      "0000010" when "00111010110101001", -- t[30121] = 2
      "0000010" when "00111010110101010", -- t[30122] = 2
      "0000010" when "00111010110101011", -- t[30123] = 2
      "0000010" when "00111010110101100", -- t[30124] = 2
      "0000010" when "00111010110101101", -- t[30125] = 2
      "0000010" when "00111010110101110", -- t[30126] = 2
      "0000010" when "00111010110101111", -- t[30127] = 2
      "0000010" when "00111010110110000", -- t[30128] = 2
      "0000010" when "00111010110110001", -- t[30129] = 2
      "0000010" when "00111010110110010", -- t[30130] = 2
      "0000010" when "00111010110110011", -- t[30131] = 2
      "0000010" when "00111010110110100", -- t[30132] = 2
      "0000010" when "00111010110110101", -- t[30133] = 2
      "0000010" when "00111010110110110", -- t[30134] = 2
      "0000010" when "00111010110110111", -- t[30135] = 2
      "0000010" when "00111010110111000", -- t[30136] = 2
      "0000010" when "00111010110111001", -- t[30137] = 2
      "0000010" when "00111010110111010", -- t[30138] = 2
      "0000010" when "00111010110111011", -- t[30139] = 2
      "0000010" when "00111010110111100", -- t[30140] = 2
      "0000010" when "00111010110111101", -- t[30141] = 2
      "0000010" when "00111010110111110", -- t[30142] = 2
      "0000010" when "00111010110111111", -- t[30143] = 2
      "0000010" when "00111010111000000", -- t[30144] = 2
      "0000010" when "00111010111000001", -- t[30145] = 2
      "0000010" when "00111010111000010", -- t[30146] = 2
      "0000010" when "00111010111000011", -- t[30147] = 2
      "0000010" when "00111010111000100", -- t[30148] = 2
      "0000010" when "00111010111000101", -- t[30149] = 2
      "0000010" when "00111010111000110", -- t[30150] = 2
      "0000010" when "00111010111000111", -- t[30151] = 2
      "0000010" when "00111010111001000", -- t[30152] = 2
      "0000010" when "00111010111001001", -- t[30153] = 2
      "0000010" when "00111010111001010", -- t[30154] = 2
      "0000010" when "00111010111001011", -- t[30155] = 2
      "0000010" when "00111010111001100", -- t[30156] = 2
      "0000010" when "00111010111001101", -- t[30157] = 2
      "0000010" when "00111010111001110", -- t[30158] = 2
      "0000010" when "00111010111001111", -- t[30159] = 2
      "0000010" when "00111010111010000", -- t[30160] = 2
      "0000010" when "00111010111010001", -- t[30161] = 2
      "0000010" when "00111010111010010", -- t[30162] = 2
      "0000010" when "00111010111010011", -- t[30163] = 2
      "0000010" when "00111010111010100", -- t[30164] = 2
      "0000010" when "00111010111010101", -- t[30165] = 2
      "0000010" when "00111010111010110", -- t[30166] = 2
      "0000010" when "00111010111010111", -- t[30167] = 2
      "0000010" when "00111010111011000", -- t[30168] = 2
      "0000010" when "00111010111011001", -- t[30169] = 2
      "0000010" when "00111010111011010", -- t[30170] = 2
      "0000010" when "00111010111011011", -- t[30171] = 2
      "0000010" when "00111010111011100", -- t[30172] = 2
      "0000010" when "00111010111011101", -- t[30173] = 2
      "0000010" when "00111010111011110", -- t[30174] = 2
      "0000010" when "00111010111011111", -- t[30175] = 2
      "0000010" when "00111010111100000", -- t[30176] = 2
      "0000010" when "00111010111100001", -- t[30177] = 2
      "0000010" when "00111010111100010", -- t[30178] = 2
      "0000010" when "00111010111100011", -- t[30179] = 2
      "0000010" when "00111010111100100", -- t[30180] = 2
      "0000010" when "00111010111100101", -- t[30181] = 2
      "0000010" when "00111010111100110", -- t[30182] = 2
      "0000010" when "00111010111100111", -- t[30183] = 2
      "0000010" when "00111010111101000", -- t[30184] = 2
      "0000010" when "00111010111101001", -- t[30185] = 2
      "0000010" when "00111010111101010", -- t[30186] = 2
      "0000010" when "00111010111101011", -- t[30187] = 2
      "0000010" when "00111010111101100", -- t[30188] = 2
      "0000010" when "00111010111101101", -- t[30189] = 2
      "0000010" when "00111010111101110", -- t[30190] = 2
      "0000010" when "00111010111101111", -- t[30191] = 2
      "0000010" when "00111010111110000", -- t[30192] = 2
      "0000010" when "00111010111110001", -- t[30193] = 2
      "0000010" when "00111010111110010", -- t[30194] = 2
      "0000010" when "00111010111110011", -- t[30195] = 2
      "0000010" when "00111010111110100", -- t[30196] = 2
      "0000010" when "00111010111110101", -- t[30197] = 2
      "0000010" when "00111010111110110", -- t[30198] = 2
      "0000010" when "00111010111110111", -- t[30199] = 2
      "0000010" when "00111010111111000", -- t[30200] = 2
      "0000010" when "00111010111111001", -- t[30201] = 2
      "0000010" when "00111010111111010", -- t[30202] = 2
      "0000010" when "00111010111111011", -- t[30203] = 2
      "0000010" when "00111010111111100", -- t[30204] = 2
      "0000010" when "00111010111111101", -- t[30205] = 2
      "0000010" when "00111010111111110", -- t[30206] = 2
      "0000010" when "00111010111111111", -- t[30207] = 2
      "0000010" when "00111011000000000", -- t[30208] = 2
      "0000010" when "00111011000000001", -- t[30209] = 2
      "0000010" when "00111011000000010", -- t[30210] = 2
      "0000010" when "00111011000000011", -- t[30211] = 2
      "0000010" when "00111011000000100", -- t[30212] = 2
      "0000010" when "00111011000000101", -- t[30213] = 2
      "0000010" when "00111011000000110", -- t[30214] = 2
      "0000010" when "00111011000000111", -- t[30215] = 2
      "0000010" when "00111011000001000", -- t[30216] = 2
      "0000010" when "00111011000001001", -- t[30217] = 2
      "0000010" when "00111011000001010", -- t[30218] = 2
      "0000010" when "00111011000001011", -- t[30219] = 2
      "0000010" when "00111011000001100", -- t[30220] = 2
      "0000010" when "00111011000001101", -- t[30221] = 2
      "0000010" when "00111011000001110", -- t[30222] = 2
      "0000010" when "00111011000001111", -- t[30223] = 2
      "0000010" when "00111011000010000", -- t[30224] = 2
      "0000010" when "00111011000010001", -- t[30225] = 2
      "0000010" when "00111011000010010", -- t[30226] = 2
      "0000010" when "00111011000010011", -- t[30227] = 2
      "0000010" when "00111011000010100", -- t[30228] = 2
      "0000010" when "00111011000010101", -- t[30229] = 2
      "0000010" when "00111011000010110", -- t[30230] = 2
      "0000010" when "00111011000010111", -- t[30231] = 2
      "0000010" when "00111011000011000", -- t[30232] = 2
      "0000010" when "00111011000011001", -- t[30233] = 2
      "0000010" when "00111011000011010", -- t[30234] = 2
      "0000010" when "00111011000011011", -- t[30235] = 2
      "0000010" when "00111011000011100", -- t[30236] = 2
      "0000010" when "00111011000011101", -- t[30237] = 2
      "0000010" when "00111011000011110", -- t[30238] = 2
      "0000010" when "00111011000011111", -- t[30239] = 2
      "0000010" when "00111011000100000", -- t[30240] = 2
      "0000010" when "00111011000100001", -- t[30241] = 2
      "0000010" when "00111011000100010", -- t[30242] = 2
      "0000010" when "00111011000100011", -- t[30243] = 2
      "0000010" when "00111011000100100", -- t[30244] = 2
      "0000010" when "00111011000100101", -- t[30245] = 2
      "0000010" when "00111011000100110", -- t[30246] = 2
      "0000010" when "00111011000100111", -- t[30247] = 2
      "0000010" when "00111011000101000", -- t[30248] = 2
      "0000010" when "00111011000101001", -- t[30249] = 2
      "0000010" when "00111011000101010", -- t[30250] = 2
      "0000010" when "00111011000101011", -- t[30251] = 2
      "0000010" when "00111011000101100", -- t[30252] = 2
      "0000010" when "00111011000101101", -- t[30253] = 2
      "0000010" when "00111011000101110", -- t[30254] = 2
      "0000010" when "00111011000101111", -- t[30255] = 2
      "0000010" when "00111011000110000", -- t[30256] = 2
      "0000010" when "00111011000110001", -- t[30257] = 2
      "0000010" when "00111011000110010", -- t[30258] = 2
      "0000010" when "00111011000110011", -- t[30259] = 2
      "0000010" when "00111011000110100", -- t[30260] = 2
      "0000010" when "00111011000110101", -- t[30261] = 2
      "0000010" when "00111011000110110", -- t[30262] = 2
      "0000010" when "00111011000110111", -- t[30263] = 2
      "0000010" when "00111011000111000", -- t[30264] = 2
      "0000010" when "00111011000111001", -- t[30265] = 2
      "0000010" when "00111011000111010", -- t[30266] = 2
      "0000010" when "00111011000111011", -- t[30267] = 2
      "0000010" when "00111011000111100", -- t[30268] = 2
      "0000010" when "00111011000111101", -- t[30269] = 2
      "0000010" when "00111011000111110", -- t[30270] = 2
      "0000010" when "00111011000111111", -- t[30271] = 2
      "0000010" when "00111011001000000", -- t[30272] = 2
      "0000010" when "00111011001000001", -- t[30273] = 2
      "0000010" when "00111011001000010", -- t[30274] = 2
      "0000010" when "00111011001000011", -- t[30275] = 2
      "0000010" when "00111011001000100", -- t[30276] = 2
      "0000010" when "00111011001000101", -- t[30277] = 2
      "0000010" when "00111011001000110", -- t[30278] = 2
      "0000010" when "00111011001000111", -- t[30279] = 2
      "0000010" when "00111011001001000", -- t[30280] = 2
      "0000010" when "00111011001001001", -- t[30281] = 2
      "0000010" when "00111011001001010", -- t[30282] = 2
      "0000010" when "00111011001001011", -- t[30283] = 2
      "0000010" when "00111011001001100", -- t[30284] = 2
      "0000010" when "00111011001001101", -- t[30285] = 2
      "0000010" when "00111011001001110", -- t[30286] = 2
      "0000010" when "00111011001001111", -- t[30287] = 2
      "0000010" when "00111011001010000", -- t[30288] = 2
      "0000010" when "00111011001010001", -- t[30289] = 2
      "0000010" when "00111011001010010", -- t[30290] = 2
      "0000010" when "00111011001010011", -- t[30291] = 2
      "0000010" when "00111011001010100", -- t[30292] = 2
      "0000010" when "00111011001010101", -- t[30293] = 2
      "0000010" when "00111011001010110", -- t[30294] = 2
      "0000010" when "00111011001010111", -- t[30295] = 2
      "0000010" when "00111011001011000", -- t[30296] = 2
      "0000010" when "00111011001011001", -- t[30297] = 2
      "0000010" when "00111011001011010", -- t[30298] = 2
      "0000010" when "00111011001011011", -- t[30299] = 2
      "0000010" when "00111011001011100", -- t[30300] = 2
      "0000010" when "00111011001011101", -- t[30301] = 2
      "0000010" when "00111011001011110", -- t[30302] = 2
      "0000010" when "00111011001011111", -- t[30303] = 2
      "0000010" when "00111011001100000", -- t[30304] = 2
      "0000010" when "00111011001100001", -- t[30305] = 2
      "0000010" when "00111011001100010", -- t[30306] = 2
      "0000010" when "00111011001100011", -- t[30307] = 2
      "0000010" when "00111011001100100", -- t[30308] = 2
      "0000010" when "00111011001100101", -- t[30309] = 2
      "0000010" when "00111011001100110", -- t[30310] = 2
      "0000010" when "00111011001100111", -- t[30311] = 2
      "0000010" when "00111011001101000", -- t[30312] = 2
      "0000010" when "00111011001101001", -- t[30313] = 2
      "0000010" when "00111011001101010", -- t[30314] = 2
      "0000010" when "00111011001101011", -- t[30315] = 2
      "0000010" when "00111011001101100", -- t[30316] = 2
      "0000010" when "00111011001101101", -- t[30317] = 2
      "0000010" when "00111011001101110", -- t[30318] = 2
      "0000010" when "00111011001101111", -- t[30319] = 2
      "0000010" when "00111011001110000", -- t[30320] = 2
      "0000010" when "00111011001110001", -- t[30321] = 2
      "0000010" when "00111011001110010", -- t[30322] = 2
      "0000010" when "00111011001110011", -- t[30323] = 2
      "0000010" when "00111011001110100", -- t[30324] = 2
      "0000010" when "00111011001110101", -- t[30325] = 2
      "0000010" when "00111011001110110", -- t[30326] = 2
      "0000010" when "00111011001110111", -- t[30327] = 2
      "0000010" when "00111011001111000", -- t[30328] = 2
      "0000010" when "00111011001111001", -- t[30329] = 2
      "0000010" when "00111011001111010", -- t[30330] = 2
      "0000010" when "00111011001111011", -- t[30331] = 2
      "0000010" when "00111011001111100", -- t[30332] = 2
      "0000010" when "00111011001111101", -- t[30333] = 2
      "0000010" when "00111011001111110", -- t[30334] = 2
      "0000010" when "00111011001111111", -- t[30335] = 2
      "0000010" when "00111011010000000", -- t[30336] = 2
      "0000010" when "00111011010000001", -- t[30337] = 2
      "0000010" when "00111011010000010", -- t[30338] = 2
      "0000010" when "00111011010000011", -- t[30339] = 2
      "0000010" when "00111011010000100", -- t[30340] = 2
      "0000010" when "00111011010000101", -- t[30341] = 2
      "0000010" when "00111011010000110", -- t[30342] = 2
      "0000010" when "00111011010000111", -- t[30343] = 2
      "0000010" when "00111011010001000", -- t[30344] = 2
      "0000010" when "00111011010001001", -- t[30345] = 2
      "0000010" when "00111011010001010", -- t[30346] = 2
      "0000010" when "00111011010001011", -- t[30347] = 2
      "0000010" when "00111011010001100", -- t[30348] = 2
      "0000010" when "00111011010001101", -- t[30349] = 2
      "0000010" when "00111011010001110", -- t[30350] = 2
      "0000010" when "00111011010001111", -- t[30351] = 2
      "0000010" when "00111011010010000", -- t[30352] = 2
      "0000010" when "00111011010010001", -- t[30353] = 2
      "0000010" when "00111011010010010", -- t[30354] = 2
      "0000010" when "00111011010010011", -- t[30355] = 2
      "0000010" when "00111011010010100", -- t[30356] = 2
      "0000010" when "00111011010010101", -- t[30357] = 2
      "0000010" when "00111011010010110", -- t[30358] = 2
      "0000010" when "00111011010010111", -- t[30359] = 2
      "0000010" when "00111011010011000", -- t[30360] = 2
      "0000010" when "00111011010011001", -- t[30361] = 2
      "0000010" when "00111011010011010", -- t[30362] = 2
      "0000010" when "00111011010011011", -- t[30363] = 2
      "0000010" when "00111011010011100", -- t[30364] = 2
      "0000010" when "00111011010011101", -- t[30365] = 2
      "0000010" when "00111011010011110", -- t[30366] = 2
      "0000010" when "00111011010011111", -- t[30367] = 2
      "0000010" when "00111011010100000", -- t[30368] = 2
      "0000010" when "00111011010100001", -- t[30369] = 2
      "0000010" when "00111011010100010", -- t[30370] = 2
      "0000010" when "00111011010100011", -- t[30371] = 2
      "0000010" when "00111011010100100", -- t[30372] = 2
      "0000010" when "00111011010100101", -- t[30373] = 2
      "0000010" when "00111011010100110", -- t[30374] = 2
      "0000010" when "00111011010100111", -- t[30375] = 2
      "0000010" when "00111011010101000", -- t[30376] = 2
      "0000010" when "00111011010101001", -- t[30377] = 2
      "0000010" when "00111011010101010", -- t[30378] = 2
      "0000010" when "00111011010101011", -- t[30379] = 2
      "0000010" when "00111011010101100", -- t[30380] = 2
      "0000010" when "00111011010101101", -- t[30381] = 2
      "0000010" when "00111011010101110", -- t[30382] = 2
      "0000010" when "00111011010101111", -- t[30383] = 2
      "0000010" when "00111011010110000", -- t[30384] = 2
      "0000010" when "00111011010110001", -- t[30385] = 2
      "0000010" when "00111011010110010", -- t[30386] = 2
      "0000010" when "00111011010110011", -- t[30387] = 2
      "0000010" when "00111011010110100", -- t[30388] = 2
      "0000010" when "00111011010110101", -- t[30389] = 2
      "0000010" when "00111011010110110", -- t[30390] = 2
      "0000010" when "00111011010110111", -- t[30391] = 2
      "0000010" when "00111011010111000", -- t[30392] = 2
      "0000010" when "00111011010111001", -- t[30393] = 2
      "0000010" when "00111011010111010", -- t[30394] = 2
      "0000010" when "00111011010111011", -- t[30395] = 2
      "0000010" when "00111011010111100", -- t[30396] = 2
      "0000010" when "00111011010111101", -- t[30397] = 2
      "0000010" when "00111011010111110", -- t[30398] = 2
      "0000010" when "00111011010111111", -- t[30399] = 2
      "0000010" when "00111011011000000", -- t[30400] = 2
      "0000010" when "00111011011000001", -- t[30401] = 2
      "0000010" when "00111011011000010", -- t[30402] = 2
      "0000010" when "00111011011000011", -- t[30403] = 2
      "0000010" when "00111011011000100", -- t[30404] = 2
      "0000010" when "00111011011000101", -- t[30405] = 2
      "0000010" when "00111011011000110", -- t[30406] = 2
      "0000010" when "00111011011000111", -- t[30407] = 2
      "0000010" when "00111011011001000", -- t[30408] = 2
      "0000010" when "00111011011001001", -- t[30409] = 2
      "0000010" when "00111011011001010", -- t[30410] = 2
      "0000010" when "00111011011001011", -- t[30411] = 2
      "0000010" when "00111011011001100", -- t[30412] = 2
      "0000010" when "00111011011001101", -- t[30413] = 2
      "0000010" when "00111011011001110", -- t[30414] = 2
      "0000010" when "00111011011001111", -- t[30415] = 2
      "0000010" when "00111011011010000", -- t[30416] = 2
      "0000010" when "00111011011010001", -- t[30417] = 2
      "0000010" when "00111011011010010", -- t[30418] = 2
      "0000010" when "00111011011010011", -- t[30419] = 2
      "0000010" when "00111011011010100", -- t[30420] = 2
      "0000010" when "00111011011010101", -- t[30421] = 2
      "0000010" when "00111011011010110", -- t[30422] = 2
      "0000010" when "00111011011010111", -- t[30423] = 2
      "0000010" when "00111011011011000", -- t[30424] = 2
      "0000010" when "00111011011011001", -- t[30425] = 2
      "0000010" when "00111011011011010", -- t[30426] = 2
      "0000010" when "00111011011011011", -- t[30427] = 2
      "0000010" when "00111011011011100", -- t[30428] = 2
      "0000010" when "00111011011011101", -- t[30429] = 2
      "0000010" when "00111011011011110", -- t[30430] = 2
      "0000010" when "00111011011011111", -- t[30431] = 2
      "0000010" when "00111011011100000", -- t[30432] = 2
      "0000010" when "00111011011100001", -- t[30433] = 2
      "0000010" when "00111011011100010", -- t[30434] = 2
      "0000010" when "00111011011100011", -- t[30435] = 2
      "0000010" when "00111011011100100", -- t[30436] = 2
      "0000010" when "00111011011100101", -- t[30437] = 2
      "0000010" when "00111011011100110", -- t[30438] = 2
      "0000010" when "00111011011100111", -- t[30439] = 2
      "0000010" when "00111011011101000", -- t[30440] = 2
      "0000010" when "00111011011101001", -- t[30441] = 2
      "0000010" when "00111011011101010", -- t[30442] = 2
      "0000010" when "00111011011101011", -- t[30443] = 2
      "0000010" when "00111011011101100", -- t[30444] = 2
      "0000010" when "00111011011101101", -- t[30445] = 2
      "0000010" when "00111011011101110", -- t[30446] = 2
      "0000010" when "00111011011101111", -- t[30447] = 2
      "0000010" when "00111011011110000", -- t[30448] = 2
      "0000010" when "00111011011110001", -- t[30449] = 2
      "0000010" when "00111011011110010", -- t[30450] = 2
      "0000010" when "00111011011110011", -- t[30451] = 2
      "0000010" when "00111011011110100", -- t[30452] = 2
      "0000010" when "00111011011110101", -- t[30453] = 2
      "0000010" when "00111011011110110", -- t[30454] = 2
      "0000010" when "00111011011110111", -- t[30455] = 2
      "0000010" when "00111011011111000", -- t[30456] = 2
      "0000010" when "00111011011111001", -- t[30457] = 2
      "0000010" when "00111011011111010", -- t[30458] = 2
      "0000010" when "00111011011111011", -- t[30459] = 2
      "0000010" when "00111011011111100", -- t[30460] = 2
      "0000010" when "00111011011111101", -- t[30461] = 2
      "0000010" when "00111011011111110", -- t[30462] = 2
      "0000010" when "00111011011111111", -- t[30463] = 2
      "0000010" when "00111011100000000", -- t[30464] = 2
      "0000010" when "00111011100000001", -- t[30465] = 2
      "0000010" when "00111011100000010", -- t[30466] = 2
      "0000010" when "00111011100000011", -- t[30467] = 2
      "0000010" when "00111011100000100", -- t[30468] = 2
      "0000010" when "00111011100000101", -- t[30469] = 2
      "0000010" when "00111011100000110", -- t[30470] = 2
      "0000010" when "00111011100000111", -- t[30471] = 2
      "0000010" when "00111011100001000", -- t[30472] = 2
      "0000010" when "00111011100001001", -- t[30473] = 2
      "0000010" when "00111011100001010", -- t[30474] = 2
      "0000010" when "00111011100001011", -- t[30475] = 2
      "0000010" when "00111011100001100", -- t[30476] = 2
      "0000010" when "00111011100001101", -- t[30477] = 2
      "0000010" when "00111011100001110", -- t[30478] = 2
      "0000010" when "00111011100001111", -- t[30479] = 2
      "0000010" when "00111011100010000", -- t[30480] = 2
      "0000010" when "00111011100010001", -- t[30481] = 2
      "0000010" when "00111011100010010", -- t[30482] = 2
      "0000010" when "00111011100010011", -- t[30483] = 2
      "0000010" when "00111011100010100", -- t[30484] = 2
      "0000010" when "00111011100010101", -- t[30485] = 2
      "0000010" when "00111011100010110", -- t[30486] = 2
      "0000010" when "00111011100010111", -- t[30487] = 2
      "0000010" when "00111011100011000", -- t[30488] = 2
      "0000010" when "00111011100011001", -- t[30489] = 2
      "0000010" when "00111011100011010", -- t[30490] = 2
      "0000010" when "00111011100011011", -- t[30491] = 2
      "0000010" when "00111011100011100", -- t[30492] = 2
      "0000010" when "00111011100011101", -- t[30493] = 2
      "0000010" when "00111011100011110", -- t[30494] = 2
      "0000010" when "00111011100011111", -- t[30495] = 2
      "0000010" when "00111011100100000", -- t[30496] = 2
      "0000010" when "00111011100100001", -- t[30497] = 2
      "0000010" when "00111011100100010", -- t[30498] = 2
      "0000010" when "00111011100100011", -- t[30499] = 2
      "0000010" when "00111011100100100", -- t[30500] = 2
      "0000010" when "00111011100100101", -- t[30501] = 2
      "0000010" when "00111011100100110", -- t[30502] = 2
      "0000010" when "00111011100100111", -- t[30503] = 2
      "0000010" when "00111011100101000", -- t[30504] = 2
      "0000010" when "00111011100101001", -- t[30505] = 2
      "0000010" when "00111011100101010", -- t[30506] = 2
      "0000010" when "00111011100101011", -- t[30507] = 2
      "0000010" when "00111011100101100", -- t[30508] = 2
      "0000010" when "00111011100101101", -- t[30509] = 2
      "0000010" when "00111011100101110", -- t[30510] = 2
      "0000010" when "00111011100101111", -- t[30511] = 2
      "0000010" when "00111011100110000", -- t[30512] = 2
      "0000010" when "00111011100110001", -- t[30513] = 2
      "0000010" when "00111011100110010", -- t[30514] = 2
      "0000010" when "00111011100110011", -- t[30515] = 2
      "0000010" when "00111011100110100", -- t[30516] = 2
      "0000010" when "00111011100110101", -- t[30517] = 2
      "0000010" when "00111011100110110", -- t[30518] = 2
      "0000010" when "00111011100110111", -- t[30519] = 2
      "0000010" when "00111011100111000", -- t[30520] = 2
      "0000010" when "00111011100111001", -- t[30521] = 2
      "0000010" when "00111011100111010", -- t[30522] = 2
      "0000010" when "00111011100111011", -- t[30523] = 2
      "0000010" when "00111011100111100", -- t[30524] = 2
      "0000010" when "00111011100111101", -- t[30525] = 2
      "0000010" when "00111011100111110", -- t[30526] = 2
      "0000010" when "00111011100111111", -- t[30527] = 2
      "0000010" when "00111011101000000", -- t[30528] = 2
      "0000010" when "00111011101000001", -- t[30529] = 2
      "0000010" when "00111011101000010", -- t[30530] = 2
      "0000010" when "00111011101000011", -- t[30531] = 2
      "0000010" when "00111011101000100", -- t[30532] = 2
      "0000010" when "00111011101000101", -- t[30533] = 2
      "0000010" when "00111011101000110", -- t[30534] = 2
      "0000010" when "00111011101000111", -- t[30535] = 2
      "0000010" when "00111011101001000", -- t[30536] = 2
      "0000010" when "00111011101001001", -- t[30537] = 2
      "0000010" when "00111011101001010", -- t[30538] = 2
      "0000010" when "00111011101001011", -- t[30539] = 2
      "0000010" when "00111011101001100", -- t[30540] = 2
      "0000010" when "00111011101001101", -- t[30541] = 2
      "0000010" when "00111011101001110", -- t[30542] = 2
      "0000010" when "00111011101001111", -- t[30543] = 2
      "0000010" when "00111011101010000", -- t[30544] = 2
      "0000010" when "00111011101010001", -- t[30545] = 2
      "0000010" when "00111011101010010", -- t[30546] = 2
      "0000010" when "00111011101010011", -- t[30547] = 2
      "0000010" when "00111011101010100", -- t[30548] = 2
      "0000010" when "00111011101010101", -- t[30549] = 2
      "0000010" when "00111011101010110", -- t[30550] = 2
      "0000010" when "00111011101010111", -- t[30551] = 2
      "0000010" when "00111011101011000", -- t[30552] = 2
      "0000010" when "00111011101011001", -- t[30553] = 2
      "0000010" when "00111011101011010", -- t[30554] = 2
      "0000010" when "00111011101011011", -- t[30555] = 2
      "0000010" when "00111011101011100", -- t[30556] = 2
      "0000010" when "00111011101011101", -- t[30557] = 2
      "0000010" when "00111011101011110", -- t[30558] = 2
      "0000010" when "00111011101011111", -- t[30559] = 2
      "0000010" when "00111011101100000", -- t[30560] = 2
      "0000010" when "00111011101100001", -- t[30561] = 2
      "0000010" when "00111011101100010", -- t[30562] = 2
      "0000010" when "00111011101100011", -- t[30563] = 2
      "0000010" when "00111011101100100", -- t[30564] = 2
      "0000010" when "00111011101100101", -- t[30565] = 2
      "0000010" when "00111011101100110", -- t[30566] = 2
      "0000010" when "00111011101100111", -- t[30567] = 2
      "0000010" when "00111011101101000", -- t[30568] = 2
      "0000010" when "00111011101101001", -- t[30569] = 2
      "0000010" when "00111011101101010", -- t[30570] = 2
      "0000010" when "00111011101101011", -- t[30571] = 2
      "0000010" when "00111011101101100", -- t[30572] = 2
      "0000010" when "00111011101101101", -- t[30573] = 2
      "0000010" when "00111011101101110", -- t[30574] = 2
      "0000010" when "00111011101101111", -- t[30575] = 2
      "0000010" when "00111011101110000", -- t[30576] = 2
      "0000010" when "00111011101110001", -- t[30577] = 2
      "0000010" when "00111011101110010", -- t[30578] = 2
      "0000010" when "00111011101110011", -- t[30579] = 2
      "0000010" when "00111011101110100", -- t[30580] = 2
      "0000010" when "00111011101110101", -- t[30581] = 2
      "0000010" when "00111011101110110", -- t[30582] = 2
      "0000010" when "00111011101110111", -- t[30583] = 2
      "0000010" when "00111011101111000", -- t[30584] = 2
      "0000010" when "00111011101111001", -- t[30585] = 2
      "0000010" when "00111011101111010", -- t[30586] = 2
      "0000010" when "00111011101111011", -- t[30587] = 2
      "0000010" when "00111011101111100", -- t[30588] = 2
      "0000010" when "00111011101111101", -- t[30589] = 2
      "0000010" when "00111011101111110", -- t[30590] = 2
      "0000010" when "00111011101111111", -- t[30591] = 2
      "0000010" when "00111011110000000", -- t[30592] = 2
      "0000010" when "00111011110000001", -- t[30593] = 2
      "0000010" when "00111011110000010", -- t[30594] = 2
      "0000010" when "00111011110000011", -- t[30595] = 2
      "0000010" when "00111011110000100", -- t[30596] = 2
      "0000010" when "00111011110000101", -- t[30597] = 2
      "0000010" when "00111011110000110", -- t[30598] = 2
      "0000010" when "00111011110000111", -- t[30599] = 2
      "0000010" when "00111011110001000", -- t[30600] = 2
      "0000010" when "00111011110001001", -- t[30601] = 2
      "0000010" when "00111011110001010", -- t[30602] = 2
      "0000010" when "00111011110001011", -- t[30603] = 2
      "0000010" when "00111011110001100", -- t[30604] = 2
      "0000010" when "00111011110001101", -- t[30605] = 2
      "0000010" when "00111011110001110", -- t[30606] = 2
      "0000010" when "00111011110001111", -- t[30607] = 2
      "0000010" when "00111011110010000", -- t[30608] = 2
      "0000010" when "00111011110010001", -- t[30609] = 2
      "0000010" when "00111011110010010", -- t[30610] = 2
      "0000010" when "00111011110010011", -- t[30611] = 2
      "0000010" when "00111011110010100", -- t[30612] = 2
      "0000010" when "00111011110010101", -- t[30613] = 2
      "0000010" when "00111011110010110", -- t[30614] = 2
      "0000010" when "00111011110010111", -- t[30615] = 2
      "0000010" when "00111011110011000", -- t[30616] = 2
      "0000010" when "00111011110011001", -- t[30617] = 2
      "0000010" when "00111011110011010", -- t[30618] = 2
      "0000010" when "00111011110011011", -- t[30619] = 2
      "0000010" when "00111011110011100", -- t[30620] = 2
      "0000010" when "00111011110011101", -- t[30621] = 2
      "0000010" when "00111011110011110", -- t[30622] = 2
      "0000010" when "00111011110011111", -- t[30623] = 2
      "0000010" when "00111011110100000", -- t[30624] = 2
      "0000010" when "00111011110100001", -- t[30625] = 2
      "0000010" when "00111011110100010", -- t[30626] = 2
      "0000010" when "00111011110100011", -- t[30627] = 2
      "0000010" when "00111011110100100", -- t[30628] = 2
      "0000010" when "00111011110100101", -- t[30629] = 2
      "0000010" when "00111011110100110", -- t[30630] = 2
      "0000010" when "00111011110100111", -- t[30631] = 2
      "0000010" when "00111011110101000", -- t[30632] = 2
      "0000010" when "00111011110101001", -- t[30633] = 2
      "0000010" when "00111011110101010", -- t[30634] = 2
      "0000010" when "00111011110101011", -- t[30635] = 2
      "0000010" when "00111011110101100", -- t[30636] = 2
      "0000010" when "00111011110101101", -- t[30637] = 2
      "0000010" when "00111011110101110", -- t[30638] = 2
      "0000010" when "00111011110101111", -- t[30639] = 2
      "0000010" when "00111011110110000", -- t[30640] = 2
      "0000010" when "00111011110110001", -- t[30641] = 2
      "0000010" when "00111011110110010", -- t[30642] = 2
      "0000010" when "00111011110110011", -- t[30643] = 2
      "0000010" when "00111011110110100", -- t[30644] = 2
      "0000010" when "00111011110110101", -- t[30645] = 2
      "0000010" when "00111011110110110", -- t[30646] = 2
      "0000010" when "00111011110110111", -- t[30647] = 2
      "0000010" when "00111011110111000", -- t[30648] = 2
      "0000010" when "00111011110111001", -- t[30649] = 2
      "0000010" when "00111011110111010", -- t[30650] = 2
      "0000010" when "00111011110111011", -- t[30651] = 2
      "0000010" when "00111011110111100", -- t[30652] = 2
      "0000010" when "00111011110111101", -- t[30653] = 2
      "0000010" when "00111011110111110", -- t[30654] = 2
      "0000010" when "00111011110111111", -- t[30655] = 2
      "0000010" when "00111011111000000", -- t[30656] = 2
      "0000010" when "00111011111000001", -- t[30657] = 2
      "0000010" when "00111011111000010", -- t[30658] = 2
      "0000010" when "00111011111000011", -- t[30659] = 2
      "0000010" when "00111011111000100", -- t[30660] = 2
      "0000010" when "00111011111000101", -- t[30661] = 2
      "0000010" when "00111011111000110", -- t[30662] = 2
      "0000010" when "00111011111000111", -- t[30663] = 2
      "0000010" when "00111011111001000", -- t[30664] = 2
      "0000010" when "00111011111001001", -- t[30665] = 2
      "0000010" when "00111011111001010", -- t[30666] = 2
      "0000010" when "00111011111001011", -- t[30667] = 2
      "0000010" when "00111011111001100", -- t[30668] = 2
      "0000010" when "00111011111001101", -- t[30669] = 2
      "0000010" when "00111011111001110", -- t[30670] = 2
      "0000010" when "00111011111001111", -- t[30671] = 2
      "0000010" when "00111011111010000", -- t[30672] = 2
      "0000010" when "00111011111010001", -- t[30673] = 2
      "0000010" when "00111011111010010", -- t[30674] = 2
      "0000010" when "00111011111010011", -- t[30675] = 2
      "0000010" when "00111011111010100", -- t[30676] = 2
      "0000010" when "00111011111010101", -- t[30677] = 2
      "0000010" when "00111011111010110", -- t[30678] = 2
      "0000010" when "00111011111010111", -- t[30679] = 2
      "0000010" when "00111011111011000", -- t[30680] = 2
      "0000010" when "00111011111011001", -- t[30681] = 2
      "0000010" when "00111011111011010", -- t[30682] = 2
      "0000010" when "00111011111011011", -- t[30683] = 2
      "0000010" when "00111011111011100", -- t[30684] = 2
      "0000010" when "00111011111011101", -- t[30685] = 2
      "0000010" when "00111011111011110", -- t[30686] = 2
      "0000010" when "00111011111011111", -- t[30687] = 2
      "0000010" when "00111011111100000", -- t[30688] = 2
      "0000010" when "00111011111100001", -- t[30689] = 2
      "0000010" when "00111011111100010", -- t[30690] = 2
      "0000010" when "00111011111100011", -- t[30691] = 2
      "0000010" when "00111011111100100", -- t[30692] = 2
      "0000010" when "00111011111100101", -- t[30693] = 2
      "0000010" when "00111011111100110", -- t[30694] = 2
      "0000010" when "00111011111100111", -- t[30695] = 2
      "0000010" when "00111011111101000", -- t[30696] = 2
      "0000010" when "00111011111101001", -- t[30697] = 2
      "0000010" when "00111011111101010", -- t[30698] = 2
      "0000010" when "00111011111101011", -- t[30699] = 2
      "0000010" when "00111011111101100", -- t[30700] = 2
      "0000010" when "00111011111101101", -- t[30701] = 2
      "0000010" when "00111011111101110", -- t[30702] = 2
      "0000010" when "00111011111101111", -- t[30703] = 2
      "0000010" when "00111011111110000", -- t[30704] = 2
      "0000010" when "00111011111110001", -- t[30705] = 2
      "0000010" when "00111011111110010", -- t[30706] = 2
      "0000010" when "00111011111110011", -- t[30707] = 2
      "0000010" when "00111011111110100", -- t[30708] = 2
      "0000010" when "00111011111110101", -- t[30709] = 2
      "0000010" when "00111011111110110", -- t[30710] = 2
      "0000010" when "00111011111110111", -- t[30711] = 2
      "0000010" when "00111011111111000", -- t[30712] = 2
      "0000010" when "00111011111111001", -- t[30713] = 2
      "0000010" when "00111011111111010", -- t[30714] = 2
      "0000010" when "00111011111111011", -- t[30715] = 2
      "0000010" when "00111011111111100", -- t[30716] = 2
      "0000010" when "00111011111111101", -- t[30717] = 2
      "0000010" when "00111011111111110", -- t[30718] = 2
      "0000010" when "00111011111111111", -- t[30719] = 2
      "0000010" when "00111100000000000", -- t[30720] = 2
      "0000010" when "00111100000000001", -- t[30721] = 2
      "0000010" when "00111100000000010", -- t[30722] = 2
      "0000010" when "00111100000000011", -- t[30723] = 2
      "0000010" when "00111100000000100", -- t[30724] = 2
      "0000010" when "00111100000000101", -- t[30725] = 2
      "0000010" when "00111100000000110", -- t[30726] = 2
      "0000010" when "00111100000000111", -- t[30727] = 2
      "0000010" when "00111100000001000", -- t[30728] = 2
      "0000010" when "00111100000001001", -- t[30729] = 2
      "0000010" when "00111100000001010", -- t[30730] = 2
      "0000010" when "00111100000001011", -- t[30731] = 2
      "0000010" when "00111100000001100", -- t[30732] = 2
      "0000010" when "00111100000001101", -- t[30733] = 2
      "0000010" when "00111100000001110", -- t[30734] = 2
      "0000010" when "00111100000001111", -- t[30735] = 2
      "0000010" when "00111100000010000", -- t[30736] = 2
      "0000010" when "00111100000010001", -- t[30737] = 2
      "0000010" when "00111100000010010", -- t[30738] = 2
      "0000010" when "00111100000010011", -- t[30739] = 2
      "0000010" when "00111100000010100", -- t[30740] = 2
      "0000010" when "00111100000010101", -- t[30741] = 2
      "0000010" when "00111100000010110", -- t[30742] = 2
      "0000010" when "00111100000010111", -- t[30743] = 2
      "0000010" when "00111100000011000", -- t[30744] = 2
      "0000010" when "00111100000011001", -- t[30745] = 2
      "0000010" when "00111100000011010", -- t[30746] = 2
      "0000010" when "00111100000011011", -- t[30747] = 2
      "0000010" when "00111100000011100", -- t[30748] = 2
      "0000010" when "00111100000011101", -- t[30749] = 2
      "0000010" when "00111100000011110", -- t[30750] = 2
      "0000010" when "00111100000011111", -- t[30751] = 2
      "0000010" when "00111100000100000", -- t[30752] = 2
      "0000010" when "00111100000100001", -- t[30753] = 2
      "0000010" when "00111100000100010", -- t[30754] = 2
      "0000010" when "00111100000100011", -- t[30755] = 2
      "0000010" when "00111100000100100", -- t[30756] = 2
      "0000010" when "00111100000100101", -- t[30757] = 2
      "0000010" when "00111100000100110", -- t[30758] = 2
      "0000010" when "00111100000100111", -- t[30759] = 2
      "0000010" when "00111100000101000", -- t[30760] = 2
      "0000010" when "00111100000101001", -- t[30761] = 2
      "0000010" when "00111100000101010", -- t[30762] = 2
      "0000010" when "00111100000101011", -- t[30763] = 2
      "0000010" when "00111100000101100", -- t[30764] = 2
      "0000010" when "00111100000101101", -- t[30765] = 2
      "0000010" when "00111100000101110", -- t[30766] = 2
      "0000010" when "00111100000101111", -- t[30767] = 2
      "0000010" when "00111100000110000", -- t[30768] = 2
      "0000010" when "00111100000110001", -- t[30769] = 2
      "0000010" when "00111100000110010", -- t[30770] = 2
      "0000010" when "00111100000110011", -- t[30771] = 2
      "0000010" when "00111100000110100", -- t[30772] = 2
      "0000010" when "00111100000110101", -- t[30773] = 2
      "0000010" when "00111100000110110", -- t[30774] = 2
      "0000010" when "00111100000110111", -- t[30775] = 2
      "0000010" when "00111100000111000", -- t[30776] = 2
      "0000010" when "00111100000111001", -- t[30777] = 2
      "0000010" when "00111100000111010", -- t[30778] = 2
      "0000010" when "00111100000111011", -- t[30779] = 2
      "0000010" when "00111100000111100", -- t[30780] = 2
      "0000010" when "00111100000111101", -- t[30781] = 2
      "0000010" when "00111100000111110", -- t[30782] = 2
      "0000010" when "00111100000111111", -- t[30783] = 2
      "0000010" when "00111100001000000", -- t[30784] = 2
      "0000010" when "00111100001000001", -- t[30785] = 2
      "0000010" when "00111100001000010", -- t[30786] = 2
      "0000010" when "00111100001000011", -- t[30787] = 2
      "0000010" when "00111100001000100", -- t[30788] = 2
      "0000010" when "00111100001000101", -- t[30789] = 2
      "0000010" when "00111100001000110", -- t[30790] = 2
      "0000010" when "00111100001000111", -- t[30791] = 2
      "0000010" when "00111100001001000", -- t[30792] = 2
      "0000010" when "00111100001001001", -- t[30793] = 2
      "0000010" when "00111100001001010", -- t[30794] = 2
      "0000010" when "00111100001001011", -- t[30795] = 2
      "0000010" when "00111100001001100", -- t[30796] = 2
      "0000010" when "00111100001001101", -- t[30797] = 2
      "0000010" when "00111100001001110", -- t[30798] = 2
      "0000010" when "00111100001001111", -- t[30799] = 2
      "0000010" when "00111100001010000", -- t[30800] = 2
      "0000010" when "00111100001010001", -- t[30801] = 2
      "0000010" when "00111100001010010", -- t[30802] = 2
      "0000010" when "00111100001010011", -- t[30803] = 2
      "0000010" when "00111100001010100", -- t[30804] = 2
      "0000010" when "00111100001010101", -- t[30805] = 2
      "0000010" when "00111100001010110", -- t[30806] = 2
      "0000010" when "00111100001010111", -- t[30807] = 2
      "0000010" when "00111100001011000", -- t[30808] = 2
      "0000010" when "00111100001011001", -- t[30809] = 2
      "0000010" when "00111100001011010", -- t[30810] = 2
      "0000010" when "00111100001011011", -- t[30811] = 2
      "0000010" when "00111100001011100", -- t[30812] = 2
      "0000010" when "00111100001011101", -- t[30813] = 2
      "0000010" when "00111100001011110", -- t[30814] = 2
      "0000010" when "00111100001011111", -- t[30815] = 2
      "0000010" when "00111100001100000", -- t[30816] = 2
      "0000010" when "00111100001100001", -- t[30817] = 2
      "0000010" when "00111100001100010", -- t[30818] = 2
      "0000010" when "00111100001100011", -- t[30819] = 2
      "0000010" when "00111100001100100", -- t[30820] = 2
      "0000010" when "00111100001100101", -- t[30821] = 2
      "0000010" when "00111100001100110", -- t[30822] = 2
      "0000010" when "00111100001100111", -- t[30823] = 2
      "0000010" when "00111100001101000", -- t[30824] = 2
      "0000010" when "00111100001101001", -- t[30825] = 2
      "0000010" when "00111100001101010", -- t[30826] = 2
      "0000010" when "00111100001101011", -- t[30827] = 2
      "0000010" when "00111100001101100", -- t[30828] = 2
      "0000010" when "00111100001101101", -- t[30829] = 2
      "0000010" when "00111100001101110", -- t[30830] = 2
      "0000010" when "00111100001101111", -- t[30831] = 2
      "0000010" when "00111100001110000", -- t[30832] = 2
      "0000010" when "00111100001110001", -- t[30833] = 2
      "0000010" when "00111100001110010", -- t[30834] = 2
      "0000010" when "00111100001110011", -- t[30835] = 2
      "0000010" when "00111100001110100", -- t[30836] = 2
      "0000010" when "00111100001110101", -- t[30837] = 2
      "0000010" when "00111100001110110", -- t[30838] = 2
      "0000010" when "00111100001110111", -- t[30839] = 2
      "0000010" when "00111100001111000", -- t[30840] = 2
      "0000010" when "00111100001111001", -- t[30841] = 2
      "0000010" when "00111100001111010", -- t[30842] = 2
      "0000010" when "00111100001111011", -- t[30843] = 2
      "0000010" when "00111100001111100", -- t[30844] = 2
      "0000010" when "00111100001111101", -- t[30845] = 2
      "0000010" when "00111100001111110", -- t[30846] = 2
      "0000010" when "00111100001111111", -- t[30847] = 2
      "0000010" when "00111100010000000", -- t[30848] = 2
      "0000010" when "00111100010000001", -- t[30849] = 2
      "0000010" when "00111100010000010", -- t[30850] = 2
      "0000010" when "00111100010000011", -- t[30851] = 2
      "0000010" when "00111100010000100", -- t[30852] = 2
      "0000010" when "00111100010000101", -- t[30853] = 2
      "0000010" when "00111100010000110", -- t[30854] = 2
      "0000010" when "00111100010000111", -- t[30855] = 2
      "0000010" when "00111100010001000", -- t[30856] = 2
      "0000010" when "00111100010001001", -- t[30857] = 2
      "0000010" when "00111100010001010", -- t[30858] = 2
      "0000010" when "00111100010001011", -- t[30859] = 2
      "0000010" when "00111100010001100", -- t[30860] = 2
      "0000010" when "00111100010001101", -- t[30861] = 2
      "0000010" when "00111100010001110", -- t[30862] = 2
      "0000010" when "00111100010001111", -- t[30863] = 2
      "0000010" when "00111100010010000", -- t[30864] = 2
      "0000010" when "00111100010010001", -- t[30865] = 2
      "0000010" when "00111100010010010", -- t[30866] = 2
      "0000010" when "00111100010010011", -- t[30867] = 2
      "0000010" when "00111100010010100", -- t[30868] = 2
      "0000010" when "00111100010010101", -- t[30869] = 2
      "0000010" when "00111100010010110", -- t[30870] = 2
      "0000010" when "00111100010010111", -- t[30871] = 2
      "0000010" when "00111100010011000", -- t[30872] = 2
      "0000010" when "00111100010011001", -- t[30873] = 2
      "0000010" when "00111100010011010", -- t[30874] = 2
      "0000010" when "00111100010011011", -- t[30875] = 2
      "0000010" when "00111100010011100", -- t[30876] = 2
      "0000010" when "00111100010011101", -- t[30877] = 2
      "0000010" when "00111100010011110", -- t[30878] = 2
      "0000010" when "00111100010011111", -- t[30879] = 2
      "0000010" when "00111100010100000", -- t[30880] = 2
      "0000010" when "00111100010100001", -- t[30881] = 2
      "0000010" when "00111100010100010", -- t[30882] = 2
      "0000010" when "00111100010100011", -- t[30883] = 2
      "0000010" when "00111100010100100", -- t[30884] = 2
      "0000010" when "00111100010100101", -- t[30885] = 2
      "0000010" when "00111100010100110", -- t[30886] = 2
      "0000010" when "00111100010100111", -- t[30887] = 2
      "0000010" when "00111100010101000", -- t[30888] = 2
      "0000010" when "00111100010101001", -- t[30889] = 2
      "0000010" when "00111100010101010", -- t[30890] = 2
      "0000010" when "00111100010101011", -- t[30891] = 2
      "0000010" when "00111100010101100", -- t[30892] = 2
      "0000010" when "00111100010101101", -- t[30893] = 2
      "0000010" when "00111100010101110", -- t[30894] = 2
      "0000010" when "00111100010101111", -- t[30895] = 2
      "0000010" when "00111100010110000", -- t[30896] = 2
      "0000010" when "00111100010110001", -- t[30897] = 2
      "0000010" when "00111100010110010", -- t[30898] = 2
      "0000010" when "00111100010110011", -- t[30899] = 2
      "0000010" when "00111100010110100", -- t[30900] = 2
      "0000010" when "00111100010110101", -- t[30901] = 2
      "0000010" when "00111100010110110", -- t[30902] = 2
      "0000010" when "00111100010110111", -- t[30903] = 2
      "0000010" when "00111100010111000", -- t[30904] = 2
      "0000010" when "00111100010111001", -- t[30905] = 2
      "0000010" when "00111100010111010", -- t[30906] = 2
      "0000010" when "00111100010111011", -- t[30907] = 2
      "0000010" when "00111100010111100", -- t[30908] = 2
      "0000010" when "00111100010111101", -- t[30909] = 2
      "0000010" when "00111100010111110", -- t[30910] = 2
      "0000010" when "00111100010111111", -- t[30911] = 2
      "0000010" when "00111100011000000", -- t[30912] = 2
      "0000010" when "00111100011000001", -- t[30913] = 2
      "0000010" when "00111100011000010", -- t[30914] = 2
      "0000010" when "00111100011000011", -- t[30915] = 2
      "0000010" when "00111100011000100", -- t[30916] = 2
      "0000010" when "00111100011000101", -- t[30917] = 2
      "0000010" when "00111100011000110", -- t[30918] = 2
      "0000010" when "00111100011000111", -- t[30919] = 2
      "0000010" when "00111100011001000", -- t[30920] = 2
      "0000010" when "00111100011001001", -- t[30921] = 2
      "0000010" when "00111100011001010", -- t[30922] = 2
      "0000010" when "00111100011001011", -- t[30923] = 2
      "0000010" when "00111100011001100", -- t[30924] = 2
      "0000010" when "00111100011001101", -- t[30925] = 2
      "0000010" when "00111100011001110", -- t[30926] = 2
      "0000010" when "00111100011001111", -- t[30927] = 2
      "0000010" when "00111100011010000", -- t[30928] = 2
      "0000010" when "00111100011010001", -- t[30929] = 2
      "0000010" when "00111100011010010", -- t[30930] = 2
      "0000010" when "00111100011010011", -- t[30931] = 2
      "0000010" when "00111100011010100", -- t[30932] = 2
      "0000010" when "00111100011010101", -- t[30933] = 2
      "0000010" when "00111100011010110", -- t[30934] = 2
      "0000010" when "00111100011010111", -- t[30935] = 2
      "0000010" when "00111100011011000", -- t[30936] = 2
      "0000010" when "00111100011011001", -- t[30937] = 2
      "0000010" when "00111100011011010", -- t[30938] = 2
      "0000010" when "00111100011011011", -- t[30939] = 2
      "0000010" when "00111100011011100", -- t[30940] = 2
      "0000010" when "00111100011011101", -- t[30941] = 2
      "0000010" when "00111100011011110", -- t[30942] = 2
      "0000010" when "00111100011011111", -- t[30943] = 2
      "0000010" when "00111100011100000", -- t[30944] = 2
      "0000010" when "00111100011100001", -- t[30945] = 2
      "0000010" when "00111100011100010", -- t[30946] = 2
      "0000010" when "00111100011100011", -- t[30947] = 2
      "0000010" when "00111100011100100", -- t[30948] = 2
      "0000010" when "00111100011100101", -- t[30949] = 2
      "0000010" when "00111100011100110", -- t[30950] = 2
      "0000010" when "00111100011100111", -- t[30951] = 2
      "0000010" when "00111100011101000", -- t[30952] = 2
      "0000010" when "00111100011101001", -- t[30953] = 2
      "0000010" when "00111100011101010", -- t[30954] = 2
      "0000010" when "00111100011101011", -- t[30955] = 2
      "0000010" when "00111100011101100", -- t[30956] = 2
      "0000010" when "00111100011101101", -- t[30957] = 2
      "0000010" when "00111100011101110", -- t[30958] = 2
      "0000010" when "00111100011101111", -- t[30959] = 2
      "0000010" when "00111100011110000", -- t[30960] = 2
      "0000010" when "00111100011110001", -- t[30961] = 2
      "0000010" when "00111100011110010", -- t[30962] = 2
      "0000010" when "00111100011110011", -- t[30963] = 2
      "0000010" when "00111100011110100", -- t[30964] = 2
      "0000010" when "00111100011110101", -- t[30965] = 2
      "0000010" when "00111100011110110", -- t[30966] = 2
      "0000010" when "00111100011110111", -- t[30967] = 2
      "0000010" when "00111100011111000", -- t[30968] = 2
      "0000010" when "00111100011111001", -- t[30969] = 2
      "0000010" when "00111100011111010", -- t[30970] = 2
      "0000010" when "00111100011111011", -- t[30971] = 2
      "0000010" when "00111100011111100", -- t[30972] = 2
      "0000010" when "00111100011111101", -- t[30973] = 2
      "0000010" when "00111100011111110", -- t[30974] = 2
      "0000010" when "00111100011111111", -- t[30975] = 2
      "0000010" when "00111100100000000", -- t[30976] = 2
      "0000010" when "00111100100000001", -- t[30977] = 2
      "0000010" when "00111100100000010", -- t[30978] = 2
      "0000010" when "00111100100000011", -- t[30979] = 2
      "0000010" when "00111100100000100", -- t[30980] = 2
      "0000010" when "00111100100000101", -- t[30981] = 2
      "0000010" when "00111100100000110", -- t[30982] = 2
      "0000010" when "00111100100000111", -- t[30983] = 2
      "0000010" when "00111100100001000", -- t[30984] = 2
      "0000010" when "00111100100001001", -- t[30985] = 2
      "0000010" when "00111100100001010", -- t[30986] = 2
      "0000010" when "00111100100001011", -- t[30987] = 2
      "0000010" when "00111100100001100", -- t[30988] = 2
      "0000010" when "00111100100001101", -- t[30989] = 2
      "0000010" when "00111100100001110", -- t[30990] = 2
      "0000010" when "00111100100001111", -- t[30991] = 2
      "0000010" when "00111100100010000", -- t[30992] = 2
      "0000010" when "00111100100010001", -- t[30993] = 2
      "0000010" when "00111100100010010", -- t[30994] = 2
      "0000010" when "00111100100010011", -- t[30995] = 2
      "0000010" when "00111100100010100", -- t[30996] = 2
      "0000010" when "00111100100010101", -- t[30997] = 2
      "0000010" when "00111100100010110", -- t[30998] = 2
      "0000010" when "00111100100010111", -- t[30999] = 2
      "0000010" when "00111100100011000", -- t[31000] = 2
      "0000010" when "00111100100011001", -- t[31001] = 2
      "0000010" when "00111100100011010", -- t[31002] = 2
      "0000010" when "00111100100011011", -- t[31003] = 2
      "0000010" when "00111100100011100", -- t[31004] = 2
      "0000010" when "00111100100011101", -- t[31005] = 2
      "0000010" when "00111100100011110", -- t[31006] = 2
      "0000010" when "00111100100011111", -- t[31007] = 2
      "0000010" when "00111100100100000", -- t[31008] = 2
      "0000010" when "00111100100100001", -- t[31009] = 2
      "0000010" when "00111100100100010", -- t[31010] = 2
      "0000010" when "00111100100100011", -- t[31011] = 2
      "0000010" when "00111100100100100", -- t[31012] = 2
      "0000010" when "00111100100100101", -- t[31013] = 2
      "0000010" when "00111100100100110", -- t[31014] = 2
      "0000010" when "00111100100100111", -- t[31015] = 2
      "0000010" when "00111100100101000", -- t[31016] = 2
      "0000010" when "00111100100101001", -- t[31017] = 2
      "0000010" when "00111100100101010", -- t[31018] = 2
      "0000010" when "00111100100101011", -- t[31019] = 2
      "0000010" when "00111100100101100", -- t[31020] = 2
      "0000010" when "00111100100101101", -- t[31021] = 2
      "0000010" when "00111100100101110", -- t[31022] = 2
      "0000010" when "00111100100101111", -- t[31023] = 2
      "0000010" when "00111100100110000", -- t[31024] = 2
      "0000010" when "00111100100110001", -- t[31025] = 2
      "0000010" when "00111100100110010", -- t[31026] = 2
      "0000010" when "00111100100110011", -- t[31027] = 2
      "0000010" when "00111100100110100", -- t[31028] = 2
      "0000010" when "00111100100110101", -- t[31029] = 2
      "0000010" when "00111100100110110", -- t[31030] = 2
      "0000010" when "00111100100110111", -- t[31031] = 2
      "0000010" when "00111100100111000", -- t[31032] = 2
      "0000010" when "00111100100111001", -- t[31033] = 2
      "0000010" when "00111100100111010", -- t[31034] = 2
      "0000010" when "00111100100111011", -- t[31035] = 2
      "0000010" when "00111100100111100", -- t[31036] = 2
      "0000010" when "00111100100111101", -- t[31037] = 2
      "0000010" when "00111100100111110", -- t[31038] = 2
      "0000010" when "00111100100111111", -- t[31039] = 2
      "0000010" when "00111100101000000", -- t[31040] = 2
      "0000010" when "00111100101000001", -- t[31041] = 2
      "0000010" when "00111100101000010", -- t[31042] = 2
      "0000010" when "00111100101000011", -- t[31043] = 2
      "0000010" when "00111100101000100", -- t[31044] = 2
      "0000010" when "00111100101000101", -- t[31045] = 2
      "0000010" when "00111100101000110", -- t[31046] = 2
      "0000010" when "00111100101000111", -- t[31047] = 2
      "0000010" when "00111100101001000", -- t[31048] = 2
      "0000010" when "00111100101001001", -- t[31049] = 2
      "0000010" when "00111100101001010", -- t[31050] = 2
      "0000010" when "00111100101001011", -- t[31051] = 2
      "0000010" when "00111100101001100", -- t[31052] = 2
      "0000010" when "00111100101001101", -- t[31053] = 2
      "0000010" when "00111100101001110", -- t[31054] = 2
      "0000010" when "00111100101001111", -- t[31055] = 2
      "0000010" when "00111100101010000", -- t[31056] = 2
      "0000010" when "00111100101010001", -- t[31057] = 2
      "0000010" when "00111100101010010", -- t[31058] = 2
      "0000010" when "00111100101010011", -- t[31059] = 2
      "0000010" when "00111100101010100", -- t[31060] = 2
      "0000010" when "00111100101010101", -- t[31061] = 2
      "0000010" when "00111100101010110", -- t[31062] = 2
      "0000010" when "00111100101010111", -- t[31063] = 2
      "0000010" when "00111100101011000", -- t[31064] = 2
      "0000010" when "00111100101011001", -- t[31065] = 2
      "0000010" when "00111100101011010", -- t[31066] = 2
      "0000010" when "00111100101011011", -- t[31067] = 2
      "0000010" when "00111100101011100", -- t[31068] = 2
      "0000010" when "00111100101011101", -- t[31069] = 2
      "0000010" when "00111100101011110", -- t[31070] = 2
      "0000010" when "00111100101011111", -- t[31071] = 2
      "0000010" when "00111100101100000", -- t[31072] = 2
      "0000011" when "00111100101100001", -- t[31073] = 3
      "0000011" when "00111100101100010", -- t[31074] = 3
      "0000011" when "00111100101100011", -- t[31075] = 3
      "0000011" when "00111100101100100", -- t[31076] = 3
      "0000011" when "00111100101100101", -- t[31077] = 3
      "0000011" when "00111100101100110", -- t[31078] = 3
      "0000011" when "00111100101100111", -- t[31079] = 3
      "0000011" when "00111100101101000", -- t[31080] = 3
      "0000011" when "00111100101101001", -- t[31081] = 3
      "0000011" when "00111100101101010", -- t[31082] = 3
      "0000011" when "00111100101101011", -- t[31083] = 3
      "0000011" when "00111100101101100", -- t[31084] = 3
      "0000011" when "00111100101101101", -- t[31085] = 3
      "0000011" when "00111100101101110", -- t[31086] = 3
      "0000011" when "00111100101101111", -- t[31087] = 3
      "0000011" when "00111100101110000", -- t[31088] = 3
      "0000011" when "00111100101110001", -- t[31089] = 3
      "0000011" when "00111100101110010", -- t[31090] = 3
      "0000011" when "00111100101110011", -- t[31091] = 3
      "0000011" when "00111100101110100", -- t[31092] = 3
      "0000011" when "00111100101110101", -- t[31093] = 3
      "0000011" when "00111100101110110", -- t[31094] = 3
      "0000011" when "00111100101110111", -- t[31095] = 3
      "0000011" when "00111100101111000", -- t[31096] = 3
      "0000011" when "00111100101111001", -- t[31097] = 3
      "0000011" when "00111100101111010", -- t[31098] = 3
      "0000011" when "00111100101111011", -- t[31099] = 3
      "0000011" when "00111100101111100", -- t[31100] = 3
      "0000011" when "00111100101111101", -- t[31101] = 3
      "0000011" when "00111100101111110", -- t[31102] = 3
      "0000011" when "00111100101111111", -- t[31103] = 3
      "0000011" when "00111100110000000", -- t[31104] = 3
      "0000011" when "00111100110000001", -- t[31105] = 3
      "0000011" when "00111100110000010", -- t[31106] = 3
      "0000011" when "00111100110000011", -- t[31107] = 3
      "0000011" when "00111100110000100", -- t[31108] = 3
      "0000011" when "00111100110000101", -- t[31109] = 3
      "0000011" when "00111100110000110", -- t[31110] = 3
      "0000011" when "00111100110000111", -- t[31111] = 3
      "0000011" when "00111100110001000", -- t[31112] = 3
      "0000011" when "00111100110001001", -- t[31113] = 3
      "0000011" when "00111100110001010", -- t[31114] = 3
      "0000011" when "00111100110001011", -- t[31115] = 3
      "0000011" when "00111100110001100", -- t[31116] = 3
      "0000011" when "00111100110001101", -- t[31117] = 3
      "0000011" when "00111100110001110", -- t[31118] = 3
      "0000011" when "00111100110001111", -- t[31119] = 3
      "0000011" when "00111100110010000", -- t[31120] = 3
      "0000011" when "00111100110010001", -- t[31121] = 3
      "0000011" when "00111100110010010", -- t[31122] = 3
      "0000011" when "00111100110010011", -- t[31123] = 3
      "0000011" when "00111100110010100", -- t[31124] = 3
      "0000011" when "00111100110010101", -- t[31125] = 3
      "0000011" when "00111100110010110", -- t[31126] = 3
      "0000011" when "00111100110010111", -- t[31127] = 3
      "0000011" when "00111100110011000", -- t[31128] = 3
      "0000011" when "00111100110011001", -- t[31129] = 3
      "0000011" when "00111100110011010", -- t[31130] = 3
      "0000011" when "00111100110011011", -- t[31131] = 3
      "0000011" when "00111100110011100", -- t[31132] = 3
      "0000011" when "00111100110011101", -- t[31133] = 3
      "0000011" when "00111100110011110", -- t[31134] = 3
      "0000011" when "00111100110011111", -- t[31135] = 3
      "0000011" when "00111100110100000", -- t[31136] = 3
      "0000011" when "00111100110100001", -- t[31137] = 3
      "0000011" when "00111100110100010", -- t[31138] = 3
      "0000011" when "00111100110100011", -- t[31139] = 3
      "0000011" when "00111100110100100", -- t[31140] = 3
      "0000011" when "00111100110100101", -- t[31141] = 3
      "0000011" when "00111100110100110", -- t[31142] = 3
      "0000011" when "00111100110100111", -- t[31143] = 3
      "0000011" when "00111100110101000", -- t[31144] = 3
      "0000011" when "00111100110101001", -- t[31145] = 3
      "0000011" when "00111100110101010", -- t[31146] = 3
      "0000011" when "00111100110101011", -- t[31147] = 3
      "0000011" when "00111100110101100", -- t[31148] = 3
      "0000011" when "00111100110101101", -- t[31149] = 3
      "0000011" when "00111100110101110", -- t[31150] = 3
      "0000011" when "00111100110101111", -- t[31151] = 3
      "0000011" when "00111100110110000", -- t[31152] = 3
      "0000011" when "00111100110110001", -- t[31153] = 3
      "0000011" when "00111100110110010", -- t[31154] = 3
      "0000011" when "00111100110110011", -- t[31155] = 3
      "0000011" when "00111100110110100", -- t[31156] = 3
      "0000011" when "00111100110110101", -- t[31157] = 3
      "0000011" when "00111100110110110", -- t[31158] = 3
      "0000011" when "00111100110110111", -- t[31159] = 3
      "0000011" when "00111100110111000", -- t[31160] = 3
      "0000011" when "00111100110111001", -- t[31161] = 3
      "0000011" when "00111100110111010", -- t[31162] = 3
      "0000011" when "00111100110111011", -- t[31163] = 3
      "0000011" when "00111100110111100", -- t[31164] = 3
      "0000011" when "00111100110111101", -- t[31165] = 3
      "0000011" when "00111100110111110", -- t[31166] = 3
      "0000011" when "00111100110111111", -- t[31167] = 3
      "0000011" when "00111100111000000", -- t[31168] = 3
      "0000011" when "00111100111000001", -- t[31169] = 3
      "0000011" when "00111100111000010", -- t[31170] = 3
      "0000011" when "00111100111000011", -- t[31171] = 3
      "0000011" when "00111100111000100", -- t[31172] = 3
      "0000011" when "00111100111000101", -- t[31173] = 3
      "0000011" when "00111100111000110", -- t[31174] = 3
      "0000011" when "00111100111000111", -- t[31175] = 3
      "0000011" when "00111100111001000", -- t[31176] = 3
      "0000011" when "00111100111001001", -- t[31177] = 3
      "0000011" when "00111100111001010", -- t[31178] = 3
      "0000011" when "00111100111001011", -- t[31179] = 3
      "0000011" when "00111100111001100", -- t[31180] = 3
      "0000011" when "00111100111001101", -- t[31181] = 3
      "0000011" when "00111100111001110", -- t[31182] = 3
      "0000011" when "00111100111001111", -- t[31183] = 3
      "0000011" when "00111100111010000", -- t[31184] = 3
      "0000011" when "00111100111010001", -- t[31185] = 3
      "0000011" when "00111100111010010", -- t[31186] = 3
      "0000011" when "00111100111010011", -- t[31187] = 3
      "0000011" when "00111100111010100", -- t[31188] = 3
      "0000011" when "00111100111010101", -- t[31189] = 3
      "0000011" when "00111100111010110", -- t[31190] = 3
      "0000011" when "00111100111010111", -- t[31191] = 3
      "0000011" when "00111100111011000", -- t[31192] = 3
      "0000011" when "00111100111011001", -- t[31193] = 3
      "0000011" when "00111100111011010", -- t[31194] = 3
      "0000011" when "00111100111011011", -- t[31195] = 3
      "0000011" when "00111100111011100", -- t[31196] = 3
      "0000011" when "00111100111011101", -- t[31197] = 3
      "0000011" when "00111100111011110", -- t[31198] = 3
      "0000011" when "00111100111011111", -- t[31199] = 3
      "0000011" when "00111100111100000", -- t[31200] = 3
      "0000011" when "00111100111100001", -- t[31201] = 3
      "0000011" when "00111100111100010", -- t[31202] = 3
      "0000011" when "00111100111100011", -- t[31203] = 3
      "0000011" when "00111100111100100", -- t[31204] = 3
      "0000011" when "00111100111100101", -- t[31205] = 3
      "0000011" when "00111100111100110", -- t[31206] = 3
      "0000011" when "00111100111100111", -- t[31207] = 3
      "0000011" when "00111100111101000", -- t[31208] = 3
      "0000011" when "00111100111101001", -- t[31209] = 3
      "0000011" when "00111100111101010", -- t[31210] = 3
      "0000011" when "00111100111101011", -- t[31211] = 3
      "0000011" when "00111100111101100", -- t[31212] = 3
      "0000011" when "00111100111101101", -- t[31213] = 3
      "0000011" when "00111100111101110", -- t[31214] = 3
      "0000011" when "00111100111101111", -- t[31215] = 3
      "0000011" when "00111100111110000", -- t[31216] = 3
      "0000011" when "00111100111110001", -- t[31217] = 3
      "0000011" when "00111100111110010", -- t[31218] = 3
      "0000011" when "00111100111110011", -- t[31219] = 3
      "0000011" when "00111100111110100", -- t[31220] = 3
      "0000011" when "00111100111110101", -- t[31221] = 3
      "0000011" when "00111100111110110", -- t[31222] = 3
      "0000011" when "00111100111110111", -- t[31223] = 3
      "0000011" when "00111100111111000", -- t[31224] = 3
      "0000011" when "00111100111111001", -- t[31225] = 3
      "0000011" when "00111100111111010", -- t[31226] = 3
      "0000011" when "00111100111111011", -- t[31227] = 3
      "0000011" when "00111100111111100", -- t[31228] = 3
      "0000011" when "00111100111111101", -- t[31229] = 3
      "0000011" when "00111100111111110", -- t[31230] = 3
      "0000011" when "00111100111111111", -- t[31231] = 3
      "0000011" when "00111101000000000", -- t[31232] = 3
      "0000011" when "00111101000000001", -- t[31233] = 3
      "0000011" when "00111101000000010", -- t[31234] = 3
      "0000011" when "00111101000000011", -- t[31235] = 3
      "0000011" when "00111101000000100", -- t[31236] = 3
      "0000011" when "00111101000000101", -- t[31237] = 3
      "0000011" when "00111101000000110", -- t[31238] = 3
      "0000011" when "00111101000000111", -- t[31239] = 3
      "0000011" when "00111101000001000", -- t[31240] = 3
      "0000011" when "00111101000001001", -- t[31241] = 3
      "0000011" when "00111101000001010", -- t[31242] = 3
      "0000011" when "00111101000001011", -- t[31243] = 3
      "0000011" when "00111101000001100", -- t[31244] = 3
      "0000011" when "00111101000001101", -- t[31245] = 3
      "0000011" when "00111101000001110", -- t[31246] = 3
      "0000011" when "00111101000001111", -- t[31247] = 3
      "0000011" when "00111101000010000", -- t[31248] = 3
      "0000011" when "00111101000010001", -- t[31249] = 3
      "0000011" when "00111101000010010", -- t[31250] = 3
      "0000011" when "00111101000010011", -- t[31251] = 3
      "0000011" when "00111101000010100", -- t[31252] = 3
      "0000011" when "00111101000010101", -- t[31253] = 3
      "0000011" when "00111101000010110", -- t[31254] = 3
      "0000011" when "00111101000010111", -- t[31255] = 3
      "0000011" when "00111101000011000", -- t[31256] = 3
      "0000011" when "00111101000011001", -- t[31257] = 3
      "0000011" when "00111101000011010", -- t[31258] = 3
      "0000011" when "00111101000011011", -- t[31259] = 3
      "0000011" when "00111101000011100", -- t[31260] = 3
      "0000011" when "00111101000011101", -- t[31261] = 3
      "0000011" when "00111101000011110", -- t[31262] = 3
      "0000011" when "00111101000011111", -- t[31263] = 3
      "0000011" when "00111101000100000", -- t[31264] = 3
      "0000011" when "00111101000100001", -- t[31265] = 3
      "0000011" when "00111101000100010", -- t[31266] = 3
      "0000011" when "00111101000100011", -- t[31267] = 3
      "0000011" when "00111101000100100", -- t[31268] = 3
      "0000011" when "00111101000100101", -- t[31269] = 3
      "0000011" when "00111101000100110", -- t[31270] = 3
      "0000011" when "00111101000100111", -- t[31271] = 3
      "0000011" when "00111101000101000", -- t[31272] = 3
      "0000011" when "00111101000101001", -- t[31273] = 3
      "0000011" when "00111101000101010", -- t[31274] = 3
      "0000011" when "00111101000101011", -- t[31275] = 3
      "0000011" when "00111101000101100", -- t[31276] = 3
      "0000011" when "00111101000101101", -- t[31277] = 3
      "0000011" when "00111101000101110", -- t[31278] = 3
      "0000011" when "00111101000101111", -- t[31279] = 3
      "0000011" when "00111101000110000", -- t[31280] = 3
      "0000011" when "00111101000110001", -- t[31281] = 3
      "0000011" when "00111101000110010", -- t[31282] = 3
      "0000011" when "00111101000110011", -- t[31283] = 3
      "0000011" when "00111101000110100", -- t[31284] = 3
      "0000011" when "00111101000110101", -- t[31285] = 3
      "0000011" when "00111101000110110", -- t[31286] = 3
      "0000011" when "00111101000110111", -- t[31287] = 3
      "0000011" when "00111101000111000", -- t[31288] = 3
      "0000011" when "00111101000111001", -- t[31289] = 3
      "0000011" when "00111101000111010", -- t[31290] = 3
      "0000011" when "00111101000111011", -- t[31291] = 3
      "0000011" when "00111101000111100", -- t[31292] = 3
      "0000011" when "00111101000111101", -- t[31293] = 3
      "0000011" when "00111101000111110", -- t[31294] = 3
      "0000011" when "00111101000111111", -- t[31295] = 3
      "0000011" when "00111101001000000", -- t[31296] = 3
      "0000011" when "00111101001000001", -- t[31297] = 3
      "0000011" when "00111101001000010", -- t[31298] = 3
      "0000011" when "00111101001000011", -- t[31299] = 3
      "0000011" when "00111101001000100", -- t[31300] = 3
      "0000011" when "00111101001000101", -- t[31301] = 3
      "0000011" when "00111101001000110", -- t[31302] = 3
      "0000011" when "00111101001000111", -- t[31303] = 3
      "0000011" when "00111101001001000", -- t[31304] = 3
      "0000011" when "00111101001001001", -- t[31305] = 3
      "0000011" when "00111101001001010", -- t[31306] = 3
      "0000011" when "00111101001001011", -- t[31307] = 3
      "0000011" when "00111101001001100", -- t[31308] = 3
      "0000011" when "00111101001001101", -- t[31309] = 3
      "0000011" when "00111101001001110", -- t[31310] = 3
      "0000011" when "00111101001001111", -- t[31311] = 3
      "0000011" when "00111101001010000", -- t[31312] = 3
      "0000011" when "00111101001010001", -- t[31313] = 3
      "0000011" when "00111101001010010", -- t[31314] = 3
      "0000011" when "00111101001010011", -- t[31315] = 3
      "0000011" when "00111101001010100", -- t[31316] = 3
      "0000011" when "00111101001010101", -- t[31317] = 3
      "0000011" when "00111101001010110", -- t[31318] = 3
      "0000011" when "00111101001010111", -- t[31319] = 3
      "0000011" when "00111101001011000", -- t[31320] = 3
      "0000011" when "00111101001011001", -- t[31321] = 3
      "0000011" when "00111101001011010", -- t[31322] = 3
      "0000011" when "00111101001011011", -- t[31323] = 3
      "0000011" when "00111101001011100", -- t[31324] = 3
      "0000011" when "00111101001011101", -- t[31325] = 3
      "0000011" when "00111101001011110", -- t[31326] = 3
      "0000011" when "00111101001011111", -- t[31327] = 3
      "0000011" when "00111101001100000", -- t[31328] = 3
      "0000011" when "00111101001100001", -- t[31329] = 3
      "0000011" when "00111101001100010", -- t[31330] = 3
      "0000011" when "00111101001100011", -- t[31331] = 3
      "0000011" when "00111101001100100", -- t[31332] = 3
      "0000011" when "00111101001100101", -- t[31333] = 3
      "0000011" when "00111101001100110", -- t[31334] = 3
      "0000011" when "00111101001100111", -- t[31335] = 3
      "0000011" when "00111101001101000", -- t[31336] = 3
      "0000011" when "00111101001101001", -- t[31337] = 3
      "0000011" when "00111101001101010", -- t[31338] = 3
      "0000011" when "00111101001101011", -- t[31339] = 3
      "0000011" when "00111101001101100", -- t[31340] = 3
      "0000011" when "00111101001101101", -- t[31341] = 3
      "0000011" when "00111101001101110", -- t[31342] = 3
      "0000011" when "00111101001101111", -- t[31343] = 3
      "0000011" when "00111101001110000", -- t[31344] = 3
      "0000011" when "00111101001110001", -- t[31345] = 3
      "0000011" when "00111101001110010", -- t[31346] = 3
      "0000011" when "00111101001110011", -- t[31347] = 3
      "0000011" when "00111101001110100", -- t[31348] = 3
      "0000011" when "00111101001110101", -- t[31349] = 3
      "0000011" when "00111101001110110", -- t[31350] = 3
      "0000011" when "00111101001110111", -- t[31351] = 3
      "0000011" when "00111101001111000", -- t[31352] = 3
      "0000011" when "00111101001111001", -- t[31353] = 3
      "0000011" when "00111101001111010", -- t[31354] = 3
      "0000011" when "00111101001111011", -- t[31355] = 3
      "0000011" when "00111101001111100", -- t[31356] = 3
      "0000011" when "00111101001111101", -- t[31357] = 3
      "0000011" when "00111101001111110", -- t[31358] = 3
      "0000011" when "00111101001111111", -- t[31359] = 3
      "0000011" when "00111101010000000", -- t[31360] = 3
      "0000011" when "00111101010000001", -- t[31361] = 3
      "0000011" when "00111101010000010", -- t[31362] = 3
      "0000011" when "00111101010000011", -- t[31363] = 3
      "0000011" when "00111101010000100", -- t[31364] = 3
      "0000011" when "00111101010000101", -- t[31365] = 3
      "0000011" when "00111101010000110", -- t[31366] = 3
      "0000011" when "00111101010000111", -- t[31367] = 3
      "0000011" when "00111101010001000", -- t[31368] = 3
      "0000011" when "00111101010001001", -- t[31369] = 3
      "0000011" when "00111101010001010", -- t[31370] = 3
      "0000011" when "00111101010001011", -- t[31371] = 3
      "0000011" when "00111101010001100", -- t[31372] = 3
      "0000011" when "00111101010001101", -- t[31373] = 3
      "0000011" when "00111101010001110", -- t[31374] = 3
      "0000011" when "00111101010001111", -- t[31375] = 3
      "0000011" when "00111101010010000", -- t[31376] = 3
      "0000011" when "00111101010010001", -- t[31377] = 3
      "0000011" when "00111101010010010", -- t[31378] = 3
      "0000011" when "00111101010010011", -- t[31379] = 3
      "0000011" when "00111101010010100", -- t[31380] = 3
      "0000011" when "00111101010010101", -- t[31381] = 3
      "0000011" when "00111101010010110", -- t[31382] = 3
      "0000011" when "00111101010010111", -- t[31383] = 3
      "0000011" when "00111101010011000", -- t[31384] = 3
      "0000011" when "00111101010011001", -- t[31385] = 3
      "0000011" when "00111101010011010", -- t[31386] = 3
      "0000011" when "00111101010011011", -- t[31387] = 3
      "0000011" when "00111101010011100", -- t[31388] = 3
      "0000011" when "00111101010011101", -- t[31389] = 3
      "0000011" when "00111101010011110", -- t[31390] = 3
      "0000011" when "00111101010011111", -- t[31391] = 3
      "0000011" when "00111101010100000", -- t[31392] = 3
      "0000011" when "00111101010100001", -- t[31393] = 3
      "0000011" when "00111101010100010", -- t[31394] = 3
      "0000011" when "00111101010100011", -- t[31395] = 3
      "0000011" when "00111101010100100", -- t[31396] = 3
      "0000011" when "00111101010100101", -- t[31397] = 3
      "0000011" when "00111101010100110", -- t[31398] = 3
      "0000011" when "00111101010100111", -- t[31399] = 3
      "0000011" when "00111101010101000", -- t[31400] = 3
      "0000011" when "00111101010101001", -- t[31401] = 3
      "0000011" when "00111101010101010", -- t[31402] = 3
      "0000011" when "00111101010101011", -- t[31403] = 3
      "0000011" when "00111101010101100", -- t[31404] = 3
      "0000011" when "00111101010101101", -- t[31405] = 3
      "0000011" when "00111101010101110", -- t[31406] = 3
      "0000011" when "00111101010101111", -- t[31407] = 3
      "0000011" when "00111101010110000", -- t[31408] = 3
      "0000011" when "00111101010110001", -- t[31409] = 3
      "0000011" when "00111101010110010", -- t[31410] = 3
      "0000011" when "00111101010110011", -- t[31411] = 3
      "0000011" when "00111101010110100", -- t[31412] = 3
      "0000011" when "00111101010110101", -- t[31413] = 3
      "0000011" when "00111101010110110", -- t[31414] = 3
      "0000011" when "00111101010110111", -- t[31415] = 3
      "0000011" when "00111101010111000", -- t[31416] = 3
      "0000011" when "00111101010111001", -- t[31417] = 3
      "0000011" when "00111101010111010", -- t[31418] = 3
      "0000011" when "00111101010111011", -- t[31419] = 3
      "0000011" when "00111101010111100", -- t[31420] = 3
      "0000011" when "00111101010111101", -- t[31421] = 3
      "0000011" when "00111101010111110", -- t[31422] = 3
      "0000011" when "00111101010111111", -- t[31423] = 3
      "0000011" when "00111101011000000", -- t[31424] = 3
      "0000011" when "00111101011000001", -- t[31425] = 3
      "0000011" when "00111101011000010", -- t[31426] = 3
      "0000011" when "00111101011000011", -- t[31427] = 3
      "0000011" when "00111101011000100", -- t[31428] = 3
      "0000011" when "00111101011000101", -- t[31429] = 3
      "0000011" when "00111101011000110", -- t[31430] = 3
      "0000011" when "00111101011000111", -- t[31431] = 3
      "0000011" when "00111101011001000", -- t[31432] = 3
      "0000011" when "00111101011001001", -- t[31433] = 3
      "0000011" when "00111101011001010", -- t[31434] = 3
      "0000011" when "00111101011001011", -- t[31435] = 3
      "0000011" when "00111101011001100", -- t[31436] = 3
      "0000011" when "00111101011001101", -- t[31437] = 3
      "0000011" when "00111101011001110", -- t[31438] = 3
      "0000011" when "00111101011001111", -- t[31439] = 3
      "0000011" when "00111101011010000", -- t[31440] = 3
      "0000011" when "00111101011010001", -- t[31441] = 3
      "0000011" when "00111101011010010", -- t[31442] = 3
      "0000011" when "00111101011010011", -- t[31443] = 3
      "0000011" when "00111101011010100", -- t[31444] = 3
      "0000011" when "00111101011010101", -- t[31445] = 3
      "0000011" when "00111101011010110", -- t[31446] = 3
      "0000011" when "00111101011010111", -- t[31447] = 3
      "0000011" when "00111101011011000", -- t[31448] = 3
      "0000011" when "00111101011011001", -- t[31449] = 3
      "0000011" when "00111101011011010", -- t[31450] = 3
      "0000011" when "00111101011011011", -- t[31451] = 3
      "0000011" when "00111101011011100", -- t[31452] = 3
      "0000011" when "00111101011011101", -- t[31453] = 3
      "0000011" when "00111101011011110", -- t[31454] = 3
      "0000011" when "00111101011011111", -- t[31455] = 3
      "0000011" when "00111101011100000", -- t[31456] = 3
      "0000011" when "00111101011100001", -- t[31457] = 3
      "0000011" when "00111101011100010", -- t[31458] = 3
      "0000011" when "00111101011100011", -- t[31459] = 3
      "0000011" when "00111101011100100", -- t[31460] = 3
      "0000011" when "00111101011100101", -- t[31461] = 3
      "0000011" when "00111101011100110", -- t[31462] = 3
      "0000011" when "00111101011100111", -- t[31463] = 3
      "0000011" when "00111101011101000", -- t[31464] = 3
      "0000011" when "00111101011101001", -- t[31465] = 3
      "0000011" when "00111101011101010", -- t[31466] = 3
      "0000011" when "00111101011101011", -- t[31467] = 3
      "0000011" when "00111101011101100", -- t[31468] = 3
      "0000011" when "00111101011101101", -- t[31469] = 3
      "0000011" when "00111101011101110", -- t[31470] = 3
      "0000011" when "00111101011101111", -- t[31471] = 3
      "0000011" when "00111101011110000", -- t[31472] = 3
      "0000011" when "00111101011110001", -- t[31473] = 3
      "0000011" when "00111101011110010", -- t[31474] = 3
      "0000011" when "00111101011110011", -- t[31475] = 3
      "0000011" when "00111101011110100", -- t[31476] = 3
      "0000011" when "00111101011110101", -- t[31477] = 3
      "0000011" when "00111101011110110", -- t[31478] = 3
      "0000011" when "00111101011110111", -- t[31479] = 3
      "0000011" when "00111101011111000", -- t[31480] = 3
      "0000011" when "00111101011111001", -- t[31481] = 3
      "0000011" when "00111101011111010", -- t[31482] = 3
      "0000011" when "00111101011111011", -- t[31483] = 3
      "0000011" when "00111101011111100", -- t[31484] = 3
      "0000011" when "00111101011111101", -- t[31485] = 3
      "0000011" when "00111101011111110", -- t[31486] = 3
      "0000011" when "00111101011111111", -- t[31487] = 3
      "0000011" when "00111101100000000", -- t[31488] = 3
      "0000011" when "00111101100000001", -- t[31489] = 3
      "0000011" when "00111101100000010", -- t[31490] = 3
      "0000011" when "00111101100000011", -- t[31491] = 3
      "0000011" when "00111101100000100", -- t[31492] = 3
      "0000011" when "00111101100000101", -- t[31493] = 3
      "0000011" when "00111101100000110", -- t[31494] = 3
      "0000011" when "00111101100000111", -- t[31495] = 3
      "0000011" when "00111101100001000", -- t[31496] = 3
      "0000011" when "00111101100001001", -- t[31497] = 3
      "0000011" when "00111101100001010", -- t[31498] = 3
      "0000011" when "00111101100001011", -- t[31499] = 3
      "0000011" when "00111101100001100", -- t[31500] = 3
      "0000011" when "00111101100001101", -- t[31501] = 3
      "0000011" when "00111101100001110", -- t[31502] = 3
      "0000011" when "00111101100001111", -- t[31503] = 3
      "0000011" when "00111101100010000", -- t[31504] = 3
      "0000011" when "00111101100010001", -- t[31505] = 3
      "0000011" when "00111101100010010", -- t[31506] = 3
      "0000011" when "00111101100010011", -- t[31507] = 3
      "0000011" when "00111101100010100", -- t[31508] = 3
      "0000011" when "00111101100010101", -- t[31509] = 3
      "0000011" when "00111101100010110", -- t[31510] = 3
      "0000011" when "00111101100010111", -- t[31511] = 3
      "0000011" when "00111101100011000", -- t[31512] = 3
      "0000011" when "00111101100011001", -- t[31513] = 3
      "0000011" when "00111101100011010", -- t[31514] = 3
      "0000011" when "00111101100011011", -- t[31515] = 3
      "0000011" when "00111101100011100", -- t[31516] = 3
      "0000011" when "00111101100011101", -- t[31517] = 3
      "0000011" when "00111101100011110", -- t[31518] = 3
      "0000011" when "00111101100011111", -- t[31519] = 3
      "0000011" when "00111101100100000", -- t[31520] = 3
      "0000011" when "00111101100100001", -- t[31521] = 3
      "0000011" when "00111101100100010", -- t[31522] = 3
      "0000011" when "00111101100100011", -- t[31523] = 3
      "0000011" when "00111101100100100", -- t[31524] = 3
      "0000011" when "00111101100100101", -- t[31525] = 3
      "0000011" when "00111101100100110", -- t[31526] = 3
      "0000011" when "00111101100100111", -- t[31527] = 3
      "0000011" when "00111101100101000", -- t[31528] = 3
      "0000011" when "00111101100101001", -- t[31529] = 3
      "0000011" when "00111101100101010", -- t[31530] = 3
      "0000011" when "00111101100101011", -- t[31531] = 3
      "0000011" when "00111101100101100", -- t[31532] = 3
      "0000011" when "00111101100101101", -- t[31533] = 3
      "0000011" when "00111101100101110", -- t[31534] = 3
      "0000011" when "00111101100101111", -- t[31535] = 3
      "0000011" when "00111101100110000", -- t[31536] = 3
      "0000011" when "00111101100110001", -- t[31537] = 3
      "0000011" when "00111101100110010", -- t[31538] = 3
      "0000011" when "00111101100110011", -- t[31539] = 3
      "0000011" when "00111101100110100", -- t[31540] = 3
      "0000011" when "00111101100110101", -- t[31541] = 3
      "0000011" when "00111101100110110", -- t[31542] = 3
      "0000011" when "00111101100110111", -- t[31543] = 3
      "0000011" when "00111101100111000", -- t[31544] = 3
      "0000011" when "00111101100111001", -- t[31545] = 3
      "0000011" when "00111101100111010", -- t[31546] = 3
      "0000011" when "00111101100111011", -- t[31547] = 3
      "0000011" when "00111101100111100", -- t[31548] = 3
      "0000011" when "00111101100111101", -- t[31549] = 3
      "0000011" when "00111101100111110", -- t[31550] = 3
      "0000011" when "00111101100111111", -- t[31551] = 3
      "0000011" when "00111101101000000", -- t[31552] = 3
      "0000011" when "00111101101000001", -- t[31553] = 3
      "0000011" when "00111101101000010", -- t[31554] = 3
      "0000011" when "00111101101000011", -- t[31555] = 3
      "0000011" when "00111101101000100", -- t[31556] = 3
      "0000011" when "00111101101000101", -- t[31557] = 3
      "0000011" when "00111101101000110", -- t[31558] = 3
      "0000011" when "00111101101000111", -- t[31559] = 3
      "0000011" when "00111101101001000", -- t[31560] = 3
      "0000011" when "00111101101001001", -- t[31561] = 3
      "0000011" when "00111101101001010", -- t[31562] = 3
      "0000011" when "00111101101001011", -- t[31563] = 3
      "0000011" when "00111101101001100", -- t[31564] = 3
      "0000011" when "00111101101001101", -- t[31565] = 3
      "0000011" when "00111101101001110", -- t[31566] = 3
      "0000011" when "00111101101001111", -- t[31567] = 3
      "0000011" when "00111101101010000", -- t[31568] = 3
      "0000011" when "00111101101010001", -- t[31569] = 3
      "0000011" when "00111101101010010", -- t[31570] = 3
      "0000011" when "00111101101010011", -- t[31571] = 3
      "0000011" when "00111101101010100", -- t[31572] = 3
      "0000011" when "00111101101010101", -- t[31573] = 3
      "0000011" when "00111101101010110", -- t[31574] = 3
      "0000011" when "00111101101010111", -- t[31575] = 3
      "0000011" when "00111101101011000", -- t[31576] = 3
      "0000011" when "00111101101011001", -- t[31577] = 3
      "0000011" when "00111101101011010", -- t[31578] = 3
      "0000011" when "00111101101011011", -- t[31579] = 3
      "0000011" when "00111101101011100", -- t[31580] = 3
      "0000011" when "00111101101011101", -- t[31581] = 3
      "0000011" when "00111101101011110", -- t[31582] = 3
      "0000011" when "00111101101011111", -- t[31583] = 3
      "0000011" when "00111101101100000", -- t[31584] = 3
      "0000011" when "00111101101100001", -- t[31585] = 3
      "0000011" when "00111101101100010", -- t[31586] = 3
      "0000011" when "00111101101100011", -- t[31587] = 3
      "0000011" when "00111101101100100", -- t[31588] = 3
      "0000011" when "00111101101100101", -- t[31589] = 3
      "0000011" when "00111101101100110", -- t[31590] = 3
      "0000011" when "00111101101100111", -- t[31591] = 3
      "0000011" when "00111101101101000", -- t[31592] = 3
      "0000011" when "00111101101101001", -- t[31593] = 3
      "0000011" when "00111101101101010", -- t[31594] = 3
      "0000011" when "00111101101101011", -- t[31595] = 3
      "0000011" when "00111101101101100", -- t[31596] = 3
      "0000011" when "00111101101101101", -- t[31597] = 3
      "0000011" when "00111101101101110", -- t[31598] = 3
      "0000011" when "00111101101101111", -- t[31599] = 3
      "0000011" when "00111101101110000", -- t[31600] = 3
      "0000011" when "00111101101110001", -- t[31601] = 3
      "0000011" when "00111101101110010", -- t[31602] = 3
      "0000011" when "00111101101110011", -- t[31603] = 3
      "0000011" when "00111101101110100", -- t[31604] = 3
      "0000011" when "00111101101110101", -- t[31605] = 3
      "0000011" when "00111101101110110", -- t[31606] = 3
      "0000011" when "00111101101110111", -- t[31607] = 3
      "0000011" when "00111101101111000", -- t[31608] = 3
      "0000011" when "00111101101111001", -- t[31609] = 3
      "0000011" when "00111101101111010", -- t[31610] = 3
      "0000011" when "00111101101111011", -- t[31611] = 3
      "0000011" when "00111101101111100", -- t[31612] = 3
      "0000011" when "00111101101111101", -- t[31613] = 3
      "0000011" when "00111101101111110", -- t[31614] = 3
      "0000011" when "00111101101111111", -- t[31615] = 3
      "0000011" when "00111101110000000", -- t[31616] = 3
      "0000011" when "00111101110000001", -- t[31617] = 3
      "0000011" when "00111101110000010", -- t[31618] = 3
      "0000011" when "00111101110000011", -- t[31619] = 3
      "0000011" when "00111101110000100", -- t[31620] = 3
      "0000011" when "00111101110000101", -- t[31621] = 3
      "0000011" when "00111101110000110", -- t[31622] = 3
      "0000011" when "00111101110000111", -- t[31623] = 3
      "0000011" when "00111101110001000", -- t[31624] = 3
      "0000011" when "00111101110001001", -- t[31625] = 3
      "0000011" when "00111101110001010", -- t[31626] = 3
      "0000011" when "00111101110001011", -- t[31627] = 3
      "0000011" when "00111101110001100", -- t[31628] = 3
      "0000011" when "00111101110001101", -- t[31629] = 3
      "0000011" when "00111101110001110", -- t[31630] = 3
      "0000011" when "00111101110001111", -- t[31631] = 3
      "0000011" when "00111101110010000", -- t[31632] = 3
      "0000011" when "00111101110010001", -- t[31633] = 3
      "0000011" when "00111101110010010", -- t[31634] = 3
      "0000011" when "00111101110010011", -- t[31635] = 3
      "0000011" when "00111101110010100", -- t[31636] = 3
      "0000011" when "00111101110010101", -- t[31637] = 3
      "0000011" when "00111101110010110", -- t[31638] = 3
      "0000011" when "00111101110010111", -- t[31639] = 3
      "0000011" when "00111101110011000", -- t[31640] = 3
      "0000011" when "00111101110011001", -- t[31641] = 3
      "0000011" when "00111101110011010", -- t[31642] = 3
      "0000011" when "00111101110011011", -- t[31643] = 3
      "0000011" when "00111101110011100", -- t[31644] = 3
      "0000011" when "00111101110011101", -- t[31645] = 3
      "0000011" when "00111101110011110", -- t[31646] = 3
      "0000011" when "00111101110011111", -- t[31647] = 3
      "0000011" when "00111101110100000", -- t[31648] = 3
      "0000011" when "00111101110100001", -- t[31649] = 3
      "0000011" when "00111101110100010", -- t[31650] = 3
      "0000011" when "00111101110100011", -- t[31651] = 3
      "0000011" when "00111101110100100", -- t[31652] = 3
      "0000011" when "00111101110100101", -- t[31653] = 3
      "0000011" when "00111101110100110", -- t[31654] = 3
      "0000011" when "00111101110100111", -- t[31655] = 3
      "0000011" when "00111101110101000", -- t[31656] = 3
      "0000011" when "00111101110101001", -- t[31657] = 3
      "0000011" when "00111101110101010", -- t[31658] = 3
      "0000011" when "00111101110101011", -- t[31659] = 3
      "0000011" when "00111101110101100", -- t[31660] = 3
      "0000011" when "00111101110101101", -- t[31661] = 3
      "0000011" when "00111101110101110", -- t[31662] = 3
      "0000011" when "00111101110101111", -- t[31663] = 3
      "0000011" when "00111101110110000", -- t[31664] = 3
      "0000011" when "00111101110110001", -- t[31665] = 3
      "0000011" when "00111101110110010", -- t[31666] = 3
      "0000011" when "00111101110110011", -- t[31667] = 3
      "0000011" when "00111101110110100", -- t[31668] = 3
      "0000011" when "00111101110110101", -- t[31669] = 3
      "0000011" when "00111101110110110", -- t[31670] = 3
      "0000011" when "00111101110110111", -- t[31671] = 3
      "0000011" when "00111101110111000", -- t[31672] = 3
      "0000011" when "00111101110111001", -- t[31673] = 3
      "0000011" when "00111101110111010", -- t[31674] = 3
      "0000011" when "00111101110111011", -- t[31675] = 3
      "0000011" when "00111101110111100", -- t[31676] = 3
      "0000011" when "00111101110111101", -- t[31677] = 3
      "0000011" when "00111101110111110", -- t[31678] = 3
      "0000011" when "00111101110111111", -- t[31679] = 3
      "0000011" when "00111101111000000", -- t[31680] = 3
      "0000011" when "00111101111000001", -- t[31681] = 3
      "0000011" when "00111101111000010", -- t[31682] = 3
      "0000011" when "00111101111000011", -- t[31683] = 3
      "0000011" when "00111101111000100", -- t[31684] = 3
      "0000011" when "00111101111000101", -- t[31685] = 3
      "0000011" when "00111101111000110", -- t[31686] = 3
      "0000011" when "00111101111000111", -- t[31687] = 3
      "0000011" when "00111101111001000", -- t[31688] = 3
      "0000011" when "00111101111001001", -- t[31689] = 3
      "0000011" when "00111101111001010", -- t[31690] = 3
      "0000011" when "00111101111001011", -- t[31691] = 3
      "0000011" when "00111101111001100", -- t[31692] = 3
      "0000011" when "00111101111001101", -- t[31693] = 3
      "0000011" when "00111101111001110", -- t[31694] = 3
      "0000011" when "00111101111001111", -- t[31695] = 3
      "0000011" when "00111101111010000", -- t[31696] = 3
      "0000011" when "00111101111010001", -- t[31697] = 3
      "0000011" when "00111101111010010", -- t[31698] = 3
      "0000011" when "00111101111010011", -- t[31699] = 3
      "0000011" when "00111101111010100", -- t[31700] = 3
      "0000011" when "00111101111010101", -- t[31701] = 3
      "0000011" when "00111101111010110", -- t[31702] = 3
      "0000011" when "00111101111010111", -- t[31703] = 3
      "0000011" when "00111101111011000", -- t[31704] = 3
      "0000011" when "00111101111011001", -- t[31705] = 3
      "0000011" when "00111101111011010", -- t[31706] = 3
      "0000011" when "00111101111011011", -- t[31707] = 3
      "0000011" when "00111101111011100", -- t[31708] = 3
      "0000011" when "00111101111011101", -- t[31709] = 3
      "0000011" when "00111101111011110", -- t[31710] = 3
      "0000011" when "00111101111011111", -- t[31711] = 3
      "0000011" when "00111101111100000", -- t[31712] = 3
      "0000011" when "00111101111100001", -- t[31713] = 3
      "0000011" when "00111101111100010", -- t[31714] = 3
      "0000011" when "00111101111100011", -- t[31715] = 3
      "0000011" when "00111101111100100", -- t[31716] = 3
      "0000011" when "00111101111100101", -- t[31717] = 3
      "0000011" when "00111101111100110", -- t[31718] = 3
      "0000011" when "00111101111100111", -- t[31719] = 3
      "0000011" when "00111101111101000", -- t[31720] = 3
      "0000011" when "00111101111101001", -- t[31721] = 3
      "0000011" when "00111101111101010", -- t[31722] = 3
      "0000011" when "00111101111101011", -- t[31723] = 3
      "0000011" when "00111101111101100", -- t[31724] = 3
      "0000011" when "00111101111101101", -- t[31725] = 3
      "0000011" when "00111101111101110", -- t[31726] = 3
      "0000011" when "00111101111101111", -- t[31727] = 3
      "0000011" when "00111101111110000", -- t[31728] = 3
      "0000011" when "00111101111110001", -- t[31729] = 3
      "0000011" when "00111101111110010", -- t[31730] = 3
      "0000011" when "00111101111110011", -- t[31731] = 3
      "0000011" when "00111101111110100", -- t[31732] = 3
      "0000011" when "00111101111110101", -- t[31733] = 3
      "0000011" when "00111101111110110", -- t[31734] = 3
      "0000011" when "00111101111110111", -- t[31735] = 3
      "0000011" when "00111101111111000", -- t[31736] = 3
      "0000011" when "00111101111111001", -- t[31737] = 3
      "0000011" when "00111101111111010", -- t[31738] = 3
      "0000011" when "00111101111111011", -- t[31739] = 3
      "0000011" when "00111101111111100", -- t[31740] = 3
      "0000011" when "00111101111111101", -- t[31741] = 3
      "0000011" when "00111101111111110", -- t[31742] = 3
      "0000011" when "00111101111111111", -- t[31743] = 3
      "0000011" when "00111110000000000", -- t[31744] = 3
      "0000011" when "00111110000000001", -- t[31745] = 3
      "0000011" when "00111110000000010", -- t[31746] = 3
      "0000011" when "00111110000000011", -- t[31747] = 3
      "0000011" when "00111110000000100", -- t[31748] = 3
      "0000011" when "00111110000000101", -- t[31749] = 3
      "0000011" when "00111110000000110", -- t[31750] = 3
      "0000011" when "00111110000000111", -- t[31751] = 3
      "0000011" when "00111110000001000", -- t[31752] = 3
      "0000011" when "00111110000001001", -- t[31753] = 3
      "0000011" when "00111110000001010", -- t[31754] = 3
      "0000011" when "00111110000001011", -- t[31755] = 3
      "0000011" when "00111110000001100", -- t[31756] = 3
      "0000011" when "00111110000001101", -- t[31757] = 3
      "0000011" when "00111110000001110", -- t[31758] = 3
      "0000011" when "00111110000001111", -- t[31759] = 3
      "0000011" when "00111110000010000", -- t[31760] = 3
      "0000011" when "00111110000010001", -- t[31761] = 3
      "0000011" when "00111110000010010", -- t[31762] = 3
      "0000011" when "00111110000010011", -- t[31763] = 3
      "0000011" when "00111110000010100", -- t[31764] = 3
      "0000011" when "00111110000010101", -- t[31765] = 3
      "0000011" when "00111110000010110", -- t[31766] = 3
      "0000011" when "00111110000010111", -- t[31767] = 3
      "0000011" when "00111110000011000", -- t[31768] = 3
      "0000011" when "00111110000011001", -- t[31769] = 3
      "0000011" when "00111110000011010", -- t[31770] = 3
      "0000011" when "00111110000011011", -- t[31771] = 3
      "0000011" when "00111110000011100", -- t[31772] = 3
      "0000011" when "00111110000011101", -- t[31773] = 3
      "0000011" when "00111110000011110", -- t[31774] = 3
      "0000011" when "00111110000011111", -- t[31775] = 3
      "0000011" when "00111110000100000", -- t[31776] = 3
      "0000011" when "00111110000100001", -- t[31777] = 3
      "0000011" when "00111110000100010", -- t[31778] = 3
      "0000011" when "00111110000100011", -- t[31779] = 3
      "0000011" when "00111110000100100", -- t[31780] = 3
      "0000011" when "00111110000100101", -- t[31781] = 3
      "0000011" when "00111110000100110", -- t[31782] = 3
      "0000011" when "00111110000100111", -- t[31783] = 3
      "0000011" when "00111110000101000", -- t[31784] = 3
      "0000011" when "00111110000101001", -- t[31785] = 3
      "0000011" when "00111110000101010", -- t[31786] = 3
      "0000011" when "00111110000101011", -- t[31787] = 3
      "0000011" when "00111110000101100", -- t[31788] = 3
      "0000011" when "00111110000101101", -- t[31789] = 3
      "0000011" when "00111110000101110", -- t[31790] = 3
      "0000011" when "00111110000101111", -- t[31791] = 3
      "0000011" when "00111110000110000", -- t[31792] = 3
      "0000011" when "00111110000110001", -- t[31793] = 3
      "0000011" when "00111110000110010", -- t[31794] = 3
      "0000011" when "00111110000110011", -- t[31795] = 3
      "0000011" when "00111110000110100", -- t[31796] = 3
      "0000011" when "00111110000110101", -- t[31797] = 3
      "0000011" when "00111110000110110", -- t[31798] = 3
      "0000011" when "00111110000110111", -- t[31799] = 3
      "0000011" when "00111110000111000", -- t[31800] = 3
      "0000011" when "00111110000111001", -- t[31801] = 3
      "0000011" when "00111110000111010", -- t[31802] = 3
      "0000011" when "00111110000111011", -- t[31803] = 3
      "0000011" when "00111110000111100", -- t[31804] = 3
      "0000011" when "00111110000111101", -- t[31805] = 3
      "0000011" when "00111110000111110", -- t[31806] = 3
      "0000011" when "00111110000111111", -- t[31807] = 3
      "0000011" when "00111110001000000", -- t[31808] = 3
      "0000011" when "00111110001000001", -- t[31809] = 3
      "0000011" when "00111110001000010", -- t[31810] = 3
      "0000011" when "00111110001000011", -- t[31811] = 3
      "0000011" when "00111110001000100", -- t[31812] = 3
      "0000011" when "00111110001000101", -- t[31813] = 3
      "0000011" when "00111110001000110", -- t[31814] = 3
      "0000011" when "00111110001000111", -- t[31815] = 3
      "0000011" when "00111110001001000", -- t[31816] = 3
      "0000011" when "00111110001001001", -- t[31817] = 3
      "0000011" when "00111110001001010", -- t[31818] = 3
      "0000011" when "00111110001001011", -- t[31819] = 3
      "0000011" when "00111110001001100", -- t[31820] = 3
      "0000011" when "00111110001001101", -- t[31821] = 3
      "0000011" when "00111110001001110", -- t[31822] = 3
      "0000011" when "00111110001001111", -- t[31823] = 3
      "0000011" when "00111110001010000", -- t[31824] = 3
      "0000011" when "00111110001010001", -- t[31825] = 3
      "0000011" when "00111110001010010", -- t[31826] = 3
      "0000011" when "00111110001010011", -- t[31827] = 3
      "0000011" when "00111110001010100", -- t[31828] = 3
      "0000011" when "00111110001010101", -- t[31829] = 3
      "0000011" when "00111110001010110", -- t[31830] = 3
      "0000011" when "00111110001010111", -- t[31831] = 3
      "0000011" when "00111110001011000", -- t[31832] = 3
      "0000011" when "00111110001011001", -- t[31833] = 3
      "0000011" when "00111110001011010", -- t[31834] = 3
      "0000011" when "00111110001011011", -- t[31835] = 3
      "0000011" when "00111110001011100", -- t[31836] = 3
      "0000011" when "00111110001011101", -- t[31837] = 3
      "0000011" when "00111110001011110", -- t[31838] = 3
      "0000011" when "00111110001011111", -- t[31839] = 3
      "0000011" when "00111110001100000", -- t[31840] = 3
      "0000011" when "00111110001100001", -- t[31841] = 3
      "0000011" when "00111110001100010", -- t[31842] = 3
      "0000011" when "00111110001100011", -- t[31843] = 3
      "0000011" when "00111110001100100", -- t[31844] = 3
      "0000011" when "00111110001100101", -- t[31845] = 3
      "0000011" when "00111110001100110", -- t[31846] = 3
      "0000011" when "00111110001100111", -- t[31847] = 3
      "0000011" when "00111110001101000", -- t[31848] = 3
      "0000011" when "00111110001101001", -- t[31849] = 3
      "0000011" when "00111110001101010", -- t[31850] = 3
      "0000011" when "00111110001101011", -- t[31851] = 3
      "0000011" when "00111110001101100", -- t[31852] = 3
      "0000011" when "00111110001101101", -- t[31853] = 3
      "0000011" when "00111110001101110", -- t[31854] = 3
      "0000011" when "00111110001101111", -- t[31855] = 3
      "0000011" when "00111110001110000", -- t[31856] = 3
      "0000011" when "00111110001110001", -- t[31857] = 3
      "0000011" when "00111110001110010", -- t[31858] = 3
      "0000011" when "00111110001110011", -- t[31859] = 3
      "0000011" when "00111110001110100", -- t[31860] = 3
      "0000011" when "00111110001110101", -- t[31861] = 3
      "0000011" when "00111110001110110", -- t[31862] = 3
      "0000011" when "00111110001110111", -- t[31863] = 3
      "0000011" when "00111110001111000", -- t[31864] = 3
      "0000011" when "00111110001111001", -- t[31865] = 3
      "0000011" when "00111110001111010", -- t[31866] = 3
      "0000011" when "00111110001111011", -- t[31867] = 3
      "0000011" when "00111110001111100", -- t[31868] = 3
      "0000011" when "00111110001111101", -- t[31869] = 3
      "0000011" when "00111110001111110", -- t[31870] = 3
      "0000011" when "00111110001111111", -- t[31871] = 3
      "0000011" when "00111110010000000", -- t[31872] = 3
      "0000011" when "00111110010000001", -- t[31873] = 3
      "0000011" when "00111110010000010", -- t[31874] = 3
      "0000011" when "00111110010000011", -- t[31875] = 3
      "0000011" when "00111110010000100", -- t[31876] = 3
      "0000011" when "00111110010000101", -- t[31877] = 3
      "0000011" when "00111110010000110", -- t[31878] = 3
      "0000011" when "00111110010000111", -- t[31879] = 3
      "0000011" when "00111110010001000", -- t[31880] = 3
      "0000011" when "00111110010001001", -- t[31881] = 3
      "0000011" when "00111110010001010", -- t[31882] = 3
      "0000011" when "00111110010001011", -- t[31883] = 3
      "0000011" when "00111110010001100", -- t[31884] = 3
      "0000011" when "00111110010001101", -- t[31885] = 3
      "0000011" when "00111110010001110", -- t[31886] = 3
      "0000011" when "00111110010001111", -- t[31887] = 3
      "0000011" when "00111110010010000", -- t[31888] = 3
      "0000011" when "00111110010010001", -- t[31889] = 3
      "0000011" when "00111110010010010", -- t[31890] = 3
      "0000011" when "00111110010010011", -- t[31891] = 3
      "0000011" when "00111110010010100", -- t[31892] = 3
      "0000011" when "00111110010010101", -- t[31893] = 3
      "0000011" when "00111110010010110", -- t[31894] = 3
      "0000011" when "00111110010010111", -- t[31895] = 3
      "0000011" when "00111110010011000", -- t[31896] = 3
      "0000011" when "00111110010011001", -- t[31897] = 3
      "0000011" when "00111110010011010", -- t[31898] = 3
      "0000011" when "00111110010011011", -- t[31899] = 3
      "0000011" when "00111110010011100", -- t[31900] = 3
      "0000011" when "00111110010011101", -- t[31901] = 3
      "0000011" when "00111110010011110", -- t[31902] = 3
      "0000011" when "00111110010011111", -- t[31903] = 3
      "0000011" when "00111110010100000", -- t[31904] = 3
      "0000011" when "00111110010100001", -- t[31905] = 3
      "0000011" when "00111110010100010", -- t[31906] = 3
      "0000011" when "00111110010100011", -- t[31907] = 3
      "0000011" when "00111110010100100", -- t[31908] = 3
      "0000011" when "00111110010100101", -- t[31909] = 3
      "0000011" when "00111110010100110", -- t[31910] = 3
      "0000011" when "00111110010100111", -- t[31911] = 3
      "0000011" when "00111110010101000", -- t[31912] = 3
      "0000011" when "00111110010101001", -- t[31913] = 3
      "0000011" when "00111110010101010", -- t[31914] = 3
      "0000011" when "00111110010101011", -- t[31915] = 3
      "0000011" when "00111110010101100", -- t[31916] = 3
      "0000011" when "00111110010101101", -- t[31917] = 3
      "0000011" when "00111110010101110", -- t[31918] = 3
      "0000011" when "00111110010101111", -- t[31919] = 3
      "0000011" when "00111110010110000", -- t[31920] = 3
      "0000011" when "00111110010110001", -- t[31921] = 3
      "0000011" when "00111110010110010", -- t[31922] = 3
      "0000011" when "00111110010110011", -- t[31923] = 3
      "0000011" when "00111110010110100", -- t[31924] = 3
      "0000011" when "00111110010110101", -- t[31925] = 3
      "0000011" when "00111110010110110", -- t[31926] = 3
      "0000011" when "00111110010110111", -- t[31927] = 3
      "0000011" when "00111110010111000", -- t[31928] = 3
      "0000011" when "00111110010111001", -- t[31929] = 3
      "0000011" when "00111110010111010", -- t[31930] = 3
      "0000011" when "00111110010111011", -- t[31931] = 3
      "0000011" when "00111110010111100", -- t[31932] = 3
      "0000011" when "00111110010111101", -- t[31933] = 3
      "0000011" when "00111110010111110", -- t[31934] = 3
      "0000011" when "00111110010111111", -- t[31935] = 3
      "0000011" when "00111110011000000", -- t[31936] = 3
      "0000011" when "00111110011000001", -- t[31937] = 3
      "0000011" when "00111110011000010", -- t[31938] = 3
      "0000011" when "00111110011000011", -- t[31939] = 3
      "0000011" when "00111110011000100", -- t[31940] = 3
      "0000011" when "00111110011000101", -- t[31941] = 3
      "0000011" when "00111110011000110", -- t[31942] = 3
      "0000011" when "00111110011000111", -- t[31943] = 3
      "0000011" when "00111110011001000", -- t[31944] = 3
      "0000011" when "00111110011001001", -- t[31945] = 3
      "0000011" when "00111110011001010", -- t[31946] = 3
      "0000011" when "00111110011001011", -- t[31947] = 3
      "0000011" when "00111110011001100", -- t[31948] = 3
      "0000011" when "00111110011001101", -- t[31949] = 3
      "0000011" when "00111110011001110", -- t[31950] = 3
      "0000011" when "00111110011001111", -- t[31951] = 3
      "0000011" when "00111110011010000", -- t[31952] = 3
      "0000011" when "00111110011010001", -- t[31953] = 3
      "0000011" when "00111110011010010", -- t[31954] = 3
      "0000011" when "00111110011010011", -- t[31955] = 3
      "0000011" when "00111110011010100", -- t[31956] = 3
      "0000011" when "00111110011010101", -- t[31957] = 3
      "0000011" when "00111110011010110", -- t[31958] = 3
      "0000011" when "00111110011010111", -- t[31959] = 3
      "0000011" when "00111110011011000", -- t[31960] = 3
      "0000011" when "00111110011011001", -- t[31961] = 3
      "0000011" when "00111110011011010", -- t[31962] = 3
      "0000011" when "00111110011011011", -- t[31963] = 3
      "0000011" when "00111110011011100", -- t[31964] = 3
      "0000011" when "00111110011011101", -- t[31965] = 3
      "0000011" when "00111110011011110", -- t[31966] = 3
      "0000011" when "00111110011011111", -- t[31967] = 3
      "0000011" when "00111110011100000", -- t[31968] = 3
      "0000011" when "00111110011100001", -- t[31969] = 3
      "0000011" when "00111110011100010", -- t[31970] = 3
      "0000011" when "00111110011100011", -- t[31971] = 3
      "0000011" when "00111110011100100", -- t[31972] = 3
      "0000011" when "00111110011100101", -- t[31973] = 3
      "0000011" when "00111110011100110", -- t[31974] = 3
      "0000011" when "00111110011100111", -- t[31975] = 3
      "0000011" when "00111110011101000", -- t[31976] = 3
      "0000011" when "00111110011101001", -- t[31977] = 3
      "0000011" when "00111110011101010", -- t[31978] = 3
      "0000011" when "00111110011101011", -- t[31979] = 3
      "0000011" when "00111110011101100", -- t[31980] = 3
      "0000011" when "00111110011101101", -- t[31981] = 3
      "0000011" when "00111110011101110", -- t[31982] = 3
      "0000011" when "00111110011101111", -- t[31983] = 3
      "0000011" when "00111110011110000", -- t[31984] = 3
      "0000011" when "00111110011110001", -- t[31985] = 3
      "0000011" when "00111110011110010", -- t[31986] = 3
      "0000011" when "00111110011110011", -- t[31987] = 3
      "0000011" when "00111110011110100", -- t[31988] = 3
      "0000011" when "00111110011110101", -- t[31989] = 3
      "0000011" when "00111110011110110", -- t[31990] = 3
      "0000011" when "00111110011110111", -- t[31991] = 3
      "0000011" when "00111110011111000", -- t[31992] = 3
      "0000011" when "00111110011111001", -- t[31993] = 3
      "0000011" when "00111110011111010", -- t[31994] = 3
      "0000011" when "00111110011111011", -- t[31995] = 3
      "0000011" when "00111110011111100", -- t[31996] = 3
      "0000011" when "00111110011111101", -- t[31997] = 3
      "0000011" when "00111110011111110", -- t[31998] = 3
      "0000011" when "00111110011111111", -- t[31999] = 3
      "0000011" when "00111110100000000", -- t[32000] = 3
      "0000011" when "00111110100000001", -- t[32001] = 3
      "0000011" when "00111110100000010", -- t[32002] = 3
      "0000011" when "00111110100000011", -- t[32003] = 3
      "0000011" when "00111110100000100", -- t[32004] = 3
      "0000011" when "00111110100000101", -- t[32005] = 3
      "0000011" when "00111110100000110", -- t[32006] = 3
      "0000011" when "00111110100000111", -- t[32007] = 3
      "0000011" when "00111110100001000", -- t[32008] = 3
      "0000011" when "00111110100001001", -- t[32009] = 3
      "0000011" when "00111110100001010", -- t[32010] = 3
      "0000011" when "00111110100001011", -- t[32011] = 3
      "0000011" when "00111110100001100", -- t[32012] = 3
      "0000011" when "00111110100001101", -- t[32013] = 3
      "0000011" when "00111110100001110", -- t[32014] = 3
      "0000011" when "00111110100001111", -- t[32015] = 3
      "0000011" when "00111110100010000", -- t[32016] = 3
      "0000011" when "00111110100010001", -- t[32017] = 3
      "0000011" when "00111110100010010", -- t[32018] = 3
      "0000011" when "00111110100010011", -- t[32019] = 3
      "0000011" when "00111110100010100", -- t[32020] = 3
      "0000011" when "00111110100010101", -- t[32021] = 3
      "0000011" when "00111110100010110", -- t[32022] = 3
      "0000011" when "00111110100010111", -- t[32023] = 3
      "0000011" when "00111110100011000", -- t[32024] = 3
      "0000011" when "00111110100011001", -- t[32025] = 3
      "0000011" when "00111110100011010", -- t[32026] = 3
      "0000011" when "00111110100011011", -- t[32027] = 3
      "0000011" when "00111110100011100", -- t[32028] = 3
      "0000011" when "00111110100011101", -- t[32029] = 3
      "0000011" when "00111110100011110", -- t[32030] = 3
      "0000011" when "00111110100011111", -- t[32031] = 3
      "0000011" when "00111110100100000", -- t[32032] = 3
      "0000011" when "00111110100100001", -- t[32033] = 3
      "0000011" when "00111110100100010", -- t[32034] = 3
      "0000011" when "00111110100100011", -- t[32035] = 3
      "0000011" when "00111110100100100", -- t[32036] = 3
      "0000011" when "00111110100100101", -- t[32037] = 3
      "0000011" when "00111110100100110", -- t[32038] = 3
      "0000011" when "00111110100100111", -- t[32039] = 3
      "0000011" when "00111110100101000", -- t[32040] = 3
      "0000011" when "00111110100101001", -- t[32041] = 3
      "0000011" when "00111110100101010", -- t[32042] = 3
      "0000011" when "00111110100101011", -- t[32043] = 3
      "0000011" when "00111110100101100", -- t[32044] = 3
      "0000011" when "00111110100101101", -- t[32045] = 3
      "0000011" when "00111110100101110", -- t[32046] = 3
      "0000011" when "00111110100101111", -- t[32047] = 3
      "0000011" when "00111110100110000", -- t[32048] = 3
      "0000011" when "00111110100110001", -- t[32049] = 3
      "0000011" when "00111110100110010", -- t[32050] = 3
      "0000011" when "00111110100110011", -- t[32051] = 3
      "0000011" when "00111110100110100", -- t[32052] = 3
      "0000011" when "00111110100110101", -- t[32053] = 3
      "0000011" when "00111110100110110", -- t[32054] = 3
      "0000011" when "00111110100110111", -- t[32055] = 3
      "0000011" when "00111110100111000", -- t[32056] = 3
      "0000011" when "00111110100111001", -- t[32057] = 3
      "0000011" when "00111110100111010", -- t[32058] = 3
      "0000011" when "00111110100111011", -- t[32059] = 3
      "0000011" when "00111110100111100", -- t[32060] = 3
      "0000011" when "00111110100111101", -- t[32061] = 3
      "0000011" when "00111110100111110", -- t[32062] = 3
      "0000011" when "00111110100111111", -- t[32063] = 3
      "0000011" when "00111110101000000", -- t[32064] = 3
      "0000011" when "00111110101000001", -- t[32065] = 3
      "0000011" when "00111110101000010", -- t[32066] = 3
      "0000011" when "00111110101000011", -- t[32067] = 3
      "0000011" when "00111110101000100", -- t[32068] = 3
      "0000011" when "00111110101000101", -- t[32069] = 3
      "0000011" when "00111110101000110", -- t[32070] = 3
      "0000011" when "00111110101000111", -- t[32071] = 3
      "0000011" when "00111110101001000", -- t[32072] = 3
      "0000011" when "00111110101001001", -- t[32073] = 3
      "0000011" when "00111110101001010", -- t[32074] = 3
      "0000011" when "00111110101001011", -- t[32075] = 3
      "0000011" when "00111110101001100", -- t[32076] = 3
      "0000011" when "00111110101001101", -- t[32077] = 3
      "0000011" when "00111110101001110", -- t[32078] = 3
      "0000011" when "00111110101001111", -- t[32079] = 3
      "0000011" when "00111110101010000", -- t[32080] = 3
      "0000011" when "00111110101010001", -- t[32081] = 3
      "0000011" when "00111110101010010", -- t[32082] = 3
      "0000011" when "00111110101010011", -- t[32083] = 3
      "0000011" when "00111110101010100", -- t[32084] = 3
      "0000011" when "00111110101010101", -- t[32085] = 3
      "0000011" when "00111110101010110", -- t[32086] = 3
      "0000011" when "00111110101010111", -- t[32087] = 3
      "0000011" when "00111110101011000", -- t[32088] = 3
      "0000011" when "00111110101011001", -- t[32089] = 3
      "0000011" when "00111110101011010", -- t[32090] = 3
      "0000011" when "00111110101011011", -- t[32091] = 3
      "0000011" when "00111110101011100", -- t[32092] = 3
      "0000011" when "00111110101011101", -- t[32093] = 3
      "0000011" when "00111110101011110", -- t[32094] = 3
      "0000011" when "00111110101011111", -- t[32095] = 3
      "0000011" when "00111110101100000", -- t[32096] = 3
      "0000011" when "00111110101100001", -- t[32097] = 3
      "0000011" when "00111110101100010", -- t[32098] = 3
      "0000011" when "00111110101100011", -- t[32099] = 3
      "0000011" when "00111110101100100", -- t[32100] = 3
      "0000011" when "00111110101100101", -- t[32101] = 3
      "0000011" when "00111110101100110", -- t[32102] = 3
      "0000011" when "00111110101100111", -- t[32103] = 3
      "0000011" when "00111110101101000", -- t[32104] = 3
      "0000011" when "00111110101101001", -- t[32105] = 3
      "0000011" when "00111110101101010", -- t[32106] = 3
      "0000011" when "00111110101101011", -- t[32107] = 3
      "0000011" when "00111110101101100", -- t[32108] = 3
      "0000011" when "00111110101101101", -- t[32109] = 3
      "0000011" when "00111110101101110", -- t[32110] = 3
      "0000011" when "00111110101101111", -- t[32111] = 3
      "0000011" when "00111110101110000", -- t[32112] = 3
      "0000011" when "00111110101110001", -- t[32113] = 3
      "0000011" when "00111110101110010", -- t[32114] = 3
      "0000011" when "00111110101110011", -- t[32115] = 3
      "0000011" when "00111110101110100", -- t[32116] = 3
      "0000011" when "00111110101110101", -- t[32117] = 3
      "0000011" when "00111110101110110", -- t[32118] = 3
      "0000011" when "00111110101110111", -- t[32119] = 3
      "0000011" when "00111110101111000", -- t[32120] = 3
      "0000011" when "00111110101111001", -- t[32121] = 3
      "0000011" when "00111110101111010", -- t[32122] = 3
      "0000011" when "00111110101111011", -- t[32123] = 3
      "0000011" when "00111110101111100", -- t[32124] = 3
      "0000011" when "00111110101111101", -- t[32125] = 3
      "0000011" when "00111110101111110", -- t[32126] = 3
      "0000011" when "00111110101111111", -- t[32127] = 3
      "0000011" when "00111110110000000", -- t[32128] = 3
      "0000011" when "00111110110000001", -- t[32129] = 3
      "0000011" when "00111110110000010", -- t[32130] = 3
      "0000011" when "00111110110000011", -- t[32131] = 3
      "0000011" when "00111110110000100", -- t[32132] = 3
      "0000011" when "00111110110000101", -- t[32133] = 3
      "0000011" when "00111110110000110", -- t[32134] = 3
      "0000011" when "00111110110000111", -- t[32135] = 3
      "0000011" when "00111110110001000", -- t[32136] = 3
      "0000011" when "00111110110001001", -- t[32137] = 3
      "0000011" when "00111110110001010", -- t[32138] = 3
      "0000011" when "00111110110001011", -- t[32139] = 3
      "0000011" when "00111110110001100", -- t[32140] = 3
      "0000011" when "00111110110001101", -- t[32141] = 3
      "0000011" when "00111110110001110", -- t[32142] = 3
      "0000011" when "00111110110001111", -- t[32143] = 3
      "0000011" when "00111110110010000", -- t[32144] = 3
      "0000011" when "00111110110010001", -- t[32145] = 3
      "0000011" when "00111110110010010", -- t[32146] = 3
      "0000011" when "00111110110010011", -- t[32147] = 3
      "0000011" when "00111110110010100", -- t[32148] = 3
      "0000011" when "00111110110010101", -- t[32149] = 3
      "0000011" when "00111110110010110", -- t[32150] = 3
      "0000011" when "00111110110010111", -- t[32151] = 3
      "0000011" when "00111110110011000", -- t[32152] = 3
      "0000011" when "00111110110011001", -- t[32153] = 3
      "0000011" when "00111110110011010", -- t[32154] = 3
      "0000011" when "00111110110011011", -- t[32155] = 3
      "0000011" when "00111110110011100", -- t[32156] = 3
      "0000011" when "00111110110011101", -- t[32157] = 3
      "0000011" when "00111110110011110", -- t[32158] = 3
      "0000011" when "00111110110011111", -- t[32159] = 3
      "0000011" when "00111110110100000", -- t[32160] = 3
      "0000011" when "00111110110100001", -- t[32161] = 3
      "0000011" when "00111110110100010", -- t[32162] = 3
      "0000011" when "00111110110100011", -- t[32163] = 3
      "0000011" when "00111110110100100", -- t[32164] = 3
      "0000011" when "00111110110100101", -- t[32165] = 3
      "0000011" when "00111110110100110", -- t[32166] = 3
      "0000011" when "00111110110100111", -- t[32167] = 3
      "0000011" when "00111110110101000", -- t[32168] = 3
      "0000011" when "00111110110101001", -- t[32169] = 3
      "0000011" when "00111110110101010", -- t[32170] = 3
      "0000011" when "00111110110101011", -- t[32171] = 3
      "0000011" when "00111110110101100", -- t[32172] = 3
      "0000011" when "00111110110101101", -- t[32173] = 3
      "0000011" when "00111110110101110", -- t[32174] = 3
      "0000011" when "00111110110101111", -- t[32175] = 3
      "0000011" when "00111110110110000", -- t[32176] = 3
      "0000011" when "00111110110110001", -- t[32177] = 3
      "0000011" when "00111110110110010", -- t[32178] = 3
      "0000011" when "00111110110110011", -- t[32179] = 3
      "0000011" when "00111110110110100", -- t[32180] = 3
      "0000011" when "00111110110110101", -- t[32181] = 3
      "0000011" when "00111110110110110", -- t[32182] = 3
      "0000011" when "00111110110110111", -- t[32183] = 3
      "0000011" when "00111110110111000", -- t[32184] = 3
      "0000011" when "00111110110111001", -- t[32185] = 3
      "0000011" when "00111110110111010", -- t[32186] = 3
      "0000011" when "00111110110111011", -- t[32187] = 3
      "0000011" when "00111110110111100", -- t[32188] = 3
      "0000011" when "00111110110111101", -- t[32189] = 3
      "0000011" when "00111110110111110", -- t[32190] = 3
      "0000011" when "00111110110111111", -- t[32191] = 3
      "0000011" when "00111110111000000", -- t[32192] = 3
      "0000011" when "00111110111000001", -- t[32193] = 3
      "0000011" when "00111110111000010", -- t[32194] = 3
      "0000011" when "00111110111000011", -- t[32195] = 3
      "0000011" when "00111110111000100", -- t[32196] = 3
      "0000011" when "00111110111000101", -- t[32197] = 3
      "0000011" when "00111110111000110", -- t[32198] = 3
      "0000011" when "00111110111000111", -- t[32199] = 3
      "0000011" when "00111110111001000", -- t[32200] = 3
      "0000011" when "00111110111001001", -- t[32201] = 3
      "0000011" when "00111110111001010", -- t[32202] = 3
      "0000011" when "00111110111001011", -- t[32203] = 3
      "0000011" when "00111110111001100", -- t[32204] = 3
      "0000011" when "00111110111001101", -- t[32205] = 3
      "0000011" when "00111110111001110", -- t[32206] = 3
      "0000011" when "00111110111001111", -- t[32207] = 3
      "0000011" when "00111110111010000", -- t[32208] = 3
      "0000011" when "00111110111010001", -- t[32209] = 3
      "0000011" when "00111110111010010", -- t[32210] = 3
      "0000011" when "00111110111010011", -- t[32211] = 3
      "0000011" when "00111110111010100", -- t[32212] = 3
      "0000011" when "00111110111010101", -- t[32213] = 3
      "0000011" when "00111110111010110", -- t[32214] = 3
      "0000011" when "00111110111010111", -- t[32215] = 3
      "0000011" when "00111110111011000", -- t[32216] = 3
      "0000011" when "00111110111011001", -- t[32217] = 3
      "0000011" when "00111110111011010", -- t[32218] = 3
      "0000011" when "00111110111011011", -- t[32219] = 3
      "0000011" when "00111110111011100", -- t[32220] = 3
      "0000011" when "00111110111011101", -- t[32221] = 3
      "0000011" when "00111110111011110", -- t[32222] = 3
      "0000011" when "00111110111011111", -- t[32223] = 3
      "0000011" when "00111110111100000", -- t[32224] = 3
      "0000011" when "00111110111100001", -- t[32225] = 3
      "0000011" when "00111110111100010", -- t[32226] = 3
      "0000011" when "00111110111100011", -- t[32227] = 3
      "0000011" when "00111110111100100", -- t[32228] = 3
      "0000011" when "00111110111100101", -- t[32229] = 3
      "0000011" when "00111110111100110", -- t[32230] = 3
      "0000011" when "00111110111100111", -- t[32231] = 3
      "0000011" when "00111110111101000", -- t[32232] = 3
      "0000011" when "00111110111101001", -- t[32233] = 3
      "0000011" when "00111110111101010", -- t[32234] = 3
      "0000011" when "00111110111101011", -- t[32235] = 3
      "0000011" when "00111110111101100", -- t[32236] = 3
      "0000011" when "00111110111101101", -- t[32237] = 3
      "0000011" when "00111110111101110", -- t[32238] = 3
      "0000011" when "00111110111101111", -- t[32239] = 3
      "0000011" when "00111110111110000", -- t[32240] = 3
      "0000011" when "00111110111110001", -- t[32241] = 3
      "0000011" when "00111110111110010", -- t[32242] = 3
      "0000011" when "00111110111110011", -- t[32243] = 3
      "0000011" when "00111110111110100", -- t[32244] = 3
      "0000011" when "00111110111110101", -- t[32245] = 3
      "0000011" when "00111110111110110", -- t[32246] = 3
      "0000011" when "00111110111110111", -- t[32247] = 3
      "0000011" when "00111110111111000", -- t[32248] = 3
      "0000011" when "00111110111111001", -- t[32249] = 3
      "0000011" when "00111110111111010", -- t[32250] = 3
      "0000011" when "00111110111111011", -- t[32251] = 3
      "0000011" when "00111110111111100", -- t[32252] = 3
      "0000011" when "00111110111111101", -- t[32253] = 3
      "0000011" when "00111110111111110", -- t[32254] = 3
      "0000011" when "00111110111111111", -- t[32255] = 3
      "0000011" when "00111111000000000", -- t[32256] = 3
      "0000011" when "00111111000000001", -- t[32257] = 3
      "0000011" when "00111111000000010", -- t[32258] = 3
      "0000011" when "00111111000000011", -- t[32259] = 3
      "0000011" when "00111111000000100", -- t[32260] = 3
      "0000011" when "00111111000000101", -- t[32261] = 3
      "0000011" when "00111111000000110", -- t[32262] = 3
      "0000011" when "00111111000000111", -- t[32263] = 3
      "0000011" when "00111111000001000", -- t[32264] = 3
      "0000011" when "00111111000001001", -- t[32265] = 3
      "0000011" when "00111111000001010", -- t[32266] = 3
      "0000011" when "00111111000001011", -- t[32267] = 3
      "0000011" when "00111111000001100", -- t[32268] = 3
      "0000011" when "00111111000001101", -- t[32269] = 3
      "0000011" when "00111111000001110", -- t[32270] = 3
      "0000011" when "00111111000001111", -- t[32271] = 3
      "0000011" when "00111111000010000", -- t[32272] = 3
      "0000011" when "00111111000010001", -- t[32273] = 3
      "0000011" when "00111111000010010", -- t[32274] = 3
      "0000011" when "00111111000010011", -- t[32275] = 3
      "0000011" when "00111111000010100", -- t[32276] = 3
      "0000011" when "00111111000010101", -- t[32277] = 3
      "0000011" when "00111111000010110", -- t[32278] = 3
      "0000011" when "00111111000010111", -- t[32279] = 3
      "0000011" when "00111111000011000", -- t[32280] = 3
      "0000011" when "00111111000011001", -- t[32281] = 3
      "0000011" when "00111111000011010", -- t[32282] = 3
      "0000011" when "00111111000011011", -- t[32283] = 3
      "0000011" when "00111111000011100", -- t[32284] = 3
      "0000011" when "00111111000011101", -- t[32285] = 3
      "0000011" when "00111111000011110", -- t[32286] = 3
      "0000011" when "00111111000011111", -- t[32287] = 3
      "0000011" when "00111111000100000", -- t[32288] = 3
      "0000011" when "00111111000100001", -- t[32289] = 3
      "0000011" when "00111111000100010", -- t[32290] = 3
      "0000011" when "00111111000100011", -- t[32291] = 3
      "0000011" when "00111111000100100", -- t[32292] = 3
      "0000011" when "00111111000100101", -- t[32293] = 3
      "0000011" when "00111111000100110", -- t[32294] = 3
      "0000011" when "00111111000100111", -- t[32295] = 3
      "0000011" when "00111111000101000", -- t[32296] = 3
      "0000011" when "00111111000101001", -- t[32297] = 3
      "0000011" when "00111111000101010", -- t[32298] = 3
      "0000011" when "00111111000101011", -- t[32299] = 3
      "0000011" when "00111111000101100", -- t[32300] = 3
      "0000011" when "00111111000101101", -- t[32301] = 3
      "0000011" when "00111111000101110", -- t[32302] = 3
      "0000011" when "00111111000101111", -- t[32303] = 3
      "0000011" when "00111111000110000", -- t[32304] = 3
      "0000011" when "00111111000110001", -- t[32305] = 3
      "0000011" when "00111111000110010", -- t[32306] = 3
      "0000011" when "00111111000110011", -- t[32307] = 3
      "0000011" when "00111111000110100", -- t[32308] = 3
      "0000011" when "00111111000110101", -- t[32309] = 3
      "0000011" when "00111111000110110", -- t[32310] = 3
      "0000011" when "00111111000110111", -- t[32311] = 3
      "0000011" when "00111111000111000", -- t[32312] = 3
      "0000011" when "00111111000111001", -- t[32313] = 3
      "0000011" when "00111111000111010", -- t[32314] = 3
      "0000011" when "00111111000111011", -- t[32315] = 3
      "0000011" when "00111111000111100", -- t[32316] = 3
      "0000011" when "00111111000111101", -- t[32317] = 3
      "0000011" when "00111111000111110", -- t[32318] = 3
      "0000011" when "00111111000111111", -- t[32319] = 3
      "0000011" when "00111111001000000", -- t[32320] = 3
      "0000011" when "00111111001000001", -- t[32321] = 3
      "0000011" when "00111111001000010", -- t[32322] = 3
      "0000011" when "00111111001000011", -- t[32323] = 3
      "0000011" when "00111111001000100", -- t[32324] = 3
      "0000011" when "00111111001000101", -- t[32325] = 3
      "0000011" when "00111111001000110", -- t[32326] = 3
      "0000011" when "00111111001000111", -- t[32327] = 3
      "0000011" when "00111111001001000", -- t[32328] = 3
      "0000011" when "00111111001001001", -- t[32329] = 3
      "0000011" when "00111111001001010", -- t[32330] = 3
      "0000011" when "00111111001001011", -- t[32331] = 3
      "0000011" when "00111111001001100", -- t[32332] = 3
      "0000011" when "00111111001001101", -- t[32333] = 3
      "0000011" when "00111111001001110", -- t[32334] = 3
      "0000011" when "00111111001001111", -- t[32335] = 3
      "0000011" when "00111111001010000", -- t[32336] = 3
      "0000011" when "00111111001010001", -- t[32337] = 3
      "0000011" when "00111111001010010", -- t[32338] = 3
      "0000011" when "00111111001010011", -- t[32339] = 3
      "0000011" when "00111111001010100", -- t[32340] = 3
      "0000011" when "00111111001010101", -- t[32341] = 3
      "0000011" when "00111111001010110", -- t[32342] = 3
      "0000011" when "00111111001010111", -- t[32343] = 3
      "0000011" when "00111111001011000", -- t[32344] = 3
      "0000011" when "00111111001011001", -- t[32345] = 3
      "0000011" when "00111111001011010", -- t[32346] = 3
      "0000011" when "00111111001011011", -- t[32347] = 3
      "0000011" when "00111111001011100", -- t[32348] = 3
      "0000011" when "00111111001011101", -- t[32349] = 3
      "0000011" when "00111111001011110", -- t[32350] = 3
      "0000011" when "00111111001011111", -- t[32351] = 3
      "0000011" when "00111111001100000", -- t[32352] = 3
      "0000011" when "00111111001100001", -- t[32353] = 3
      "0000011" when "00111111001100010", -- t[32354] = 3
      "0000011" when "00111111001100011", -- t[32355] = 3
      "0000011" when "00111111001100100", -- t[32356] = 3
      "0000011" when "00111111001100101", -- t[32357] = 3
      "0000011" when "00111111001100110", -- t[32358] = 3
      "0000011" when "00111111001100111", -- t[32359] = 3
      "0000011" when "00111111001101000", -- t[32360] = 3
      "0000011" when "00111111001101001", -- t[32361] = 3
      "0000011" when "00111111001101010", -- t[32362] = 3
      "0000011" when "00111111001101011", -- t[32363] = 3
      "0000011" when "00111111001101100", -- t[32364] = 3
      "0000011" when "00111111001101101", -- t[32365] = 3
      "0000011" when "00111111001101110", -- t[32366] = 3
      "0000011" when "00111111001101111", -- t[32367] = 3
      "0000011" when "00111111001110000", -- t[32368] = 3
      "0000011" when "00111111001110001", -- t[32369] = 3
      "0000011" when "00111111001110010", -- t[32370] = 3
      "0000011" when "00111111001110011", -- t[32371] = 3
      "0000011" when "00111111001110100", -- t[32372] = 3
      "0000011" when "00111111001110101", -- t[32373] = 3
      "0000011" when "00111111001110110", -- t[32374] = 3
      "0000011" when "00111111001110111", -- t[32375] = 3
      "0000011" when "00111111001111000", -- t[32376] = 3
      "0000011" when "00111111001111001", -- t[32377] = 3
      "0000011" when "00111111001111010", -- t[32378] = 3
      "0000011" when "00111111001111011", -- t[32379] = 3
      "0000011" when "00111111001111100", -- t[32380] = 3
      "0000011" when "00111111001111101", -- t[32381] = 3
      "0000011" when "00111111001111110", -- t[32382] = 3
      "0000011" when "00111111001111111", -- t[32383] = 3
      "0000011" when "00111111010000000", -- t[32384] = 3
      "0000011" when "00111111010000001", -- t[32385] = 3
      "0000011" when "00111111010000010", -- t[32386] = 3
      "0000011" when "00111111010000011", -- t[32387] = 3
      "0000011" when "00111111010000100", -- t[32388] = 3
      "0000011" when "00111111010000101", -- t[32389] = 3
      "0000011" when "00111111010000110", -- t[32390] = 3
      "0000011" when "00111111010000111", -- t[32391] = 3
      "0000011" when "00111111010001000", -- t[32392] = 3
      "0000011" when "00111111010001001", -- t[32393] = 3
      "0000011" when "00111111010001010", -- t[32394] = 3
      "0000011" when "00111111010001011", -- t[32395] = 3
      "0000011" when "00111111010001100", -- t[32396] = 3
      "0000011" when "00111111010001101", -- t[32397] = 3
      "0000011" when "00111111010001110", -- t[32398] = 3
      "0000011" when "00111111010001111", -- t[32399] = 3
      "0000011" when "00111111010010000", -- t[32400] = 3
      "0000011" when "00111111010010001", -- t[32401] = 3
      "0000011" when "00111111010010010", -- t[32402] = 3
      "0000011" when "00111111010010011", -- t[32403] = 3
      "0000011" when "00111111010010100", -- t[32404] = 3
      "0000011" when "00111111010010101", -- t[32405] = 3
      "0000011" when "00111111010010110", -- t[32406] = 3
      "0000011" when "00111111010010111", -- t[32407] = 3
      "0000011" when "00111111010011000", -- t[32408] = 3
      "0000011" when "00111111010011001", -- t[32409] = 3
      "0000011" when "00111111010011010", -- t[32410] = 3
      "0000011" when "00111111010011011", -- t[32411] = 3
      "0000011" when "00111111010011100", -- t[32412] = 3
      "0000011" when "00111111010011101", -- t[32413] = 3
      "0000011" when "00111111010011110", -- t[32414] = 3
      "0000011" when "00111111010011111", -- t[32415] = 3
      "0000011" when "00111111010100000", -- t[32416] = 3
      "0000011" when "00111111010100001", -- t[32417] = 3
      "0000011" when "00111111010100010", -- t[32418] = 3
      "0000011" when "00111111010100011", -- t[32419] = 3
      "0000011" when "00111111010100100", -- t[32420] = 3
      "0000011" when "00111111010100101", -- t[32421] = 3
      "0000011" when "00111111010100110", -- t[32422] = 3
      "0000011" when "00111111010100111", -- t[32423] = 3
      "0000011" when "00111111010101000", -- t[32424] = 3
      "0000011" when "00111111010101001", -- t[32425] = 3
      "0000011" when "00111111010101010", -- t[32426] = 3
      "0000011" when "00111111010101011", -- t[32427] = 3
      "0000011" when "00111111010101100", -- t[32428] = 3
      "0000011" when "00111111010101101", -- t[32429] = 3
      "0000011" when "00111111010101110", -- t[32430] = 3
      "0000011" when "00111111010101111", -- t[32431] = 3
      "0000011" when "00111111010110000", -- t[32432] = 3
      "0000011" when "00111111010110001", -- t[32433] = 3
      "0000011" when "00111111010110010", -- t[32434] = 3
      "0000011" when "00111111010110011", -- t[32435] = 3
      "0000011" when "00111111010110100", -- t[32436] = 3
      "0000011" when "00111111010110101", -- t[32437] = 3
      "0000011" when "00111111010110110", -- t[32438] = 3
      "0000011" when "00111111010110111", -- t[32439] = 3
      "0000011" when "00111111010111000", -- t[32440] = 3
      "0000011" when "00111111010111001", -- t[32441] = 3
      "0000011" when "00111111010111010", -- t[32442] = 3
      "0000011" when "00111111010111011", -- t[32443] = 3
      "0000011" when "00111111010111100", -- t[32444] = 3
      "0000011" when "00111111010111101", -- t[32445] = 3
      "0000011" when "00111111010111110", -- t[32446] = 3
      "0000011" when "00111111010111111", -- t[32447] = 3
      "0000011" when "00111111011000000", -- t[32448] = 3
      "0000011" when "00111111011000001", -- t[32449] = 3
      "0000011" when "00111111011000010", -- t[32450] = 3
      "0000011" when "00111111011000011", -- t[32451] = 3
      "0000011" when "00111111011000100", -- t[32452] = 3
      "0000011" when "00111111011000101", -- t[32453] = 3
      "0000011" when "00111111011000110", -- t[32454] = 3
      "0000011" when "00111111011000111", -- t[32455] = 3
      "0000011" when "00111111011001000", -- t[32456] = 3
      "0000011" when "00111111011001001", -- t[32457] = 3
      "0000011" when "00111111011001010", -- t[32458] = 3
      "0000011" when "00111111011001011", -- t[32459] = 3
      "0000011" when "00111111011001100", -- t[32460] = 3
      "0000011" when "00111111011001101", -- t[32461] = 3
      "0000011" when "00111111011001110", -- t[32462] = 3
      "0000011" when "00111111011001111", -- t[32463] = 3
      "0000011" when "00111111011010000", -- t[32464] = 3
      "0000011" when "00111111011010001", -- t[32465] = 3
      "0000011" when "00111111011010010", -- t[32466] = 3
      "0000011" when "00111111011010011", -- t[32467] = 3
      "0000011" when "00111111011010100", -- t[32468] = 3
      "0000011" when "00111111011010101", -- t[32469] = 3
      "0000011" when "00111111011010110", -- t[32470] = 3
      "0000011" when "00111111011010111", -- t[32471] = 3
      "0000011" when "00111111011011000", -- t[32472] = 3
      "0000011" when "00111111011011001", -- t[32473] = 3
      "0000011" when "00111111011011010", -- t[32474] = 3
      "0000011" when "00111111011011011", -- t[32475] = 3
      "0000011" when "00111111011011100", -- t[32476] = 3
      "0000011" when "00111111011011101", -- t[32477] = 3
      "0000011" when "00111111011011110", -- t[32478] = 3
      "0000011" when "00111111011011111", -- t[32479] = 3
      "0000011" when "00111111011100000", -- t[32480] = 3
      "0000011" when "00111111011100001", -- t[32481] = 3
      "0000011" when "00111111011100010", -- t[32482] = 3
      "0000011" when "00111111011100011", -- t[32483] = 3
      "0000011" when "00111111011100100", -- t[32484] = 3
      "0000011" when "00111111011100101", -- t[32485] = 3
      "0000011" when "00111111011100110", -- t[32486] = 3
      "0000011" when "00111111011100111", -- t[32487] = 3
      "0000011" when "00111111011101000", -- t[32488] = 3
      "0000011" when "00111111011101001", -- t[32489] = 3
      "0000011" when "00111111011101010", -- t[32490] = 3
      "0000011" when "00111111011101011", -- t[32491] = 3
      "0000011" when "00111111011101100", -- t[32492] = 3
      "0000011" when "00111111011101101", -- t[32493] = 3
      "0000011" when "00111111011101110", -- t[32494] = 3
      "0000011" when "00111111011101111", -- t[32495] = 3
      "0000011" when "00111111011110000", -- t[32496] = 3
      "0000011" when "00111111011110001", -- t[32497] = 3
      "0000011" when "00111111011110010", -- t[32498] = 3
      "0000011" when "00111111011110011", -- t[32499] = 3
      "0000011" when "00111111011110100", -- t[32500] = 3
      "0000011" when "00111111011110101", -- t[32501] = 3
      "0000011" when "00111111011110110", -- t[32502] = 3
      "0000011" when "00111111011110111", -- t[32503] = 3
      "0000011" when "00111111011111000", -- t[32504] = 3
      "0000011" when "00111111011111001", -- t[32505] = 3
      "0000011" when "00111111011111010", -- t[32506] = 3
      "0000011" when "00111111011111011", -- t[32507] = 3
      "0000011" when "00111111011111100", -- t[32508] = 3
      "0000011" when "00111111011111101", -- t[32509] = 3
      "0000011" when "00111111011111110", -- t[32510] = 3
      "0000011" when "00111111011111111", -- t[32511] = 3
      "0000011" when "00111111100000000", -- t[32512] = 3
      "0000011" when "00111111100000001", -- t[32513] = 3
      "0000011" when "00111111100000010", -- t[32514] = 3
      "0000011" when "00111111100000011", -- t[32515] = 3
      "0000011" when "00111111100000100", -- t[32516] = 3
      "0000011" when "00111111100000101", -- t[32517] = 3
      "0000011" when "00111111100000110", -- t[32518] = 3
      "0000011" when "00111111100000111", -- t[32519] = 3
      "0000011" when "00111111100001000", -- t[32520] = 3
      "0000011" when "00111111100001001", -- t[32521] = 3
      "0000011" when "00111111100001010", -- t[32522] = 3
      "0000011" when "00111111100001011", -- t[32523] = 3
      "0000011" when "00111111100001100", -- t[32524] = 3
      "0000011" when "00111111100001101", -- t[32525] = 3
      "0000011" when "00111111100001110", -- t[32526] = 3
      "0000011" when "00111111100001111", -- t[32527] = 3
      "0000011" when "00111111100010000", -- t[32528] = 3
      "0000011" when "00111111100010001", -- t[32529] = 3
      "0000011" when "00111111100010010", -- t[32530] = 3
      "0000011" when "00111111100010011", -- t[32531] = 3
      "0000011" when "00111111100010100", -- t[32532] = 3
      "0000011" when "00111111100010101", -- t[32533] = 3
      "0000011" when "00111111100010110", -- t[32534] = 3
      "0000011" when "00111111100010111", -- t[32535] = 3
      "0000011" when "00111111100011000", -- t[32536] = 3
      "0000011" when "00111111100011001", -- t[32537] = 3
      "0000011" when "00111111100011010", -- t[32538] = 3
      "0000011" when "00111111100011011", -- t[32539] = 3
      "0000011" when "00111111100011100", -- t[32540] = 3
      "0000011" when "00111111100011101", -- t[32541] = 3
      "0000011" when "00111111100011110", -- t[32542] = 3
      "0000011" when "00111111100011111", -- t[32543] = 3
      "0000011" when "00111111100100000", -- t[32544] = 3
      "0000011" when "00111111100100001", -- t[32545] = 3
      "0000011" when "00111111100100010", -- t[32546] = 3
      "0000011" when "00111111100100011", -- t[32547] = 3
      "0000011" when "00111111100100100", -- t[32548] = 3
      "0000011" when "00111111100100101", -- t[32549] = 3
      "0000011" when "00111111100100110", -- t[32550] = 3
      "0000011" when "00111111100100111", -- t[32551] = 3
      "0000011" when "00111111100101000", -- t[32552] = 3
      "0000011" when "00111111100101001", -- t[32553] = 3
      "0000011" when "00111111100101010", -- t[32554] = 3
      "0000011" when "00111111100101011", -- t[32555] = 3
      "0000011" when "00111111100101100", -- t[32556] = 3
      "0000011" when "00111111100101101", -- t[32557] = 3
      "0000011" when "00111111100101110", -- t[32558] = 3
      "0000011" when "00111111100101111", -- t[32559] = 3
      "0000011" when "00111111100110000", -- t[32560] = 3
      "0000011" when "00111111100110001", -- t[32561] = 3
      "0000011" when "00111111100110010", -- t[32562] = 3
      "0000011" when "00111111100110011", -- t[32563] = 3
      "0000011" when "00111111100110100", -- t[32564] = 3
      "0000011" when "00111111100110101", -- t[32565] = 3
      "0000011" when "00111111100110110", -- t[32566] = 3
      "0000011" when "00111111100110111", -- t[32567] = 3
      "0000011" when "00111111100111000", -- t[32568] = 3
      "0000011" when "00111111100111001", -- t[32569] = 3
      "0000011" when "00111111100111010", -- t[32570] = 3
      "0000011" when "00111111100111011", -- t[32571] = 3
      "0000011" when "00111111100111100", -- t[32572] = 3
      "0000011" when "00111111100111101", -- t[32573] = 3
      "0000011" when "00111111100111110", -- t[32574] = 3
      "0000011" when "00111111100111111", -- t[32575] = 3
      "0000011" when "00111111101000000", -- t[32576] = 3
      "0000011" when "00111111101000001", -- t[32577] = 3
      "0000011" when "00111111101000010", -- t[32578] = 3
      "0000011" when "00111111101000011", -- t[32579] = 3
      "0000011" when "00111111101000100", -- t[32580] = 3
      "0000011" when "00111111101000101", -- t[32581] = 3
      "0000011" when "00111111101000110", -- t[32582] = 3
      "0000011" when "00111111101000111", -- t[32583] = 3
      "0000011" when "00111111101001000", -- t[32584] = 3
      "0000011" when "00111111101001001", -- t[32585] = 3
      "0000011" when "00111111101001010", -- t[32586] = 3
      "0000011" when "00111111101001011", -- t[32587] = 3
      "0000011" when "00111111101001100", -- t[32588] = 3
      "0000011" when "00111111101001101", -- t[32589] = 3
      "0000011" when "00111111101001110", -- t[32590] = 3
      "0000011" when "00111111101001111", -- t[32591] = 3
      "0000011" when "00111111101010000", -- t[32592] = 3
      "0000011" when "00111111101010001", -- t[32593] = 3
      "0000011" when "00111111101010010", -- t[32594] = 3
      "0000011" when "00111111101010011", -- t[32595] = 3
      "0000011" when "00111111101010100", -- t[32596] = 3
      "0000011" when "00111111101010101", -- t[32597] = 3
      "0000011" when "00111111101010110", -- t[32598] = 3
      "0000011" when "00111111101010111", -- t[32599] = 3
      "0000011" when "00111111101011000", -- t[32600] = 3
      "0000011" when "00111111101011001", -- t[32601] = 3
      "0000011" when "00111111101011010", -- t[32602] = 3
      "0000011" when "00111111101011011", -- t[32603] = 3
      "0000011" when "00111111101011100", -- t[32604] = 3
      "0000011" when "00111111101011101", -- t[32605] = 3
      "0000011" when "00111111101011110", -- t[32606] = 3
      "0000011" when "00111111101011111", -- t[32607] = 3
      "0000011" when "00111111101100000", -- t[32608] = 3
      "0000011" when "00111111101100001", -- t[32609] = 3
      "0000011" when "00111111101100010", -- t[32610] = 3
      "0000011" when "00111111101100011", -- t[32611] = 3
      "0000011" when "00111111101100100", -- t[32612] = 3
      "0000011" when "00111111101100101", -- t[32613] = 3
      "0000011" when "00111111101100110", -- t[32614] = 3
      "0000011" when "00111111101100111", -- t[32615] = 3
      "0000011" when "00111111101101000", -- t[32616] = 3
      "0000011" when "00111111101101001", -- t[32617] = 3
      "0000011" when "00111111101101010", -- t[32618] = 3
      "0000011" when "00111111101101011", -- t[32619] = 3
      "0000011" when "00111111101101100", -- t[32620] = 3
      "0000011" when "00111111101101101", -- t[32621] = 3
      "0000011" when "00111111101101110", -- t[32622] = 3
      "0000011" when "00111111101101111", -- t[32623] = 3
      "0000011" when "00111111101110000", -- t[32624] = 3
      "0000011" when "00111111101110001", -- t[32625] = 3
      "0000011" when "00111111101110010", -- t[32626] = 3
      "0000011" when "00111111101110011", -- t[32627] = 3
      "0000011" when "00111111101110100", -- t[32628] = 3
      "0000011" when "00111111101110101", -- t[32629] = 3
      "0000011" when "00111111101110110", -- t[32630] = 3
      "0000011" when "00111111101110111", -- t[32631] = 3
      "0000011" when "00111111101111000", -- t[32632] = 3
      "0000011" when "00111111101111001", -- t[32633] = 3
      "0000011" when "00111111101111010", -- t[32634] = 3
      "0000011" when "00111111101111011", -- t[32635] = 3
      "0000011" when "00111111101111100", -- t[32636] = 3
      "0000011" when "00111111101111101", -- t[32637] = 3
      "0000011" when "00111111101111110", -- t[32638] = 3
      "0000011" when "00111111101111111", -- t[32639] = 3
      "0000011" when "00111111110000000", -- t[32640] = 3
      "0000011" when "00111111110000001", -- t[32641] = 3
      "0000011" when "00111111110000010", -- t[32642] = 3
      "0000011" when "00111111110000011", -- t[32643] = 3
      "0000011" when "00111111110000100", -- t[32644] = 3
      "0000011" when "00111111110000101", -- t[32645] = 3
      "0000011" when "00111111110000110", -- t[32646] = 3
      "0000011" when "00111111110000111", -- t[32647] = 3
      "0000011" when "00111111110001000", -- t[32648] = 3
      "0000011" when "00111111110001001", -- t[32649] = 3
      "0000011" when "00111111110001010", -- t[32650] = 3
      "0000011" when "00111111110001011", -- t[32651] = 3
      "0000011" when "00111111110001100", -- t[32652] = 3
      "0000011" when "00111111110001101", -- t[32653] = 3
      "0000011" when "00111111110001110", -- t[32654] = 3
      "0000011" when "00111111110001111", -- t[32655] = 3
      "0000011" when "00111111110010000", -- t[32656] = 3
      "0000011" when "00111111110010001", -- t[32657] = 3
      "0000011" when "00111111110010010", -- t[32658] = 3
      "0000011" when "00111111110010011", -- t[32659] = 3
      "0000011" when "00111111110010100", -- t[32660] = 3
      "0000011" when "00111111110010101", -- t[32661] = 3
      "0000011" when "00111111110010110", -- t[32662] = 3
      "0000011" when "00111111110010111", -- t[32663] = 3
      "0000011" when "00111111110011000", -- t[32664] = 3
      "0000011" when "00111111110011001", -- t[32665] = 3
      "0000011" when "00111111110011010", -- t[32666] = 3
      "0000011" when "00111111110011011", -- t[32667] = 3
      "0000011" when "00111111110011100", -- t[32668] = 3
      "0000011" when "00111111110011101", -- t[32669] = 3
      "0000011" when "00111111110011110", -- t[32670] = 3
      "0000011" when "00111111110011111", -- t[32671] = 3
      "0000011" when "00111111110100000", -- t[32672] = 3
      "0000011" when "00111111110100001", -- t[32673] = 3
      "0000011" when "00111111110100010", -- t[32674] = 3
      "0000011" when "00111111110100011", -- t[32675] = 3
      "0000011" when "00111111110100100", -- t[32676] = 3
      "0000011" when "00111111110100101", -- t[32677] = 3
      "0000011" when "00111111110100110", -- t[32678] = 3
      "0000011" when "00111111110100111", -- t[32679] = 3
      "0000011" when "00111111110101000", -- t[32680] = 3
      "0000011" when "00111111110101001", -- t[32681] = 3
      "0000011" when "00111111110101010", -- t[32682] = 3
      "0000011" when "00111111110101011", -- t[32683] = 3
      "0000011" when "00111111110101100", -- t[32684] = 3
      "0000011" when "00111111110101101", -- t[32685] = 3
      "0000011" when "00111111110101110", -- t[32686] = 3
      "0000011" when "00111111110101111", -- t[32687] = 3
      "0000011" when "00111111110110000", -- t[32688] = 3
      "0000011" when "00111111110110001", -- t[32689] = 3
      "0000011" when "00111111110110010", -- t[32690] = 3
      "0000011" when "00111111110110011", -- t[32691] = 3
      "0000011" when "00111111110110100", -- t[32692] = 3
      "0000011" when "00111111110110101", -- t[32693] = 3
      "0000011" when "00111111110110110", -- t[32694] = 3
      "0000011" when "00111111110110111", -- t[32695] = 3
      "0000011" when "00111111110111000", -- t[32696] = 3
      "0000011" when "00111111110111001", -- t[32697] = 3
      "0000011" when "00111111110111010", -- t[32698] = 3
      "0000011" when "00111111110111011", -- t[32699] = 3
      "0000011" when "00111111110111100", -- t[32700] = 3
      "0000011" when "00111111110111101", -- t[32701] = 3
      "0000011" when "00111111110111110", -- t[32702] = 3
      "0000011" when "00111111110111111", -- t[32703] = 3
      "0000011" when "00111111111000000", -- t[32704] = 3
      "0000011" when "00111111111000001", -- t[32705] = 3
      "0000011" when "00111111111000010", -- t[32706] = 3
      "0000011" when "00111111111000011", -- t[32707] = 3
      "0000011" when "00111111111000100", -- t[32708] = 3
      "0000011" when "00111111111000101", -- t[32709] = 3
      "0000011" when "00111111111000110", -- t[32710] = 3
      "0000011" when "00111111111000111", -- t[32711] = 3
      "0000011" when "00111111111001000", -- t[32712] = 3
      "0000011" when "00111111111001001", -- t[32713] = 3
      "0000011" when "00111111111001010", -- t[32714] = 3
      "0000011" when "00111111111001011", -- t[32715] = 3
      "0000011" when "00111111111001100", -- t[32716] = 3
      "0000011" when "00111111111001101", -- t[32717] = 3
      "0000011" when "00111111111001110", -- t[32718] = 3
      "0000011" when "00111111111001111", -- t[32719] = 3
      "0000011" when "00111111111010000", -- t[32720] = 3
      "0000011" when "00111111111010001", -- t[32721] = 3
      "0000011" when "00111111111010010", -- t[32722] = 3
      "0000011" when "00111111111010011", -- t[32723] = 3
      "0000011" when "00111111111010100", -- t[32724] = 3
      "0000011" when "00111111111010101", -- t[32725] = 3
      "0000011" when "00111111111010110", -- t[32726] = 3
      "0000011" when "00111111111010111", -- t[32727] = 3
      "0000011" when "00111111111011000", -- t[32728] = 3
      "0000011" when "00111111111011001", -- t[32729] = 3
      "0000011" when "00111111111011010", -- t[32730] = 3
      "0000011" when "00111111111011011", -- t[32731] = 3
      "0000011" when "00111111111011100", -- t[32732] = 3
      "0000011" when "00111111111011101", -- t[32733] = 3
      "0000011" when "00111111111011110", -- t[32734] = 3
      "0000011" when "00111111111011111", -- t[32735] = 3
      "0000011" when "00111111111100000", -- t[32736] = 3
      "0000011" when "00111111111100001", -- t[32737] = 3
      "0000011" when "00111111111100010", -- t[32738] = 3
      "0000011" when "00111111111100011", -- t[32739] = 3
      "0000011" when "00111111111100100", -- t[32740] = 3
      "0000011" when "00111111111100101", -- t[32741] = 3
      "0000011" when "00111111111100110", -- t[32742] = 3
      "0000011" when "00111111111100111", -- t[32743] = 3
      "0000011" when "00111111111101000", -- t[32744] = 3
      "0000011" when "00111111111101001", -- t[32745] = 3
      "0000011" when "00111111111101010", -- t[32746] = 3
      "0000011" when "00111111111101011", -- t[32747] = 3
      "0000011" when "00111111111101100", -- t[32748] = 3
      "0000011" when "00111111111101101", -- t[32749] = 3
      "0000011" when "00111111111101110", -- t[32750] = 3
      "0000011" when "00111111111101111", -- t[32751] = 3
      "0000011" when "00111111111110000", -- t[32752] = 3
      "0000011" when "00111111111110001", -- t[32753] = 3
      "0000011" when "00111111111110010", -- t[32754] = 3
      "0000011" when "00111111111110011", -- t[32755] = 3
      "0000011" when "00111111111110100", -- t[32756] = 3
      "0000011" when "00111111111110101", -- t[32757] = 3
      "0000011" when "00111111111110110", -- t[32758] = 3
      "0000011" when "00111111111110111", -- t[32759] = 3
      "0000011" when "00111111111111000", -- t[32760] = 3
      "0000011" when "00111111111111001", -- t[32761] = 3
      "0000011" when "00111111111111010", -- t[32762] = 3
      "0000011" when "00111111111111011", -- t[32763] = 3
      "0000011" when "00111111111111100", -- t[32764] = 3
      "0000011" when "00111111111111101", -- t[32765] = 3
      "0000011" when "00111111111111110", -- t[32766] = 3
      "0000011" when "00111111111111111", -- t[32767] = 3
      "0000011" when "01000000000000000", -- t[32768] = 3
      "0000011" when "01000000000000001", -- t[32769] = 3
      "0000011" when "01000000000000010", -- t[32770] = 3
      "0000011" when "01000000000000011", -- t[32771] = 3
      "0000011" when "01000000000000100", -- t[32772] = 3
      "0000011" when "01000000000000101", -- t[32773] = 3
      "0000011" when "01000000000000110", -- t[32774] = 3
      "0000011" when "01000000000000111", -- t[32775] = 3
      "0000011" when "01000000000001000", -- t[32776] = 3
      "0000011" when "01000000000001001", -- t[32777] = 3
      "0000011" when "01000000000001010", -- t[32778] = 3
      "0000011" when "01000000000001011", -- t[32779] = 3
      "0000011" when "01000000000001100", -- t[32780] = 3
      "0000011" when "01000000000001101", -- t[32781] = 3
      "0000011" when "01000000000001110", -- t[32782] = 3
      "0000011" when "01000000000001111", -- t[32783] = 3
      "0000011" when "01000000000010000", -- t[32784] = 3
      "0000011" when "01000000000010001", -- t[32785] = 3
      "0000011" when "01000000000010010", -- t[32786] = 3
      "0000011" when "01000000000010011", -- t[32787] = 3
      "0000011" when "01000000000010100", -- t[32788] = 3
      "0000011" when "01000000000010101", -- t[32789] = 3
      "0000011" when "01000000000010110", -- t[32790] = 3
      "0000011" when "01000000000010111", -- t[32791] = 3
      "0000011" when "01000000000011000", -- t[32792] = 3
      "0000011" when "01000000000011001", -- t[32793] = 3
      "0000011" when "01000000000011010", -- t[32794] = 3
      "0000011" when "01000000000011011", -- t[32795] = 3
      "0000011" when "01000000000011100", -- t[32796] = 3
      "0000011" when "01000000000011101", -- t[32797] = 3
      "0000011" when "01000000000011110", -- t[32798] = 3
      "0000011" when "01000000000011111", -- t[32799] = 3
      "0000011" when "01000000000100000", -- t[32800] = 3
      "0000011" when "01000000000100001", -- t[32801] = 3
      "0000011" when "01000000000100010", -- t[32802] = 3
      "0000011" when "01000000000100011", -- t[32803] = 3
      "0000011" when "01000000000100100", -- t[32804] = 3
      "0000011" when "01000000000100101", -- t[32805] = 3
      "0000011" when "01000000000100110", -- t[32806] = 3
      "0000011" when "01000000000100111", -- t[32807] = 3
      "0000011" when "01000000000101000", -- t[32808] = 3
      "0000011" when "01000000000101001", -- t[32809] = 3
      "0000011" when "01000000000101010", -- t[32810] = 3
      "0000011" when "01000000000101011", -- t[32811] = 3
      "0000011" when "01000000000101100", -- t[32812] = 3
      "0000011" when "01000000000101101", -- t[32813] = 3
      "0000011" when "01000000000101110", -- t[32814] = 3
      "0000011" when "01000000000101111", -- t[32815] = 3
      "0000011" when "01000000000110000", -- t[32816] = 3
      "0000011" when "01000000000110001", -- t[32817] = 3
      "0000011" when "01000000000110010", -- t[32818] = 3
      "0000011" when "01000000000110011", -- t[32819] = 3
      "0000011" when "01000000000110100", -- t[32820] = 3
      "0000011" when "01000000000110101", -- t[32821] = 3
      "0000011" when "01000000000110110", -- t[32822] = 3
      "0000011" when "01000000000110111", -- t[32823] = 3
      "0000011" when "01000000000111000", -- t[32824] = 3
      "0000011" when "01000000000111001", -- t[32825] = 3
      "0000011" when "01000000000111010", -- t[32826] = 3
      "0000011" when "01000000000111011", -- t[32827] = 3
      "0000011" when "01000000000111100", -- t[32828] = 3
      "0000011" when "01000000000111101", -- t[32829] = 3
      "0000011" when "01000000000111110", -- t[32830] = 3
      "0000011" when "01000000000111111", -- t[32831] = 3
      "0000011" when "01000000001000000", -- t[32832] = 3
      "0000011" when "01000000001000001", -- t[32833] = 3
      "0000011" when "01000000001000010", -- t[32834] = 3
      "0000011" when "01000000001000011", -- t[32835] = 3
      "0000011" when "01000000001000100", -- t[32836] = 3
      "0000011" when "01000000001000101", -- t[32837] = 3
      "0000011" when "01000000001000110", -- t[32838] = 3
      "0000011" when "01000000001000111", -- t[32839] = 3
      "0000011" when "01000000001001000", -- t[32840] = 3
      "0000011" when "01000000001001001", -- t[32841] = 3
      "0000011" when "01000000001001010", -- t[32842] = 3
      "0000011" when "01000000001001011", -- t[32843] = 3
      "0000011" when "01000000001001100", -- t[32844] = 3
      "0000011" when "01000000001001101", -- t[32845] = 3
      "0000011" when "01000000001001110", -- t[32846] = 3
      "0000011" when "01000000001001111", -- t[32847] = 3
      "0000011" when "01000000001010000", -- t[32848] = 3
      "0000011" when "01000000001010001", -- t[32849] = 3
      "0000011" when "01000000001010010", -- t[32850] = 3
      "0000011" when "01000000001010011", -- t[32851] = 3
      "0000011" when "01000000001010100", -- t[32852] = 3
      "0000011" when "01000000001010101", -- t[32853] = 3
      "0000011" when "01000000001010110", -- t[32854] = 3
      "0000011" when "01000000001010111", -- t[32855] = 3
      "0000011" when "01000000001011000", -- t[32856] = 3
      "0000011" when "01000000001011001", -- t[32857] = 3
      "0000011" when "01000000001011010", -- t[32858] = 3
      "0000011" when "01000000001011011", -- t[32859] = 3
      "0000011" when "01000000001011100", -- t[32860] = 3
      "0000011" when "01000000001011101", -- t[32861] = 3
      "0000011" when "01000000001011110", -- t[32862] = 3
      "0000011" when "01000000001011111", -- t[32863] = 3
      "0000011" when "01000000001100000", -- t[32864] = 3
      "0000011" when "01000000001100001", -- t[32865] = 3
      "0000011" when "01000000001100010", -- t[32866] = 3
      "0000011" when "01000000001100011", -- t[32867] = 3
      "0000011" when "01000000001100100", -- t[32868] = 3
      "0000011" when "01000000001100101", -- t[32869] = 3
      "0000011" when "01000000001100110", -- t[32870] = 3
      "0000011" when "01000000001100111", -- t[32871] = 3
      "0000011" when "01000000001101000", -- t[32872] = 3
      "0000011" when "01000000001101001", -- t[32873] = 3
      "0000011" when "01000000001101010", -- t[32874] = 3
      "0000011" when "01000000001101011", -- t[32875] = 3
      "0000011" when "01000000001101100", -- t[32876] = 3
      "0000011" when "01000000001101101", -- t[32877] = 3
      "0000011" when "01000000001101110", -- t[32878] = 3
      "0000011" when "01000000001101111", -- t[32879] = 3
      "0000011" when "01000000001110000", -- t[32880] = 3
      "0000011" when "01000000001110001", -- t[32881] = 3
      "0000011" when "01000000001110010", -- t[32882] = 3
      "0000011" when "01000000001110011", -- t[32883] = 3
      "0000011" when "01000000001110100", -- t[32884] = 3
      "0000011" when "01000000001110101", -- t[32885] = 3
      "0000011" when "01000000001110110", -- t[32886] = 3
      "0000011" when "01000000001110111", -- t[32887] = 3
      "0000011" when "01000000001111000", -- t[32888] = 3
      "0000011" when "01000000001111001", -- t[32889] = 3
      "0000011" when "01000000001111010", -- t[32890] = 3
      "0000011" when "01000000001111011", -- t[32891] = 3
      "0000011" when "01000000001111100", -- t[32892] = 3
      "0000011" when "01000000001111101", -- t[32893] = 3
      "0000011" when "01000000001111110", -- t[32894] = 3
      "0000011" when "01000000001111111", -- t[32895] = 3
      "0000011" when "01000000010000000", -- t[32896] = 3
      "0000011" when "01000000010000001", -- t[32897] = 3
      "0000011" when "01000000010000010", -- t[32898] = 3
      "0000011" when "01000000010000011", -- t[32899] = 3
      "0000011" when "01000000010000100", -- t[32900] = 3
      "0000011" when "01000000010000101", -- t[32901] = 3
      "0000011" when "01000000010000110", -- t[32902] = 3
      "0000011" when "01000000010000111", -- t[32903] = 3
      "0000011" when "01000000010001000", -- t[32904] = 3
      "0000011" when "01000000010001001", -- t[32905] = 3
      "0000011" when "01000000010001010", -- t[32906] = 3
      "0000011" when "01000000010001011", -- t[32907] = 3
      "0000011" when "01000000010001100", -- t[32908] = 3
      "0000011" when "01000000010001101", -- t[32909] = 3
      "0000011" when "01000000010001110", -- t[32910] = 3
      "0000011" when "01000000010001111", -- t[32911] = 3
      "0000011" when "01000000010010000", -- t[32912] = 3
      "0000011" when "01000000010010001", -- t[32913] = 3
      "0000011" when "01000000010010010", -- t[32914] = 3
      "0000011" when "01000000010010011", -- t[32915] = 3
      "0000011" when "01000000010010100", -- t[32916] = 3
      "0000011" when "01000000010010101", -- t[32917] = 3
      "0000011" when "01000000010010110", -- t[32918] = 3
      "0000011" when "01000000010010111", -- t[32919] = 3
      "0000011" when "01000000010011000", -- t[32920] = 3
      "0000011" when "01000000010011001", -- t[32921] = 3
      "0000011" when "01000000010011010", -- t[32922] = 3
      "0000011" when "01000000010011011", -- t[32923] = 3
      "0000011" when "01000000010011100", -- t[32924] = 3
      "0000011" when "01000000010011101", -- t[32925] = 3
      "0000011" when "01000000010011110", -- t[32926] = 3
      "0000011" when "01000000010011111", -- t[32927] = 3
      "0000011" when "01000000010100000", -- t[32928] = 3
      "0000011" when "01000000010100001", -- t[32929] = 3
      "0000011" when "01000000010100010", -- t[32930] = 3
      "0000011" when "01000000010100011", -- t[32931] = 3
      "0000011" when "01000000010100100", -- t[32932] = 3
      "0000011" when "01000000010100101", -- t[32933] = 3
      "0000011" when "01000000010100110", -- t[32934] = 3
      "0000011" when "01000000010100111", -- t[32935] = 3
      "0000011" when "01000000010101000", -- t[32936] = 3
      "0000011" when "01000000010101001", -- t[32937] = 3
      "0000011" when "01000000010101010", -- t[32938] = 3
      "0000011" when "01000000010101011", -- t[32939] = 3
      "0000011" when "01000000010101100", -- t[32940] = 3
      "0000011" when "01000000010101101", -- t[32941] = 3
      "0000011" when "01000000010101110", -- t[32942] = 3
      "0000011" when "01000000010101111", -- t[32943] = 3
      "0000011" when "01000000010110000", -- t[32944] = 3
      "0000011" when "01000000010110001", -- t[32945] = 3
      "0000011" when "01000000010110010", -- t[32946] = 3
      "0000011" when "01000000010110011", -- t[32947] = 3
      "0000011" when "01000000010110100", -- t[32948] = 3
      "0000011" when "01000000010110101", -- t[32949] = 3
      "0000011" when "01000000010110110", -- t[32950] = 3
      "0000011" when "01000000010110111", -- t[32951] = 3
      "0000011" when "01000000010111000", -- t[32952] = 3
      "0000011" when "01000000010111001", -- t[32953] = 3
      "0000011" when "01000000010111010", -- t[32954] = 3
      "0000011" when "01000000010111011", -- t[32955] = 3
      "0000011" when "01000000010111100", -- t[32956] = 3
      "0000011" when "01000000010111101", -- t[32957] = 3
      "0000011" when "01000000010111110", -- t[32958] = 3
      "0000011" when "01000000010111111", -- t[32959] = 3
      "0000011" when "01000000011000000", -- t[32960] = 3
      "0000011" when "01000000011000001", -- t[32961] = 3
      "0000011" when "01000000011000010", -- t[32962] = 3
      "0000011" when "01000000011000011", -- t[32963] = 3
      "0000011" when "01000000011000100", -- t[32964] = 3
      "0000011" when "01000000011000101", -- t[32965] = 3
      "0000011" when "01000000011000110", -- t[32966] = 3
      "0000011" when "01000000011000111", -- t[32967] = 3
      "0000011" when "01000000011001000", -- t[32968] = 3
      "0000011" when "01000000011001001", -- t[32969] = 3
      "0000011" when "01000000011001010", -- t[32970] = 3
      "0000011" when "01000000011001011", -- t[32971] = 3
      "0000011" when "01000000011001100", -- t[32972] = 3
      "0000011" when "01000000011001101", -- t[32973] = 3
      "0000011" when "01000000011001110", -- t[32974] = 3
      "0000011" when "01000000011001111", -- t[32975] = 3
      "0000011" when "01000000011010000", -- t[32976] = 3
      "0000011" when "01000000011010001", -- t[32977] = 3
      "0000011" when "01000000011010010", -- t[32978] = 3
      "0000011" when "01000000011010011", -- t[32979] = 3
      "0000011" when "01000000011010100", -- t[32980] = 3
      "0000011" when "01000000011010101", -- t[32981] = 3
      "0000011" when "01000000011010110", -- t[32982] = 3
      "0000011" when "01000000011010111", -- t[32983] = 3
      "0000011" when "01000000011011000", -- t[32984] = 3
      "0000011" when "01000000011011001", -- t[32985] = 3
      "0000011" when "01000000011011010", -- t[32986] = 3
      "0000011" when "01000000011011011", -- t[32987] = 3
      "0000011" when "01000000011011100", -- t[32988] = 3
      "0000011" when "01000000011011101", -- t[32989] = 3
      "0000011" when "01000000011011110", -- t[32990] = 3
      "0000011" when "01000000011011111", -- t[32991] = 3
      "0000011" when "01000000011100000", -- t[32992] = 3
      "0000011" when "01000000011100001", -- t[32993] = 3
      "0000011" when "01000000011100010", -- t[32994] = 3
      "0000011" when "01000000011100011", -- t[32995] = 3
      "0000011" when "01000000011100100", -- t[32996] = 3
      "0000011" when "01000000011100101", -- t[32997] = 3
      "0000011" when "01000000011100110", -- t[32998] = 3
      "0000011" when "01000000011100111", -- t[32999] = 3
      "0000011" when "01000000011101000", -- t[33000] = 3
      "0000011" when "01000000011101001", -- t[33001] = 3
      "0000011" when "01000000011101010", -- t[33002] = 3
      "0000011" when "01000000011101011", -- t[33003] = 3
      "0000011" when "01000000011101100", -- t[33004] = 3
      "0000011" when "01000000011101101", -- t[33005] = 3
      "0000011" when "01000000011101110", -- t[33006] = 3
      "0000011" when "01000000011101111", -- t[33007] = 3
      "0000011" when "01000000011110000", -- t[33008] = 3
      "0000011" when "01000000011110001", -- t[33009] = 3
      "0000011" when "01000000011110010", -- t[33010] = 3
      "0000011" when "01000000011110011", -- t[33011] = 3
      "0000011" when "01000000011110100", -- t[33012] = 3
      "0000011" when "01000000011110101", -- t[33013] = 3
      "0000011" when "01000000011110110", -- t[33014] = 3
      "0000011" when "01000000011110111", -- t[33015] = 3
      "0000011" when "01000000011111000", -- t[33016] = 3
      "0000011" when "01000000011111001", -- t[33017] = 3
      "0000011" when "01000000011111010", -- t[33018] = 3
      "0000011" when "01000000011111011", -- t[33019] = 3
      "0000011" when "01000000011111100", -- t[33020] = 3
      "0000011" when "01000000011111101", -- t[33021] = 3
      "0000011" when "01000000011111110", -- t[33022] = 3
      "0000011" when "01000000011111111", -- t[33023] = 3
      "0000011" when "01000000100000000", -- t[33024] = 3
      "0000011" when "01000000100000001", -- t[33025] = 3
      "0000011" when "01000000100000010", -- t[33026] = 3
      "0000011" when "01000000100000011", -- t[33027] = 3
      "0000011" when "01000000100000100", -- t[33028] = 3
      "0000011" when "01000000100000101", -- t[33029] = 3
      "0000011" when "01000000100000110", -- t[33030] = 3
      "0000011" when "01000000100000111", -- t[33031] = 3
      "0000011" when "01000000100001000", -- t[33032] = 3
      "0000011" when "01000000100001001", -- t[33033] = 3
      "0000011" when "01000000100001010", -- t[33034] = 3
      "0000011" when "01000000100001011", -- t[33035] = 3
      "0000011" when "01000000100001100", -- t[33036] = 3
      "0000011" when "01000000100001101", -- t[33037] = 3
      "0000011" when "01000000100001110", -- t[33038] = 3
      "0000011" when "01000000100001111", -- t[33039] = 3
      "0000011" when "01000000100010000", -- t[33040] = 3
      "0000011" when "01000000100010001", -- t[33041] = 3
      "0000011" when "01000000100010010", -- t[33042] = 3
      "0000011" when "01000000100010011", -- t[33043] = 3
      "0000011" when "01000000100010100", -- t[33044] = 3
      "0000011" when "01000000100010101", -- t[33045] = 3
      "0000011" when "01000000100010110", -- t[33046] = 3
      "0000011" when "01000000100010111", -- t[33047] = 3
      "0000011" when "01000000100011000", -- t[33048] = 3
      "0000011" when "01000000100011001", -- t[33049] = 3
      "0000011" when "01000000100011010", -- t[33050] = 3
      "0000011" when "01000000100011011", -- t[33051] = 3
      "0000011" when "01000000100011100", -- t[33052] = 3
      "0000011" when "01000000100011101", -- t[33053] = 3
      "0000011" when "01000000100011110", -- t[33054] = 3
      "0000011" when "01000000100011111", -- t[33055] = 3
      "0000011" when "01000000100100000", -- t[33056] = 3
      "0000011" when "01000000100100001", -- t[33057] = 3
      "0000011" when "01000000100100010", -- t[33058] = 3
      "0000011" when "01000000100100011", -- t[33059] = 3
      "0000011" when "01000000100100100", -- t[33060] = 3
      "0000011" when "01000000100100101", -- t[33061] = 3
      "0000011" when "01000000100100110", -- t[33062] = 3
      "0000011" when "01000000100100111", -- t[33063] = 3
      "0000011" when "01000000100101000", -- t[33064] = 3
      "0000011" when "01000000100101001", -- t[33065] = 3
      "0000011" when "01000000100101010", -- t[33066] = 3
      "0000011" when "01000000100101011", -- t[33067] = 3
      "0000011" when "01000000100101100", -- t[33068] = 3
      "0000011" when "01000000100101101", -- t[33069] = 3
      "0000011" when "01000000100101110", -- t[33070] = 3
      "0000011" when "01000000100101111", -- t[33071] = 3
      "0000011" when "01000000100110000", -- t[33072] = 3
      "0000011" when "01000000100110001", -- t[33073] = 3
      "0000011" when "01000000100110010", -- t[33074] = 3
      "0000011" when "01000000100110011", -- t[33075] = 3
      "0000011" when "01000000100110100", -- t[33076] = 3
      "0000011" when "01000000100110101", -- t[33077] = 3
      "0000011" when "01000000100110110", -- t[33078] = 3
      "0000011" when "01000000100110111", -- t[33079] = 3
      "0000011" when "01000000100111000", -- t[33080] = 3
      "0000011" when "01000000100111001", -- t[33081] = 3
      "0000011" when "01000000100111010", -- t[33082] = 3
      "0000011" when "01000000100111011", -- t[33083] = 3
      "0000011" when "01000000100111100", -- t[33084] = 3
      "0000011" when "01000000100111101", -- t[33085] = 3
      "0000011" when "01000000100111110", -- t[33086] = 3
      "0000011" when "01000000100111111", -- t[33087] = 3
      "0000011" when "01000000101000000", -- t[33088] = 3
      "0000011" when "01000000101000001", -- t[33089] = 3
      "0000011" when "01000000101000010", -- t[33090] = 3
      "0000011" when "01000000101000011", -- t[33091] = 3
      "0000011" when "01000000101000100", -- t[33092] = 3
      "0000011" when "01000000101000101", -- t[33093] = 3
      "0000011" when "01000000101000110", -- t[33094] = 3
      "0000011" when "01000000101000111", -- t[33095] = 3
      "0000011" when "01000000101001000", -- t[33096] = 3
      "0000011" when "01000000101001001", -- t[33097] = 3
      "0000011" when "01000000101001010", -- t[33098] = 3
      "0000011" when "01000000101001011", -- t[33099] = 3
      "0000011" when "01000000101001100", -- t[33100] = 3
      "0000011" when "01000000101001101", -- t[33101] = 3
      "0000011" when "01000000101001110", -- t[33102] = 3
      "0000011" when "01000000101001111", -- t[33103] = 3
      "0000011" when "01000000101010000", -- t[33104] = 3
      "0000011" when "01000000101010001", -- t[33105] = 3
      "0000011" when "01000000101010010", -- t[33106] = 3
      "0000011" when "01000000101010011", -- t[33107] = 3
      "0000011" when "01000000101010100", -- t[33108] = 3
      "0000011" when "01000000101010101", -- t[33109] = 3
      "0000011" when "01000000101010110", -- t[33110] = 3
      "0000011" when "01000000101010111", -- t[33111] = 3
      "0000011" when "01000000101011000", -- t[33112] = 3
      "0000011" when "01000000101011001", -- t[33113] = 3
      "0000011" when "01000000101011010", -- t[33114] = 3
      "0000011" when "01000000101011011", -- t[33115] = 3
      "0000011" when "01000000101011100", -- t[33116] = 3
      "0000011" when "01000000101011101", -- t[33117] = 3
      "0000011" when "01000000101011110", -- t[33118] = 3
      "0000011" when "01000000101011111", -- t[33119] = 3
      "0000011" when "01000000101100000", -- t[33120] = 3
      "0000011" when "01000000101100001", -- t[33121] = 3
      "0000011" when "01000000101100010", -- t[33122] = 3
      "0000011" when "01000000101100011", -- t[33123] = 3
      "0000011" when "01000000101100100", -- t[33124] = 3
      "0000011" when "01000000101100101", -- t[33125] = 3
      "0000011" when "01000000101100110", -- t[33126] = 3
      "0000011" when "01000000101100111", -- t[33127] = 3
      "0000011" when "01000000101101000", -- t[33128] = 3
      "0000011" when "01000000101101001", -- t[33129] = 3
      "0000011" when "01000000101101010", -- t[33130] = 3
      "0000011" when "01000000101101011", -- t[33131] = 3
      "0000011" when "01000000101101100", -- t[33132] = 3
      "0000011" when "01000000101101101", -- t[33133] = 3
      "0000011" when "01000000101101110", -- t[33134] = 3
      "0000011" when "01000000101101111", -- t[33135] = 3
      "0000011" when "01000000101110000", -- t[33136] = 3
      "0000011" when "01000000101110001", -- t[33137] = 3
      "0000011" when "01000000101110010", -- t[33138] = 3
      "0000011" when "01000000101110011", -- t[33139] = 3
      "0000011" when "01000000101110100", -- t[33140] = 3
      "0000011" when "01000000101110101", -- t[33141] = 3
      "0000011" when "01000000101110110", -- t[33142] = 3
      "0000011" when "01000000101110111", -- t[33143] = 3
      "0000011" when "01000000101111000", -- t[33144] = 3
      "0000011" when "01000000101111001", -- t[33145] = 3
      "0000011" when "01000000101111010", -- t[33146] = 3
      "0000011" when "01000000101111011", -- t[33147] = 3
      "0000011" when "01000000101111100", -- t[33148] = 3
      "0000011" when "01000000101111101", -- t[33149] = 3
      "0000011" when "01000000101111110", -- t[33150] = 3
      "0000011" when "01000000101111111", -- t[33151] = 3
      "0000011" when "01000000110000000", -- t[33152] = 3
      "0000011" when "01000000110000001", -- t[33153] = 3
      "0000011" when "01000000110000010", -- t[33154] = 3
      "0000011" when "01000000110000011", -- t[33155] = 3
      "0000011" when "01000000110000100", -- t[33156] = 3
      "0000011" when "01000000110000101", -- t[33157] = 3
      "0000011" when "01000000110000110", -- t[33158] = 3
      "0000011" when "01000000110000111", -- t[33159] = 3
      "0000011" when "01000000110001000", -- t[33160] = 3
      "0000011" when "01000000110001001", -- t[33161] = 3
      "0000011" when "01000000110001010", -- t[33162] = 3
      "0000011" when "01000000110001011", -- t[33163] = 3
      "0000011" when "01000000110001100", -- t[33164] = 3
      "0000011" when "01000000110001101", -- t[33165] = 3
      "0000011" when "01000000110001110", -- t[33166] = 3
      "0000011" when "01000000110001111", -- t[33167] = 3
      "0000011" when "01000000110010000", -- t[33168] = 3
      "0000011" when "01000000110010001", -- t[33169] = 3
      "0000011" when "01000000110010010", -- t[33170] = 3
      "0000011" when "01000000110010011", -- t[33171] = 3
      "0000011" when "01000000110010100", -- t[33172] = 3
      "0000011" when "01000000110010101", -- t[33173] = 3
      "0000011" when "01000000110010110", -- t[33174] = 3
      "0000011" when "01000000110010111", -- t[33175] = 3
      "0000011" when "01000000110011000", -- t[33176] = 3
      "0000011" when "01000000110011001", -- t[33177] = 3
      "0000011" when "01000000110011010", -- t[33178] = 3
      "0000011" when "01000000110011011", -- t[33179] = 3
      "0000011" when "01000000110011100", -- t[33180] = 3
      "0000011" when "01000000110011101", -- t[33181] = 3
      "0000011" when "01000000110011110", -- t[33182] = 3
      "0000011" when "01000000110011111", -- t[33183] = 3
      "0000011" when "01000000110100000", -- t[33184] = 3
      "0000011" when "01000000110100001", -- t[33185] = 3
      "0000011" when "01000000110100010", -- t[33186] = 3
      "0000011" when "01000000110100011", -- t[33187] = 3
      "0000011" when "01000000110100100", -- t[33188] = 3
      "0000011" when "01000000110100101", -- t[33189] = 3
      "0000011" when "01000000110100110", -- t[33190] = 3
      "0000011" when "01000000110100111", -- t[33191] = 3
      "0000011" when "01000000110101000", -- t[33192] = 3
      "0000011" when "01000000110101001", -- t[33193] = 3
      "0000011" when "01000000110101010", -- t[33194] = 3
      "0000011" when "01000000110101011", -- t[33195] = 3
      "0000011" when "01000000110101100", -- t[33196] = 3
      "0000011" when "01000000110101101", -- t[33197] = 3
      "0000011" when "01000000110101110", -- t[33198] = 3
      "0000011" when "01000000110101111", -- t[33199] = 3
      "0000011" when "01000000110110000", -- t[33200] = 3
      "0000011" when "01000000110110001", -- t[33201] = 3
      "0000011" when "01000000110110010", -- t[33202] = 3
      "0000011" when "01000000110110011", -- t[33203] = 3
      "0000011" when "01000000110110100", -- t[33204] = 3
      "0000011" when "01000000110110101", -- t[33205] = 3
      "0000011" when "01000000110110110", -- t[33206] = 3
      "0000011" when "01000000110110111", -- t[33207] = 3
      "0000011" when "01000000110111000", -- t[33208] = 3
      "0000011" when "01000000110111001", -- t[33209] = 3
      "0000011" when "01000000110111010", -- t[33210] = 3
      "0000011" when "01000000110111011", -- t[33211] = 3
      "0000011" when "01000000110111100", -- t[33212] = 3
      "0000011" when "01000000110111101", -- t[33213] = 3
      "0000011" when "01000000110111110", -- t[33214] = 3
      "0000011" when "01000000110111111", -- t[33215] = 3
      "0000011" when "01000000111000000", -- t[33216] = 3
      "0000011" when "01000000111000001", -- t[33217] = 3
      "0000011" when "01000000111000010", -- t[33218] = 3
      "0000011" when "01000000111000011", -- t[33219] = 3
      "0000011" when "01000000111000100", -- t[33220] = 3
      "0000011" when "01000000111000101", -- t[33221] = 3
      "0000011" when "01000000111000110", -- t[33222] = 3
      "0000011" when "01000000111000111", -- t[33223] = 3
      "0000011" when "01000000111001000", -- t[33224] = 3
      "0000011" when "01000000111001001", -- t[33225] = 3
      "0000011" when "01000000111001010", -- t[33226] = 3
      "0000011" when "01000000111001011", -- t[33227] = 3
      "0000011" when "01000000111001100", -- t[33228] = 3
      "0000011" when "01000000111001101", -- t[33229] = 3
      "0000011" when "01000000111001110", -- t[33230] = 3
      "0000011" when "01000000111001111", -- t[33231] = 3
      "0000011" when "01000000111010000", -- t[33232] = 3
      "0000011" when "01000000111010001", -- t[33233] = 3
      "0000011" when "01000000111010010", -- t[33234] = 3
      "0000011" when "01000000111010011", -- t[33235] = 3
      "0000011" when "01000000111010100", -- t[33236] = 3
      "0000011" when "01000000111010101", -- t[33237] = 3
      "0000011" when "01000000111010110", -- t[33238] = 3
      "0000011" when "01000000111010111", -- t[33239] = 3
      "0000011" when "01000000111011000", -- t[33240] = 3
      "0000011" when "01000000111011001", -- t[33241] = 3
      "0000011" when "01000000111011010", -- t[33242] = 3
      "0000011" when "01000000111011011", -- t[33243] = 3
      "0000011" when "01000000111011100", -- t[33244] = 3
      "0000011" when "01000000111011101", -- t[33245] = 3
      "0000011" when "01000000111011110", -- t[33246] = 3
      "0000011" when "01000000111011111", -- t[33247] = 3
      "0000011" when "01000000111100000", -- t[33248] = 3
      "0000011" when "01000000111100001", -- t[33249] = 3
      "0000011" when "01000000111100010", -- t[33250] = 3
      "0000011" when "01000000111100011", -- t[33251] = 3
      "0000011" when "01000000111100100", -- t[33252] = 3
      "0000011" when "01000000111100101", -- t[33253] = 3
      "0000011" when "01000000111100110", -- t[33254] = 3
      "0000011" when "01000000111100111", -- t[33255] = 3
      "0000011" when "01000000111101000", -- t[33256] = 3
      "0000011" when "01000000111101001", -- t[33257] = 3
      "0000011" when "01000000111101010", -- t[33258] = 3
      "0000011" when "01000000111101011", -- t[33259] = 3
      "0000011" when "01000000111101100", -- t[33260] = 3
      "0000011" when "01000000111101101", -- t[33261] = 3
      "0000011" when "01000000111101110", -- t[33262] = 3
      "0000011" when "01000000111101111", -- t[33263] = 3
      "0000011" when "01000000111110000", -- t[33264] = 3
      "0000011" when "01000000111110001", -- t[33265] = 3
      "0000011" when "01000000111110010", -- t[33266] = 3
      "0000011" when "01000000111110011", -- t[33267] = 3
      "0000011" when "01000000111110100", -- t[33268] = 3
      "0000011" when "01000000111110101", -- t[33269] = 3
      "0000011" when "01000000111110110", -- t[33270] = 3
      "0000011" when "01000000111110111", -- t[33271] = 3
      "0000011" when "01000000111111000", -- t[33272] = 3
      "0000011" when "01000000111111001", -- t[33273] = 3
      "0000011" when "01000000111111010", -- t[33274] = 3
      "0000011" when "01000000111111011", -- t[33275] = 3
      "0000011" when "01000000111111100", -- t[33276] = 3
      "0000011" when "01000000111111101", -- t[33277] = 3
      "0000011" when "01000000111111110", -- t[33278] = 3
      "0000011" when "01000000111111111", -- t[33279] = 3
      "0000011" when "01000001000000000", -- t[33280] = 3
      "0000011" when "01000001000000001", -- t[33281] = 3
      "0000011" when "01000001000000010", -- t[33282] = 3
      "0000011" when "01000001000000011", -- t[33283] = 3
      "0000011" when "01000001000000100", -- t[33284] = 3
      "0000011" when "01000001000000101", -- t[33285] = 3
      "0000011" when "01000001000000110", -- t[33286] = 3
      "0000011" when "01000001000000111", -- t[33287] = 3
      "0000011" when "01000001000001000", -- t[33288] = 3
      "0000011" when "01000001000001001", -- t[33289] = 3
      "0000011" when "01000001000001010", -- t[33290] = 3
      "0000011" when "01000001000001011", -- t[33291] = 3
      "0000011" when "01000001000001100", -- t[33292] = 3
      "0000011" when "01000001000001101", -- t[33293] = 3
      "0000011" when "01000001000001110", -- t[33294] = 3
      "0000011" when "01000001000001111", -- t[33295] = 3
      "0000011" when "01000001000010000", -- t[33296] = 3
      "0000011" when "01000001000010001", -- t[33297] = 3
      "0000011" when "01000001000010010", -- t[33298] = 3
      "0000011" when "01000001000010011", -- t[33299] = 3
      "0000011" when "01000001000010100", -- t[33300] = 3
      "0000011" when "01000001000010101", -- t[33301] = 3
      "0000011" when "01000001000010110", -- t[33302] = 3
      "0000011" when "01000001000010111", -- t[33303] = 3
      "0000011" when "01000001000011000", -- t[33304] = 3
      "0000011" when "01000001000011001", -- t[33305] = 3
      "0000011" when "01000001000011010", -- t[33306] = 3
      "0000011" when "01000001000011011", -- t[33307] = 3
      "0000011" when "01000001000011100", -- t[33308] = 3
      "0000011" when "01000001000011101", -- t[33309] = 3
      "0000011" when "01000001000011110", -- t[33310] = 3
      "0000011" when "01000001000011111", -- t[33311] = 3
      "0000011" when "01000001000100000", -- t[33312] = 3
      "0000011" when "01000001000100001", -- t[33313] = 3
      "0000011" when "01000001000100010", -- t[33314] = 3
      "0000011" when "01000001000100011", -- t[33315] = 3
      "0000011" when "01000001000100100", -- t[33316] = 3
      "0000011" when "01000001000100101", -- t[33317] = 3
      "0000011" when "01000001000100110", -- t[33318] = 3
      "0000011" when "01000001000100111", -- t[33319] = 3
      "0000011" when "01000001000101000", -- t[33320] = 3
      "0000011" when "01000001000101001", -- t[33321] = 3
      "0000011" when "01000001000101010", -- t[33322] = 3
      "0000011" when "01000001000101011", -- t[33323] = 3
      "0000011" when "01000001000101100", -- t[33324] = 3
      "0000011" when "01000001000101101", -- t[33325] = 3
      "0000011" when "01000001000101110", -- t[33326] = 3
      "0000011" when "01000001000101111", -- t[33327] = 3
      "0000011" when "01000001000110000", -- t[33328] = 3
      "0000011" when "01000001000110001", -- t[33329] = 3
      "0000011" when "01000001000110010", -- t[33330] = 3
      "0000011" when "01000001000110011", -- t[33331] = 3
      "0000011" when "01000001000110100", -- t[33332] = 3
      "0000011" when "01000001000110101", -- t[33333] = 3
      "0000011" when "01000001000110110", -- t[33334] = 3
      "0000011" when "01000001000110111", -- t[33335] = 3
      "0000011" when "01000001000111000", -- t[33336] = 3
      "0000011" when "01000001000111001", -- t[33337] = 3
      "0000011" when "01000001000111010", -- t[33338] = 3
      "0000011" when "01000001000111011", -- t[33339] = 3
      "0000011" when "01000001000111100", -- t[33340] = 3
      "0000011" when "01000001000111101", -- t[33341] = 3
      "0000011" when "01000001000111110", -- t[33342] = 3
      "0000011" when "01000001000111111", -- t[33343] = 3
      "0000011" when "01000001001000000", -- t[33344] = 3
      "0000011" when "01000001001000001", -- t[33345] = 3
      "0000011" when "01000001001000010", -- t[33346] = 3
      "0000011" when "01000001001000011", -- t[33347] = 3
      "0000011" when "01000001001000100", -- t[33348] = 3
      "0000011" when "01000001001000101", -- t[33349] = 3
      "0000011" when "01000001001000110", -- t[33350] = 3
      "0000011" when "01000001001000111", -- t[33351] = 3
      "0000011" when "01000001001001000", -- t[33352] = 3
      "0000011" when "01000001001001001", -- t[33353] = 3
      "0000011" when "01000001001001010", -- t[33354] = 3
      "0000011" when "01000001001001011", -- t[33355] = 3
      "0000011" when "01000001001001100", -- t[33356] = 3
      "0000011" when "01000001001001101", -- t[33357] = 3
      "0000011" when "01000001001001110", -- t[33358] = 3
      "0000011" when "01000001001001111", -- t[33359] = 3
      "0000011" when "01000001001010000", -- t[33360] = 3
      "0000011" when "01000001001010001", -- t[33361] = 3
      "0000011" when "01000001001010010", -- t[33362] = 3
      "0000011" when "01000001001010011", -- t[33363] = 3
      "0000011" when "01000001001010100", -- t[33364] = 3
      "0000011" when "01000001001010101", -- t[33365] = 3
      "0000011" when "01000001001010110", -- t[33366] = 3
      "0000011" when "01000001001010111", -- t[33367] = 3
      "0000011" when "01000001001011000", -- t[33368] = 3
      "0000011" when "01000001001011001", -- t[33369] = 3
      "0000011" when "01000001001011010", -- t[33370] = 3
      "0000011" when "01000001001011011", -- t[33371] = 3
      "0000011" when "01000001001011100", -- t[33372] = 3
      "0000011" when "01000001001011101", -- t[33373] = 3
      "0000011" when "01000001001011110", -- t[33374] = 3
      "0000011" when "01000001001011111", -- t[33375] = 3
      "0000011" when "01000001001100000", -- t[33376] = 3
      "0000011" when "01000001001100001", -- t[33377] = 3
      "0000011" when "01000001001100010", -- t[33378] = 3
      "0000011" when "01000001001100011", -- t[33379] = 3
      "0000011" when "01000001001100100", -- t[33380] = 3
      "0000011" when "01000001001100101", -- t[33381] = 3
      "0000011" when "01000001001100110", -- t[33382] = 3
      "0000011" when "01000001001100111", -- t[33383] = 3
      "0000011" when "01000001001101000", -- t[33384] = 3
      "0000011" when "01000001001101001", -- t[33385] = 3
      "0000011" when "01000001001101010", -- t[33386] = 3
      "0000011" when "01000001001101011", -- t[33387] = 3
      "0000011" when "01000001001101100", -- t[33388] = 3
      "0000011" when "01000001001101101", -- t[33389] = 3
      "0000011" when "01000001001101110", -- t[33390] = 3
      "0000011" when "01000001001101111", -- t[33391] = 3
      "0000011" when "01000001001110000", -- t[33392] = 3
      "0000011" when "01000001001110001", -- t[33393] = 3
      "0000011" when "01000001001110010", -- t[33394] = 3
      "0000011" when "01000001001110011", -- t[33395] = 3
      "0000011" when "01000001001110100", -- t[33396] = 3
      "0000011" when "01000001001110101", -- t[33397] = 3
      "0000011" when "01000001001110110", -- t[33398] = 3
      "0000011" when "01000001001110111", -- t[33399] = 3
      "0000011" when "01000001001111000", -- t[33400] = 3
      "0000011" when "01000001001111001", -- t[33401] = 3
      "0000011" when "01000001001111010", -- t[33402] = 3
      "0000011" when "01000001001111011", -- t[33403] = 3
      "0000011" when "01000001001111100", -- t[33404] = 3
      "0000011" when "01000001001111101", -- t[33405] = 3
      "0000011" when "01000001001111110", -- t[33406] = 3
      "0000011" when "01000001001111111", -- t[33407] = 3
      "0000011" when "01000001010000000", -- t[33408] = 3
      "0000011" when "01000001010000001", -- t[33409] = 3
      "0000011" when "01000001010000010", -- t[33410] = 3
      "0000011" when "01000001010000011", -- t[33411] = 3
      "0000011" when "01000001010000100", -- t[33412] = 3
      "0000011" when "01000001010000101", -- t[33413] = 3
      "0000011" when "01000001010000110", -- t[33414] = 3
      "0000011" when "01000001010000111", -- t[33415] = 3
      "0000011" when "01000001010001000", -- t[33416] = 3
      "0000011" when "01000001010001001", -- t[33417] = 3
      "0000011" when "01000001010001010", -- t[33418] = 3
      "0000011" when "01000001010001011", -- t[33419] = 3
      "0000011" when "01000001010001100", -- t[33420] = 3
      "0000011" when "01000001010001101", -- t[33421] = 3
      "0000011" when "01000001010001110", -- t[33422] = 3
      "0000011" when "01000001010001111", -- t[33423] = 3
      "0000011" when "01000001010010000", -- t[33424] = 3
      "0000011" when "01000001010010001", -- t[33425] = 3
      "0000011" when "01000001010010010", -- t[33426] = 3
      "0000011" when "01000001010010011", -- t[33427] = 3
      "0000011" when "01000001010010100", -- t[33428] = 3
      "0000011" when "01000001010010101", -- t[33429] = 3
      "0000011" when "01000001010010110", -- t[33430] = 3
      "0000011" when "01000001010010111", -- t[33431] = 3
      "0000011" when "01000001010011000", -- t[33432] = 3
      "0000011" when "01000001010011001", -- t[33433] = 3
      "0000011" when "01000001010011010", -- t[33434] = 3
      "0000011" when "01000001010011011", -- t[33435] = 3
      "0000011" when "01000001010011100", -- t[33436] = 3
      "0000011" when "01000001010011101", -- t[33437] = 3
      "0000011" when "01000001010011110", -- t[33438] = 3
      "0000011" when "01000001010011111", -- t[33439] = 3
      "0000011" when "01000001010100000", -- t[33440] = 3
      "0000011" when "01000001010100001", -- t[33441] = 3
      "0000011" when "01000001010100010", -- t[33442] = 3
      "0000011" when "01000001010100011", -- t[33443] = 3
      "0000011" when "01000001010100100", -- t[33444] = 3
      "0000011" when "01000001010100101", -- t[33445] = 3
      "0000011" when "01000001010100110", -- t[33446] = 3
      "0000011" when "01000001010100111", -- t[33447] = 3
      "0000011" when "01000001010101000", -- t[33448] = 3
      "0000011" when "01000001010101001", -- t[33449] = 3
      "0000011" when "01000001010101010", -- t[33450] = 3
      "0000011" when "01000001010101011", -- t[33451] = 3
      "0000011" when "01000001010101100", -- t[33452] = 3
      "0000011" when "01000001010101101", -- t[33453] = 3
      "0000011" when "01000001010101110", -- t[33454] = 3
      "0000011" when "01000001010101111", -- t[33455] = 3
      "0000011" when "01000001010110000", -- t[33456] = 3
      "0000011" when "01000001010110001", -- t[33457] = 3
      "0000011" when "01000001010110010", -- t[33458] = 3
      "0000011" when "01000001010110011", -- t[33459] = 3
      "0000011" when "01000001010110100", -- t[33460] = 3
      "0000011" when "01000001010110101", -- t[33461] = 3
      "0000011" when "01000001010110110", -- t[33462] = 3
      "0000011" when "01000001010110111", -- t[33463] = 3
      "0000011" when "01000001010111000", -- t[33464] = 3
      "0000011" when "01000001010111001", -- t[33465] = 3
      "0000011" when "01000001010111010", -- t[33466] = 3
      "0000011" when "01000001010111011", -- t[33467] = 3
      "0000011" when "01000001010111100", -- t[33468] = 3
      "0000011" when "01000001010111101", -- t[33469] = 3
      "0000011" when "01000001010111110", -- t[33470] = 3
      "0000011" when "01000001010111111", -- t[33471] = 3
      "0000011" when "01000001011000000", -- t[33472] = 3
      "0000011" when "01000001011000001", -- t[33473] = 3
      "0000011" when "01000001011000010", -- t[33474] = 3
      "0000011" when "01000001011000011", -- t[33475] = 3
      "0000011" when "01000001011000100", -- t[33476] = 3
      "0000011" when "01000001011000101", -- t[33477] = 3
      "0000011" when "01000001011000110", -- t[33478] = 3
      "0000011" when "01000001011000111", -- t[33479] = 3
      "0000011" when "01000001011001000", -- t[33480] = 3
      "0000011" when "01000001011001001", -- t[33481] = 3
      "0000011" when "01000001011001010", -- t[33482] = 3
      "0000011" when "01000001011001011", -- t[33483] = 3
      "0000011" when "01000001011001100", -- t[33484] = 3
      "0000011" when "01000001011001101", -- t[33485] = 3
      "0000011" when "01000001011001110", -- t[33486] = 3
      "0000011" when "01000001011001111", -- t[33487] = 3
      "0000011" when "01000001011010000", -- t[33488] = 3
      "0000011" when "01000001011010001", -- t[33489] = 3
      "0000011" when "01000001011010010", -- t[33490] = 3
      "0000011" when "01000001011010011", -- t[33491] = 3
      "0000011" when "01000001011010100", -- t[33492] = 3
      "0000011" when "01000001011010101", -- t[33493] = 3
      "0000011" when "01000001011010110", -- t[33494] = 3
      "0000011" when "01000001011010111", -- t[33495] = 3
      "0000011" when "01000001011011000", -- t[33496] = 3
      "0000011" when "01000001011011001", -- t[33497] = 3
      "0000011" when "01000001011011010", -- t[33498] = 3
      "0000011" when "01000001011011011", -- t[33499] = 3
      "0000011" when "01000001011011100", -- t[33500] = 3
      "0000011" when "01000001011011101", -- t[33501] = 3
      "0000011" when "01000001011011110", -- t[33502] = 3
      "0000011" when "01000001011011111", -- t[33503] = 3
      "0000011" when "01000001011100000", -- t[33504] = 3
      "0000011" when "01000001011100001", -- t[33505] = 3
      "0000011" when "01000001011100010", -- t[33506] = 3
      "0000011" when "01000001011100011", -- t[33507] = 3
      "0000011" when "01000001011100100", -- t[33508] = 3
      "0000011" when "01000001011100101", -- t[33509] = 3
      "0000011" when "01000001011100110", -- t[33510] = 3
      "0000011" when "01000001011100111", -- t[33511] = 3
      "0000011" when "01000001011101000", -- t[33512] = 3
      "0000011" when "01000001011101001", -- t[33513] = 3
      "0000011" when "01000001011101010", -- t[33514] = 3
      "0000011" when "01000001011101011", -- t[33515] = 3
      "0000011" when "01000001011101100", -- t[33516] = 3
      "0000011" when "01000001011101101", -- t[33517] = 3
      "0000011" when "01000001011101110", -- t[33518] = 3
      "0000011" when "01000001011101111", -- t[33519] = 3
      "0000011" when "01000001011110000", -- t[33520] = 3
      "0000011" when "01000001011110001", -- t[33521] = 3
      "0000011" when "01000001011110010", -- t[33522] = 3
      "0000011" when "01000001011110011", -- t[33523] = 3
      "0000011" when "01000001011110100", -- t[33524] = 3
      "0000011" when "01000001011110101", -- t[33525] = 3
      "0000011" when "01000001011110110", -- t[33526] = 3
      "0000011" when "01000001011110111", -- t[33527] = 3
      "0000011" when "01000001011111000", -- t[33528] = 3
      "0000011" when "01000001011111001", -- t[33529] = 3
      "0000011" when "01000001011111010", -- t[33530] = 3
      "0000011" when "01000001011111011", -- t[33531] = 3
      "0000011" when "01000001011111100", -- t[33532] = 3
      "0000011" when "01000001011111101", -- t[33533] = 3
      "0000011" when "01000001011111110", -- t[33534] = 3
      "0000011" when "01000001011111111", -- t[33535] = 3
      "0000011" when "01000001100000000", -- t[33536] = 3
      "0000011" when "01000001100000001", -- t[33537] = 3
      "0000011" when "01000001100000010", -- t[33538] = 3
      "0000011" when "01000001100000011", -- t[33539] = 3
      "0000011" when "01000001100000100", -- t[33540] = 3
      "0000011" when "01000001100000101", -- t[33541] = 3
      "0000011" when "01000001100000110", -- t[33542] = 3
      "0000011" when "01000001100000111", -- t[33543] = 3
      "0000011" when "01000001100001000", -- t[33544] = 3
      "0000011" when "01000001100001001", -- t[33545] = 3
      "0000011" when "01000001100001010", -- t[33546] = 3
      "0000011" when "01000001100001011", -- t[33547] = 3
      "0000011" when "01000001100001100", -- t[33548] = 3
      "0000011" when "01000001100001101", -- t[33549] = 3
      "0000011" when "01000001100001110", -- t[33550] = 3
      "0000011" when "01000001100001111", -- t[33551] = 3
      "0000011" when "01000001100010000", -- t[33552] = 3
      "0000011" when "01000001100010001", -- t[33553] = 3
      "0000011" when "01000001100010010", -- t[33554] = 3
      "0000011" when "01000001100010011", -- t[33555] = 3
      "0000011" when "01000001100010100", -- t[33556] = 3
      "0000011" when "01000001100010101", -- t[33557] = 3
      "0000011" when "01000001100010110", -- t[33558] = 3
      "0000011" when "01000001100010111", -- t[33559] = 3
      "0000011" when "01000001100011000", -- t[33560] = 3
      "0000011" when "01000001100011001", -- t[33561] = 3
      "0000011" when "01000001100011010", -- t[33562] = 3
      "0000011" when "01000001100011011", -- t[33563] = 3
      "0000011" when "01000001100011100", -- t[33564] = 3
      "0000011" when "01000001100011101", -- t[33565] = 3
      "0000011" when "01000001100011110", -- t[33566] = 3
      "0000011" when "01000001100011111", -- t[33567] = 3
      "0000011" when "01000001100100000", -- t[33568] = 3
      "0000011" when "01000001100100001", -- t[33569] = 3
      "0000011" when "01000001100100010", -- t[33570] = 3
      "0000011" when "01000001100100011", -- t[33571] = 3
      "0000011" when "01000001100100100", -- t[33572] = 3
      "0000011" when "01000001100100101", -- t[33573] = 3
      "0000011" when "01000001100100110", -- t[33574] = 3
      "0000011" when "01000001100100111", -- t[33575] = 3
      "0000011" when "01000001100101000", -- t[33576] = 3
      "0000011" when "01000001100101001", -- t[33577] = 3
      "0000011" when "01000001100101010", -- t[33578] = 3
      "0000011" when "01000001100101011", -- t[33579] = 3
      "0000011" when "01000001100101100", -- t[33580] = 3
      "0000011" when "01000001100101101", -- t[33581] = 3
      "0000011" when "01000001100101110", -- t[33582] = 3
      "0000011" when "01000001100101111", -- t[33583] = 3
      "0000011" when "01000001100110000", -- t[33584] = 3
      "0000011" when "01000001100110001", -- t[33585] = 3
      "0000011" when "01000001100110010", -- t[33586] = 3
      "0000011" when "01000001100110011", -- t[33587] = 3
      "0000011" when "01000001100110100", -- t[33588] = 3
      "0000011" when "01000001100110101", -- t[33589] = 3
      "0000011" when "01000001100110110", -- t[33590] = 3
      "0000011" when "01000001100110111", -- t[33591] = 3
      "0000011" when "01000001100111000", -- t[33592] = 3
      "0000011" when "01000001100111001", -- t[33593] = 3
      "0000011" when "01000001100111010", -- t[33594] = 3
      "0000011" when "01000001100111011", -- t[33595] = 3
      "0000011" when "01000001100111100", -- t[33596] = 3
      "0000011" when "01000001100111101", -- t[33597] = 3
      "0000011" when "01000001100111110", -- t[33598] = 3
      "0000011" when "01000001100111111", -- t[33599] = 3
      "0000011" when "01000001101000000", -- t[33600] = 3
      "0000011" when "01000001101000001", -- t[33601] = 3
      "0000011" when "01000001101000010", -- t[33602] = 3
      "0000011" when "01000001101000011", -- t[33603] = 3
      "0000011" when "01000001101000100", -- t[33604] = 3
      "0000011" when "01000001101000101", -- t[33605] = 3
      "0000011" when "01000001101000110", -- t[33606] = 3
      "0000011" when "01000001101000111", -- t[33607] = 3
      "0000011" when "01000001101001000", -- t[33608] = 3
      "0000011" when "01000001101001001", -- t[33609] = 3
      "0000011" when "01000001101001010", -- t[33610] = 3
      "0000011" when "01000001101001011", -- t[33611] = 3
      "0000011" when "01000001101001100", -- t[33612] = 3
      "0000011" when "01000001101001101", -- t[33613] = 3
      "0000011" when "01000001101001110", -- t[33614] = 3
      "0000011" when "01000001101001111", -- t[33615] = 3
      "0000011" when "01000001101010000", -- t[33616] = 3
      "0000011" when "01000001101010001", -- t[33617] = 3
      "0000011" when "01000001101010010", -- t[33618] = 3
      "0000011" when "01000001101010011", -- t[33619] = 3
      "0000011" when "01000001101010100", -- t[33620] = 3
      "0000011" when "01000001101010101", -- t[33621] = 3
      "0000011" when "01000001101010110", -- t[33622] = 3
      "0000011" when "01000001101010111", -- t[33623] = 3
      "0000011" when "01000001101011000", -- t[33624] = 3
      "0000011" when "01000001101011001", -- t[33625] = 3
      "0000011" when "01000001101011010", -- t[33626] = 3
      "0000011" when "01000001101011011", -- t[33627] = 3
      "0000011" when "01000001101011100", -- t[33628] = 3
      "0000011" when "01000001101011101", -- t[33629] = 3
      "0000011" when "01000001101011110", -- t[33630] = 3
      "0000011" when "01000001101011111", -- t[33631] = 3
      "0000011" when "01000001101100000", -- t[33632] = 3
      "0000011" when "01000001101100001", -- t[33633] = 3
      "0000011" when "01000001101100010", -- t[33634] = 3
      "0000011" when "01000001101100011", -- t[33635] = 3
      "0000011" when "01000001101100100", -- t[33636] = 3
      "0000011" when "01000001101100101", -- t[33637] = 3
      "0000011" when "01000001101100110", -- t[33638] = 3
      "0000011" when "01000001101100111", -- t[33639] = 3
      "0000011" when "01000001101101000", -- t[33640] = 3
      "0000011" when "01000001101101001", -- t[33641] = 3
      "0000011" when "01000001101101010", -- t[33642] = 3
      "0000011" when "01000001101101011", -- t[33643] = 3
      "0000011" when "01000001101101100", -- t[33644] = 3
      "0000011" when "01000001101101101", -- t[33645] = 3
      "0000011" when "01000001101101110", -- t[33646] = 3
      "0000011" when "01000001101101111", -- t[33647] = 3
      "0000011" when "01000001101110000", -- t[33648] = 3
      "0000011" when "01000001101110001", -- t[33649] = 3
      "0000011" when "01000001101110010", -- t[33650] = 3
      "0000011" when "01000001101110011", -- t[33651] = 3
      "0000011" when "01000001101110100", -- t[33652] = 3
      "0000011" when "01000001101110101", -- t[33653] = 3
      "0000011" when "01000001101110110", -- t[33654] = 3
      "0000011" when "01000001101110111", -- t[33655] = 3
      "0000011" when "01000001101111000", -- t[33656] = 3
      "0000011" when "01000001101111001", -- t[33657] = 3
      "0000011" when "01000001101111010", -- t[33658] = 3
      "0000011" when "01000001101111011", -- t[33659] = 3
      "0000011" when "01000001101111100", -- t[33660] = 3
      "0000011" when "01000001101111101", -- t[33661] = 3
      "0000011" when "01000001101111110", -- t[33662] = 3
      "0000011" when "01000001101111111", -- t[33663] = 3
      "0000011" when "01000001110000000", -- t[33664] = 3
      "0000011" when "01000001110000001", -- t[33665] = 3
      "0000011" when "01000001110000010", -- t[33666] = 3
      "0000011" when "01000001110000011", -- t[33667] = 3
      "0000011" when "01000001110000100", -- t[33668] = 3
      "0000011" when "01000001110000101", -- t[33669] = 3
      "0000011" when "01000001110000110", -- t[33670] = 3
      "0000011" when "01000001110000111", -- t[33671] = 3
      "0000011" when "01000001110001000", -- t[33672] = 3
      "0000011" when "01000001110001001", -- t[33673] = 3
      "0000011" when "01000001110001010", -- t[33674] = 3
      "0000011" when "01000001110001011", -- t[33675] = 3
      "0000011" when "01000001110001100", -- t[33676] = 3
      "0000011" when "01000001110001101", -- t[33677] = 3
      "0000011" when "01000001110001110", -- t[33678] = 3
      "0000011" when "01000001110001111", -- t[33679] = 3
      "0000011" when "01000001110010000", -- t[33680] = 3
      "0000011" when "01000001110010001", -- t[33681] = 3
      "0000011" when "01000001110010010", -- t[33682] = 3
      "0000011" when "01000001110010011", -- t[33683] = 3
      "0000011" when "01000001110010100", -- t[33684] = 3
      "0000011" when "01000001110010101", -- t[33685] = 3
      "0000011" when "01000001110010110", -- t[33686] = 3
      "0000011" when "01000001110010111", -- t[33687] = 3
      "0000011" when "01000001110011000", -- t[33688] = 3
      "0000011" when "01000001110011001", -- t[33689] = 3
      "0000011" when "01000001110011010", -- t[33690] = 3
      "0000011" when "01000001110011011", -- t[33691] = 3
      "0000011" when "01000001110011100", -- t[33692] = 3
      "0000011" when "01000001110011101", -- t[33693] = 3
      "0000011" when "01000001110011110", -- t[33694] = 3
      "0000011" when "01000001110011111", -- t[33695] = 3
      "0000011" when "01000001110100000", -- t[33696] = 3
      "0000011" when "01000001110100001", -- t[33697] = 3
      "0000011" when "01000001110100010", -- t[33698] = 3
      "0000011" when "01000001110100011", -- t[33699] = 3
      "0000011" when "01000001110100100", -- t[33700] = 3
      "0000011" when "01000001110100101", -- t[33701] = 3
      "0000011" when "01000001110100110", -- t[33702] = 3
      "0000011" when "01000001110100111", -- t[33703] = 3
      "0000011" when "01000001110101000", -- t[33704] = 3
      "0000011" when "01000001110101001", -- t[33705] = 3
      "0000011" when "01000001110101010", -- t[33706] = 3
      "0000011" when "01000001110101011", -- t[33707] = 3
      "0000011" when "01000001110101100", -- t[33708] = 3
      "0000011" when "01000001110101101", -- t[33709] = 3
      "0000011" when "01000001110101110", -- t[33710] = 3
      "0000011" when "01000001110101111", -- t[33711] = 3
      "0000011" when "01000001110110000", -- t[33712] = 3
      "0000011" when "01000001110110001", -- t[33713] = 3
      "0000011" when "01000001110110010", -- t[33714] = 3
      "0000011" when "01000001110110011", -- t[33715] = 3
      "0000011" when "01000001110110100", -- t[33716] = 3
      "0000011" when "01000001110110101", -- t[33717] = 3
      "0000011" when "01000001110110110", -- t[33718] = 3
      "0000011" when "01000001110110111", -- t[33719] = 3
      "0000011" when "01000001110111000", -- t[33720] = 3
      "0000011" when "01000001110111001", -- t[33721] = 3
      "0000011" when "01000001110111010", -- t[33722] = 3
      "0000011" when "01000001110111011", -- t[33723] = 3
      "0000011" when "01000001110111100", -- t[33724] = 3
      "0000011" when "01000001110111101", -- t[33725] = 3
      "0000011" when "01000001110111110", -- t[33726] = 3
      "0000011" when "01000001110111111", -- t[33727] = 3
      "0000011" when "01000001111000000", -- t[33728] = 3
      "0000011" when "01000001111000001", -- t[33729] = 3
      "0000011" when "01000001111000010", -- t[33730] = 3
      "0000011" when "01000001111000011", -- t[33731] = 3
      "0000011" when "01000001111000100", -- t[33732] = 3
      "0000011" when "01000001111000101", -- t[33733] = 3
      "0000011" when "01000001111000110", -- t[33734] = 3
      "0000011" when "01000001111000111", -- t[33735] = 3
      "0000011" when "01000001111001000", -- t[33736] = 3
      "0000011" when "01000001111001001", -- t[33737] = 3
      "0000011" when "01000001111001010", -- t[33738] = 3
      "0000011" when "01000001111001011", -- t[33739] = 3
      "0000011" when "01000001111001100", -- t[33740] = 3
      "0000011" when "01000001111001101", -- t[33741] = 3
      "0000011" when "01000001111001110", -- t[33742] = 3
      "0000011" when "01000001111001111", -- t[33743] = 3
      "0000011" when "01000001111010000", -- t[33744] = 3
      "0000011" when "01000001111010001", -- t[33745] = 3
      "0000011" when "01000001111010010", -- t[33746] = 3
      "0000011" when "01000001111010011", -- t[33747] = 3
      "0000011" when "01000001111010100", -- t[33748] = 3
      "0000011" when "01000001111010101", -- t[33749] = 3
      "0000011" when "01000001111010110", -- t[33750] = 3
      "0000011" when "01000001111010111", -- t[33751] = 3
      "0000011" when "01000001111011000", -- t[33752] = 3
      "0000011" when "01000001111011001", -- t[33753] = 3
      "0000011" when "01000001111011010", -- t[33754] = 3
      "0000011" when "01000001111011011", -- t[33755] = 3
      "0000011" when "01000001111011100", -- t[33756] = 3
      "0000011" when "01000001111011101", -- t[33757] = 3
      "0000011" when "01000001111011110", -- t[33758] = 3
      "0000011" when "01000001111011111", -- t[33759] = 3
      "0000011" when "01000001111100000", -- t[33760] = 3
      "0000011" when "01000001111100001", -- t[33761] = 3
      "0000011" when "01000001111100010", -- t[33762] = 3
      "0000011" when "01000001111100011", -- t[33763] = 3
      "0000011" when "01000001111100100", -- t[33764] = 3
      "0000011" when "01000001111100101", -- t[33765] = 3
      "0000011" when "01000001111100110", -- t[33766] = 3
      "0000011" when "01000001111100111", -- t[33767] = 3
      "0000011" when "01000001111101000", -- t[33768] = 3
      "0000011" when "01000001111101001", -- t[33769] = 3
      "0000011" when "01000001111101010", -- t[33770] = 3
      "0000011" when "01000001111101011", -- t[33771] = 3
      "0000011" when "01000001111101100", -- t[33772] = 3
      "0000011" when "01000001111101101", -- t[33773] = 3
      "0000011" when "01000001111101110", -- t[33774] = 3
      "0000011" when "01000001111101111", -- t[33775] = 3
      "0000011" when "01000001111110000", -- t[33776] = 3
      "0000011" when "01000001111110001", -- t[33777] = 3
      "0000011" when "01000001111110010", -- t[33778] = 3
      "0000011" when "01000001111110011", -- t[33779] = 3
      "0000011" when "01000001111110100", -- t[33780] = 3
      "0000011" when "01000001111110101", -- t[33781] = 3
      "0000011" when "01000001111110110", -- t[33782] = 3
      "0000011" when "01000001111110111", -- t[33783] = 3
      "0000011" when "01000001111111000", -- t[33784] = 3
      "0000011" when "01000001111111001", -- t[33785] = 3
      "0000011" when "01000001111111010", -- t[33786] = 3
      "0000011" when "01000001111111011", -- t[33787] = 3
      "0000011" when "01000001111111100", -- t[33788] = 3
      "0000011" when "01000001111111101", -- t[33789] = 3
      "0000011" when "01000001111111110", -- t[33790] = 3
      "0000011" when "01000001111111111", -- t[33791] = 3
      "0000011" when "01000010000000000", -- t[33792] = 3
      "0000011" when "01000010000000001", -- t[33793] = 3
      "0000011" when "01000010000000010", -- t[33794] = 3
      "0000011" when "01000010000000011", -- t[33795] = 3
      "0000011" when "01000010000000100", -- t[33796] = 3
      "0000011" when "01000010000000101", -- t[33797] = 3
      "0000011" when "01000010000000110", -- t[33798] = 3
      "0000011" when "01000010000000111", -- t[33799] = 3
      "0000011" when "01000010000001000", -- t[33800] = 3
      "0000011" when "01000010000001001", -- t[33801] = 3
      "0000011" when "01000010000001010", -- t[33802] = 3
      "0000011" when "01000010000001011", -- t[33803] = 3
      "0000011" when "01000010000001100", -- t[33804] = 3
      "0000011" when "01000010000001101", -- t[33805] = 3
      "0000011" when "01000010000001110", -- t[33806] = 3
      "0000011" when "01000010000001111", -- t[33807] = 3
      "0000011" when "01000010000010000", -- t[33808] = 3
      "0000011" when "01000010000010001", -- t[33809] = 3
      "0000011" when "01000010000010010", -- t[33810] = 3
      "0000011" when "01000010000010011", -- t[33811] = 3
      "0000011" when "01000010000010100", -- t[33812] = 3
      "0000011" when "01000010000010101", -- t[33813] = 3
      "0000011" when "01000010000010110", -- t[33814] = 3
      "0000011" when "01000010000010111", -- t[33815] = 3
      "0000011" when "01000010000011000", -- t[33816] = 3
      "0000011" when "01000010000011001", -- t[33817] = 3
      "0000011" when "01000010000011010", -- t[33818] = 3
      "0000011" when "01000010000011011", -- t[33819] = 3
      "0000011" when "01000010000011100", -- t[33820] = 3
      "0000011" when "01000010000011101", -- t[33821] = 3
      "0000011" when "01000010000011110", -- t[33822] = 3
      "0000011" when "01000010000011111", -- t[33823] = 3
      "0000011" when "01000010000100000", -- t[33824] = 3
      "0000011" when "01000010000100001", -- t[33825] = 3
      "0000011" when "01000010000100010", -- t[33826] = 3
      "0000011" when "01000010000100011", -- t[33827] = 3
      "0000011" when "01000010000100100", -- t[33828] = 3
      "0000011" when "01000010000100101", -- t[33829] = 3
      "0000011" when "01000010000100110", -- t[33830] = 3
      "0000011" when "01000010000100111", -- t[33831] = 3
      "0000011" when "01000010000101000", -- t[33832] = 3
      "0000011" when "01000010000101001", -- t[33833] = 3
      "0000011" when "01000010000101010", -- t[33834] = 3
      "0000011" when "01000010000101011", -- t[33835] = 3
      "0000011" when "01000010000101100", -- t[33836] = 3
      "0000011" when "01000010000101101", -- t[33837] = 3
      "0000011" when "01000010000101110", -- t[33838] = 3
      "0000011" when "01000010000101111", -- t[33839] = 3
      "0000011" when "01000010000110000", -- t[33840] = 3
      "0000011" when "01000010000110001", -- t[33841] = 3
      "0000011" when "01000010000110010", -- t[33842] = 3
      "0000011" when "01000010000110011", -- t[33843] = 3
      "0000011" when "01000010000110100", -- t[33844] = 3
      "0000011" when "01000010000110101", -- t[33845] = 3
      "0000011" when "01000010000110110", -- t[33846] = 3
      "0000011" when "01000010000110111", -- t[33847] = 3
      "0000011" when "01000010000111000", -- t[33848] = 3
      "0000011" when "01000010000111001", -- t[33849] = 3
      "0000011" when "01000010000111010", -- t[33850] = 3
      "0000011" when "01000010000111011", -- t[33851] = 3
      "0000011" when "01000010000111100", -- t[33852] = 3
      "0000011" when "01000010000111101", -- t[33853] = 3
      "0000011" when "01000010000111110", -- t[33854] = 3
      "0000011" when "01000010000111111", -- t[33855] = 3
      "0000011" when "01000010001000000", -- t[33856] = 3
      "0000011" when "01000010001000001", -- t[33857] = 3
      "0000011" when "01000010001000010", -- t[33858] = 3
      "0000011" when "01000010001000011", -- t[33859] = 3
      "0000011" when "01000010001000100", -- t[33860] = 3
      "0000011" when "01000010001000101", -- t[33861] = 3
      "0000011" when "01000010001000110", -- t[33862] = 3
      "0000011" when "01000010001000111", -- t[33863] = 3
      "0000011" when "01000010001001000", -- t[33864] = 3
      "0000011" when "01000010001001001", -- t[33865] = 3
      "0000011" when "01000010001001010", -- t[33866] = 3
      "0000011" when "01000010001001011", -- t[33867] = 3
      "0000011" when "01000010001001100", -- t[33868] = 3
      "0000011" when "01000010001001101", -- t[33869] = 3
      "0000011" when "01000010001001110", -- t[33870] = 3
      "0000011" when "01000010001001111", -- t[33871] = 3
      "0000011" when "01000010001010000", -- t[33872] = 3
      "0000011" when "01000010001010001", -- t[33873] = 3
      "0000011" when "01000010001010010", -- t[33874] = 3
      "0000011" when "01000010001010011", -- t[33875] = 3
      "0000011" when "01000010001010100", -- t[33876] = 3
      "0000011" when "01000010001010101", -- t[33877] = 3
      "0000011" when "01000010001010110", -- t[33878] = 3
      "0000011" when "01000010001010111", -- t[33879] = 3
      "0000011" when "01000010001011000", -- t[33880] = 3
      "0000011" when "01000010001011001", -- t[33881] = 3
      "0000011" when "01000010001011010", -- t[33882] = 3
      "0000011" when "01000010001011011", -- t[33883] = 3
      "0000011" when "01000010001011100", -- t[33884] = 3
      "0000011" when "01000010001011101", -- t[33885] = 3
      "0000011" when "01000010001011110", -- t[33886] = 3
      "0000011" when "01000010001011111", -- t[33887] = 3
      "0000011" when "01000010001100000", -- t[33888] = 3
      "0000011" when "01000010001100001", -- t[33889] = 3
      "0000011" when "01000010001100010", -- t[33890] = 3
      "0000011" when "01000010001100011", -- t[33891] = 3
      "0000011" when "01000010001100100", -- t[33892] = 3
      "0000011" when "01000010001100101", -- t[33893] = 3
      "0000011" when "01000010001100110", -- t[33894] = 3
      "0000011" when "01000010001100111", -- t[33895] = 3
      "0000011" when "01000010001101000", -- t[33896] = 3
      "0000011" when "01000010001101001", -- t[33897] = 3
      "0000011" when "01000010001101010", -- t[33898] = 3
      "0000011" when "01000010001101011", -- t[33899] = 3
      "0000011" when "01000010001101100", -- t[33900] = 3
      "0000011" when "01000010001101101", -- t[33901] = 3
      "0000011" when "01000010001101110", -- t[33902] = 3
      "0000011" when "01000010001101111", -- t[33903] = 3
      "0000011" when "01000010001110000", -- t[33904] = 3
      "0000011" when "01000010001110001", -- t[33905] = 3
      "0000011" when "01000010001110010", -- t[33906] = 3
      "0000011" when "01000010001110011", -- t[33907] = 3
      "0000011" when "01000010001110100", -- t[33908] = 3
      "0000011" when "01000010001110101", -- t[33909] = 3
      "0000011" when "01000010001110110", -- t[33910] = 3
      "0000011" when "01000010001110111", -- t[33911] = 3
      "0000011" when "01000010001111000", -- t[33912] = 3
      "0000011" when "01000010001111001", -- t[33913] = 3
      "0000011" when "01000010001111010", -- t[33914] = 3
      "0000011" when "01000010001111011", -- t[33915] = 3
      "0000011" when "01000010001111100", -- t[33916] = 3
      "0000011" when "01000010001111101", -- t[33917] = 3
      "0000011" when "01000010001111110", -- t[33918] = 3
      "0000011" when "01000010001111111", -- t[33919] = 3
      "0000011" when "01000010010000000", -- t[33920] = 3
      "0000011" when "01000010010000001", -- t[33921] = 3
      "0000011" when "01000010010000010", -- t[33922] = 3
      "0000011" when "01000010010000011", -- t[33923] = 3
      "0000011" when "01000010010000100", -- t[33924] = 3
      "0000011" when "01000010010000101", -- t[33925] = 3
      "0000011" when "01000010010000110", -- t[33926] = 3
      "0000011" when "01000010010000111", -- t[33927] = 3
      "0000011" when "01000010010001000", -- t[33928] = 3
      "0000011" when "01000010010001001", -- t[33929] = 3
      "0000011" when "01000010010001010", -- t[33930] = 3
      "0000011" when "01000010010001011", -- t[33931] = 3
      "0000011" when "01000010010001100", -- t[33932] = 3
      "0000011" when "01000010010001101", -- t[33933] = 3
      "0000011" when "01000010010001110", -- t[33934] = 3
      "0000011" when "01000010010001111", -- t[33935] = 3
      "0000011" when "01000010010010000", -- t[33936] = 3
      "0000011" when "01000010010010001", -- t[33937] = 3
      "0000011" when "01000010010010010", -- t[33938] = 3
      "0000011" when "01000010010010011", -- t[33939] = 3
      "0000011" when "01000010010010100", -- t[33940] = 3
      "0000011" when "01000010010010101", -- t[33941] = 3
      "0000011" when "01000010010010110", -- t[33942] = 3
      "0000011" when "01000010010010111", -- t[33943] = 3
      "0000011" when "01000010010011000", -- t[33944] = 3
      "0000011" when "01000010010011001", -- t[33945] = 3
      "0000011" when "01000010010011010", -- t[33946] = 3
      "0000011" when "01000010010011011", -- t[33947] = 3
      "0000011" when "01000010010011100", -- t[33948] = 3
      "0000011" when "01000010010011101", -- t[33949] = 3
      "0000011" when "01000010010011110", -- t[33950] = 3
      "0000011" when "01000010010011111", -- t[33951] = 3
      "0000011" when "01000010010100000", -- t[33952] = 3
      "0000011" when "01000010010100001", -- t[33953] = 3
      "0000011" when "01000010010100010", -- t[33954] = 3
      "0000011" when "01000010010100011", -- t[33955] = 3
      "0000011" when "01000010010100100", -- t[33956] = 3
      "0000011" when "01000010010100101", -- t[33957] = 3
      "0000011" when "01000010010100110", -- t[33958] = 3
      "0000011" when "01000010010100111", -- t[33959] = 3
      "0000011" when "01000010010101000", -- t[33960] = 3
      "0000011" when "01000010010101001", -- t[33961] = 3
      "0000011" when "01000010010101010", -- t[33962] = 3
      "0000011" when "01000010010101011", -- t[33963] = 3
      "0000011" when "01000010010101100", -- t[33964] = 3
      "0000011" when "01000010010101101", -- t[33965] = 3
      "0000011" when "01000010010101110", -- t[33966] = 3
      "0000011" when "01000010010101111", -- t[33967] = 3
      "0000011" when "01000010010110000", -- t[33968] = 3
      "0000011" when "01000010010110001", -- t[33969] = 3
      "0000011" when "01000010010110010", -- t[33970] = 3
      "0000011" when "01000010010110011", -- t[33971] = 3
      "0000011" when "01000010010110100", -- t[33972] = 3
      "0000011" when "01000010010110101", -- t[33973] = 3
      "0000011" when "01000010010110110", -- t[33974] = 3
      "0000011" when "01000010010110111", -- t[33975] = 3
      "0000011" when "01000010010111000", -- t[33976] = 3
      "0000011" when "01000010010111001", -- t[33977] = 3
      "0000011" when "01000010010111010", -- t[33978] = 3
      "0000011" when "01000010010111011", -- t[33979] = 3
      "0000011" when "01000010010111100", -- t[33980] = 3
      "0000011" when "01000010010111101", -- t[33981] = 3
      "0000011" when "01000010010111110", -- t[33982] = 3
      "0000011" when "01000010010111111", -- t[33983] = 3
      "0000011" when "01000010011000000", -- t[33984] = 3
      "0000011" when "01000010011000001", -- t[33985] = 3
      "0000011" when "01000010011000010", -- t[33986] = 3
      "0000011" when "01000010011000011", -- t[33987] = 3
      "0000011" when "01000010011000100", -- t[33988] = 3
      "0000011" when "01000010011000101", -- t[33989] = 3
      "0000011" when "01000010011000110", -- t[33990] = 3
      "0000011" when "01000010011000111", -- t[33991] = 3
      "0000011" when "01000010011001000", -- t[33992] = 3
      "0000011" when "01000010011001001", -- t[33993] = 3
      "0000011" when "01000010011001010", -- t[33994] = 3
      "0000011" when "01000010011001011", -- t[33995] = 3
      "0000011" when "01000010011001100", -- t[33996] = 3
      "0000011" when "01000010011001101", -- t[33997] = 3
      "0000011" when "01000010011001110", -- t[33998] = 3
      "0000011" when "01000010011001111", -- t[33999] = 3
      "0000011" when "01000010011010000", -- t[34000] = 3
      "0000011" when "01000010011010001", -- t[34001] = 3
      "0000011" when "01000010011010010", -- t[34002] = 3
      "0000011" when "01000010011010011", -- t[34003] = 3
      "0000011" when "01000010011010100", -- t[34004] = 3
      "0000011" when "01000010011010101", -- t[34005] = 3
      "0000011" when "01000010011010110", -- t[34006] = 3
      "0000011" when "01000010011010111", -- t[34007] = 3
      "0000011" when "01000010011011000", -- t[34008] = 3
      "0000011" when "01000010011011001", -- t[34009] = 3
      "0000011" when "01000010011011010", -- t[34010] = 3
      "0000011" when "01000010011011011", -- t[34011] = 3
      "0000011" when "01000010011011100", -- t[34012] = 3
      "0000011" when "01000010011011101", -- t[34013] = 3
      "0000011" when "01000010011011110", -- t[34014] = 3
      "0000011" when "01000010011011111", -- t[34015] = 3
      "0000011" when "01000010011100000", -- t[34016] = 3
      "0000011" when "01000010011100001", -- t[34017] = 3
      "0000011" when "01000010011100010", -- t[34018] = 3
      "0000011" when "01000010011100011", -- t[34019] = 3
      "0000011" when "01000010011100100", -- t[34020] = 3
      "0000011" when "01000010011100101", -- t[34021] = 3
      "0000011" when "01000010011100110", -- t[34022] = 3
      "0000011" when "01000010011100111", -- t[34023] = 3
      "0000011" when "01000010011101000", -- t[34024] = 3
      "0000011" when "01000010011101001", -- t[34025] = 3
      "0000011" when "01000010011101010", -- t[34026] = 3
      "0000011" when "01000010011101011", -- t[34027] = 3
      "0000011" when "01000010011101100", -- t[34028] = 3
      "0000011" when "01000010011101101", -- t[34029] = 3
      "0000011" when "01000010011101110", -- t[34030] = 3
      "0000011" when "01000010011101111", -- t[34031] = 3
      "0000011" when "01000010011110000", -- t[34032] = 3
      "0000011" when "01000010011110001", -- t[34033] = 3
      "0000011" when "01000010011110010", -- t[34034] = 3
      "0000011" when "01000010011110011", -- t[34035] = 3
      "0000011" when "01000010011110100", -- t[34036] = 3
      "0000011" when "01000010011110101", -- t[34037] = 3
      "0000011" when "01000010011110110", -- t[34038] = 3
      "0000011" when "01000010011110111", -- t[34039] = 3
      "0000011" when "01000010011111000", -- t[34040] = 3
      "0000011" when "01000010011111001", -- t[34041] = 3
      "0000011" when "01000010011111010", -- t[34042] = 3
      "0000011" when "01000010011111011", -- t[34043] = 3
      "0000011" when "01000010011111100", -- t[34044] = 3
      "0000011" when "01000010011111101", -- t[34045] = 3
      "0000011" when "01000010011111110", -- t[34046] = 3
      "0000011" when "01000010011111111", -- t[34047] = 3
      "0000011" when "01000010100000000", -- t[34048] = 3
      "0000011" when "01000010100000001", -- t[34049] = 3
      "0000011" when "01000010100000010", -- t[34050] = 3
      "0000011" when "01000010100000011", -- t[34051] = 3
      "0000011" when "01000010100000100", -- t[34052] = 3
      "0000011" when "01000010100000101", -- t[34053] = 3
      "0000011" when "01000010100000110", -- t[34054] = 3
      "0000011" when "01000010100000111", -- t[34055] = 3
      "0000011" when "01000010100001000", -- t[34056] = 3
      "0000011" when "01000010100001001", -- t[34057] = 3
      "0000011" when "01000010100001010", -- t[34058] = 3
      "0000011" when "01000010100001011", -- t[34059] = 3
      "0000011" when "01000010100001100", -- t[34060] = 3
      "0000011" when "01000010100001101", -- t[34061] = 3
      "0000011" when "01000010100001110", -- t[34062] = 3
      "0000011" when "01000010100001111", -- t[34063] = 3
      "0000011" when "01000010100010000", -- t[34064] = 3
      "0000011" when "01000010100010001", -- t[34065] = 3
      "0000011" when "01000010100010010", -- t[34066] = 3
      "0000011" when "01000010100010011", -- t[34067] = 3
      "0000011" when "01000010100010100", -- t[34068] = 3
      "0000011" when "01000010100010101", -- t[34069] = 3
      "0000011" when "01000010100010110", -- t[34070] = 3
      "0000011" when "01000010100010111", -- t[34071] = 3
      "0000011" when "01000010100011000", -- t[34072] = 3
      "0000011" when "01000010100011001", -- t[34073] = 3
      "0000011" when "01000010100011010", -- t[34074] = 3
      "0000011" when "01000010100011011", -- t[34075] = 3
      "0000011" when "01000010100011100", -- t[34076] = 3
      "0000011" when "01000010100011101", -- t[34077] = 3
      "0000011" when "01000010100011110", -- t[34078] = 3
      "0000011" when "01000010100011111", -- t[34079] = 3
      "0000011" when "01000010100100000", -- t[34080] = 3
      "0000011" when "01000010100100001", -- t[34081] = 3
      "0000011" when "01000010100100010", -- t[34082] = 3
      "0000011" when "01000010100100011", -- t[34083] = 3
      "0000011" when "01000010100100100", -- t[34084] = 3
      "0000011" when "01000010100100101", -- t[34085] = 3
      "0000011" when "01000010100100110", -- t[34086] = 3
      "0000011" when "01000010100100111", -- t[34087] = 3
      "0000011" when "01000010100101000", -- t[34088] = 3
      "0000011" when "01000010100101001", -- t[34089] = 3
      "0000011" when "01000010100101010", -- t[34090] = 3
      "0000011" when "01000010100101011", -- t[34091] = 3
      "0000011" when "01000010100101100", -- t[34092] = 3
      "0000011" when "01000010100101101", -- t[34093] = 3
      "0000011" when "01000010100101110", -- t[34094] = 3
      "0000011" when "01000010100101111", -- t[34095] = 3
      "0000011" when "01000010100110000", -- t[34096] = 3
      "0000011" when "01000010100110001", -- t[34097] = 3
      "0000011" when "01000010100110010", -- t[34098] = 3
      "0000011" when "01000010100110011", -- t[34099] = 3
      "0000011" when "01000010100110100", -- t[34100] = 3
      "0000011" when "01000010100110101", -- t[34101] = 3
      "0000011" when "01000010100110110", -- t[34102] = 3
      "0000011" when "01000010100110111", -- t[34103] = 3
      "0000011" when "01000010100111000", -- t[34104] = 3
      "0000011" when "01000010100111001", -- t[34105] = 3
      "0000011" when "01000010100111010", -- t[34106] = 3
      "0000011" when "01000010100111011", -- t[34107] = 3
      "0000011" when "01000010100111100", -- t[34108] = 3
      "0000011" when "01000010100111101", -- t[34109] = 3
      "0000011" when "01000010100111110", -- t[34110] = 3
      "0000011" when "01000010100111111", -- t[34111] = 3
      "0000011" when "01000010101000000", -- t[34112] = 3
      "0000011" when "01000010101000001", -- t[34113] = 3
      "0000011" when "01000010101000010", -- t[34114] = 3
      "0000011" when "01000010101000011", -- t[34115] = 3
      "0000011" when "01000010101000100", -- t[34116] = 3
      "0000011" when "01000010101000101", -- t[34117] = 3
      "0000011" when "01000010101000110", -- t[34118] = 3
      "0000011" when "01000010101000111", -- t[34119] = 3
      "0000011" when "01000010101001000", -- t[34120] = 3
      "0000011" when "01000010101001001", -- t[34121] = 3
      "0000011" when "01000010101001010", -- t[34122] = 3
      "0000011" when "01000010101001011", -- t[34123] = 3
      "0000011" when "01000010101001100", -- t[34124] = 3
      "0000011" when "01000010101001101", -- t[34125] = 3
      "0000011" when "01000010101001110", -- t[34126] = 3
      "0000011" when "01000010101001111", -- t[34127] = 3
      "0000011" when "01000010101010000", -- t[34128] = 3
      "0000011" when "01000010101010001", -- t[34129] = 3
      "0000011" when "01000010101010010", -- t[34130] = 3
      "0000011" when "01000010101010011", -- t[34131] = 3
      "0000011" when "01000010101010100", -- t[34132] = 3
      "0000011" when "01000010101010101", -- t[34133] = 3
      "0000011" when "01000010101010110", -- t[34134] = 3
      "0000011" when "01000010101010111", -- t[34135] = 3
      "0000011" when "01000010101011000", -- t[34136] = 3
      "0000011" when "01000010101011001", -- t[34137] = 3
      "0000011" when "01000010101011010", -- t[34138] = 3
      "0000011" when "01000010101011011", -- t[34139] = 3
      "0000011" when "01000010101011100", -- t[34140] = 3
      "0000011" when "01000010101011101", -- t[34141] = 3
      "0000011" when "01000010101011110", -- t[34142] = 3
      "0000011" when "01000010101011111", -- t[34143] = 3
      "0000011" when "01000010101100000", -- t[34144] = 3
      "0000011" when "01000010101100001", -- t[34145] = 3
      "0000011" when "01000010101100010", -- t[34146] = 3
      "0000011" when "01000010101100011", -- t[34147] = 3
      "0000011" when "01000010101100100", -- t[34148] = 3
      "0000011" when "01000010101100101", -- t[34149] = 3
      "0000011" when "01000010101100110", -- t[34150] = 3
      "0000011" when "01000010101100111", -- t[34151] = 3
      "0000011" when "01000010101101000", -- t[34152] = 3
      "0000011" when "01000010101101001", -- t[34153] = 3
      "0000011" when "01000010101101010", -- t[34154] = 3
      "0000011" when "01000010101101011", -- t[34155] = 3
      "0000011" when "01000010101101100", -- t[34156] = 3
      "0000011" when "01000010101101101", -- t[34157] = 3
      "0000011" when "01000010101101110", -- t[34158] = 3
      "0000011" when "01000010101101111", -- t[34159] = 3
      "0000011" when "01000010101110000", -- t[34160] = 3
      "0000011" when "01000010101110001", -- t[34161] = 3
      "0000011" when "01000010101110010", -- t[34162] = 3
      "0000011" when "01000010101110011", -- t[34163] = 3
      "0000011" when "01000010101110100", -- t[34164] = 3
      "0000011" when "01000010101110101", -- t[34165] = 3
      "0000011" when "01000010101110110", -- t[34166] = 3
      "0000011" when "01000010101110111", -- t[34167] = 3
      "0000011" when "01000010101111000", -- t[34168] = 3
      "0000011" when "01000010101111001", -- t[34169] = 3
      "0000011" when "01000010101111010", -- t[34170] = 3
      "0000011" when "01000010101111011", -- t[34171] = 3
      "0000011" when "01000010101111100", -- t[34172] = 3
      "0000011" when "01000010101111101", -- t[34173] = 3
      "0000011" when "01000010101111110", -- t[34174] = 3
      "0000011" when "01000010101111111", -- t[34175] = 3
      "0000011" when "01000010110000000", -- t[34176] = 3
      "0000011" when "01000010110000001", -- t[34177] = 3
      "0000011" when "01000010110000010", -- t[34178] = 3
      "0000011" when "01000010110000011", -- t[34179] = 3
      "0000011" when "01000010110000100", -- t[34180] = 3
      "0000011" when "01000010110000101", -- t[34181] = 3
      "0000011" when "01000010110000110", -- t[34182] = 3
      "0000011" when "01000010110000111", -- t[34183] = 3
      "0000011" when "01000010110001000", -- t[34184] = 3
      "0000011" when "01000010110001001", -- t[34185] = 3
      "0000011" when "01000010110001010", -- t[34186] = 3
      "0000011" when "01000010110001011", -- t[34187] = 3
      "0000011" when "01000010110001100", -- t[34188] = 3
      "0000011" when "01000010110001101", -- t[34189] = 3
      "0000011" when "01000010110001110", -- t[34190] = 3
      "0000011" when "01000010110001111", -- t[34191] = 3
      "0000011" when "01000010110010000", -- t[34192] = 3
      "0000011" when "01000010110010001", -- t[34193] = 3
      "0000011" when "01000010110010010", -- t[34194] = 3
      "0000011" when "01000010110010011", -- t[34195] = 3
      "0000011" when "01000010110010100", -- t[34196] = 3
      "0000011" when "01000010110010101", -- t[34197] = 3
      "0000011" when "01000010110010110", -- t[34198] = 3
      "0000011" when "01000010110010111", -- t[34199] = 3
      "0000011" when "01000010110011000", -- t[34200] = 3
      "0000011" when "01000010110011001", -- t[34201] = 3
      "0000011" when "01000010110011010", -- t[34202] = 3
      "0000011" when "01000010110011011", -- t[34203] = 3
      "0000011" when "01000010110011100", -- t[34204] = 3
      "0000011" when "01000010110011101", -- t[34205] = 3
      "0000011" when "01000010110011110", -- t[34206] = 3
      "0000011" when "01000010110011111", -- t[34207] = 3
      "0000011" when "01000010110100000", -- t[34208] = 3
      "0000011" when "01000010110100001", -- t[34209] = 3
      "0000011" when "01000010110100010", -- t[34210] = 3
      "0000011" when "01000010110100011", -- t[34211] = 3
      "0000011" when "01000010110100100", -- t[34212] = 3
      "0000011" when "01000010110100101", -- t[34213] = 3
      "0000011" when "01000010110100110", -- t[34214] = 3
      "0000011" when "01000010110100111", -- t[34215] = 3
      "0000011" when "01000010110101000", -- t[34216] = 3
      "0000011" when "01000010110101001", -- t[34217] = 3
      "0000011" when "01000010110101010", -- t[34218] = 3
      "0000011" when "01000010110101011", -- t[34219] = 3
      "0000011" when "01000010110101100", -- t[34220] = 3
      "0000011" when "01000010110101101", -- t[34221] = 3
      "0000011" when "01000010110101110", -- t[34222] = 3
      "0000011" when "01000010110101111", -- t[34223] = 3
      "0000011" when "01000010110110000", -- t[34224] = 3
      "0000011" when "01000010110110001", -- t[34225] = 3
      "0000011" when "01000010110110010", -- t[34226] = 3
      "0000011" when "01000010110110011", -- t[34227] = 3
      "0000011" when "01000010110110100", -- t[34228] = 3
      "0000011" when "01000010110110101", -- t[34229] = 3
      "0000011" when "01000010110110110", -- t[34230] = 3
      "0000011" when "01000010110110111", -- t[34231] = 3
      "0000011" when "01000010110111000", -- t[34232] = 3
      "0000011" when "01000010110111001", -- t[34233] = 3
      "0000011" when "01000010110111010", -- t[34234] = 3
      "0000011" when "01000010110111011", -- t[34235] = 3
      "0000011" when "01000010110111100", -- t[34236] = 3
      "0000011" when "01000010110111101", -- t[34237] = 3
      "0000011" when "01000010110111110", -- t[34238] = 3
      "0000011" when "01000010110111111", -- t[34239] = 3
      "0000011" when "01000010111000000", -- t[34240] = 3
      "0000011" when "01000010111000001", -- t[34241] = 3
      "0000011" when "01000010111000010", -- t[34242] = 3
      "0000011" when "01000010111000011", -- t[34243] = 3
      "0000011" when "01000010111000100", -- t[34244] = 3
      "0000011" when "01000010111000101", -- t[34245] = 3
      "0000011" when "01000010111000110", -- t[34246] = 3
      "0000011" when "01000010111000111", -- t[34247] = 3
      "0000011" when "01000010111001000", -- t[34248] = 3
      "0000011" when "01000010111001001", -- t[34249] = 3
      "0000011" when "01000010111001010", -- t[34250] = 3
      "0000011" when "01000010111001011", -- t[34251] = 3
      "0000011" when "01000010111001100", -- t[34252] = 3
      "0000011" when "01000010111001101", -- t[34253] = 3
      "0000011" when "01000010111001110", -- t[34254] = 3
      "0000011" when "01000010111001111", -- t[34255] = 3
      "0000011" when "01000010111010000", -- t[34256] = 3
      "0000011" when "01000010111010001", -- t[34257] = 3
      "0000011" when "01000010111010010", -- t[34258] = 3
      "0000011" when "01000010111010011", -- t[34259] = 3
      "0000011" when "01000010111010100", -- t[34260] = 3
      "0000011" when "01000010111010101", -- t[34261] = 3
      "0000011" when "01000010111010110", -- t[34262] = 3
      "0000011" when "01000010111010111", -- t[34263] = 3
      "0000011" when "01000010111011000", -- t[34264] = 3
      "0000011" when "01000010111011001", -- t[34265] = 3
      "0000011" when "01000010111011010", -- t[34266] = 3
      "0000011" when "01000010111011011", -- t[34267] = 3
      "0000011" when "01000010111011100", -- t[34268] = 3
      "0000011" when "01000010111011101", -- t[34269] = 3
      "0000011" when "01000010111011110", -- t[34270] = 3
      "0000011" when "01000010111011111", -- t[34271] = 3
      "0000011" when "01000010111100000", -- t[34272] = 3
      "0000011" when "01000010111100001", -- t[34273] = 3
      "0000011" when "01000010111100010", -- t[34274] = 3
      "0000011" when "01000010111100011", -- t[34275] = 3
      "0000011" when "01000010111100100", -- t[34276] = 3
      "0000011" when "01000010111100101", -- t[34277] = 3
      "0000011" when "01000010111100110", -- t[34278] = 3
      "0000011" when "01000010111100111", -- t[34279] = 3
      "0000011" when "01000010111101000", -- t[34280] = 3
      "0000011" when "01000010111101001", -- t[34281] = 3
      "0000011" when "01000010111101010", -- t[34282] = 3
      "0000011" when "01000010111101011", -- t[34283] = 3
      "0000011" when "01000010111101100", -- t[34284] = 3
      "0000011" when "01000010111101101", -- t[34285] = 3
      "0000011" when "01000010111101110", -- t[34286] = 3
      "0000011" when "01000010111101111", -- t[34287] = 3
      "0000011" when "01000010111110000", -- t[34288] = 3
      "0000011" when "01000010111110001", -- t[34289] = 3
      "0000011" when "01000010111110010", -- t[34290] = 3
      "0000011" when "01000010111110011", -- t[34291] = 3
      "0000011" when "01000010111110100", -- t[34292] = 3
      "0000011" when "01000010111110101", -- t[34293] = 3
      "0000011" when "01000010111110110", -- t[34294] = 3
      "0000011" when "01000010111110111", -- t[34295] = 3
      "0000011" when "01000010111111000", -- t[34296] = 3
      "0000011" when "01000010111111001", -- t[34297] = 3
      "0000011" when "01000010111111010", -- t[34298] = 3
      "0000011" when "01000010111111011", -- t[34299] = 3
      "0000011" when "01000010111111100", -- t[34300] = 3
      "0000011" when "01000010111111101", -- t[34301] = 3
      "0000011" when "01000010111111110", -- t[34302] = 3
      "0000011" when "01000010111111111", -- t[34303] = 3
      "0000011" when "01000011000000000", -- t[34304] = 3
      "0000011" when "01000011000000001", -- t[34305] = 3
      "0000011" when "01000011000000010", -- t[34306] = 3
      "0000011" when "01000011000000011", -- t[34307] = 3
      "0000011" when "01000011000000100", -- t[34308] = 3
      "0000011" when "01000011000000101", -- t[34309] = 3
      "0000011" when "01000011000000110", -- t[34310] = 3
      "0000011" when "01000011000000111", -- t[34311] = 3
      "0000011" when "01000011000001000", -- t[34312] = 3
      "0000011" when "01000011000001001", -- t[34313] = 3
      "0000011" when "01000011000001010", -- t[34314] = 3
      "0000011" when "01000011000001011", -- t[34315] = 3
      "0000011" when "01000011000001100", -- t[34316] = 3
      "0000011" when "01000011000001101", -- t[34317] = 3
      "0000011" when "01000011000001110", -- t[34318] = 3
      "0000011" when "01000011000001111", -- t[34319] = 3
      "0000011" when "01000011000010000", -- t[34320] = 3
      "0000011" when "01000011000010001", -- t[34321] = 3
      "0000011" when "01000011000010010", -- t[34322] = 3
      "0000011" when "01000011000010011", -- t[34323] = 3
      "0000011" when "01000011000010100", -- t[34324] = 3
      "0000011" when "01000011000010101", -- t[34325] = 3
      "0000011" when "01000011000010110", -- t[34326] = 3
      "0000011" when "01000011000010111", -- t[34327] = 3
      "0000011" when "01000011000011000", -- t[34328] = 3
      "0000011" when "01000011000011001", -- t[34329] = 3
      "0000011" when "01000011000011010", -- t[34330] = 3
      "0000011" when "01000011000011011", -- t[34331] = 3
      "0000011" when "01000011000011100", -- t[34332] = 3
      "0000011" when "01000011000011101", -- t[34333] = 3
      "0000011" when "01000011000011110", -- t[34334] = 3
      "0000011" when "01000011000011111", -- t[34335] = 3
      "0000011" when "01000011000100000", -- t[34336] = 3
      "0000011" when "01000011000100001", -- t[34337] = 3
      "0000011" when "01000011000100010", -- t[34338] = 3
      "0000011" when "01000011000100011", -- t[34339] = 3
      "0000011" when "01000011000100100", -- t[34340] = 3
      "0000011" when "01000011000100101", -- t[34341] = 3
      "0000011" when "01000011000100110", -- t[34342] = 3
      "0000011" when "01000011000100111", -- t[34343] = 3
      "0000011" when "01000011000101000", -- t[34344] = 3
      "0000011" when "01000011000101001", -- t[34345] = 3
      "0000011" when "01000011000101010", -- t[34346] = 3
      "0000011" when "01000011000101011", -- t[34347] = 3
      "0000011" when "01000011000101100", -- t[34348] = 3
      "0000011" when "01000011000101101", -- t[34349] = 3
      "0000011" when "01000011000101110", -- t[34350] = 3
      "0000011" when "01000011000101111", -- t[34351] = 3
      "0000011" when "01000011000110000", -- t[34352] = 3
      "0000011" when "01000011000110001", -- t[34353] = 3
      "0000011" when "01000011000110010", -- t[34354] = 3
      "0000011" when "01000011000110011", -- t[34355] = 3
      "0000011" when "01000011000110100", -- t[34356] = 3
      "0000011" when "01000011000110101", -- t[34357] = 3
      "0000011" when "01000011000110110", -- t[34358] = 3
      "0000011" when "01000011000110111", -- t[34359] = 3
      "0000011" when "01000011000111000", -- t[34360] = 3
      "0000011" when "01000011000111001", -- t[34361] = 3
      "0000011" when "01000011000111010", -- t[34362] = 3
      "0000011" when "01000011000111011", -- t[34363] = 3
      "0000011" when "01000011000111100", -- t[34364] = 3
      "0000011" when "01000011000111101", -- t[34365] = 3
      "0000011" when "01000011000111110", -- t[34366] = 3
      "0000011" when "01000011000111111", -- t[34367] = 3
      "0000011" when "01000011001000000", -- t[34368] = 3
      "0000011" when "01000011001000001", -- t[34369] = 3
      "0000011" when "01000011001000010", -- t[34370] = 3
      "0000011" when "01000011001000011", -- t[34371] = 3
      "0000011" when "01000011001000100", -- t[34372] = 3
      "0000011" when "01000011001000101", -- t[34373] = 3
      "0000011" when "01000011001000110", -- t[34374] = 3
      "0000011" when "01000011001000111", -- t[34375] = 3
      "0000011" when "01000011001001000", -- t[34376] = 3
      "0000011" when "01000011001001001", -- t[34377] = 3
      "0000011" when "01000011001001010", -- t[34378] = 3
      "0000011" when "01000011001001011", -- t[34379] = 3
      "0000011" when "01000011001001100", -- t[34380] = 3
      "0000011" when "01000011001001101", -- t[34381] = 3
      "0000011" when "01000011001001110", -- t[34382] = 3
      "0000011" when "01000011001001111", -- t[34383] = 3
      "0000011" when "01000011001010000", -- t[34384] = 3
      "0000011" when "01000011001010001", -- t[34385] = 3
      "0000011" when "01000011001010010", -- t[34386] = 3
      "0000011" when "01000011001010011", -- t[34387] = 3
      "0000011" when "01000011001010100", -- t[34388] = 3
      "0000011" when "01000011001010101", -- t[34389] = 3
      "0000011" when "01000011001010110", -- t[34390] = 3
      "0000011" when "01000011001010111", -- t[34391] = 3
      "0000011" when "01000011001011000", -- t[34392] = 3
      "0000011" when "01000011001011001", -- t[34393] = 3
      "0000011" when "01000011001011010", -- t[34394] = 3
      "0000011" when "01000011001011011", -- t[34395] = 3
      "0000011" when "01000011001011100", -- t[34396] = 3
      "0000011" when "01000011001011101", -- t[34397] = 3
      "0000011" when "01000011001011110", -- t[34398] = 3
      "0000011" when "01000011001011111", -- t[34399] = 3
      "0000011" when "01000011001100000", -- t[34400] = 3
      "0000011" when "01000011001100001", -- t[34401] = 3
      "0000011" when "01000011001100010", -- t[34402] = 3
      "0000011" when "01000011001100011", -- t[34403] = 3
      "0000011" when "01000011001100100", -- t[34404] = 3
      "0000011" when "01000011001100101", -- t[34405] = 3
      "0000011" when "01000011001100110", -- t[34406] = 3
      "0000011" when "01000011001100111", -- t[34407] = 3
      "0000011" when "01000011001101000", -- t[34408] = 3
      "0000011" when "01000011001101001", -- t[34409] = 3
      "0000011" when "01000011001101010", -- t[34410] = 3
      "0000011" when "01000011001101011", -- t[34411] = 3
      "0000011" when "01000011001101100", -- t[34412] = 3
      "0000011" when "01000011001101101", -- t[34413] = 3
      "0000011" when "01000011001101110", -- t[34414] = 3
      "0000011" when "01000011001101111", -- t[34415] = 3
      "0000011" when "01000011001110000", -- t[34416] = 3
      "0000011" when "01000011001110001", -- t[34417] = 3
      "0000011" when "01000011001110010", -- t[34418] = 3
      "0000011" when "01000011001110011", -- t[34419] = 3
      "0000011" when "01000011001110100", -- t[34420] = 3
      "0000011" when "01000011001110101", -- t[34421] = 3
      "0000011" when "01000011001110110", -- t[34422] = 3
      "0000011" when "01000011001110111", -- t[34423] = 3
      "0000011" when "01000011001111000", -- t[34424] = 3
      "0000011" when "01000011001111001", -- t[34425] = 3
      "0000011" when "01000011001111010", -- t[34426] = 3
      "0000011" when "01000011001111011", -- t[34427] = 3
      "0000011" when "01000011001111100", -- t[34428] = 3
      "0000011" when "01000011001111101", -- t[34429] = 3
      "0000011" when "01000011001111110", -- t[34430] = 3
      "0000011" when "01000011001111111", -- t[34431] = 3
      "0000011" when "01000011010000000", -- t[34432] = 3
      "0000011" when "01000011010000001", -- t[34433] = 3
      "0000011" when "01000011010000010", -- t[34434] = 3
      "0000011" when "01000011010000011", -- t[34435] = 3
      "0000011" when "01000011010000100", -- t[34436] = 3
      "0000011" when "01000011010000101", -- t[34437] = 3
      "0000011" when "01000011010000110", -- t[34438] = 3
      "0000011" when "01000011010000111", -- t[34439] = 3
      "0000011" when "01000011010001000", -- t[34440] = 3
      "0000011" when "01000011010001001", -- t[34441] = 3
      "0000011" when "01000011010001010", -- t[34442] = 3
      "0000011" when "01000011010001011", -- t[34443] = 3
      "0000011" when "01000011010001100", -- t[34444] = 3
      "0000011" when "01000011010001101", -- t[34445] = 3
      "0000011" when "01000011010001110", -- t[34446] = 3
      "0000011" when "01000011010001111", -- t[34447] = 3
      "0000011" when "01000011010010000", -- t[34448] = 3
      "0000011" when "01000011010010001", -- t[34449] = 3
      "0000011" when "01000011010010010", -- t[34450] = 3
      "0000011" when "01000011010010011", -- t[34451] = 3
      "0000011" when "01000011010010100", -- t[34452] = 3
      "0000011" when "01000011010010101", -- t[34453] = 3
      "0000011" when "01000011010010110", -- t[34454] = 3
      "0000011" when "01000011010010111", -- t[34455] = 3
      "0000011" when "01000011010011000", -- t[34456] = 3
      "0000011" when "01000011010011001", -- t[34457] = 3
      "0000011" when "01000011010011010", -- t[34458] = 3
      "0000011" when "01000011010011011", -- t[34459] = 3
      "0000011" when "01000011010011100", -- t[34460] = 3
      "0000011" when "01000011010011101", -- t[34461] = 3
      "0000011" when "01000011010011110", -- t[34462] = 3
      "0000011" when "01000011010011111", -- t[34463] = 3
      "0000011" when "01000011010100000", -- t[34464] = 3
      "0000011" when "01000011010100001", -- t[34465] = 3
      "0000011" when "01000011010100010", -- t[34466] = 3
      "0000011" when "01000011010100011", -- t[34467] = 3
      "0000011" when "01000011010100100", -- t[34468] = 3
      "0000011" when "01000011010100101", -- t[34469] = 3
      "0000011" when "01000011010100110", -- t[34470] = 3
      "0000011" when "01000011010100111", -- t[34471] = 3
      "0000011" when "01000011010101000", -- t[34472] = 3
      "0000011" when "01000011010101001", -- t[34473] = 3
      "0000011" when "01000011010101010", -- t[34474] = 3
      "0000011" when "01000011010101011", -- t[34475] = 3
      "0000011" when "01000011010101100", -- t[34476] = 3
      "0000011" when "01000011010101101", -- t[34477] = 3
      "0000011" when "01000011010101110", -- t[34478] = 3
      "0000011" when "01000011010101111", -- t[34479] = 3
      "0000011" when "01000011010110000", -- t[34480] = 3
      "0000011" when "01000011010110001", -- t[34481] = 3
      "0000011" when "01000011010110010", -- t[34482] = 3
      "0000011" when "01000011010110011", -- t[34483] = 3
      "0000011" when "01000011010110100", -- t[34484] = 3
      "0000011" when "01000011010110101", -- t[34485] = 3
      "0000011" when "01000011010110110", -- t[34486] = 3
      "0000011" when "01000011010110111", -- t[34487] = 3
      "0000011" when "01000011010111000", -- t[34488] = 3
      "0000011" when "01000011010111001", -- t[34489] = 3
      "0000011" when "01000011010111010", -- t[34490] = 3
      "0000011" when "01000011010111011", -- t[34491] = 3
      "0000011" when "01000011010111100", -- t[34492] = 3
      "0000011" when "01000011010111101", -- t[34493] = 3
      "0000011" when "01000011010111110", -- t[34494] = 3
      "0000011" when "01000011010111111", -- t[34495] = 3
      "0000011" when "01000011011000000", -- t[34496] = 3
      "0000011" when "01000011011000001", -- t[34497] = 3
      "0000011" when "01000011011000010", -- t[34498] = 3
      "0000011" when "01000011011000011", -- t[34499] = 3
      "0000011" when "01000011011000100", -- t[34500] = 3
      "0000011" when "01000011011000101", -- t[34501] = 3
      "0000011" when "01000011011000110", -- t[34502] = 3
      "0000011" when "01000011011000111", -- t[34503] = 3
      "0000011" when "01000011011001000", -- t[34504] = 3
      "0000011" when "01000011011001001", -- t[34505] = 3
      "0000011" when "01000011011001010", -- t[34506] = 3
      "0000011" when "01000011011001011", -- t[34507] = 3
      "0000011" when "01000011011001100", -- t[34508] = 3
      "0000011" when "01000011011001101", -- t[34509] = 3
      "0000011" when "01000011011001110", -- t[34510] = 3
      "0000011" when "01000011011001111", -- t[34511] = 3
      "0000011" when "01000011011010000", -- t[34512] = 3
      "0000011" when "01000011011010001", -- t[34513] = 3
      "0000011" when "01000011011010010", -- t[34514] = 3
      "0000011" when "01000011011010011", -- t[34515] = 3
      "0000011" when "01000011011010100", -- t[34516] = 3
      "0000011" when "01000011011010101", -- t[34517] = 3
      "0000011" when "01000011011010110", -- t[34518] = 3
      "0000011" when "01000011011010111", -- t[34519] = 3
      "0000011" when "01000011011011000", -- t[34520] = 3
      "0000011" when "01000011011011001", -- t[34521] = 3
      "0000011" when "01000011011011010", -- t[34522] = 3
      "0000011" when "01000011011011011", -- t[34523] = 3
      "0000011" when "01000011011011100", -- t[34524] = 3
      "0000011" when "01000011011011101", -- t[34525] = 3
      "0000011" when "01000011011011110", -- t[34526] = 3
      "0000011" when "01000011011011111", -- t[34527] = 3
      "0000011" when "01000011011100000", -- t[34528] = 3
      "0000011" when "01000011011100001", -- t[34529] = 3
      "0000011" when "01000011011100010", -- t[34530] = 3
      "0000011" when "01000011011100011", -- t[34531] = 3
      "0000011" when "01000011011100100", -- t[34532] = 3
      "0000011" when "01000011011100101", -- t[34533] = 3
      "0000011" when "01000011011100110", -- t[34534] = 3
      "0000011" when "01000011011100111", -- t[34535] = 3
      "0000011" when "01000011011101000", -- t[34536] = 3
      "0000011" when "01000011011101001", -- t[34537] = 3
      "0000011" when "01000011011101010", -- t[34538] = 3
      "0000011" when "01000011011101011", -- t[34539] = 3
      "0000011" when "01000011011101100", -- t[34540] = 3
      "0000011" when "01000011011101101", -- t[34541] = 3
      "0000011" when "01000011011101110", -- t[34542] = 3
      "0000011" when "01000011011101111", -- t[34543] = 3
      "0000011" when "01000011011110000", -- t[34544] = 3
      "0000011" when "01000011011110001", -- t[34545] = 3
      "0000011" when "01000011011110010", -- t[34546] = 3
      "0000011" when "01000011011110011", -- t[34547] = 3
      "0000011" when "01000011011110100", -- t[34548] = 3
      "0000011" when "01000011011110101", -- t[34549] = 3
      "0000011" when "01000011011110110", -- t[34550] = 3
      "0000011" when "01000011011110111", -- t[34551] = 3
      "0000011" when "01000011011111000", -- t[34552] = 3
      "0000011" when "01000011011111001", -- t[34553] = 3
      "0000011" when "01000011011111010", -- t[34554] = 3
      "0000011" when "01000011011111011", -- t[34555] = 3
      "0000011" when "01000011011111100", -- t[34556] = 3
      "0000011" when "01000011011111101", -- t[34557] = 3
      "0000011" when "01000011011111110", -- t[34558] = 3
      "0000011" when "01000011011111111", -- t[34559] = 3
      "0000011" when "01000011100000000", -- t[34560] = 3
      "0000011" when "01000011100000001", -- t[34561] = 3
      "0000011" when "01000011100000010", -- t[34562] = 3
      "0000011" when "01000011100000011", -- t[34563] = 3
      "0000011" when "01000011100000100", -- t[34564] = 3
      "0000011" when "01000011100000101", -- t[34565] = 3
      "0000011" when "01000011100000110", -- t[34566] = 3
      "0000011" when "01000011100000111", -- t[34567] = 3
      "0000011" when "01000011100001000", -- t[34568] = 3
      "0000011" when "01000011100001001", -- t[34569] = 3
      "0000011" when "01000011100001010", -- t[34570] = 3
      "0000011" when "01000011100001011", -- t[34571] = 3
      "0000011" when "01000011100001100", -- t[34572] = 3
      "0000011" when "01000011100001101", -- t[34573] = 3
      "0000011" when "01000011100001110", -- t[34574] = 3
      "0000011" when "01000011100001111", -- t[34575] = 3
      "0000011" when "01000011100010000", -- t[34576] = 3
      "0000011" when "01000011100010001", -- t[34577] = 3
      "0000011" when "01000011100010010", -- t[34578] = 3
      "0000011" when "01000011100010011", -- t[34579] = 3
      "0000011" when "01000011100010100", -- t[34580] = 3
      "0000011" when "01000011100010101", -- t[34581] = 3
      "0000011" when "01000011100010110", -- t[34582] = 3
      "0000011" when "01000011100010111", -- t[34583] = 3
      "0000011" when "01000011100011000", -- t[34584] = 3
      "0000011" when "01000011100011001", -- t[34585] = 3
      "0000011" when "01000011100011010", -- t[34586] = 3
      "0000011" when "01000011100011011", -- t[34587] = 3
      "0000011" when "01000011100011100", -- t[34588] = 3
      "0000011" when "01000011100011101", -- t[34589] = 3
      "0000011" when "01000011100011110", -- t[34590] = 3
      "0000011" when "01000011100011111", -- t[34591] = 3
      "0000011" when "01000011100100000", -- t[34592] = 3
      "0000011" when "01000011100100001", -- t[34593] = 3
      "0000011" when "01000011100100010", -- t[34594] = 3
      "0000011" when "01000011100100011", -- t[34595] = 3
      "0000011" when "01000011100100100", -- t[34596] = 3
      "0000011" when "01000011100100101", -- t[34597] = 3
      "0000011" when "01000011100100110", -- t[34598] = 3
      "0000011" when "01000011100100111", -- t[34599] = 3
      "0000011" when "01000011100101000", -- t[34600] = 3
      "0000011" when "01000011100101001", -- t[34601] = 3
      "0000011" when "01000011100101010", -- t[34602] = 3
      "0000011" when "01000011100101011", -- t[34603] = 3
      "0000011" when "01000011100101100", -- t[34604] = 3
      "0000011" when "01000011100101101", -- t[34605] = 3
      "0000011" when "01000011100101110", -- t[34606] = 3
      "0000011" when "01000011100101111", -- t[34607] = 3
      "0000011" when "01000011100110000", -- t[34608] = 3
      "0000011" when "01000011100110001", -- t[34609] = 3
      "0000011" when "01000011100110010", -- t[34610] = 3
      "0000011" when "01000011100110011", -- t[34611] = 3
      "0000011" when "01000011100110100", -- t[34612] = 3
      "0000011" when "01000011100110101", -- t[34613] = 3
      "0000011" when "01000011100110110", -- t[34614] = 3
      "0000011" when "01000011100110111", -- t[34615] = 3
      "0000011" when "01000011100111000", -- t[34616] = 3
      "0000011" when "01000011100111001", -- t[34617] = 3
      "0000011" when "01000011100111010", -- t[34618] = 3
      "0000011" when "01000011100111011", -- t[34619] = 3
      "0000011" when "01000011100111100", -- t[34620] = 3
      "0000011" when "01000011100111101", -- t[34621] = 3
      "0000011" when "01000011100111110", -- t[34622] = 3
      "0000011" when "01000011100111111", -- t[34623] = 3
      "0000011" when "01000011101000000", -- t[34624] = 3
      "0000011" when "01000011101000001", -- t[34625] = 3
      "0000011" when "01000011101000010", -- t[34626] = 3
      "0000011" when "01000011101000011", -- t[34627] = 3
      "0000011" when "01000011101000100", -- t[34628] = 3
      "0000011" when "01000011101000101", -- t[34629] = 3
      "0000011" when "01000011101000110", -- t[34630] = 3
      "0000011" when "01000011101000111", -- t[34631] = 3
      "0000011" when "01000011101001000", -- t[34632] = 3
      "0000011" when "01000011101001001", -- t[34633] = 3
      "0000011" when "01000011101001010", -- t[34634] = 3
      "0000011" when "01000011101001011", -- t[34635] = 3
      "0000011" when "01000011101001100", -- t[34636] = 3
      "0000011" when "01000011101001101", -- t[34637] = 3
      "0000011" when "01000011101001110", -- t[34638] = 3
      "0000011" when "01000011101001111", -- t[34639] = 3
      "0000011" when "01000011101010000", -- t[34640] = 3
      "0000011" when "01000011101010001", -- t[34641] = 3
      "0000011" when "01000011101010010", -- t[34642] = 3
      "0000011" when "01000011101010011", -- t[34643] = 3
      "0000011" when "01000011101010100", -- t[34644] = 3
      "0000011" when "01000011101010101", -- t[34645] = 3
      "0000011" when "01000011101010110", -- t[34646] = 3
      "0000011" when "01000011101010111", -- t[34647] = 3
      "0000011" when "01000011101011000", -- t[34648] = 3
      "0000011" when "01000011101011001", -- t[34649] = 3
      "0000011" when "01000011101011010", -- t[34650] = 3
      "0000011" when "01000011101011011", -- t[34651] = 3
      "0000011" when "01000011101011100", -- t[34652] = 3
      "0000011" when "01000011101011101", -- t[34653] = 3
      "0000011" when "01000011101011110", -- t[34654] = 3
      "0000011" when "01000011101011111", -- t[34655] = 3
      "0000011" when "01000011101100000", -- t[34656] = 3
      "0000011" when "01000011101100001", -- t[34657] = 3
      "0000011" when "01000011101100010", -- t[34658] = 3
      "0000011" when "01000011101100011", -- t[34659] = 3
      "0000011" when "01000011101100100", -- t[34660] = 3
      "0000011" when "01000011101100101", -- t[34661] = 3
      "0000011" when "01000011101100110", -- t[34662] = 3
      "0000011" when "01000011101100111", -- t[34663] = 3
      "0000011" when "01000011101101000", -- t[34664] = 3
      "0000011" when "01000011101101001", -- t[34665] = 3
      "0000011" when "01000011101101010", -- t[34666] = 3
      "0000011" when "01000011101101011", -- t[34667] = 3
      "0000011" when "01000011101101100", -- t[34668] = 3
      "0000011" when "01000011101101101", -- t[34669] = 3
      "0000011" when "01000011101101110", -- t[34670] = 3
      "0000011" when "01000011101101111", -- t[34671] = 3
      "0000011" when "01000011101110000", -- t[34672] = 3
      "0000011" when "01000011101110001", -- t[34673] = 3
      "0000011" when "01000011101110010", -- t[34674] = 3
      "0000011" when "01000011101110011", -- t[34675] = 3
      "0000011" when "01000011101110100", -- t[34676] = 3
      "0000011" when "01000011101110101", -- t[34677] = 3
      "0000011" when "01000011101110110", -- t[34678] = 3
      "0000011" when "01000011101110111", -- t[34679] = 3
      "0000011" when "01000011101111000", -- t[34680] = 3
      "0000011" when "01000011101111001", -- t[34681] = 3
      "0000011" when "01000011101111010", -- t[34682] = 3
      "0000011" when "01000011101111011", -- t[34683] = 3
      "0000011" when "01000011101111100", -- t[34684] = 3
      "0000011" when "01000011101111101", -- t[34685] = 3
      "0000011" when "01000011101111110", -- t[34686] = 3
      "0000011" when "01000011101111111", -- t[34687] = 3
      "0000011" when "01000011110000000", -- t[34688] = 3
      "0000011" when "01000011110000001", -- t[34689] = 3
      "0000011" when "01000011110000010", -- t[34690] = 3
      "0000011" when "01000011110000011", -- t[34691] = 3
      "0000011" when "01000011110000100", -- t[34692] = 3
      "0000011" when "01000011110000101", -- t[34693] = 3
      "0000011" when "01000011110000110", -- t[34694] = 3
      "0000011" when "01000011110000111", -- t[34695] = 3
      "0000011" when "01000011110001000", -- t[34696] = 3
      "0000011" when "01000011110001001", -- t[34697] = 3
      "0000011" when "01000011110001010", -- t[34698] = 3
      "0000011" when "01000011110001011", -- t[34699] = 3
      "0000011" when "01000011110001100", -- t[34700] = 3
      "0000011" when "01000011110001101", -- t[34701] = 3
      "0000011" when "01000011110001110", -- t[34702] = 3
      "0000011" when "01000011110001111", -- t[34703] = 3
      "0000011" when "01000011110010000", -- t[34704] = 3
      "0000011" when "01000011110010001", -- t[34705] = 3
      "0000011" when "01000011110010010", -- t[34706] = 3
      "0000011" when "01000011110010011", -- t[34707] = 3
      "0000011" when "01000011110010100", -- t[34708] = 3
      "0000011" when "01000011110010101", -- t[34709] = 3
      "0000011" when "01000011110010110", -- t[34710] = 3
      "0000011" when "01000011110010111", -- t[34711] = 3
      "0000011" when "01000011110011000", -- t[34712] = 3
      "0000011" when "01000011110011001", -- t[34713] = 3
      "0000011" when "01000011110011010", -- t[34714] = 3
      "0000011" when "01000011110011011", -- t[34715] = 3
      "0000011" when "01000011110011100", -- t[34716] = 3
      "0000011" when "01000011110011101", -- t[34717] = 3
      "0000011" when "01000011110011110", -- t[34718] = 3
      "0000011" when "01000011110011111", -- t[34719] = 3
      "0000011" when "01000011110100000", -- t[34720] = 3
      "0000011" when "01000011110100001", -- t[34721] = 3
      "0000011" when "01000011110100010", -- t[34722] = 3
      "0000011" when "01000011110100011", -- t[34723] = 3
      "0000011" when "01000011110100100", -- t[34724] = 3
      "0000011" when "01000011110100101", -- t[34725] = 3
      "0000011" when "01000011110100110", -- t[34726] = 3
      "0000011" when "01000011110100111", -- t[34727] = 3
      "0000011" when "01000011110101000", -- t[34728] = 3
      "0000011" when "01000011110101001", -- t[34729] = 3
      "0000011" when "01000011110101010", -- t[34730] = 3
      "0000011" when "01000011110101011", -- t[34731] = 3
      "0000011" when "01000011110101100", -- t[34732] = 3
      "0000011" when "01000011110101101", -- t[34733] = 3
      "0000011" when "01000011110101110", -- t[34734] = 3
      "0000011" when "01000011110101111", -- t[34735] = 3
      "0000011" when "01000011110110000", -- t[34736] = 3
      "0000011" when "01000011110110001", -- t[34737] = 3
      "0000011" when "01000011110110010", -- t[34738] = 3
      "0000011" when "01000011110110011", -- t[34739] = 3
      "0000011" when "01000011110110100", -- t[34740] = 3
      "0000011" when "01000011110110101", -- t[34741] = 3
      "0000011" when "01000011110110110", -- t[34742] = 3
      "0000011" when "01000011110110111", -- t[34743] = 3
      "0000011" when "01000011110111000", -- t[34744] = 3
      "0000011" when "01000011110111001", -- t[34745] = 3
      "0000011" when "01000011110111010", -- t[34746] = 3
      "0000011" when "01000011110111011", -- t[34747] = 3
      "0000011" when "01000011110111100", -- t[34748] = 3
      "0000011" when "01000011110111101", -- t[34749] = 3
      "0000011" when "01000011110111110", -- t[34750] = 3
      "0000011" when "01000011110111111", -- t[34751] = 3
      "0000011" when "01000011111000000", -- t[34752] = 3
      "0000011" when "01000011111000001", -- t[34753] = 3
      "0000011" when "01000011111000010", -- t[34754] = 3
      "0000011" when "01000011111000011", -- t[34755] = 3
      "0000011" when "01000011111000100", -- t[34756] = 3
      "0000011" when "01000011111000101", -- t[34757] = 3
      "0000011" when "01000011111000110", -- t[34758] = 3
      "0000011" when "01000011111000111", -- t[34759] = 3
      "0000011" when "01000011111001000", -- t[34760] = 3
      "0000011" when "01000011111001001", -- t[34761] = 3
      "0000011" when "01000011111001010", -- t[34762] = 3
      "0000011" when "01000011111001011", -- t[34763] = 3
      "0000011" when "01000011111001100", -- t[34764] = 3
      "0000011" when "01000011111001101", -- t[34765] = 3
      "0000011" when "01000011111001110", -- t[34766] = 3
      "0000011" when "01000011111001111", -- t[34767] = 3
      "0000011" when "01000011111010000", -- t[34768] = 3
      "0000011" when "01000011111010001", -- t[34769] = 3
      "0000011" when "01000011111010010", -- t[34770] = 3
      "0000011" when "01000011111010011", -- t[34771] = 3
      "0000011" when "01000011111010100", -- t[34772] = 3
      "0000011" when "01000011111010101", -- t[34773] = 3
      "0000011" when "01000011111010110", -- t[34774] = 3
      "0000011" when "01000011111010111", -- t[34775] = 3
      "0000011" when "01000011111011000", -- t[34776] = 3
      "0000011" when "01000011111011001", -- t[34777] = 3
      "0000011" when "01000011111011010", -- t[34778] = 3
      "0000011" when "01000011111011011", -- t[34779] = 3
      "0000011" when "01000011111011100", -- t[34780] = 3
      "0000011" when "01000011111011101", -- t[34781] = 3
      "0000011" when "01000011111011110", -- t[34782] = 3
      "0000011" when "01000011111011111", -- t[34783] = 3
      "0000011" when "01000011111100000", -- t[34784] = 3
      "0000011" when "01000011111100001", -- t[34785] = 3
      "0000011" when "01000011111100010", -- t[34786] = 3
      "0000011" when "01000011111100011", -- t[34787] = 3
      "0000011" when "01000011111100100", -- t[34788] = 3
      "0000011" when "01000011111100101", -- t[34789] = 3
      "0000011" when "01000011111100110", -- t[34790] = 3
      "0000011" when "01000011111100111", -- t[34791] = 3
      "0000011" when "01000011111101000", -- t[34792] = 3
      "0000011" when "01000011111101001", -- t[34793] = 3
      "0000011" when "01000011111101010", -- t[34794] = 3
      "0000011" when "01000011111101011", -- t[34795] = 3
      "0000011" when "01000011111101100", -- t[34796] = 3
      "0000011" when "01000011111101101", -- t[34797] = 3
      "0000011" when "01000011111101110", -- t[34798] = 3
      "0000011" when "01000011111101111", -- t[34799] = 3
      "0000011" when "01000011111110000", -- t[34800] = 3
      "0000011" when "01000011111110001", -- t[34801] = 3
      "0000011" when "01000011111110010", -- t[34802] = 3
      "0000011" when "01000011111110011", -- t[34803] = 3
      "0000011" when "01000011111110100", -- t[34804] = 3
      "0000011" when "01000011111110101", -- t[34805] = 3
      "0000011" when "01000011111110110", -- t[34806] = 3
      "0000011" when "01000011111110111", -- t[34807] = 3
      "0000011" when "01000011111111000", -- t[34808] = 3
      "0000011" when "01000011111111001", -- t[34809] = 3
      "0000011" when "01000011111111010", -- t[34810] = 3
      "0000011" when "01000011111111011", -- t[34811] = 3
      "0000011" when "01000011111111100", -- t[34812] = 3
      "0000011" when "01000011111111101", -- t[34813] = 3
      "0000011" when "01000011111111110", -- t[34814] = 3
      "0000011" when "01000011111111111", -- t[34815] = 3
      "0000011" when "01000100000000000", -- t[34816] = 3
      "0000011" when "01000100000000001", -- t[34817] = 3
      "0000011" when "01000100000000010", -- t[34818] = 3
      "0000011" when "01000100000000011", -- t[34819] = 3
      "0000011" when "01000100000000100", -- t[34820] = 3
      "0000011" when "01000100000000101", -- t[34821] = 3
      "0000011" when "01000100000000110", -- t[34822] = 3
      "0000011" when "01000100000000111", -- t[34823] = 3
      "0000011" when "01000100000001000", -- t[34824] = 3
      "0000011" when "01000100000001001", -- t[34825] = 3
      "0000011" when "01000100000001010", -- t[34826] = 3
      "0000011" when "01000100000001011", -- t[34827] = 3
      "0000011" when "01000100000001100", -- t[34828] = 3
      "0000011" when "01000100000001101", -- t[34829] = 3
      "0000011" when "01000100000001110", -- t[34830] = 3
      "0000011" when "01000100000001111", -- t[34831] = 3
      "0000011" when "01000100000010000", -- t[34832] = 3
      "0000011" when "01000100000010001", -- t[34833] = 3
      "0000011" when "01000100000010010", -- t[34834] = 3
      "0000011" when "01000100000010011", -- t[34835] = 3
      "0000011" when "01000100000010100", -- t[34836] = 3
      "0000011" when "01000100000010101", -- t[34837] = 3
      "0000011" when "01000100000010110", -- t[34838] = 3
      "0000011" when "01000100000010111", -- t[34839] = 3
      "0000011" when "01000100000011000", -- t[34840] = 3
      "0000011" when "01000100000011001", -- t[34841] = 3
      "0000011" when "01000100000011010", -- t[34842] = 3
      "0000011" when "01000100000011011", -- t[34843] = 3
      "0000011" when "01000100000011100", -- t[34844] = 3
      "0000011" when "01000100000011101", -- t[34845] = 3
      "0000011" when "01000100000011110", -- t[34846] = 3
      "0000011" when "01000100000011111", -- t[34847] = 3
      "0000011" when "01000100000100000", -- t[34848] = 3
      "0000011" when "01000100000100001", -- t[34849] = 3
      "0000011" when "01000100000100010", -- t[34850] = 3
      "0000011" when "01000100000100011", -- t[34851] = 3
      "0000011" when "01000100000100100", -- t[34852] = 3
      "0000011" when "01000100000100101", -- t[34853] = 3
      "0000011" when "01000100000100110", -- t[34854] = 3
      "0000011" when "01000100000100111", -- t[34855] = 3
      "0000011" when "01000100000101000", -- t[34856] = 3
      "0000011" when "01000100000101001", -- t[34857] = 3
      "0000011" when "01000100000101010", -- t[34858] = 3
      "0000011" when "01000100000101011", -- t[34859] = 3
      "0000011" when "01000100000101100", -- t[34860] = 3
      "0000011" when "01000100000101101", -- t[34861] = 3
      "0000011" when "01000100000101110", -- t[34862] = 3
      "0000011" when "01000100000101111", -- t[34863] = 3
      "0000011" when "01000100000110000", -- t[34864] = 3
      "0000011" when "01000100000110001", -- t[34865] = 3
      "0000011" when "01000100000110010", -- t[34866] = 3
      "0000011" when "01000100000110011", -- t[34867] = 3
      "0000011" when "01000100000110100", -- t[34868] = 3
      "0000011" when "01000100000110101", -- t[34869] = 3
      "0000011" when "01000100000110110", -- t[34870] = 3
      "0000011" when "01000100000110111", -- t[34871] = 3
      "0000011" when "01000100000111000", -- t[34872] = 3
      "0000011" when "01000100000111001", -- t[34873] = 3
      "0000011" when "01000100000111010", -- t[34874] = 3
      "0000011" when "01000100000111011", -- t[34875] = 3
      "0000011" when "01000100000111100", -- t[34876] = 3
      "0000011" when "01000100000111101", -- t[34877] = 3
      "0000011" when "01000100000111110", -- t[34878] = 3
      "0000011" when "01000100000111111", -- t[34879] = 3
      "0000011" when "01000100001000000", -- t[34880] = 3
      "0000011" when "01000100001000001", -- t[34881] = 3
      "0000011" when "01000100001000010", -- t[34882] = 3
      "0000011" when "01000100001000011", -- t[34883] = 3
      "0000011" when "01000100001000100", -- t[34884] = 3
      "0000011" when "01000100001000101", -- t[34885] = 3
      "0000011" when "01000100001000110", -- t[34886] = 3
      "0000011" when "01000100001000111", -- t[34887] = 3
      "0000011" when "01000100001001000", -- t[34888] = 3
      "0000011" when "01000100001001001", -- t[34889] = 3
      "0000011" when "01000100001001010", -- t[34890] = 3
      "0000011" when "01000100001001011", -- t[34891] = 3
      "0000011" when "01000100001001100", -- t[34892] = 3
      "0000011" when "01000100001001101", -- t[34893] = 3
      "0000011" when "01000100001001110", -- t[34894] = 3
      "0000011" when "01000100001001111", -- t[34895] = 3
      "0000011" when "01000100001010000", -- t[34896] = 3
      "0000011" when "01000100001010001", -- t[34897] = 3
      "0000011" when "01000100001010010", -- t[34898] = 3
      "0000011" when "01000100001010011", -- t[34899] = 3
      "0000011" when "01000100001010100", -- t[34900] = 3
      "0000011" when "01000100001010101", -- t[34901] = 3
      "0000011" when "01000100001010110", -- t[34902] = 3
      "0000011" when "01000100001010111", -- t[34903] = 3
      "0000011" when "01000100001011000", -- t[34904] = 3
      "0000011" when "01000100001011001", -- t[34905] = 3
      "0000011" when "01000100001011010", -- t[34906] = 3
      "0000011" when "01000100001011011", -- t[34907] = 3
      "0000011" when "01000100001011100", -- t[34908] = 3
      "0000011" when "01000100001011101", -- t[34909] = 3
      "0000011" when "01000100001011110", -- t[34910] = 3
      "0000011" when "01000100001011111", -- t[34911] = 3
      "0000011" when "01000100001100000", -- t[34912] = 3
      "0000011" when "01000100001100001", -- t[34913] = 3
      "0000011" when "01000100001100010", -- t[34914] = 3
      "0000011" when "01000100001100011", -- t[34915] = 3
      "0000011" when "01000100001100100", -- t[34916] = 3
      "0000011" when "01000100001100101", -- t[34917] = 3
      "0000011" when "01000100001100110", -- t[34918] = 3
      "0000011" when "01000100001100111", -- t[34919] = 3
      "0000011" when "01000100001101000", -- t[34920] = 3
      "0000011" when "01000100001101001", -- t[34921] = 3
      "0000011" when "01000100001101010", -- t[34922] = 3
      "0000011" when "01000100001101011", -- t[34923] = 3
      "0000011" when "01000100001101100", -- t[34924] = 3
      "0000011" when "01000100001101101", -- t[34925] = 3
      "0000011" when "01000100001101110", -- t[34926] = 3
      "0000011" when "01000100001101111", -- t[34927] = 3
      "0000011" when "01000100001110000", -- t[34928] = 3
      "0000011" when "01000100001110001", -- t[34929] = 3
      "0000011" when "01000100001110010", -- t[34930] = 3
      "0000011" when "01000100001110011", -- t[34931] = 3
      "0000011" when "01000100001110100", -- t[34932] = 3
      "0000011" when "01000100001110101", -- t[34933] = 3
      "0000011" when "01000100001110110", -- t[34934] = 3
      "0000011" when "01000100001110111", -- t[34935] = 3
      "0000011" when "01000100001111000", -- t[34936] = 3
      "0000011" when "01000100001111001", -- t[34937] = 3
      "0000011" when "01000100001111010", -- t[34938] = 3
      "0000011" when "01000100001111011", -- t[34939] = 3
      "0000011" when "01000100001111100", -- t[34940] = 3
      "0000011" when "01000100001111101", -- t[34941] = 3
      "0000011" when "01000100001111110", -- t[34942] = 3
      "0000011" when "01000100001111111", -- t[34943] = 3
      "0000011" when "01000100010000000", -- t[34944] = 3
      "0000011" when "01000100010000001", -- t[34945] = 3
      "0000011" when "01000100010000010", -- t[34946] = 3
      "0000011" when "01000100010000011", -- t[34947] = 3
      "0000011" when "01000100010000100", -- t[34948] = 3
      "0000011" when "01000100010000101", -- t[34949] = 3
      "0000011" when "01000100010000110", -- t[34950] = 3
      "0000011" when "01000100010000111", -- t[34951] = 3
      "0000011" when "01000100010001000", -- t[34952] = 3
      "0000011" when "01000100010001001", -- t[34953] = 3
      "0000011" when "01000100010001010", -- t[34954] = 3
      "0000011" when "01000100010001011", -- t[34955] = 3
      "0000011" when "01000100010001100", -- t[34956] = 3
      "0000011" when "01000100010001101", -- t[34957] = 3
      "0000011" when "01000100010001110", -- t[34958] = 3
      "0000011" when "01000100010001111", -- t[34959] = 3
      "0000011" when "01000100010010000", -- t[34960] = 3
      "0000011" when "01000100010010001", -- t[34961] = 3
      "0000011" when "01000100010010010", -- t[34962] = 3
      "0000011" when "01000100010010011", -- t[34963] = 3
      "0000011" when "01000100010010100", -- t[34964] = 3
      "0000011" when "01000100010010101", -- t[34965] = 3
      "0000011" when "01000100010010110", -- t[34966] = 3
      "0000011" when "01000100010010111", -- t[34967] = 3
      "0000011" when "01000100010011000", -- t[34968] = 3
      "0000011" when "01000100010011001", -- t[34969] = 3
      "0000011" when "01000100010011010", -- t[34970] = 3
      "0000011" when "01000100010011011", -- t[34971] = 3
      "0000011" when "01000100010011100", -- t[34972] = 3
      "0000011" when "01000100010011101", -- t[34973] = 3
      "0000011" when "01000100010011110", -- t[34974] = 3
      "0000011" when "01000100010011111", -- t[34975] = 3
      "0000011" when "01000100010100000", -- t[34976] = 3
      "0000011" when "01000100010100001", -- t[34977] = 3
      "0000011" when "01000100010100010", -- t[34978] = 3
      "0000011" when "01000100010100011", -- t[34979] = 3
      "0000011" when "01000100010100100", -- t[34980] = 3
      "0000011" when "01000100010100101", -- t[34981] = 3
      "0000011" when "01000100010100110", -- t[34982] = 3
      "0000011" when "01000100010100111", -- t[34983] = 3
      "0000011" when "01000100010101000", -- t[34984] = 3
      "0000011" when "01000100010101001", -- t[34985] = 3
      "0000011" when "01000100010101010", -- t[34986] = 3
      "0000011" when "01000100010101011", -- t[34987] = 3
      "0000011" when "01000100010101100", -- t[34988] = 3
      "0000011" when "01000100010101101", -- t[34989] = 3
      "0000011" when "01000100010101110", -- t[34990] = 3
      "0000011" when "01000100010101111", -- t[34991] = 3
      "0000011" when "01000100010110000", -- t[34992] = 3
      "0000011" when "01000100010110001", -- t[34993] = 3
      "0000011" when "01000100010110010", -- t[34994] = 3
      "0000011" when "01000100010110011", -- t[34995] = 3
      "0000011" when "01000100010110100", -- t[34996] = 3
      "0000011" when "01000100010110101", -- t[34997] = 3
      "0000011" when "01000100010110110", -- t[34998] = 3
      "0000011" when "01000100010110111", -- t[34999] = 3
      "0000011" when "01000100010111000", -- t[35000] = 3
      "0000011" when "01000100010111001", -- t[35001] = 3
      "0000011" when "01000100010111010", -- t[35002] = 3
      "0000011" when "01000100010111011", -- t[35003] = 3
      "0000011" when "01000100010111100", -- t[35004] = 3
      "0000011" when "01000100010111101", -- t[35005] = 3
      "0000011" when "01000100010111110", -- t[35006] = 3
      "0000011" when "01000100010111111", -- t[35007] = 3
      "0000011" when "01000100011000000", -- t[35008] = 3
      "0000011" when "01000100011000001", -- t[35009] = 3
      "0000011" when "01000100011000010", -- t[35010] = 3
      "0000011" when "01000100011000011", -- t[35011] = 3
      "0000011" when "01000100011000100", -- t[35012] = 3
      "0000011" when "01000100011000101", -- t[35013] = 3
      "0000011" when "01000100011000110", -- t[35014] = 3
      "0000011" when "01000100011000111", -- t[35015] = 3
      "0000011" when "01000100011001000", -- t[35016] = 3
      "0000011" when "01000100011001001", -- t[35017] = 3
      "0000011" when "01000100011001010", -- t[35018] = 3
      "0000011" when "01000100011001011", -- t[35019] = 3
      "0000011" when "01000100011001100", -- t[35020] = 3
      "0000011" when "01000100011001101", -- t[35021] = 3
      "0000011" when "01000100011001110", -- t[35022] = 3
      "0000011" when "01000100011001111", -- t[35023] = 3
      "0000011" when "01000100011010000", -- t[35024] = 3
      "0000011" when "01000100011010001", -- t[35025] = 3
      "0000011" when "01000100011010010", -- t[35026] = 3
      "0000011" when "01000100011010011", -- t[35027] = 3
      "0000011" when "01000100011010100", -- t[35028] = 3
      "0000011" when "01000100011010101", -- t[35029] = 3
      "0000011" when "01000100011010110", -- t[35030] = 3
      "0000011" when "01000100011010111", -- t[35031] = 3
      "0000011" when "01000100011011000", -- t[35032] = 3
      "0000011" when "01000100011011001", -- t[35033] = 3
      "0000011" when "01000100011011010", -- t[35034] = 3
      "0000011" when "01000100011011011", -- t[35035] = 3
      "0000011" when "01000100011011100", -- t[35036] = 3
      "0000011" when "01000100011011101", -- t[35037] = 3
      "0000011" when "01000100011011110", -- t[35038] = 3
      "0000011" when "01000100011011111", -- t[35039] = 3
      "0000011" when "01000100011100000", -- t[35040] = 3
      "0000011" when "01000100011100001", -- t[35041] = 3
      "0000011" when "01000100011100010", -- t[35042] = 3
      "0000011" when "01000100011100011", -- t[35043] = 3
      "0000011" when "01000100011100100", -- t[35044] = 3
      "0000011" when "01000100011100101", -- t[35045] = 3
      "0000011" when "01000100011100110", -- t[35046] = 3
      "0000011" when "01000100011100111", -- t[35047] = 3
      "0000011" when "01000100011101000", -- t[35048] = 3
      "0000100" when "01000100011101001", -- t[35049] = 4
      "0000100" when "01000100011101010", -- t[35050] = 4
      "0000100" when "01000100011101011", -- t[35051] = 4
      "0000100" when "01000100011101100", -- t[35052] = 4
      "0000100" when "01000100011101101", -- t[35053] = 4
      "0000100" when "01000100011101110", -- t[35054] = 4
      "0000100" when "01000100011101111", -- t[35055] = 4
      "0000100" when "01000100011110000", -- t[35056] = 4
      "0000100" when "01000100011110001", -- t[35057] = 4
      "0000100" when "01000100011110010", -- t[35058] = 4
      "0000100" when "01000100011110011", -- t[35059] = 4
      "0000100" when "01000100011110100", -- t[35060] = 4
      "0000100" when "01000100011110101", -- t[35061] = 4
      "0000100" when "01000100011110110", -- t[35062] = 4
      "0000100" when "01000100011110111", -- t[35063] = 4
      "0000100" when "01000100011111000", -- t[35064] = 4
      "0000100" when "01000100011111001", -- t[35065] = 4
      "0000100" when "01000100011111010", -- t[35066] = 4
      "0000100" when "01000100011111011", -- t[35067] = 4
      "0000100" when "01000100011111100", -- t[35068] = 4
      "0000100" when "01000100011111101", -- t[35069] = 4
      "0000100" when "01000100011111110", -- t[35070] = 4
      "0000100" when "01000100011111111", -- t[35071] = 4
      "0000100" when "01000100100000000", -- t[35072] = 4
      "0000100" when "01000100100000001", -- t[35073] = 4
      "0000100" when "01000100100000010", -- t[35074] = 4
      "0000100" when "01000100100000011", -- t[35075] = 4
      "0000100" when "01000100100000100", -- t[35076] = 4
      "0000100" when "01000100100000101", -- t[35077] = 4
      "0000100" when "01000100100000110", -- t[35078] = 4
      "0000100" when "01000100100000111", -- t[35079] = 4
      "0000100" when "01000100100001000", -- t[35080] = 4
      "0000100" when "01000100100001001", -- t[35081] = 4
      "0000100" when "01000100100001010", -- t[35082] = 4
      "0000100" when "01000100100001011", -- t[35083] = 4
      "0000100" when "01000100100001100", -- t[35084] = 4
      "0000100" when "01000100100001101", -- t[35085] = 4
      "0000100" when "01000100100001110", -- t[35086] = 4
      "0000100" when "01000100100001111", -- t[35087] = 4
      "0000100" when "01000100100010000", -- t[35088] = 4
      "0000100" when "01000100100010001", -- t[35089] = 4
      "0000100" when "01000100100010010", -- t[35090] = 4
      "0000100" when "01000100100010011", -- t[35091] = 4
      "0000100" when "01000100100010100", -- t[35092] = 4
      "0000100" when "01000100100010101", -- t[35093] = 4
      "0000100" when "01000100100010110", -- t[35094] = 4
      "0000100" when "01000100100010111", -- t[35095] = 4
      "0000100" when "01000100100011000", -- t[35096] = 4
      "0000100" when "01000100100011001", -- t[35097] = 4
      "0000100" when "01000100100011010", -- t[35098] = 4
      "0000100" when "01000100100011011", -- t[35099] = 4
      "0000100" when "01000100100011100", -- t[35100] = 4
      "0000100" when "01000100100011101", -- t[35101] = 4
      "0000100" when "01000100100011110", -- t[35102] = 4
      "0000100" when "01000100100011111", -- t[35103] = 4
      "0000100" when "01000100100100000", -- t[35104] = 4
      "0000100" when "01000100100100001", -- t[35105] = 4
      "0000100" when "01000100100100010", -- t[35106] = 4
      "0000100" when "01000100100100011", -- t[35107] = 4
      "0000100" when "01000100100100100", -- t[35108] = 4
      "0000100" when "01000100100100101", -- t[35109] = 4
      "0000100" when "01000100100100110", -- t[35110] = 4
      "0000100" when "01000100100100111", -- t[35111] = 4
      "0000100" when "01000100100101000", -- t[35112] = 4
      "0000100" when "01000100100101001", -- t[35113] = 4
      "0000100" when "01000100100101010", -- t[35114] = 4
      "0000100" when "01000100100101011", -- t[35115] = 4
      "0000100" when "01000100100101100", -- t[35116] = 4
      "0000100" when "01000100100101101", -- t[35117] = 4
      "0000100" when "01000100100101110", -- t[35118] = 4
      "0000100" when "01000100100101111", -- t[35119] = 4
      "0000100" when "01000100100110000", -- t[35120] = 4
      "0000100" when "01000100100110001", -- t[35121] = 4
      "0000100" when "01000100100110010", -- t[35122] = 4
      "0000100" when "01000100100110011", -- t[35123] = 4
      "0000100" when "01000100100110100", -- t[35124] = 4
      "0000100" when "01000100100110101", -- t[35125] = 4
      "0000100" when "01000100100110110", -- t[35126] = 4
      "0000100" when "01000100100110111", -- t[35127] = 4
      "0000100" when "01000100100111000", -- t[35128] = 4
      "0000100" when "01000100100111001", -- t[35129] = 4
      "0000100" when "01000100100111010", -- t[35130] = 4
      "0000100" when "01000100100111011", -- t[35131] = 4
      "0000100" when "01000100100111100", -- t[35132] = 4
      "0000100" when "01000100100111101", -- t[35133] = 4
      "0000100" when "01000100100111110", -- t[35134] = 4
      "0000100" when "01000100100111111", -- t[35135] = 4
      "0000100" when "01000100101000000", -- t[35136] = 4
      "0000100" when "01000100101000001", -- t[35137] = 4
      "0000100" when "01000100101000010", -- t[35138] = 4
      "0000100" when "01000100101000011", -- t[35139] = 4
      "0000100" when "01000100101000100", -- t[35140] = 4
      "0000100" when "01000100101000101", -- t[35141] = 4
      "0000100" when "01000100101000110", -- t[35142] = 4
      "0000100" when "01000100101000111", -- t[35143] = 4
      "0000100" when "01000100101001000", -- t[35144] = 4
      "0000100" when "01000100101001001", -- t[35145] = 4
      "0000100" when "01000100101001010", -- t[35146] = 4
      "0000100" when "01000100101001011", -- t[35147] = 4
      "0000100" when "01000100101001100", -- t[35148] = 4
      "0000100" when "01000100101001101", -- t[35149] = 4
      "0000100" when "01000100101001110", -- t[35150] = 4
      "0000100" when "01000100101001111", -- t[35151] = 4
      "0000100" when "01000100101010000", -- t[35152] = 4
      "0000100" when "01000100101010001", -- t[35153] = 4
      "0000100" when "01000100101010010", -- t[35154] = 4
      "0000100" when "01000100101010011", -- t[35155] = 4
      "0000100" when "01000100101010100", -- t[35156] = 4
      "0000100" when "01000100101010101", -- t[35157] = 4
      "0000100" when "01000100101010110", -- t[35158] = 4
      "0000100" when "01000100101010111", -- t[35159] = 4
      "0000100" when "01000100101011000", -- t[35160] = 4
      "0000100" when "01000100101011001", -- t[35161] = 4
      "0000100" when "01000100101011010", -- t[35162] = 4
      "0000100" when "01000100101011011", -- t[35163] = 4
      "0000100" when "01000100101011100", -- t[35164] = 4
      "0000100" when "01000100101011101", -- t[35165] = 4
      "0000100" when "01000100101011110", -- t[35166] = 4
      "0000100" when "01000100101011111", -- t[35167] = 4
      "0000100" when "01000100101100000", -- t[35168] = 4
      "0000100" when "01000100101100001", -- t[35169] = 4
      "0000100" when "01000100101100010", -- t[35170] = 4
      "0000100" when "01000100101100011", -- t[35171] = 4
      "0000100" when "01000100101100100", -- t[35172] = 4
      "0000100" when "01000100101100101", -- t[35173] = 4
      "0000100" when "01000100101100110", -- t[35174] = 4
      "0000100" when "01000100101100111", -- t[35175] = 4
      "0000100" when "01000100101101000", -- t[35176] = 4
      "0000100" when "01000100101101001", -- t[35177] = 4
      "0000100" when "01000100101101010", -- t[35178] = 4
      "0000100" when "01000100101101011", -- t[35179] = 4
      "0000100" when "01000100101101100", -- t[35180] = 4
      "0000100" when "01000100101101101", -- t[35181] = 4
      "0000100" when "01000100101101110", -- t[35182] = 4
      "0000100" when "01000100101101111", -- t[35183] = 4
      "0000100" when "01000100101110000", -- t[35184] = 4
      "0000100" when "01000100101110001", -- t[35185] = 4
      "0000100" when "01000100101110010", -- t[35186] = 4
      "0000100" when "01000100101110011", -- t[35187] = 4
      "0000100" when "01000100101110100", -- t[35188] = 4
      "0000100" when "01000100101110101", -- t[35189] = 4
      "0000100" when "01000100101110110", -- t[35190] = 4
      "0000100" when "01000100101110111", -- t[35191] = 4
      "0000100" when "01000100101111000", -- t[35192] = 4
      "0000100" when "01000100101111001", -- t[35193] = 4
      "0000100" when "01000100101111010", -- t[35194] = 4
      "0000100" when "01000100101111011", -- t[35195] = 4
      "0000100" when "01000100101111100", -- t[35196] = 4
      "0000100" when "01000100101111101", -- t[35197] = 4
      "0000100" when "01000100101111110", -- t[35198] = 4
      "0000100" when "01000100101111111", -- t[35199] = 4
      "0000100" when "01000100110000000", -- t[35200] = 4
      "0000100" when "01000100110000001", -- t[35201] = 4
      "0000100" when "01000100110000010", -- t[35202] = 4
      "0000100" when "01000100110000011", -- t[35203] = 4
      "0000100" when "01000100110000100", -- t[35204] = 4
      "0000100" when "01000100110000101", -- t[35205] = 4
      "0000100" when "01000100110000110", -- t[35206] = 4
      "0000100" when "01000100110000111", -- t[35207] = 4
      "0000100" when "01000100110001000", -- t[35208] = 4
      "0000100" when "01000100110001001", -- t[35209] = 4
      "0000100" when "01000100110001010", -- t[35210] = 4
      "0000100" when "01000100110001011", -- t[35211] = 4
      "0000100" when "01000100110001100", -- t[35212] = 4
      "0000100" when "01000100110001101", -- t[35213] = 4
      "0000100" when "01000100110001110", -- t[35214] = 4
      "0000100" when "01000100110001111", -- t[35215] = 4
      "0000100" when "01000100110010000", -- t[35216] = 4
      "0000100" when "01000100110010001", -- t[35217] = 4
      "0000100" when "01000100110010010", -- t[35218] = 4
      "0000100" when "01000100110010011", -- t[35219] = 4
      "0000100" when "01000100110010100", -- t[35220] = 4
      "0000100" when "01000100110010101", -- t[35221] = 4
      "0000100" when "01000100110010110", -- t[35222] = 4
      "0000100" when "01000100110010111", -- t[35223] = 4
      "0000100" when "01000100110011000", -- t[35224] = 4
      "0000100" when "01000100110011001", -- t[35225] = 4
      "0000100" when "01000100110011010", -- t[35226] = 4
      "0000100" when "01000100110011011", -- t[35227] = 4
      "0000100" when "01000100110011100", -- t[35228] = 4
      "0000100" when "01000100110011101", -- t[35229] = 4
      "0000100" when "01000100110011110", -- t[35230] = 4
      "0000100" when "01000100110011111", -- t[35231] = 4
      "0000100" when "01000100110100000", -- t[35232] = 4
      "0000100" when "01000100110100001", -- t[35233] = 4
      "0000100" when "01000100110100010", -- t[35234] = 4
      "0000100" when "01000100110100011", -- t[35235] = 4
      "0000100" when "01000100110100100", -- t[35236] = 4
      "0000100" when "01000100110100101", -- t[35237] = 4
      "0000100" when "01000100110100110", -- t[35238] = 4
      "0000100" when "01000100110100111", -- t[35239] = 4
      "0000100" when "01000100110101000", -- t[35240] = 4
      "0000100" when "01000100110101001", -- t[35241] = 4
      "0000100" when "01000100110101010", -- t[35242] = 4
      "0000100" when "01000100110101011", -- t[35243] = 4
      "0000100" when "01000100110101100", -- t[35244] = 4
      "0000100" when "01000100110101101", -- t[35245] = 4
      "0000100" when "01000100110101110", -- t[35246] = 4
      "0000100" when "01000100110101111", -- t[35247] = 4
      "0000100" when "01000100110110000", -- t[35248] = 4
      "0000100" when "01000100110110001", -- t[35249] = 4
      "0000100" when "01000100110110010", -- t[35250] = 4
      "0000100" when "01000100110110011", -- t[35251] = 4
      "0000100" when "01000100110110100", -- t[35252] = 4
      "0000100" when "01000100110110101", -- t[35253] = 4
      "0000100" when "01000100110110110", -- t[35254] = 4
      "0000100" when "01000100110110111", -- t[35255] = 4
      "0000100" when "01000100110111000", -- t[35256] = 4
      "0000100" when "01000100110111001", -- t[35257] = 4
      "0000100" when "01000100110111010", -- t[35258] = 4
      "0000100" when "01000100110111011", -- t[35259] = 4
      "0000100" when "01000100110111100", -- t[35260] = 4
      "0000100" when "01000100110111101", -- t[35261] = 4
      "0000100" when "01000100110111110", -- t[35262] = 4
      "0000100" when "01000100110111111", -- t[35263] = 4
      "0000100" when "01000100111000000", -- t[35264] = 4
      "0000100" when "01000100111000001", -- t[35265] = 4
      "0000100" when "01000100111000010", -- t[35266] = 4
      "0000100" when "01000100111000011", -- t[35267] = 4
      "0000100" when "01000100111000100", -- t[35268] = 4
      "0000100" when "01000100111000101", -- t[35269] = 4
      "0000100" when "01000100111000110", -- t[35270] = 4
      "0000100" when "01000100111000111", -- t[35271] = 4
      "0000100" when "01000100111001000", -- t[35272] = 4
      "0000100" when "01000100111001001", -- t[35273] = 4
      "0000100" when "01000100111001010", -- t[35274] = 4
      "0000100" when "01000100111001011", -- t[35275] = 4
      "0000100" when "01000100111001100", -- t[35276] = 4
      "0000100" when "01000100111001101", -- t[35277] = 4
      "0000100" when "01000100111001110", -- t[35278] = 4
      "0000100" when "01000100111001111", -- t[35279] = 4
      "0000100" when "01000100111010000", -- t[35280] = 4
      "0000100" when "01000100111010001", -- t[35281] = 4
      "0000100" when "01000100111010010", -- t[35282] = 4
      "0000100" when "01000100111010011", -- t[35283] = 4
      "0000100" when "01000100111010100", -- t[35284] = 4
      "0000100" when "01000100111010101", -- t[35285] = 4
      "0000100" when "01000100111010110", -- t[35286] = 4
      "0000100" when "01000100111010111", -- t[35287] = 4
      "0000100" when "01000100111011000", -- t[35288] = 4
      "0000100" when "01000100111011001", -- t[35289] = 4
      "0000100" when "01000100111011010", -- t[35290] = 4
      "0000100" when "01000100111011011", -- t[35291] = 4
      "0000100" when "01000100111011100", -- t[35292] = 4
      "0000100" when "01000100111011101", -- t[35293] = 4
      "0000100" when "01000100111011110", -- t[35294] = 4
      "0000100" when "01000100111011111", -- t[35295] = 4
      "0000100" when "01000100111100000", -- t[35296] = 4
      "0000100" when "01000100111100001", -- t[35297] = 4
      "0000100" when "01000100111100010", -- t[35298] = 4
      "0000100" when "01000100111100011", -- t[35299] = 4
      "0000100" when "01000100111100100", -- t[35300] = 4
      "0000100" when "01000100111100101", -- t[35301] = 4
      "0000100" when "01000100111100110", -- t[35302] = 4
      "0000100" when "01000100111100111", -- t[35303] = 4
      "0000100" when "01000100111101000", -- t[35304] = 4
      "0000100" when "01000100111101001", -- t[35305] = 4
      "0000100" when "01000100111101010", -- t[35306] = 4
      "0000100" when "01000100111101011", -- t[35307] = 4
      "0000100" when "01000100111101100", -- t[35308] = 4
      "0000100" when "01000100111101101", -- t[35309] = 4
      "0000100" when "01000100111101110", -- t[35310] = 4
      "0000100" when "01000100111101111", -- t[35311] = 4
      "0000100" when "01000100111110000", -- t[35312] = 4
      "0000100" when "01000100111110001", -- t[35313] = 4
      "0000100" when "01000100111110010", -- t[35314] = 4
      "0000100" when "01000100111110011", -- t[35315] = 4
      "0000100" when "01000100111110100", -- t[35316] = 4
      "0000100" when "01000100111110101", -- t[35317] = 4
      "0000100" when "01000100111110110", -- t[35318] = 4
      "0000100" when "01000100111110111", -- t[35319] = 4
      "0000100" when "01000100111111000", -- t[35320] = 4
      "0000100" when "01000100111111001", -- t[35321] = 4
      "0000100" when "01000100111111010", -- t[35322] = 4
      "0000100" when "01000100111111011", -- t[35323] = 4
      "0000100" when "01000100111111100", -- t[35324] = 4
      "0000100" when "01000100111111101", -- t[35325] = 4
      "0000100" when "01000100111111110", -- t[35326] = 4
      "0000100" when "01000100111111111", -- t[35327] = 4
      "0000100" when "01000101000000000", -- t[35328] = 4
      "0000100" when "01000101000000001", -- t[35329] = 4
      "0000100" when "01000101000000010", -- t[35330] = 4
      "0000100" when "01000101000000011", -- t[35331] = 4
      "0000100" when "01000101000000100", -- t[35332] = 4
      "0000100" when "01000101000000101", -- t[35333] = 4
      "0000100" when "01000101000000110", -- t[35334] = 4
      "0000100" when "01000101000000111", -- t[35335] = 4
      "0000100" when "01000101000001000", -- t[35336] = 4
      "0000100" when "01000101000001001", -- t[35337] = 4
      "0000100" when "01000101000001010", -- t[35338] = 4
      "0000100" when "01000101000001011", -- t[35339] = 4
      "0000100" when "01000101000001100", -- t[35340] = 4
      "0000100" when "01000101000001101", -- t[35341] = 4
      "0000100" when "01000101000001110", -- t[35342] = 4
      "0000100" when "01000101000001111", -- t[35343] = 4
      "0000100" when "01000101000010000", -- t[35344] = 4
      "0000100" when "01000101000010001", -- t[35345] = 4
      "0000100" when "01000101000010010", -- t[35346] = 4
      "0000100" when "01000101000010011", -- t[35347] = 4
      "0000100" when "01000101000010100", -- t[35348] = 4
      "0000100" when "01000101000010101", -- t[35349] = 4
      "0000100" when "01000101000010110", -- t[35350] = 4
      "0000100" when "01000101000010111", -- t[35351] = 4
      "0000100" when "01000101000011000", -- t[35352] = 4
      "0000100" when "01000101000011001", -- t[35353] = 4
      "0000100" when "01000101000011010", -- t[35354] = 4
      "0000100" when "01000101000011011", -- t[35355] = 4
      "0000100" when "01000101000011100", -- t[35356] = 4
      "0000100" when "01000101000011101", -- t[35357] = 4
      "0000100" when "01000101000011110", -- t[35358] = 4
      "0000100" when "01000101000011111", -- t[35359] = 4
      "0000100" when "01000101000100000", -- t[35360] = 4
      "0000100" when "01000101000100001", -- t[35361] = 4
      "0000100" when "01000101000100010", -- t[35362] = 4
      "0000100" when "01000101000100011", -- t[35363] = 4
      "0000100" when "01000101000100100", -- t[35364] = 4
      "0000100" when "01000101000100101", -- t[35365] = 4
      "0000100" when "01000101000100110", -- t[35366] = 4
      "0000100" when "01000101000100111", -- t[35367] = 4
      "0000100" when "01000101000101000", -- t[35368] = 4
      "0000100" when "01000101000101001", -- t[35369] = 4
      "0000100" when "01000101000101010", -- t[35370] = 4
      "0000100" when "01000101000101011", -- t[35371] = 4
      "0000100" when "01000101000101100", -- t[35372] = 4
      "0000100" when "01000101000101101", -- t[35373] = 4
      "0000100" when "01000101000101110", -- t[35374] = 4
      "0000100" when "01000101000101111", -- t[35375] = 4
      "0000100" when "01000101000110000", -- t[35376] = 4
      "0000100" when "01000101000110001", -- t[35377] = 4
      "0000100" when "01000101000110010", -- t[35378] = 4
      "0000100" when "01000101000110011", -- t[35379] = 4
      "0000100" when "01000101000110100", -- t[35380] = 4
      "0000100" when "01000101000110101", -- t[35381] = 4
      "0000100" when "01000101000110110", -- t[35382] = 4
      "0000100" when "01000101000110111", -- t[35383] = 4
      "0000100" when "01000101000111000", -- t[35384] = 4
      "0000100" when "01000101000111001", -- t[35385] = 4
      "0000100" when "01000101000111010", -- t[35386] = 4
      "0000100" when "01000101000111011", -- t[35387] = 4
      "0000100" when "01000101000111100", -- t[35388] = 4
      "0000100" when "01000101000111101", -- t[35389] = 4
      "0000100" when "01000101000111110", -- t[35390] = 4
      "0000100" when "01000101000111111", -- t[35391] = 4
      "0000100" when "01000101001000000", -- t[35392] = 4
      "0000100" when "01000101001000001", -- t[35393] = 4
      "0000100" when "01000101001000010", -- t[35394] = 4
      "0000100" when "01000101001000011", -- t[35395] = 4
      "0000100" when "01000101001000100", -- t[35396] = 4
      "0000100" when "01000101001000101", -- t[35397] = 4
      "0000100" when "01000101001000110", -- t[35398] = 4
      "0000100" when "01000101001000111", -- t[35399] = 4
      "0000100" when "01000101001001000", -- t[35400] = 4
      "0000100" when "01000101001001001", -- t[35401] = 4
      "0000100" when "01000101001001010", -- t[35402] = 4
      "0000100" when "01000101001001011", -- t[35403] = 4
      "0000100" when "01000101001001100", -- t[35404] = 4
      "0000100" when "01000101001001101", -- t[35405] = 4
      "0000100" when "01000101001001110", -- t[35406] = 4
      "0000100" when "01000101001001111", -- t[35407] = 4
      "0000100" when "01000101001010000", -- t[35408] = 4
      "0000100" when "01000101001010001", -- t[35409] = 4
      "0000100" when "01000101001010010", -- t[35410] = 4
      "0000100" when "01000101001010011", -- t[35411] = 4
      "0000100" when "01000101001010100", -- t[35412] = 4
      "0000100" when "01000101001010101", -- t[35413] = 4
      "0000100" when "01000101001010110", -- t[35414] = 4
      "0000100" when "01000101001010111", -- t[35415] = 4
      "0000100" when "01000101001011000", -- t[35416] = 4
      "0000100" when "01000101001011001", -- t[35417] = 4
      "0000100" when "01000101001011010", -- t[35418] = 4
      "0000100" when "01000101001011011", -- t[35419] = 4
      "0000100" when "01000101001011100", -- t[35420] = 4
      "0000100" when "01000101001011101", -- t[35421] = 4
      "0000100" when "01000101001011110", -- t[35422] = 4
      "0000100" when "01000101001011111", -- t[35423] = 4
      "0000100" when "01000101001100000", -- t[35424] = 4
      "0000100" when "01000101001100001", -- t[35425] = 4
      "0000100" when "01000101001100010", -- t[35426] = 4
      "0000100" when "01000101001100011", -- t[35427] = 4
      "0000100" when "01000101001100100", -- t[35428] = 4
      "0000100" when "01000101001100101", -- t[35429] = 4
      "0000100" when "01000101001100110", -- t[35430] = 4
      "0000100" when "01000101001100111", -- t[35431] = 4
      "0000100" when "01000101001101000", -- t[35432] = 4
      "0000100" when "01000101001101001", -- t[35433] = 4
      "0000100" when "01000101001101010", -- t[35434] = 4
      "0000100" when "01000101001101011", -- t[35435] = 4
      "0000100" when "01000101001101100", -- t[35436] = 4
      "0000100" when "01000101001101101", -- t[35437] = 4
      "0000100" when "01000101001101110", -- t[35438] = 4
      "0000100" when "01000101001101111", -- t[35439] = 4
      "0000100" when "01000101001110000", -- t[35440] = 4
      "0000100" when "01000101001110001", -- t[35441] = 4
      "0000100" when "01000101001110010", -- t[35442] = 4
      "0000100" when "01000101001110011", -- t[35443] = 4
      "0000100" when "01000101001110100", -- t[35444] = 4
      "0000100" when "01000101001110101", -- t[35445] = 4
      "0000100" when "01000101001110110", -- t[35446] = 4
      "0000100" when "01000101001110111", -- t[35447] = 4
      "0000100" when "01000101001111000", -- t[35448] = 4
      "0000100" when "01000101001111001", -- t[35449] = 4
      "0000100" when "01000101001111010", -- t[35450] = 4
      "0000100" when "01000101001111011", -- t[35451] = 4
      "0000100" when "01000101001111100", -- t[35452] = 4
      "0000100" when "01000101001111101", -- t[35453] = 4
      "0000100" when "01000101001111110", -- t[35454] = 4
      "0000100" when "01000101001111111", -- t[35455] = 4
      "0000100" when "01000101010000000", -- t[35456] = 4
      "0000100" when "01000101010000001", -- t[35457] = 4
      "0000100" when "01000101010000010", -- t[35458] = 4
      "0000100" when "01000101010000011", -- t[35459] = 4
      "0000100" when "01000101010000100", -- t[35460] = 4
      "0000100" when "01000101010000101", -- t[35461] = 4
      "0000100" when "01000101010000110", -- t[35462] = 4
      "0000100" when "01000101010000111", -- t[35463] = 4
      "0000100" when "01000101010001000", -- t[35464] = 4
      "0000100" when "01000101010001001", -- t[35465] = 4
      "0000100" when "01000101010001010", -- t[35466] = 4
      "0000100" when "01000101010001011", -- t[35467] = 4
      "0000100" when "01000101010001100", -- t[35468] = 4
      "0000100" when "01000101010001101", -- t[35469] = 4
      "0000100" when "01000101010001110", -- t[35470] = 4
      "0000100" when "01000101010001111", -- t[35471] = 4
      "0000100" when "01000101010010000", -- t[35472] = 4
      "0000100" when "01000101010010001", -- t[35473] = 4
      "0000100" when "01000101010010010", -- t[35474] = 4
      "0000100" when "01000101010010011", -- t[35475] = 4
      "0000100" when "01000101010010100", -- t[35476] = 4
      "0000100" when "01000101010010101", -- t[35477] = 4
      "0000100" when "01000101010010110", -- t[35478] = 4
      "0000100" when "01000101010010111", -- t[35479] = 4
      "0000100" when "01000101010011000", -- t[35480] = 4
      "0000100" when "01000101010011001", -- t[35481] = 4
      "0000100" when "01000101010011010", -- t[35482] = 4
      "0000100" when "01000101010011011", -- t[35483] = 4
      "0000100" when "01000101010011100", -- t[35484] = 4
      "0000100" when "01000101010011101", -- t[35485] = 4
      "0000100" when "01000101010011110", -- t[35486] = 4
      "0000100" when "01000101010011111", -- t[35487] = 4
      "0000100" when "01000101010100000", -- t[35488] = 4
      "0000100" when "01000101010100001", -- t[35489] = 4
      "0000100" when "01000101010100010", -- t[35490] = 4
      "0000100" when "01000101010100011", -- t[35491] = 4
      "0000100" when "01000101010100100", -- t[35492] = 4
      "0000100" when "01000101010100101", -- t[35493] = 4
      "0000100" when "01000101010100110", -- t[35494] = 4
      "0000100" when "01000101010100111", -- t[35495] = 4
      "0000100" when "01000101010101000", -- t[35496] = 4
      "0000100" when "01000101010101001", -- t[35497] = 4
      "0000100" when "01000101010101010", -- t[35498] = 4
      "0000100" when "01000101010101011", -- t[35499] = 4
      "0000100" when "01000101010101100", -- t[35500] = 4
      "0000100" when "01000101010101101", -- t[35501] = 4
      "0000100" when "01000101010101110", -- t[35502] = 4
      "0000100" when "01000101010101111", -- t[35503] = 4
      "0000100" when "01000101010110000", -- t[35504] = 4
      "0000100" when "01000101010110001", -- t[35505] = 4
      "0000100" when "01000101010110010", -- t[35506] = 4
      "0000100" when "01000101010110011", -- t[35507] = 4
      "0000100" when "01000101010110100", -- t[35508] = 4
      "0000100" when "01000101010110101", -- t[35509] = 4
      "0000100" when "01000101010110110", -- t[35510] = 4
      "0000100" when "01000101010110111", -- t[35511] = 4
      "0000100" when "01000101010111000", -- t[35512] = 4
      "0000100" when "01000101010111001", -- t[35513] = 4
      "0000100" when "01000101010111010", -- t[35514] = 4
      "0000100" when "01000101010111011", -- t[35515] = 4
      "0000100" when "01000101010111100", -- t[35516] = 4
      "0000100" when "01000101010111101", -- t[35517] = 4
      "0000100" when "01000101010111110", -- t[35518] = 4
      "0000100" when "01000101010111111", -- t[35519] = 4
      "0000100" when "01000101011000000", -- t[35520] = 4
      "0000100" when "01000101011000001", -- t[35521] = 4
      "0000100" when "01000101011000010", -- t[35522] = 4
      "0000100" when "01000101011000011", -- t[35523] = 4
      "0000100" when "01000101011000100", -- t[35524] = 4
      "0000100" when "01000101011000101", -- t[35525] = 4
      "0000100" when "01000101011000110", -- t[35526] = 4
      "0000100" when "01000101011000111", -- t[35527] = 4
      "0000100" when "01000101011001000", -- t[35528] = 4
      "0000100" when "01000101011001001", -- t[35529] = 4
      "0000100" when "01000101011001010", -- t[35530] = 4
      "0000100" when "01000101011001011", -- t[35531] = 4
      "0000100" when "01000101011001100", -- t[35532] = 4
      "0000100" when "01000101011001101", -- t[35533] = 4
      "0000100" when "01000101011001110", -- t[35534] = 4
      "0000100" when "01000101011001111", -- t[35535] = 4
      "0000100" when "01000101011010000", -- t[35536] = 4
      "0000100" when "01000101011010001", -- t[35537] = 4
      "0000100" when "01000101011010010", -- t[35538] = 4
      "0000100" when "01000101011010011", -- t[35539] = 4
      "0000100" when "01000101011010100", -- t[35540] = 4
      "0000100" when "01000101011010101", -- t[35541] = 4
      "0000100" when "01000101011010110", -- t[35542] = 4
      "0000100" when "01000101011010111", -- t[35543] = 4
      "0000100" when "01000101011011000", -- t[35544] = 4
      "0000100" when "01000101011011001", -- t[35545] = 4
      "0000100" when "01000101011011010", -- t[35546] = 4
      "0000100" when "01000101011011011", -- t[35547] = 4
      "0000100" when "01000101011011100", -- t[35548] = 4
      "0000100" when "01000101011011101", -- t[35549] = 4
      "0000100" when "01000101011011110", -- t[35550] = 4
      "0000100" when "01000101011011111", -- t[35551] = 4
      "0000100" when "01000101011100000", -- t[35552] = 4
      "0000100" when "01000101011100001", -- t[35553] = 4
      "0000100" when "01000101011100010", -- t[35554] = 4
      "0000100" when "01000101011100011", -- t[35555] = 4
      "0000100" when "01000101011100100", -- t[35556] = 4
      "0000100" when "01000101011100101", -- t[35557] = 4
      "0000100" when "01000101011100110", -- t[35558] = 4
      "0000100" when "01000101011100111", -- t[35559] = 4
      "0000100" when "01000101011101000", -- t[35560] = 4
      "0000100" when "01000101011101001", -- t[35561] = 4
      "0000100" when "01000101011101010", -- t[35562] = 4
      "0000100" when "01000101011101011", -- t[35563] = 4
      "0000100" when "01000101011101100", -- t[35564] = 4
      "0000100" when "01000101011101101", -- t[35565] = 4
      "0000100" when "01000101011101110", -- t[35566] = 4
      "0000100" when "01000101011101111", -- t[35567] = 4
      "0000100" when "01000101011110000", -- t[35568] = 4
      "0000100" when "01000101011110001", -- t[35569] = 4
      "0000100" when "01000101011110010", -- t[35570] = 4
      "0000100" when "01000101011110011", -- t[35571] = 4
      "0000100" when "01000101011110100", -- t[35572] = 4
      "0000100" when "01000101011110101", -- t[35573] = 4
      "0000100" when "01000101011110110", -- t[35574] = 4
      "0000100" when "01000101011110111", -- t[35575] = 4
      "0000100" when "01000101011111000", -- t[35576] = 4
      "0000100" when "01000101011111001", -- t[35577] = 4
      "0000100" when "01000101011111010", -- t[35578] = 4
      "0000100" when "01000101011111011", -- t[35579] = 4
      "0000100" when "01000101011111100", -- t[35580] = 4
      "0000100" when "01000101011111101", -- t[35581] = 4
      "0000100" when "01000101011111110", -- t[35582] = 4
      "0000100" when "01000101011111111", -- t[35583] = 4
      "0000100" when "01000101100000000", -- t[35584] = 4
      "0000100" when "01000101100000001", -- t[35585] = 4
      "0000100" when "01000101100000010", -- t[35586] = 4
      "0000100" when "01000101100000011", -- t[35587] = 4
      "0000100" when "01000101100000100", -- t[35588] = 4
      "0000100" when "01000101100000101", -- t[35589] = 4
      "0000100" when "01000101100000110", -- t[35590] = 4
      "0000100" when "01000101100000111", -- t[35591] = 4
      "0000100" when "01000101100001000", -- t[35592] = 4
      "0000100" when "01000101100001001", -- t[35593] = 4
      "0000100" when "01000101100001010", -- t[35594] = 4
      "0000100" when "01000101100001011", -- t[35595] = 4
      "0000100" when "01000101100001100", -- t[35596] = 4
      "0000100" when "01000101100001101", -- t[35597] = 4
      "0000100" when "01000101100001110", -- t[35598] = 4
      "0000100" when "01000101100001111", -- t[35599] = 4
      "0000100" when "01000101100010000", -- t[35600] = 4
      "0000100" when "01000101100010001", -- t[35601] = 4
      "0000100" when "01000101100010010", -- t[35602] = 4
      "0000100" when "01000101100010011", -- t[35603] = 4
      "0000100" when "01000101100010100", -- t[35604] = 4
      "0000100" when "01000101100010101", -- t[35605] = 4
      "0000100" when "01000101100010110", -- t[35606] = 4
      "0000100" when "01000101100010111", -- t[35607] = 4
      "0000100" when "01000101100011000", -- t[35608] = 4
      "0000100" when "01000101100011001", -- t[35609] = 4
      "0000100" when "01000101100011010", -- t[35610] = 4
      "0000100" when "01000101100011011", -- t[35611] = 4
      "0000100" when "01000101100011100", -- t[35612] = 4
      "0000100" when "01000101100011101", -- t[35613] = 4
      "0000100" when "01000101100011110", -- t[35614] = 4
      "0000100" when "01000101100011111", -- t[35615] = 4
      "0000100" when "01000101100100000", -- t[35616] = 4
      "0000100" when "01000101100100001", -- t[35617] = 4
      "0000100" when "01000101100100010", -- t[35618] = 4
      "0000100" when "01000101100100011", -- t[35619] = 4
      "0000100" when "01000101100100100", -- t[35620] = 4
      "0000100" when "01000101100100101", -- t[35621] = 4
      "0000100" when "01000101100100110", -- t[35622] = 4
      "0000100" when "01000101100100111", -- t[35623] = 4
      "0000100" when "01000101100101000", -- t[35624] = 4
      "0000100" when "01000101100101001", -- t[35625] = 4
      "0000100" when "01000101100101010", -- t[35626] = 4
      "0000100" when "01000101100101011", -- t[35627] = 4
      "0000100" when "01000101100101100", -- t[35628] = 4
      "0000100" when "01000101100101101", -- t[35629] = 4
      "0000100" when "01000101100101110", -- t[35630] = 4
      "0000100" when "01000101100101111", -- t[35631] = 4
      "0000100" when "01000101100110000", -- t[35632] = 4
      "0000100" when "01000101100110001", -- t[35633] = 4
      "0000100" when "01000101100110010", -- t[35634] = 4
      "0000100" when "01000101100110011", -- t[35635] = 4
      "0000100" when "01000101100110100", -- t[35636] = 4
      "0000100" when "01000101100110101", -- t[35637] = 4
      "0000100" when "01000101100110110", -- t[35638] = 4
      "0000100" when "01000101100110111", -- t[35639] = 4
      "0000100" when "01000101100111000", -- t[35640] = 4
      "0000100" when "01000101100111001", -- t[35641] = 4
      "0000100" when "01000101100111010", -- t[35642] = 4
      "0000100" when "01000101100111011", -- t[35643] = 4
      "0000100" when "01000101100111100", -- t[35644] = 4
      "0000100" when "01000101100111101", -- t[35645] = 4
      "0000100" when "01000101100111110", -- t[35646] = 4
      "0000100" when "01000101100111111", -- t[35647] = 4
      "0000100" when "01000101101000000", -- t[35648] = 4
      "0000100" when "01000101101000001", -- t[35649] = 4
      "0000100" when "01000101101000010", -- t[35650] = 4
      "0000100" when "01000101101000011", -- t[35651] = 4
      "0000100" when "01000101101000100", -- t[35652] = 4
      "0000100" when "01000101101000101", -- t[35653] = 4
      "0000100" when "01000101101000110", -- t[35654] = 4
      "0000100" when "01000101101000111", -- t[35655] = 4
      "0000100" when "01000101101001000", -- t[35656] = 4
      "0000100" when "01000101101001001", -- t[35657] = 4
      "0000100" when "01000101101001010", -- t[35658] = 4
      "0000100" when "01000101101001011", -- t[35659] = 4
      "0000100" when "01000101101001100", -- t[35660] = 4
      "0000100" when "01000101101001101", -- t[35661] = 4
      "0000100" when "01000101101001110", -- t[35662] = 4
      "0000100" when "01000101101001111", -- t[35663] = 4
      "0000100" when "01000101101010000", -- t[35664] = 4
      "0000100" when "01000101101010001", -- t[35665] = 4
      "0000100" when "01000101101010010", -- t[35666] = 4
      "0000100" when "01000101101010011", -- t[35667] = 4
      "0000100" when "01000101101010100", -- t[35668] = 4
      "0000100" when "01000101101010101", -- t[35669] = 4
      "0000100" when "01000101101010110", -- t[35670] = 4
      "0000100" when "01000101101010111", -- t[35671] = 4
      "0000100" when "01000101101011000", -- t[35672] = 4
      "0000100" when "01000101101011001", -- t[35673] = 4
      "0000100" when "01000101101011010", -- t[35674] = 4
      "0000100" when "01000101101011011", -- t[35675] = 4
      "0000100" when "01000101101011100", -- t[35676] = 4
      "0000100" when "01000101101011101", -- t[35677] = 4
      "0000100" when "01000101101011110", -- t[35678] = 4
      "0000100" when "01000101101011111", -- t[35679] = 4
      "0000100" when "01000101101100000", -- t[35680] = 4
      "0000100" when "01000101101100001", -- t[35681] = 4
      "0000100" when "01000101101100010", -- t[35682] = 4
      "0000100" when "01000101101100011", -- t[35683] = 4
      "0000100" when "01000101101100100", -- t[35684] = 4
      "0000100" when "01000101101100101", -- t[35685] = 4
      "0000100" when "01000101101100110", -- t[35686] = 4
      "0000100" when "01000101101100111", -- t[35687] = 4
      "0000100" when "01000101101101000", -- t[35688] = 4
      "0000100" when "01000101101101001", -- t[35689] = 4
      "0000100" when "01000101101101010", -- t[35690] = 4
      "0000100" when "01000101101101011", -- t[35691] = 4
      "0000100" when "01000101101101100", -- t[35692] = 4
      "0000100" when "01000101101101101", -- t[35693] = 4
      "0000100" when "01000101101101110", -- t[35694] = 4
      "0000100" when "01000101101101111", -- t[35695] = 4
      "0000100" when "01000101101110000", -- t[35696] = 4
      "0000100" when "01000101101110001", -- t[35697] = 4
      "0000100" when "01000101101110010", -- t[35698] = 4
      "0000100" when "01000101101110011", -- t[35699] = 4
      "0000100" when "01000101101110100", -- t[35700] = 4
      "0000100" when "01000101101110101", -- t[35701] = 4
      "0000100" when "01000101101110110", -- t[35702] = 4
      "0000100" when "01000101101110111", -- t[35703] = 4
      "0000100" when "01000101101111000", -- t[35704] = 4
      "0000100" when "01000101101111001", -- t[35705] = 4
      "0000100" when "01000101101111010", -- t[35706] = 4
      "0000100" when "01000101101111011", -- t[35707] = 4
      "0000100" when "01000101101111100", -- t[35708] = 4
      "0000100" when "01000101101111101", -- t[35709] = 4
      "0000100" when "01000101101111110", -- t[35710] = 4
      "0000100" when "01000101101111111", -- t[35711] = 4
      "0000100" when "01000101110000000", -- t[35712] = 4
      "0000100" when "01000101110000001", -- t[35713] = 4
      "0000100" when "01000101110000010", -- t[35714] = 4
      "0000100" when "01000101110000011", -- t[35715] = 4
      "0000100" when "01000101110000100", -- t[35716] = 4
      "0000100" when "01000101110000101", -- t[35717] = 4
      "0000100" when "01000101110000110", -- t[35718] = 4
      "0000100" when "01000101110000111", -- t[35719] = 4
      "0000100" when "01000101110001000", -- t[35720] = 4
      "0000100" when "01000101110001001", -- t[35721] = 4
      "0000100" when "01000101110001010", -- t[35722] = 4
      "0000100" when "01000101110001011", -- t[35723] = 4
      "0000100" when "01000101110001100", -- t[35724] = 4
      "0000100" when "01000101110001101", -- t[35725] = 4
      "0000100" when "01000101110001110", -- t[35726] = 4
      "0000100" when "01000101110001111", -- t[35727] = 4
      "0000100" when "01000101110010000", -- t[35728] = 4
      "0000100" when "01000101110010001", -- t[35729] = 4
      "0000100" when "01000101110010010", -- t[35730] = 4
      "0000100" when "01000101110010011", -- t[35731] = 4
      "0000100" when "01000101110010100", -- t[35732] = 4
      "0000100" when "01000101110010101", -- t[35733] = 4
      "0000100" when "01000101110010110", -- t[35734] = 4
      "0000100" when "01000101110010111", -- t[35735] = 4
      "0000100" when "01000101110011000", -- t[35736] = 4
      "0000100" when "01000101110011001", -- t[35737] = 4
      "0000100" when "01000101110011010", -- t[35738] = 4
      "0000100" when "01000101110011011", -- t[35739] = 4
      "0000100" when "01000101110011100", -- t[35740] = 4
      "0000100" when "01000101110011101", -- t[35741] = 4
      "0000100" when "01000101110011110", -- t[35742] = 4
      "0000100" when "01000101110011111", -- t[35743] = 4
      "0000100" when "01000101110100000", -- t[35744] = 4
      "0000100" when "01000101110100001", -- t[35745] = 4
      "0000100" when "01000101110100010", -- t[35746] = 4
      "0000100" when "01000101110100011", -- t[35747] = 4
      "0000100" when "01000101110100100", -- t[35748] = 4
      "0000100" when "01000101110100101", -- t[35749] = 4
      "0000100" when "01000101110100110", -- t[35750] = 4
      "0000100" when "01000101110100111", -- t[35751] = 4
      "0000100" when "01000101110101000", -- t[35752] = 4
      "0000100" when "01000101110101001", -- t[35753] = 4
      "0000100" when "01000101110101010", -- t[35754] = 4
      "0000100" when "01000101110101011", -- t[35755] = 4
      "0000100" when "01000101110101100", -- t[35756] = 4
      "0000100" when "01000101110101101", -- t[35757] = 4
      "0000100" when "01000101110101110", -- t[35758] = 4
      "0000100" when "01000101110101111", -- t[35759] = 4
      "0000100" when "01000101110110000", -- t[35760] = 4
      "0000100" when "01000101110110001", -- t[35761] = 4
      "0000100" when "01000101110110010", -- t[35762] = 4
      "0000100" when "01000101110110011", -- t[35763] = 4
      "0000100" when "01000101110110100", -- t[35764] = 4
      "0000100" when "01000101110110101", -- t[35765] = 4
      "0000100" when "01000101110110110", -- t[35766] = 4
      "0000100" when "01000101110110111", -- t[35767] = 4
      "0000100" when "01000101110111000", -- t[35768] = 4
      "0000100" when "01000101110111001", -- t[35769] = 4
      "0000100" when "01000101110111010", -- t[35770] = 4
      "0000100" when "01000101110111011", -- t[35771] = 4
      "0000100" when "01000101110111100", -- t[35772] = 4
      "0000100" when "01000101110111101", -- t[35773] = 4
      "0000100" when "01000101110111110", -- t[35774] = 4
      "0000100" when "01000101110111111", -- t[35775] = 4
      "0000100" when "01000101111000000", -- t[35776] = 4
      "0000100" when "01000101111000001", -- t[35777] = 4
      "0000100" when "01000101111000010", -- t[35778] = 4
      "0000100" when "01000101111000011", -- t[35779] = 4
      "0000100" when "01000101111000100", -- t[35780] = 4
      "0000100" when "01000101111000101", -- t[35781] = 4
      "0000100" when "01000101111000110", -- t[35782] = 4
      "0000100" when "01000101111000111", -- t[35783] = 4
      "0000100" when "01000101111001000", -- t[35784] = 4
      "0000100" when "01000101111001001", -- t[35785] = 4
      "0000100" when "01000101111001010", -- t[35786] = 4
      "0000100" when "01000101111001011", -- t[35787] = 4
      "0000100" when "01000101111001100", -- t[35788] = 4
      "0000100" when "01000101111001101", -- t[35789] = 4
      "0000100" when "01000101111001110", -- t[35790] = 4
      "0000100" when "01000101111001111", -- t[35791] = 4
      "0000100" when "01000101111010000", -- t[35792] = 4
      "0000100" when "01000101111010001", -- t[35793] = 4
      "0000100" when "01000101111010010", -- t[35794] = 4
      "0000100" when "01000101111010011", -- t[35795] = 4
      "0000100" when "01000101111010100", -- t[35796] = 4
      "0000100" when "01000101111010101", -- t[35797] = 4
      "0000100" when "01000101111010110", -- t[35798] = 4
      "0000100" when "01000101111010111", -- t[35799] = 4
      "0000100" when "01000101111011000", -- t[35800] = 4
      "0000100" when "01000101111011001", -- t[35801] = 4
      "0000100" when "01000101111011010", -- t[35802] = 4
      "0000100" when "01000101111011011", -- t[35803] = 4
      "0000100" when "01000101111011100", -- t[35804] = 4
      "0000100" when "01000101111011101", -- t[35805] = 4
      "0000100" when "01000101111011110", -- t[35806] = 4
      "0000100" when "01000101111011111", -- t[35807] = 4
      "0000100" when "01000101111100000", -- t[35808] = 4
      "0000100" when "01000101111100001", -- t[35809] = 4
      "0000100" when "01000101111100010", -- t[35810] = 4
      "0000100" when "01000101111100011", -- t[35811] = 4
      "0000100" when "01000101111100100", -- t[35812] = 4
      "0000100" when "01000101111100101", -- t[35813] = 4
      "0000100" when "01000101111100110", -- t[35814] = 4
      "0000100" when "01000101111100111", -- t[35815] = 4
      "0000100" when "01000101111101000", -- t[35816] = 4
      "0000100" when "01000101111101001", -- t[35817] = 4
      "0000100" when "01000101111101010", -- t[35818] = 4
      "0000100" when "01000101111101011", -- t[35819] = 4
      "0000100" when "01000101111101100", -- t[35820] = 4
      "0000100" when "01000101111101101", -- t[35821] = 4
      "0000100" when "01000101111101110", -- t[35822] = 4
      "0000100" when "01000101111101111", -- t[35823] = 4
      "0000100" when "01000101111110000", -- t[35824] = 4
      "0000100" when "01000101111110001", -- t[35825] = 4
      "0000100" when "01000101111110010", -- t[35826] = 4
      "0000100" when "01000101111110011", -- t[35827] = 4
      "0000100" when "01000101111110100", -- t[35828] = 4
      "0000100" when "01000101111110101", -- t[35829] = 4
      "0000100" when "01000101111110110", -- t[35830] = 4
      "0000100" when "01000101111110111", -- t[35831] = 4
      "0000100" when "01000101111111000", -- t[35832] = 4
      "0000100" when "01000101111111001", -- t[35833] = 4
      "0000100" when "01000101111111010", -- t[35834] = 4
      "0000100" when "01000101111111011", -- t[35835] = 4
      "0000100" when "01000101111111100", -- t[35836] = 4
      "0000100" when "01000101111111101", -- t[35837] = 4
      "0000100" when "01000101111111110", -- t[35838] = 4
      "0000100" when "01000101111111111", -- t[35839] = 4
      "0000100" when "01000110000000000", -- t[35840] = 4
      "0000100" when "01000110000000001", -- t[35841] = 4
      "0000100" when "01000110000000010", -- t[35842] = 4
      "0000100" when "01000110000000011", -- t[35843] = 4
      "0000100" when "01000110000000100", -- t[35844] = 4
      "0000100" when "01000110000000101", -- t[35845] = 4
      "0000100" when "01000110000000110", -- t[35846] = 4
      "0000100" when "01000110000000111", -- t[35847] = 4
      "0000100" when "01000110000001000", -- t[35848] = 4
      "0000100" when "01000110000001001", -- t[35849] = 4
      "0000100" when "01000110000001010", -- t[35850] = 4
      "0000100" when "01000110000001011", -- t[35851] = 4
      "0000100" when "01000110000001100", -- t[35852] = 4
      "0000100" when "01000110000001101", -- t[35853] = 4
      "0000100" when "01000110000001110", -- t[35854] = 4
      "0000100" when "01000110000001111", -- t[35855] = 4
      "0000100" when "01000110000010000", -- t[35856] = 4
      "0000100" when "01000110000010001", -- t[35857] = 4
      "0000100" when "01000110000010010", -- t[35858] = 4
      "0000100" when "01000110000010011", -- t[35859] = 4
      "0000100" when "01000110000010100", -- t[35860] = 4
      "0000100" when "01000110000010101", -- t[35861] = 4
      "0000100" when "01000110000010110", -- t[35862] = 4
      "0000100" when "01000110000010111", -- t[35863] = 4
      "0000100" when "01000110000011000", -- t[35864] = 4
      "0000100" when "01000110000011001", -- t[35865] = 4
      "0000100" when "01000110000011010", -- t[35866] = 4
      "0000100" when "01000110000011011", -- t[35867] = 4
      "0000100" when "01000110000011100", -- t[35868] = 4
      "0000100" when "01000110000011101", -- t[35869] = 4
      "0000100" when "01000110000011110", -- t[35870] = 4
      "0000100" when "01000110000011111", -- t[35871] = 4
      "0000100" when "01000110000100000", -- t[35872] = 4
      "0000100" when "01000110000100001", -- t[35873] = 4
      "0000100" when "01000110000100010", -- t[35874] = 4
      "0000100" when "01000110000100011", -- t[35875] = 4
      "0000100" when "01000110000100100", -- t[35876] = 4
      "0000100" when "01000110000100101", -- t[35877] = 4
      "0000100" when "01000110000100110", -- t[35878] = 4
      "0000100" when "01000110000100111", -- t[35879] = 4
      "0000100" when "01000110000101000", -- t[35880] = 4
      "0000100" when "01000110000101001", -- t[35881] = 4
      "0000100" when "01000110000101010", -- t[35882] = 4
      "0000100" when "01000110000101011", -- t[35883] = 4
      "0000100" when "01000110000101100", -- t[35884] = 4
      "0000100" when "01000110000101101", -- t[35885] = 4
      "0000100" when "01000110000101110", -- t[35886] = 4
      "0000100" when "01000110000101111", -- t[35887] = 4
      "0000100" when "01000110000110000", -- t[35888] = 4
      "0000100" when "01000110000110001", -- t[35889] = 4
      "0000100" when "01000110000110010", -- t[35890] = 4
      "0000100" when "01000110000110011", -- t[35891] = 4
      "0000100" when "01000110000110100", -- t[35892] = 4
      "0000100" when "01000110000110101", -- t[35893] = 4
      "0000100" when "01000110000110110", -- t[35894] = 4
      "0000100" when "01000110000110111", -- t[35895] = 4
      "0000100" when "01000110000111000", -- t[35896] = 4
      "0000100" when "01000110000111001", -- t[35897] = 4
      "0000100" when "01000110000111010", -- t[35898] = 4
      "0000100" when "01000110000111011", -- t[35899] = 4
      "0000100" when "01000110000111100", -- t[35900] = 4
      "0000100" when "01000110000111101", -- t[35901] = 4
      "0000100" when "01000110000111110", -- t[35902] = 4
      "0000100" when "01000110000111111", -- t[35903] = 4
      "0000100" when "01000110001000000", -- t[35904] = 4
      "0000100" when "01000110001000001", -- t[35905] = 4
      "0000100" when "01000110001000010", -- t[35906] = 4
      "0000100" when "01000110001000011", -- t[35907] = 4
      "0000100" when "01000110001000100", -- t[35908] = 4
      "0000100" when "01000110001000101", -- t[35909] = 4
      "0000100" when "01000110001000110", -- t[35910] = 4
      "0000100" when "01000110001000111", -- t[35911] = 4
      "0000100" when "01000110001001000", -- t[35912] = 4
      "0000100" when "01000110001001001", -- t[35913] = 4
      "0000100" when "01000110001001010", -- t[35914] = 4
      "0000100" when "01000110001001011", -- t[35915] = 4
      "0000100" when "01000110001001100", -- t[35916] = 4
      "0000100" when "01000110001001101", -- t[35917] = 4
      "0000100" when "01000110001001110", -- t[35918] = 4
      "0000100" when "01000110001001111", -- t[35919] = 4
      "0000100" when "01000110001010000", -- t[35920] = 4
      "0000100" when "01000110001010001", -- t[35921] = 4
      "0000100" when "01000110001010010", -- t[35922] = 4
      "0000100" when "01000110001010011", -- t[35923] = 4
      "0000100" when "01000110001010100", -- t[35924] = 4
      "0000100" when "01000110001010101", -- t[35925] = 4
      "0000100" when "01000110001010110", -- t[35926] = 4
      "0000100" when "01000110001010111", -- t[35927] = 4
      "0000100" when "01000110001011000", -- t[35928] = 4
      "0000100" when "01000110001011001", -- t[35929] = 4
      "0000100" when "01000110001011010", -- t[35930] = 4
      "0000100" when "01000110001011011", -- t[35931] = 4
      "0000100" when "01000110001011100", -- t[35932] = 4
      "0000100" when "01000110001011101", -- t[35933] = 4
      "0000100" when "01000110001011110", -- t[35934] = 4
      "0000100" when "01000110001011111", -- t[35935] = 4
      "0000100" when "01000110001100000", -- t[35936] = 4
      "0000100" when "01000110001100001", -- t[35937] = 4
      "0000100" when "01000110001100010", -- t[35938] = 4
      "0000100" when "01000110001100011", -- t[35939] = 4
      "0000100" when "01000110001100100", -- t[35940] = 4
      "0000100" when "01000110001100101", -- t[35941] = 4
      "0000100" when "01000110001100110", -- t[35942] = 4
      "0000100" when "01000110001100111", -- t[35943] = 4
      "0000100" when "01000110001101000", -- t[35944] = 4
      "0000100" when "01000110001101001", -- t[35945] = 4
      "0000100" when "01000110001101010", -- t[35946] = 4
      "0000100" when "01000110001101011", -- t[35947] = 4
      "0000100" when "01000110001101100", -- t[35948] = 4
      "0000100" when "01000110001101101", -- t[35949] = 4
      "0000100" when "01000110001101110", -- t[35950] = 4
      "0000100" when "01000110001101111", -- t[35951] = 4
      "0000100" when "01000110001110000", -- t[35952] = 4
      "0000100" when "01000110001110001", -- t[35953] = 4
      "0000100" when "01000110001110010", -- t[35954] = 4
      "0000100" when "01000110001110011", -- t[35955] = 4
      "0000100" when "01000110001110100", -- t[35956] = 4
      "0000100" when "01000110001110101", -- t[35957] = 4
      "0000100" when "01000110001110110", -- t[35958] = 4
      "0000100" when "01000110001110111", -- t[35959] = 4
      "0000100" when "01000110001111000", -- t[35960] = 4
      "0000100" when "01000110001111001", -- t[35961] = 4
      "0000100" when "01000110001111010", -- t[35962] = 4
      "0000100" when "01000110001111011", -- t[35963] = 4
      "0000100" when "01000110001111100", -- t[35964] = 4
      "0000100" when "01000110001111101", -- t[35965] = 4
      "0000100" when "01000110001111110", -- t[35966] = 4
      "0000100" when "01000110001111111", -- t[35967] = 4
      "0000100" when "01000110010000000", -- t[35968] = 4
      "0000100" when "01000110010000001", -- t[35969] = 4
      "0000100" when "01000110010000010", -- t[35970] = 4
      "0000100" when "01000110010000011", -- t[35971] = 4
      "0000100" when "01000110010000100", -- t[35972] = 4
      "0000100" when "01000110010000101", -- t[35973] = 4
      "0000100" when "01000110010000110", -- t[35974] = 4
      "0000100" when "01000110010000111", -- t[35975] = 4
      "0000100" when "01000110010001000", -- t[35976] = 4
      "0000100" when "01000110010001001", -- t[35977] = 4
      "0000100" when "01000110010001010", -- t[35978] = 4
      "0000100" when "01000110010001011", -- t[35979] = 4
      "0000100" when "01000110010001100", -- t[35980] = 4
      "0000100" when "01000110010001101", -- t[35981] = 4
      "0000100" when "01000110010001110", -- t[35982] = 4
      "0000100" when "01000110010001111", -- t[35983] = 4
      "0000100" when "01000110010010000", -- t[35984] = 4
      "0000100" when "01000110010010001", -- t[35985] = 4
      "0000100" when "01000110010010010", -- t[35986] = 4
      "0000100" when "01000110010010011", -- t[35987] = 4
      "0000100" when "01000110010010100", -- t[35988] = 4
      "0000100" when "01000110010010101", -- t[35989] = 4
      "0000100" when "01000110010010110", -- t[35990] = 4
      "0000100" when "01000110010010111", -- t[35991] = 4
      "0000100" when "01000110010011000", -- t[35992] = 4
      "0000100" when "01000110010011001", -- t[35993] = 4
      "0000100" when "01000110010011010", -- t[35994] = 4
      "0000100" when "01000110010011011", -- t[35995] = 4
      "0000100" when "01000110010011100", -- t[35996] = 4
      "0000100" when "01000110010011101", -- t[35997] = 4
      "0000100" when "01000110010011110", -- t[35998] = 4
      "0000100" when "01000110010011111", -- t[35999] = 4
      "0000100" when "01000110010100000", -- t[36000] = 4
      "0000100" when "01000110010100001", -- t[36001] = 4
      "0000100" when "01000110010100010", -- t[36002] = 4
      "0000100" when "01000110010100011", -- t[36003] = 4
      "0000100" when "01000110010100100", -- t[36004] = 4
      "0000100" when "01000110010100101", -- t[36005] = 4
      "0000100" when "01000110010100110", -- t[36006] = 4
      "0000100" when "01000110010100111", -- t[36007] = 4
      "0000100" when "01000110010101000", -- t[36008] = 4
      "0000100" when "01000110010101001", -- t[36009] = 4
      "0000100" when "01000110010101010", -- t[36010] = 4
      "0000100" when "01000110010101011", -- t[36011] = 4
      "0000100" when "01000110010101100", -- t[36012] = 4
      "0000100" when "01000110010101101", -- t[36013] = 4
      "0000100" when "01000110010101110", -- t[36014] = 4
      "0000100" when "01000110010101111", -- t[36015] = 4
      "0000100" when "01000110010110000", -- t[36016] = 4
      "0000100" when "01000110010110001", -- t[36017] = 4
      "0000100" when "01000110010110010", -- t[36018] = 4
      "0000100" when "01000110010110011", -- t[36019] = 4
      "0000100" when "01000110010110100", -- t[36020] = 4
      "0000100" when "01000110010110101", -- t[36021] = 4
      "0000100" when "01000110010110110", -- t[36022] = 4
      "0000100" when "01000110010110111", -- t[36023] = 4
      "0000100" when "01000110010111000", -- t[36024] = 4
      "0000100" when "01000110010111001", -- t[36025] = 4
      "0000100" when "01000110010111010", -- t[36026] = 4
      "0000100" when "01000110010111011", -- t[36027] = 4
      "0000100" when "01000110010111100", -- t[36028] = 4
      "0000100" when "01000110010111101", -- t[36029] = 4
      "0000100" when "01000110010111110", -- t[36030] = 4
      "0000100" when "01000110010111111", -- t[36031] = 4
      "0000100" when "01000110011000000", -- t[36032] = 4
      "0000100" when "01000110011000001", -- t[36033] = 4
      "0000100" when "01000110011000010", -- t[36034] = 4
      "0000100" when "01000110011000011", -- t[36035] = 4
      "0000100" when "01000110011000100", -- t[36036] = 4
      "0000100" when "01000110011000101", -- t[36037] = 4
      "0000100" when "01000110011000110", -- t[36038] = 4
      "0000100" when "01000110011000111", -- t[36039] = 4
      "0000100" when "01000110011001000", -- t[36040] = 4
      "0000100" when "01000110011001001", -- t[36041] = 4
      "0000100" when "01000110011001010", -- t[36042] = 4
      "0000100" when "01000110011001011", -- t[36043] = 4
      "0000100" when "01000110011001100", -- t[36044] = 4
      "0000100" when "01000110011001101", -- t[36045] = 4
      "0000100" when "01000110011001110", -- t[36046] = 4
      "0000100" when "01000110011001111", -- t[36047] = 4
      "0000100" when "01000110011010000", -- t[36048] = 4
      "0000100" when "01000110011010001", -- t[36049] = 4
      "0000100" when "01000110011010010", -- t[36050] = 4
      "0000100" when "01000110011010011", -- t[36051] = 4
      "0000100" when "01000110011010100", -- t[36052] = 4
      "0000100" when "01000110011010101", -- t[36053] = 4
      "0000100" when "01000110011010110", -- t[36054] = 4
      "0000100" when "01000110011010111", -- t[36055] = 4
      "0000100" when "01000110011011000", -- t[36056] = 4
      "0000100" when "01000110011011001", -- t[36057] = 4
      "0000100" when "01000110011011010", -- t[36058] = 4
      "0000100" when "01000110011011011", -- t[36059] = 4
      "0000100" when "01000110011011100", -- t[36060] = 4
      "0000100" when "01000110011011101", -- t[36061] = 4
      "0000100" when "01000110011011110", -- t[36062] = 4
      "0000100" when "01000110011011111", -- t[36063] = 4
      "0000100" when "01000110011100000", -- t[36064] = 4
      "0000100" when "01000110011100001", -- t[36065] = 4
      "0000100" when "01000110011100010", -- t[36066] = 4
      "0000100" when "01000110011100011", -- t[36067] = 4
      "0000100" when "01000110011100100", -- t[36068] = 4
      "0000100" when "01000110011100101", -- t[36069] = 4
      "0000100" when "01000110011100110", -- t[36070] = 4
      "0000100" when "01000110011100111", -- t[36071] = 4
      "0000100" when "01000110011101000", -- t[36072] = 4
      "0000100" when "01000110011101001", -- t[36073] = 4
      "0000100" when "01000110011101010", -- t[36074] = 4
      "0000100" when "01000110011101011", -- t[36075] = 4
      "0000100" when "01000110011101100", -- t[36076] = 4
      "0000100" when "01000110011101101", -- t[36077] = 4
      "0000100" when "01000110011101110", -- t[36078] = 4
      "0000100" when "01000110011101111", -- t[36079] = 4
      "0000100" when "01000110011110000", -- t[36080] = 4
      "0000100" when "01000110011110001", -- t[36081] = 4
      "0000100" when "01000110011110010", -- t[36082] = 4
      "0000100" when "01000110011110011", -- t[36083] = 4
      "0000100" when "01000110011110100", -- t[36084] = 4
      "0000100" when "01000110011110101", -- t[36085] = 4
      "0000100" when "01000110011110110", -- t[36086] = 4
      "0000100" when "01000110011110111", -- t[36087] = 4
      "0000100" when "01000110011111000", -- t[36088] = 4
      "0000100" when "01000110011111001", -- t[36089] = 4
      "0000100" when "01000110011111010", -- t[36090] = 4
      "0000100" when "01000110011111011", -- t[36091] = 4
      "0000100" when "01000110011111100", -- t[36092] = 4
      "0000100" when "01000110011111101", -- t[36093] = 4
      "0000100" when "01000110011111110", -- t[36094] = 4
      "0000100" when "01000110011111111", -- t[36095] = 4
      "0000100" when "01000110100000000", -- t[36096] = 4
      "0000100" when "01000110100000001", -- t[36097] = 4
      "0000100" when "01000110100000010", -- t[36098] = 4
      "0000100" when "01000110100000011", -- t[36099] = 4
      "0000100" when "01000110100000100", -- t[36100] = 4
      "0000100" when "01000110100000101", -- t[36101] = 4
      "0000100" when "01000110100000110", -- t[36102] = 4
      "0000100" when "01000110100000111", -- t[36103] = 4
      "0000100" when "01000110100001000", -- t[36104] = 4
      "0000100" when "01000110100001001", -- t[36105] = 4
      "0000100" when "01000110100001010", -- t[36106] = 4
      "0000100" when "01000110100001011", -- t[36107] = 4
      "0000100" when "01000110100001100", -- t[36108] = 4
      "0000100" when "01000110100001101", -- t[36109] = 4
      "0000100" when "01000110100001110", -- t[36110] = 4
      "0000100" when "01000110100001111", -- t[36111] = 4
      "0000100" when "01000110100010000", -- t[36112] = 4
      "0000100" when "01000110100010001", -- t[36113] = 4
      "0000100" when "01000110100010010", -- t[36114] = 4
      "0000100" when "01000110100010011", -- t[36115] = 4
      "0000100" when "01000110100010100", -- t[36116] = 4
      "0000100" when "01000110100010101", -- t[36117] = 4
      "0000100" when "01000110100010110", -- t[36118] = 4
      "0000100" when "01000110100010111", -- t[36119] = 4
      "0000100" when "01000110100011000", -- t[36120] = 4
      "0000100" when "01000110100011001", -- t[36121] = 4
      "0000100" when "01000110100011010", -- t[36122] = 4
      "0000100" when "01000110100011011", -- t[36123] = 4
      "0000100" when "01000110100011100", -- t[36124] = 4
      "0000100" when "01000110100011101", -- t[36125] = 4
      "0000100" when "01000110100011110", -- t[36126] = 4
      "0000100" when "01000110100011111", -- t[36127] = 4
      "0000100" when "01000110100100000", -- t[36128] = 4
      "0000100" when "01000110100100001", -- t[36129] = 4
      "0000100" when "01000110100100010", -- t[36130] = 4
      "0000100" when "01000110100100011", -- t[36131] = 4
      "0000100" when "01000110100100100", -- t[36132] = 4
      "0000100" when "01000110100100101", -- t[36133] = 4
      "0000100" when "01000110100100110", -- t[36134] = 4
      "0000100" when "01000110100100111", -- t[36135] = 4
      "0000100" when "01000110100101000", -- t[36136] = 4
      "0000100" when "01000110100101001", -- t[36137] = 4
      "0000100" when "01000110100101010", -- t[36138] = 4
      "0000100" when "01000110100101011", -- t[36139] = 4
      "0000100" when "01000110100101100", -- t[36140] = 4
      "0000100" when "01000110100101101", -- t[36141] = 4
      "0000100" when "01000110100101110", -- t[36142] = 4
      "0000100" when "01000110100101111", -- t[36143] = 4
      "0000100" when "01000110100110000", -- t[36144] = 4
      "0000100" when "01000110100110001", -- t[36145] = 4
      "0000100" when "01000110100110010", -- t[36146] = 4
      "0000100" when "01000110100110011", -- t[36147] = 4
      "0000100" when "01000110100110100", -- t[36148] = 4
      "0000100" when "01000110100110101", -- t[36149] = 4
      "0000100" when "01000110100110110", -- t[36150] = 4
      "0000100" when "01000110100110111", -- t[36151] = 4
      "0000100" when "01000110100111000", -- t[36152] = 4
      "0000100" when "01000110100111001", -- t[36153] = 4
      "0000100" when "01000110100111010", -- t[36154] = 4
      "0000100" when "01000110100111011", -- t[36155] = 4
      "0000100" when "01000110100111100", -- t[36156] = 4
      "0000100" when "01000110100111101", -- t[36157] = 4
      "0000100" when "01000110100111110", -- t[36158] = 4
      "0000100" when "01000110100111111", -- t[36159] = 4
      "0000100" when "01000110101000000", -- t[36160] = 4
      "0000100" when "01000110101000001", -- t[36161] = 4
      "0000100" when "01000110101000010", -- t[36162] = 4
      "0000100" when "01000110101000011", -- t[36163] = 4
      "0000100" when "01000110101000100", -- t[36164] = 4
      "0000100" when "01000110101000101", -- t[36165] = 4
      "0000100" when "01000110101000110", -- t[36166] = 4
      "0000100" when "01000110101000111", -- t[36167] = 4
      "0000100" when "01000110101001000", -- t[36168] = 4
      "0000100" when "01000110101001001", -- t[36169] = 4
      "0000100" when "01000110101001010", -- t[36170] = 4
      "0000100" when "01000110101001011", -- t[36171] = 4
      "0000100" when "01000110101001100", -- t[36172] = 4
      "0000100" when "01000110101001101", -- t[36173] = 4
      "0000100" when "01000110101001110", -- t[36174] = 4
      "0000100" when "01000110101001111", -- t[36175] = 4
      "0000100" when "01000110101010000", -- t[36176] = 4
      "0000100" when "01000110101010001", -- t[36177] = 4
      "0000100" when "01000110101010010", -- t[36178] = 4
      "0000100" when "01000110101010011", -- t[36179] = 4
      "0000100" when "01000110101010100", -- t[36180] = 4
      "0000100" when "01000110101010101", -- t[36181] = 4
      "0000100" when "01000110101010110", -- t[36182] = 4
      "0000100" when "01000110101010111", -- t[36183] = 4
      "0000100" when "01000110101011000", -- t[36184] = 4
      "0000100" when "01000110101011001", -- t[36185] = 4
      "0000100" when "01000110101011010", -- t[36186] = 4
      "0000100" when "01000110101011011", -- t[36187] = 4
      "0000100" when "01000110101011100", -- t[36188] = 4
      "0000100" when "01000110101011101", -- t[36189] = 4
      "0000100" when "01000110101011110", -- t[36190] = 4
      "0000100" when "01000110101011111", -- t[36191] = 4
      "0000100" when "01000110101100000", -- t[36192] = 4
      "0000100" when "01000110101100001", -- t[36193] = 4
      "0000100" when "01000110101100010", -- t[36194] = 4
      "0000100" when "01000110101100011", -- t[36195] = 4
      "0000100" when "01000110101100100", -- t[36196] = 4
      "0000100" when "01000110101100101", -- t[36197] = 4
      "0000100" when "01000110101100110", -- t[36198] = 4
      "0000100" when "01000110101100111", -- t[36199] = 4
      "0000100" when "01000110101101000", -- t[36200] = 4
      "0000100" when "01000110101101001", -- t[36201] = 4
      "0000100" when "01000110101101010", -- t[36202] = 4
      "0000100" when "01000110101101011", -- t[36203] = 4
      "0000100" when "01000110101101100", -- t[36204] = 4
      "0000100" when "01000110101101101", -- t[36205] = 4
      "0000100" when "01000110101101110", -- t[36206] = 4
      "0000100" when "01000110101101111", -- t[36207] = 4
      "0000100" when "01000110101110000", -- t[36208] = 4
      "0000100" when "01000110101110001", -- t[36209] = 4
      "0000100" when "01000110101110010", -- t[36210] = 4
      "0000100" when "01000110101110011", -- t[36211] = 4
      "0000100" when "01000110101110100", -- t[36212] = 4
      "0000100" when "01000110101110101", -- t[36213] = 4
      "0000100" when "01000110101110110", -- t[36214] = 4
      "0000100" when "01000110101110111", -- t[36215] = 4
      "0000100" when "01000110101111000", -- t[36216] = 4
      "0000100" when "01000110101111001", -- t[36217] = 4
      "0000100" when "01000110101111010", -- t[36218] = 4
      "0000100" when "01000110101111011", -- t[36219] = 4
      "0000100" when "01000110101111100", -- t[36220] = 4
      "0000100" when "01000110101111101", -- t[36221] = 4
      "0000100" when "01000110101111110", -- t[36222] = 4
      "0000100" when "01000110101111111", -- t[36223] = 4
      "0000100" when "01000110110000000", -- t[36224] = 4
      "0000100" when "01000110110000001", -- t[36225] = 4
      "0000100" when "01000110110000010", -- t[36226] = 4
      "0000100" when "01000110110000011", -- t[36227] = 4
      "0000100" when "01000110110000100", -- t[36228] = 4
      "0000100" when "01000110110000101", -- t[36229] = 4
      "0000100" when "01000110110000110", -- t[36230] = 4
      "0000100" when "01000110110000111", -- t[36231] = 4
      "0000100" when "01000110110001000", -- t[36232] = 4
      "0000100" when "01000110110001001", -- t[36233] = 4
      "0000100" when "01000110110001010", -- t[36234] = 4
      "0000100" when "01000110110001011", -- t[36235] = 4
      "0000100" when "01000110110001100", -- t[36236] = 4
      "0000100" when "01000110110001101", -- t[36237] = 4
      "0000100" when "01000110110001110", -- t[36238] = 4
      "0000100" when "01000110110001111", -- t[36239] = 4
      "0000100" when "01000110110010000", -- t[36240] = 4
      "0000100" when "01000110110010001", -- t[36241] = 4
      "0000100" when "01000110110010010", -- t[36242] = 4
      "0000100" when "01000110110010011", -- t[36243] = 4
      "0000100" when "01000110110010100", -- t[36244] = 4
      "0000100" when "01000110110010101", -- t[36245] = 4
      "0000100" when "01000110110010110", -- t[36246] = 4
      "0000100" when "01000110110010111", -- t[36247] = 4
      "0000100" when "01000110110011000", -- t[36248] = 4
      "0000100" when "01000110110011001", -- t[36249] = 4
      "0000100" when "01000110110011010", -- t[36250] = 4
      "0000100" when "01000110110011011", -- t[36251] = 4
      "0000100" when "01000110110011100", -- t[36252] = 4
      "0000100" when "01000110110011101", -- t[36253] = 4
      "0000100" when "01000110110011110", -- t[36254] = 4
      "0000100" when "01000110110011111", -- t[36255] = 4
      "0000100" when "01000110110100000", -- t[36256] = 4
      "0000100" when "01000110110100001", -- t[36257] = 4
      "0000100" when "01000110110100010", -- t[36258] = 4
      "0000100" when "01000110110100011", -- t[36259] = 4
      "0000100" when "01000110110100100", -- t[36260] = 4
      "0000100" when "01000110110100101", -- t[36261] = 4
      "0000100" when "01000110110100110", -- t[36262] = 4
      "0000100" when "01000110110100111", -- t[36263] = 4
      "0000100" when "01000110110101000", -- t[36264] = 4
      "0000100" when "01000110110101001", -- t[36265] = 4
      "0000100" when "01000110110101010", -- t[36266] = 4
      "0000100" when "01000110110101011", -- t[36267] = 4
      "0000100" when "01000110110101100", -- t[36268] = 4
      "0000100" when "01000110110101101", -- t[36269] = 4
      "0000100" when "01000110110101110", -- t[36270] = 4
      "0000100" when "01000110110101111", -- t[36271] = 4
      "0000100" when "01000110110110000", -- t[36272] = 4
      "0000100" when "01000110110110001", -- t[36273] = 4
      "0000100" when "01000110110110010", -- t[36274] = 4
      "0000100" when "01000110110110011", -- t[36275] = 4
      "0000100" when "01000110110110100", -- t[36276] = 4
      "0000100" when "01000110110110101", -- t[36277] = 4
      "0000100" when "01000110110110110", -- t[36278] = 4
      "0000100" when "01000110110110111", -- t[36279] = 4
      "0000100" when "01000110110111000", -- t[36280] = 4
      "0000100" when "01000110110111001", -- t[36281] = 4
      "0000100" when "01000110110111010", -- t[36282] = 4
      "0000100" when "01000110110111011", -- t[36283] = 4
      "0000100" when "01000110110111100", -- t[36284] = 4
      "0000100" when "01000110110111101", -- t[36285] = 4
      "0000100" when "01000110110111110", -- t[36286] = 4
      "0000100" when "01000110110111111", -- t[36287] = 4
      "0000100" when "01000110111000000", -- t[36288] = 4
      "0000100" when "01000110111000001", -- t[36289] = 4
      "0000100" when "01000110111000010", -- t[36290] = 4
      "0000100" when "01000110111000011", -- t[36291] = 4
      "0000100" when "01000110111000100", -- t[36292] = 4
      "0000100" when "01000110111000101", -- t[36293] = 4
      "0000100" when "01000110111000110", -- t[36294] = 4
      "0000100" when "01000110111000111", -- t[36295] = 4
      "0000100" when "01000110111001000", -- t[36296] = 4
      "0000100" when "01000110111001001", -- t[36297] = 4
      "0000100" when "01000110111001010", -- t[36298] = 4
      "0000100" when "01000110111001011", -- t[36299] = 4
      "0000100" when "01000110111001100", -- t[36300] = 4
      "0000100" when "01000110111001101", -- t[36301] = 4
      "0000100" when "01000110111001110", -- t[36302] = 4
      "0000100" when "01000110111001111", -- t[36303] = 4
      "0000100" when "01000110111010000", -- t[36304] = 4
      "0000100" when "01000110111010001", -- t[36305] = 4
      "0000100" when "01000110111010010", -- t[36306] = 4
      "0000100" when "01000110111010011", -- t[36307] = 4
      "0000100" when "01000110111010100", -- t[36308] = 4
      "0000100" when "01000110111010101", -- t[36309] = 4
      "0000100" when "01000110111010110", -- t[36310] = 4
      "0000100" when "01000110111010111", -- t[36311] = 4
      "0000100" when "01000110111011000", -- t[36312] = 4
      "0000100" when "01000110111011001", -- t[36313] = 4
      "0000100" when "01000110111011010", -- t[36314] = 4
      "0000100" when "01000110111011011", -- t[36315] = 4
      "0000100" when "01000110111011100", -- t[36316] = 4
      "0000100" when "01000110111011101", -- t[36317] = 4
      "0000100" when "01000110111011110", -- t[36318] = 4
      "0000100" when "01000110111011111", -- t[36319] = 4
      "0000100" when "01000110111100000", -- t[36320] = 4
      "0000100" when "01000110111100001", -- t[36321] = 4
      "0000100" when "01000110111100010", -- t[36322] = 4
      "0000100" when "01000110111100011", -- t[36323] = 4
      "0000100" when "01000110111100100", -- t[36324] = 4
      "0000100" when "01000110111100101", -- t[36325] = 4
      "0000100" when "01000110111100110", -- t[36326] = 4
      "0000100" when "01000110111100111", -- t[36327] = 4
      "0000100" when "01000110111101000", -- t[36328] = 4
      "0000100" when "01000110111101001", -- t[36329] = 4
      "0000100" when "01000110111101010", -- t[36330] = 4
      "0000100" when "01000110111101011", -- t[36331] = 4
      "0000100" when "01000110111101100", -- t[36332] = 4
      "0000100" when "01000110111101101", -- t[36333] = 4
      "0000100" when "01000110111101110", -- t[36334] = 4
      "0000100" when "01000110111101111", -- t[36335] = 4
      "0000100" when "01000110111110000", -- t[36336] = 4
      "0000100" when "01000110111110001", -- t[36337] = 4
      "0000100" when "01000110111110010", -- t[36338] = 4
      "0000100" when "01000110111110011", -- t[36339] = 4
      "0000100" when "01000110111110100", -- t[36340] = 4
      "0000100" when "01000110111110101", -- t[36341] = 4
      "0000100" when "01000110111110110", -- t[36342] = 4
      "0000100" when "01000110111110111", -- t[36343] = 4
      "0000100" when "01000110111111000", -- t[36344] = 4
      "0000100" when "01000110111111001", -- t[36345] = 4
      "0000100" when "01000110111111010", -- t[36346] = 4
      "0000100" when "01000110111111011", -- t[36347] = 4
      "0000100" when "01000110111111100", -- t[36348] = 4
      "0000100" when "01000110111111101", -- t[36349] = 4
      "0000100" when "01000110111111110", -- t[36350] = 4
      "0000100" when "01000110111111111", -- t[36351] = 4
      "0000100" when "01000111000000000", -- t[36352] = 4
      "0000100" when "01000111000000001", -- t[36353] = 4
      "0000100" when "01000111000000010", -- t[36354] = 4
      "0000100" when "01000111000000011", -- t[36355] = 4
      "0000100" when "01000111000000100", -- t[36356] = 4
      "0000100" when "01000111000000101", -- t[36357] = 4
      "0000100" when "01000111000000110", -- t[36358] = 4
      "0000100" when "01000111000000111", -- t[36359] = 4
      "0000100" when "01000111000001000", -- t[36360] = 4
      "0000100" when "01000111000001001", -- t[36361] = 4
      "0000100" when "01000111000001010", -- t[36362] = 4
      "0000100" when "01000111000001011", -- t[36363] = 4
      "0000100" when "01000111000001100", -- t[36364] = 4
      "0000100" when "01000111000001101", -- t[36365] = 4
      "0000100" when "01000111000001110", -- t[36366] = 4
      "0000100" when "01000111000001111", -- t[36367] = 4
      "0000100" when "01000111000010000", -- t[36368] = 4
      "0000100" when "01000111000010001", -- t[36369] = 4
      "0000100" when "01000111000010010", -- t[36370] = 4
      "0000100" when "01000111000010011", -- t[36371] = 4
      "0000100" when "01000111000010100", -- t[36372] = 4
      "0000100" when "01000111000010101", -- t[36373] = 4
      "0000100" when "01000111000010110", -- t[36374] = 4
      "0000100" when "01000111000010111", -- t[36375] = 4
      "0000100" when "01000111000011000", -- t[36376] = 4
      "0000100" when "01000111000011001", -- t[36377] = 4
      "0000100" when "01000111000011010", -- t[36378] = 4
      "0000100" when "01000111000011011", -- t[36379] = 4
      "0000100" when "01000111000011100", -- t[36380] = 4
      "0000100" when "01000111000011101", -- t[36381] = 4
      "0000100" when "01000111000011110", -- t[36382] = 4
      "0000100" when "01000111000011111", -- t[36383] = 4
      "0000100" when "01000111000100000", -- t[36384] = 4
      "0000100" when "01000111000100001", -- t[36385] = 4
      "0000100" when "01000111000100010", -- t[36386] = 4
      "0000100" when "01000111000100011", -- t[36387] = 4
      "0000100" when "01000111000100100", -- t[36388] = 4
      "0000100" when "01000111000100101", -- t[36389] = 4
      "0000100" when "01000111000100110", -- t[36390] = 4
      "0000100" when "01000111000100111", -- t[36391] = 4
      "0000100" when "01000111000101000", -- t[36392] = 4
      "0000100" when "01000111000101001", -- t[36393] = 4
      "0000100" when "01000111000101010", -- t[36394] = 4
      "0000100" when "01000111000101011", -- t[36395] = 4
      "0000100" when "01000111000101100", -- t[36396] = 4
      "0000100" when "01000111000101101", -- t[36397] = 4
      "0000100" when "01000111000101110", -- t[36398] = 4
      "0000100" when "01000111000101111", -- t[36399] = 4
      "0000100" when "01000111000110000", -- t[36400] = 4
      "0000100" when "01000111000110001", -- t[36401] = 4
      "0000100" when "01000111000110010", -- t[36402] = 4
      "0000100" when "01000111000110011", -- t[36403] = 4
      "0000100" when "01000111000110100", -- t[36404] = 4
      "0000100" when "01000111000110101", -- t[36405] = 4
      "0000100" when "01000111000110110", -- t[36406] = 4
      "0000100" when "01000111000110111", -- t[36407] = 4
      "0000100" when "01000111000111000", -- t[36408] = 4
      "0000100" when "01000111000111001", -- t[36409] = 4
      "0000100" when "01000111000111010", -- t[36410] = 4
      "0000100" when "01000111000111011", -- t[36411] = 4
      "0000100" when "01000111000111100", -- t[36412] = 4
      "0000100" when "01000111000111101", -- t[36413] = 4
      "0000100" when "01000111000111110", -- t[36414] = 4
      "0000100" when "01000111000111111", -- t[36415] = 4
      "0000100" when "01000111001000000", -- t[36416] = 4
      "0000100" when "01000111001000001", -- t[36417] = 4
      "0000100" when "01000111001000010", -- t[36418] = 4
      "0000100" when "01000111001000011", -- t[36419] = 4
      "0000100" when "01000111001000100", -- t[36420] = 4
      "0000100" when "01000111001000101", -- t[36421] = 4
      "0000100" when "01000111001000110", -- t[36422] = 4
      "0000100" when "01000111001000111", -- t[36423] = 4
      "0000100" when "01000111001001000", -- t[36424] = 4
      "0000100" when "01000111001001001", -- t[36425] = 4
      "0000100" when "01000111001001010", -- t[36426] = 4
      "0000100" when "01000111001001011", -- t[36427] = 4
      "0000100" when "01000111001001100", -- t[36428] = 4
      "0000100" when "01000111001001101", -- t[36429] = 4
      "0000100" when "01000111001001110", -- t[36430] = 4
      "0000100" when "01000111001001111", -- t[36431] = 4
      "0000100" when "01000111001010000", -- t[36432] = 4
      "0000100" when "01000111001010001", -- t[36433] = 4
      "0000100" when "01000111001010010", -- t[36434] = 4
      "0000100" when "01000111001010011", -- t[36435] = 4
      "0000100" when "01000111001010100", -- t[36436] = 4
      "0000100" when "01000111001010101", -- t[36437] = 4
      "0000100" when "01000111001010110", -- t[36438] = 4
      "0000100" when "01000111001010111", -- t[36439] = 4
      "0000100" when "01000111001011000", -- t[36440] = 4
      "0000100" when "01000111001011001", -- t[36441] = 4
      "0000100" when "01000111001011010", -- t[36442] = 4
      "0000100" when "01000111001011011", -- t[36443] = 4
      "0000100" when "01000111001011100", -- t[36444] = 4
      "0000100" when "01000111001011101", -- t[36445] = 4
      "0000100" when "01000111001011110", -- t[36446] = 4
      "0000100" when "01000111001011111", -- t[36447] = 4
      "0000100" when "01000111001100000", -- t[36448] = 4
      "0000100" when "01000111001100001", -- t[36449] = 4
      "0000100" when "01000111001100010", -- t[36450] = 4
      "0000100" when "01000111001100011", -- t[36451] = 4
      "0000100" when "01000111001100100", -- t[36452] = 4
      "0000100" when "01000111001100101", -- t[36453] = 4
      "0000100" when "01000111001100110", -- t[36454] = 4
      "0000100" when "01000111001100111", -- t[36455] = 4
      "0000100" when "01000111001101000", -- t[36456] = 4
      "0000100" when "01000111001101001", -- t[36457] = 4
      "0000100" when "01000111001101010", -- t[36458] = 4
      "0000100" when "01000111001101011", -- t[36459] = 4
      "0000100" when "01000111001101100", -- t[36460] = 4
      "0000100" when "01000111001101101", -- t[36461] = 4
      "0000100" when "01000111001101110", -- t[36462] = 4
      "0000100" when "01000111001101111", -- t[36463] = 4
      "0000100" when "01000111001110000", -- t[36464] = 4
      "0000100" when "01000111001110001", -- t[36465] = 4
      "0000100" when "01000111001110010", -- t[36466] = 4
      "0000100" when "01000111001110011", -- t[36467] = 4
      "0000100" when "01000111001110100", -- t[36468] = 4
      "0000100" when "01000111001110101", -- t[36469] = 4
      "0000100" when "01000111001110110", -- t[36470] = 4
      "0000100" when "01000111001110111", -- t[36471] = 4
      "0000100" when "01000111001111000", -- t[36472] = 4
      "0000100" when "01000111001111001", -- t[36473] = 4
      "0000100" when "01000111001111010", -- t[36474] = 4
      "0000100" when "01000111001111011", -- t[36475] = 4
      "0000100" when "01000111001111100", -- t[36476] = 4
      "0000100" when "01000111001111101", -- t[36477] = 4
      "0000100" when "01000111001111110", -- t[36478] = 4
      "0000100" when "01000111001111111", -- t[36479] = 4
      "0000100" when "01000111010000000", -- t[36480] = 4
      "0000100" when "01000111010000001", -- t[36481] = 4
      "0000100" when "01000111010000010", -- t[36482] = 4
      "0000100" when "01000111010000011", -- t[36483] = 4
      "0000100" when "01000111010000100", -- t[36484] = 4
      "0000100" when "01000111010000101", -- t[36485] = 4
      "0000100" when "01000111010000110", -- t[36486] = 4
      "0000100" when "01000111010000111", -- t[36487] = 4
      "0000100" when "01000111010001000", -- t[36488] = 4
      "0000100" when "01000111010001001", -- t[36489] = 4
      "0000100" when "01000111010001010", -- t[36490] = 4
      "0000100" when "01000111010001011", -- t[36491] = 4
      "0000100" when "01000111010001100", -- t[36492] = 4
      "0000100" when "01000111010001101", -- t[36493] = 4
      "0000100" when "01000111010001110", -- t[36494] = 4
      "0000100" when "01000111010001111", -- t[36495] = 4
      "0000100" when "01000111010010000", -- t[36496] = 4
      "0000100" when "01000111010010001", -- t[36497] = 4
      "0000100" when "01000111010010010", -- t[36498] = 4
      "0000100" when "01000111010010011", -- t[36499] = 4
      "0000100" when "01000111010010100", -- t[36500] = 4
      "0000100" when "01000111010010101", -- t[36501] = 4
      "0000100" when "01000111010010110", -- t[36502] = 4
      "0000100" when "01000111010010111", -- t[36503] = 4
      "0000100" when "01000111010011000", -- t[36504] = 4
      "0000100" when "01000111010011001", -- t[36505] = 4
      "0000100" when "01000111010011010", -- t[36506] = 4
      "0000100" when "01000111010011011", -- t[36507] = 4
      "0000100" when "01000111010011100", -- t[36508] = 4
      "0000100" when "01000111010011101", -- t[36509] = 4
      "0000100" when "01000111010011110", -- t[36510] = 4
      "0000100" when "01000111010011111", -- t[36511] = 4
      "0000100" when "01000111010100000", -- t[36512] = 4
      "0000100" when "01000111010100001", -- t[36513] = 4
      "0000100" when "01000111010100010", -- t[36514] = 4
      "0000100" when "01000111010100011", -- t[36515] = 4
      "0000100" when "01000111010100100", -- t[36516] = 4
      "0000100" when "01000111010100101", -- t[36517] = 4
      "0000100" when "01000111010100110", -- t[36518] = 4
      "0000100" when "01000111010100111", -- t[36519] = 4
      "0000100" when "01000111010101000", -- t[36520] = 4
      "0000100" when "01000111010101001", -- t[36521] = 4
      "0000100" when "01000111010101010", -- t[36522] = 4
      "0000100" when "01000111010101011", -- t[36523] = 4
      "0000100" when "01000111010101100", -- t[36524] = 4
      "0000100" when "01000111010101101", -- t[36525] = 4
      "0000100" when "01000111010101110", -- t[36526] = 4
      "0000100" when "01000111010101111", -- t[36527] = 4
      "0000100" when "01000111010110000", -- t[36528] = 4
      "0000100" when "01000111010110001", -- t[36529] = 4
      "0000100" when "01000111010110010", -- t[36530] = 4
      "0000100" when "01000111010110011", -- t[36531] = 4
      "0000100" when "01000111010110100", -- t[36532] = 4
      "0000100" when "01000111010110101", -- t[36533] = 4
      "0000100" when "01000111010110110", -- t[36534] = 4
      "0000100" when "01000111010110111", -- t[36535] = 4
      "0000100" when "01000111010111000", -- t[36536] = 4
      "0000100" when "01000111010111001", -- t[36537] = 4
      "0000100" when "01000111010111010", -- t[36538] = 4
      "0000100" when "01000111010111011", -- t[36539] = 4
      "0000100" when "01000111010111100", -- t[36540] = 4
      "0000100" when "01000111010111101", -- t[36541] = 4
      "0000100" when "01000111010111110", -- t[36542] = 4
      "0000100" when "01000111010111111", -- t[36543] = 4
      "0000100" when "01000111011000000", -- t[36544] = 4
      "0000100" when "01000111011000001", -- t[36545] = 4
      "0000100" when "01000111011000010", -- t[36546] = 4
      "0000100" when "01000111011000011", -- t[36547] = 4
      "0000100" when "01000111011000100", -- t[36548] = 4
      "0000100" when "01000111011000101", -- t[36549] = 4
      "0000100" when "01000111011000110", -- t[36550] = 4
      "0000100" when "01000111011000111", -- t[36551] = 4
      "0000100" when "01000111011001000", -- t[36552] = 4
      "0000100" when "01000111011001001", -- t[36553] = 4
      "0000100" when "01000111011001010", -- t[36554] = 4
      "0000100" when "01000111011001011", -- t[36555] = 4
      "0000100" when "01000111011001100", -- t[36556] = 4
      "0000100" when "01000111011001101", -- t[36557] = 4
      "0000100" when "01000111011001110", -- t[36558] = 4
      "0000100" when "01000111011001111", -- t[36559] = 4
      "0000100" when "01000111011010000", -- t[36560] = 4
      "0000100" when "01000111011010001", -- t[36561] = 4
      "0000100" when "01000111011010010", -- t[36562] = 4
      "0000100" when "01000111011010011", -- t[36563] = 4
      "0000100" when "01000111011010100", -- t[36564] = 4
      "0000100" when "01000111011010101", -- t[36565] = 4
      "0000100" when "01000111011010110", -- t[36566] = 4
      "0000100" when "01000111011010111", -- t[36567] = 4
      "0000100" when "01000111011011000", -- t[36568] = 4
      "0000100" when "01000111011011001", -- t[36569] = 4
      "0000100" when "01000111011011010", -- t[36570] = 4
      "0000100" when "01000111011011011", -- t[36571] = 4
      "0000100" when "01000111011011100", -- t[36572] = 4
      "0000100" when "01000111011011101", -- t[36573] = 4
      "0000100" when "01000111011011110", -- t[36574] = 4
      "0000100" when "01000111011011111", -- t[36575] = 4
      "0000100" when "01000111011100000", -- t[36576] = 4
      "0000100" when "01000111011100001", -- t[36577] = 4
      "0000100" when "01000111011100010", -- t[36578] = 4
      "0000100" when "01000111011100011", -- t[36579] = 4
      "0000100" when "01000111011100100", -- t[36580] = 4
      "0000100" when "01000111011100101", -- t[36581] = 4
      "0000100" when "01000111011100110", -- t[36582] = 4
      "0000100" when "01000111011100111", -- t[36583] = 4
      "0000100" when "01000111011101000", -- t[36584] = 4
      "0000100" when "01000111011101001", -- t[36585] = 4
      "0000100" when "01000111011101010", -- t[36586] = 4
      "0000100" when "01000111011101011", -- t[36587] = 4
      "0000100" when "01000111011101100", -- t[36588] = 4
      "0000100" when "01000111011101101", -- t[36589] = 4
      "0000100" when "01000111011101110", -- t[36590] = 4
      "0000100" when "01000111011101111", -- t[36591] = 4
      "0000100" when "01000111011110000", -- t[36592] = 4
      "0000100" when "01000111011110001", -- t[36593] = 4
      "0000100" when "01000111011110010", -- t[36594] = 4
      "0000100" when "01000111011110011", -- t[36595] = 4
      "0000100" when "01000111011110100", -- t[36596] = 4
      "0000100" when "01000111011110101", -- t[36597] = 4
      "0000100" when "01000111011110110", -- t[36598] = 4
      "0000100" when "01000111011110111", -- t[36599] = 4
      "0000100" when "01000111011111000", -- t[36600] = 4
      "0000100" when "01000111011111001", -- t[36601] = 4
      "0000100" when "01000111011111010", -- t[36602] = 4
      "0000100" when "01000111011111011", -- t[36603] = 4
      "0000100" when "01000111011111100", -- t[36604] = 4
      "0000100" when "01000111011111101", -- t[36605] = 4
      "0000100" when "01000111011111110", -- t[36606] = 4
      "0000100" when "01000111011111111", -- t[36607] = 4
      "0000100" when "01000111100000000", -- t[36608] = 4
      "0000100" when "01000111100000001", -- t[36609] = 4
      "0000100" when "01000111100000010", -- t[36610] = 4
      "0000100" when "01000111100000011", -- t[36611] = 4
      "0000100" when "01000111100000100", -- t[36612] = 4
      "0000100" when "01000111100000101", -- t[36613] = 4
      "0000100" when "01000111100000110", -- t[36614] = 4
      "0000100" when "01000111100000111", -- t[36615] = 4
      "0000100" when "01000111100001000", -- t[36616] = 4
      "0000100" when "01000111100001001", -- t[36617] = 4
      "0000100" when "01000111100001010", -- t[36618] = 4
      "0000100" when "01000111100001011", -- t[36619] = 4
      "0000100" when "01000111100001100", -- t[36620] = 4
      "0000100" when "01000111100001101", -- t[36621] = 4
      "0000100" when "01000111100001110", -- t[36622] = 4
      "0000100" when "01000111100001111", -- t[36623] = 4
      "0000100" when "01000111100010000", -- t[36624] = 4
      "0000100" when "01000111100010001", -- t[36625] = 4
      "0000100" when "01000111100010010", -- t[36626] = 4
      "0000100" when "01000111100010011", -- t[36627] = 4
      "0000100" when "01000111100010100", -- t[36628] = 4
      "0000100" when "01000111100010101", -- t[36629] = 4
      "0000100" when "01000111100010110", -- t[36630] = 4
      "0000100" when "01000111100010111", -- t[36631] = 4
      "0000100" when "01000111100011000", -- t[36632] = 4
      "0000100" when "01000111100011001", -- t[36633] = 4
      "0000100" when "01000111100011010", -- t[36634] = 4
      "0000100" when "01000111100011011", -- t[36635] = 4
      "0000100" when "01000111100011100", -- t[36636] = 4
      "0000100" when "01000111100011101", -- t[36637] = 4
      "0000100" when "01000111100011110", -- t[36638] = 4
      "0000100" when "01000111100011111", -- t[36639] = 4
      "0000100" when "01000111100100000", -- t[36640] = 4
      "0000100" when "01000111100100001", -- t[36641] = 4
      "0000100" when "01000111100100010", -- t[36642] = 4
      "0000100" when "01000111100100011", -- t[36643] = 4
      "0000100" when "01000111100100100", -- t[36644] = 4
      "0000100" when "01000111100100101", -- t[36645] = 4
      "0000100" when "01000111100100110", -- t[36646] = 4
      "0000100" when "01000111100100111", -- t[36647] = 4
      "0000100" when "01000111100101000", -- t[36648] = 4
      "0000100" when "01000111100101001", -- t[36649] = 4
      "0000100" when "01000111100101010", -- t[36650] = 4
      "0000100" when "01000111100101011", -- t[36651] = 4
      "0000100" when "01000111100101100", -- t[36652] = 4
      "0000100" when "01000111100101101", -- t[36653] = 4
      "0000100" when "01000111100101110", -- t[36654] = 4
      "0000100" when "01000111100101111", -- t[36655] = 4
      "0000100" when "01000111100110000", -- t[36656] = 4
      "0000100" when "01000111100110001", -- t[36657] = 4
      "0000100" when "01000111100110010", -- t[36658] = 4
      "0000100" when "01000111100110011", -- t[36659] = 4
      "0000100" when "01000111100110100", -- t[36660] = 4
      "0000100" when "01000111100110101", -- t[36661] = 4
      "0000100" when "01000111100110110", -- t[36662] = 4
      "0000100" when "01000111100110111", -- t[36663] = 4
      "0000100" when "01000111100111000", -- t[36664] = 4
      "0000100" when "01000111100111001", -- t[36665] = 4
      "0000100" when "01000111100111010", -- t[36666] = 4
      "0000100" when "01000111100111011", -- t[36667] = 4
      "0000100" when "01000111100111100", -- t[36668] = 4
      "0000100" when "01000111100111101", -- t[36669] = 4
      "0000100" when "01000111100111110", -- t[36670] = 4
      "0000100" when "01000111100111111", -- t[36671] = 4
      "0000100" when "01000111101000000", -- t[36672] = 4
      "0000100" when "01000111101000001", -- t[36673] = 4
      "0000100" when "01000111101000010", -- t[36674] = 4
      "0000100" when "01000111101000011", -- t[36675] = 4
      "0000100" when "01000111101000100", -- t[36676] = 4
      "0000100" when "01000111101000101", -- t[36677] = 4
      "0000100" when "01000111101000110", -- t[36678] = 4
      "0000100" when "01000111101000111", -- t[36679] = 4
      "0000100" when "01000111101001000", -- t[36680] = 4
      "0000100" when "01000111101001001", -- t[36681] = 4
      "0000100" when "01000111101001010", -- t[36682] = 4
      "0000100" when "01000111101001011", -- t[36683] = 4
      "0000100" when "01000111101001100", -- t[36684] = 4
      "0000100" when "01000111101001101", -- t[36685] = 4
      "0000100" when "01000111101001110", -- t[36686] = 4
      "0000100" when "01000111101001111", -- t[36687] = 4
      "0000100" when "01000111101010000", -- t[36688] = 4
      "0000100" when "01000111101010001", -- t[36689] = 4
      "0000100" when "01000111101010010", -- t[36690] = 4
      "0000100" when "01000111101010011", -- t[36691] = 4
      "0000100" when "01000111101010100", -- t[36692] = 4
      "0000100" when "01000111101010101", -- t[36693] = 4
      "0000100" when "01000111101010110", -- t[36694] = 4
      "0000100" when "01000111101010111", -- t[36695] = 4
      "0000100" when "01000111101011000", -- t[36696] = 4
      "0000100" when "01000111101011001", -- t[36697] = 4
      "0000100" when "01000111101011010", -- t[36698] = 4
      "0000100" when "01000111101011011", -- t[36699] = 4
      "0000100" when "01000111101011100", -- t[36700] = 4
      "0000100" when "01000111101011101", -- t[36701] = 4
      "0000100" when "01000111101011110", -- t[36702] = 4
      "0000100" when "01000111101011111", -- t[36703] = 4
      "0000100" when "01000111101100000", -- t[36704] = 4
      "0000100" when "01000111101100001", -- t[36705] = 4
      "0000100" when "01000111101100010", -- t[36706] = 4
      "0000100" when "01000111101100011", -- t[36707] = 4
      "0000100" when "01000111101100100", -- t[36708] = 4
      "0000100" when "01000111101100101", -- t[36709] = 4
      "0000100" when "01000111101100110", -- t[36710] = 4
      "0000100" when "01000111101100111", -- t[36711] = 4
      "0000100" when "01000111101101000", -- t[36712] = 4
      "0000100" when "01000111101101001", -- t[36713] = 4
      "0000100" when "01000111101101010", -- t[36714] = 4
      "0000100" when "01000111101101011", -- t[36715] = 4
      "0000100" when "01000111101101100", -- t[36716] = 4
      "0000100" when "01000111101101101", -- t[36717] = 4
      "0000100" when "01000111101101110", -- t[36718] = 4
      "0000100" when "01000111101101111", -- t[36719] = 4
      "0000100" when "01000111101110000", -- t[36720] = 4
      "0000100" when "01000111101110001", -- t[36721] = 4
      "0000100" when "01000111101110010", -- t[36722] = 4
      "0000100" when "01000111101110011", -- t[36723] = 4
      "0000100" when "01000111101110100", -- t[36724] = 4
      "0000100" when "01000111101110101", -- t[36725] = 4
      "0000100" when "01000111101110110", -- t[36726] = 4
      "0000100" when "01000111101110111", -- t[36727] = 4
      "0000100" when "01000111101111000", -- t[36728] = 4
      "0000100" when "01000111101111001", -- t[36729] = 4
      "0000100" when "01000111101111010", -- t[36730] = 4
      "0000100" when "01000111101111011", -- t[36731] = 4
      "0000100" when "01000111101111100", -- t[36732] = 4
      "0000100" when "01000111101111101", -- t[36733] = 4
      "0000100" when "01000111101111110", -- t[36734] = 4
      "0000100" when "01000111101111111", -- t[36735] = 4
      "0000100" when "01000111110000000", -- t[36736] = 4
      "0000100" when "01000111110000001", -- t[36737] = 4
      "0000100" when "01000111110000010", -- t[36738] = 4
      "0000100" when "01000111110000011", -- t[36739] = 4
      "0000100" when "01000111110000100", -- t[36740] = 4
      "0000100" when "01000111110000101", -- t[36741] = 4
      "0000100" when "01000111110000110", -- t[36742] = 4
      "0000100" when "01000111110000111", -- t[36743] = 4
      "0000100" when "01000111110001000", -- t[36744] = 4
      "0000100" when "01000111110001001", -- t[36745] = 4
      "0000100" when "01000111110001010", -- t[36746] = 4
      "0000100" when "01000111110001011", -- t[36747] = 4
      "0000100" when "01000111110001100", -- t[36748] = 4
      "0000100" when "01000111110001101", -- t[36749] = 4
      "0000100" when "01000111110001110", -- t[36750] = 4
      "0000100" when "01000111110001111", -- t[36751] = 4
      "0000100" when "01000111110010000", -- t[36752] = 4
      "0000100" when "01000111110010001", -- t[36753] = 4
      "0000100" when "01000111110010010", -- t[36754] = 4
      "0000100" when "01000111110010011", -- t[36755] = 4
      "0000100" when "01000111110010100", -- t[36756] = 4
      "0000100" when "01000111110010101", -- t[36757] = 4
      "0000100" when "01000111110010110", -- t[36758] = 4
      "0000100" when "01000111110010111", -- t[36759] = 4
      "0000100" when "01000111110011000", -- t[36760] = 4
      "0000100" when "01000111110011001", -- t[36761] = 4
      "0000100" when "01000111110011010", -- t[36762] = 4
      "0000100" when "01000111110011011", -- t[36763] = 4
      "0000100" when "01000111110011100", -- t[36764] = 4
      "0000100" when "01000111110011101", -- t[36765] = 4
      "0000100" when "01000111110011110", -- t[36766] = 4
      "0000100" when "01000111110011111", -- t[36767] = 4
      "0000100" when "01000111110100000", -- t[36768] = 4
      "0000100" when "01000111110100001", -- t[36769] = 4
      "0000100" when "01000111110100010", -- t[36770] = 4
      "0000100" when "01000111110100011", -- t[36771] = 4
      "0000100" when "01000111110100100", -- t[36772] = 4
      "0000100" when "01000111110100101", -- t[36773] = 4
      "0000100" when "01000111110100110", -- t[36774] = 4
      "0000100" when "01000111110100111", -- t[36775] = 4
      "0000100" when "01000111110101000", -- t[36776] = 4
      "0000100" when "01000111110101001", -- t[36777] = 4
      "0000100" when "01000111110101010", -- t[36778] = 4
      "0000100" when "01000111110101011", -- t[36779] = 4
      "0000100" when "01000111110101100", -- t[36780] = 4
      "0000100" when "01000111110101101", -- t[36781] = 4
      "0000100" when "01000111110101110", -- t[36782] = 4
      "0000100" when "01000111110101111", -- t[36783] = 4
      "0000100" when "01000111110110000", -- t[36784] = 4
      "0000100" when "01000111110110001", -- t[36785] = 4
      "0000100" when "01000111110110010", -- t[36786] = 4
      "0000100" when "01000111110110011", -- t[36787] = 4
      "0000100" when "01000111110110100", -- t[36788] = 4
      "0000100" when "01000111110110101", -- t[36789] = 4
      "0000100" when "01000111110110110", -- t[36790] = 4
      "0000100" when "01000111110110111", -- t[36791] = 4
      "0000100" when "01000111110111000", -- t[36792] = 4
      "0000100" when "01000111110111001", -- t[36793] = 4
      "0000100" when "01000111110111010", -- t[36794] = 4
      "0000100" when "01000111110111011", -- t[36795] = 4
      "0000100" when "01000111110111100", -- t[36796] = 4
      "0000100" when "01000111110111101", -- t[36797] = 4
      "0000100" when "01000111110111110", -- t[36798] = 4
      "0000100" when "01000111110111111", -- t[36799] = 4
      "0000100" when "01000111111000000", -- t[36800] = 4
      "0000100" when "01000111111000001", -- t[36801] = 4
      "0000100" when "01000111111000010", -- t[36802] = 4
      "0000100" when "01000111111000011", -- t[36803] = 4
      "0000100" when "01000111111000100", -- t[36804] = 4
      "0000100" when "01000111111000101", -- t[36805] = 4
      "0000100" when "01000111111000110", -- t[36806] = 4
      "0000100" when "01000111111000111", -- t[36807] = 4
      "0000100" when "01000111111001000", -- t[36808] = 4
      "0000100" when "01000111111001001", -- t[36809] = 4
      "0000100" when "01000111111001010", -- t[36810] = 4
      "0000100" when "01000111111001011", -- t[36811] = 4
      "0000100" when "01000111111001100", -- t[36812] = 4
      "0000100" when "01000111111001101", -- t[36813] = 4
      "0000100" when "01000111111001110", -- t[36814] = 4
      "0000100" when "01000111111001111", -- t[36815] = 4
      "0000100" when "01000111111010000", -- t[36816] = 4
      "0000100" when "01000111111010001", -- t[36817] = 4
      "0000100" when "01000111111010010", -- t[36818] = 4
      "0000100" when "01000111111010011", -- t[36819] = 4
      "0000100" when "01000111111010100", -- t[36820] = 4
      "0000100" when "01000111111010101", -- t[36821] = 4
      "0000100" when "01000111111010110", -- t[36822] = 4
      "0000100" when "01000111111010111", -- t[36823] = 4
      "0000100" when "01000111111011000", -- t[36824] = 4
      "0000100" when "01000111111011001", -- t[36825] = 4
      "0000100" when "01000111111011010", -- t[36826] = 4
      "0000100" when "01000111111011011", -- t[36827] = 4
      "0000100" when "01000111111011100", -- t[36828] = 4
      "0000100" when "01000111111011101", -- t[36829] = 4
      "0000100" when "01000111111011110", -- t[36830] = 4
      "0000100" when "01000111111011111", -- t[36831] = 4
      "0000100" when "01000111111100000", -- t[36832] = 4
      "0000100" when "01000111111100001", -- t[36833] = 4
      "0000100" when "01000111111100010", -- t[36834] = 4
      "0000100" when "01000111111100011", -- t[36835] = 4
      "0000100" when "01000111111100100", -- t[36836] = 4
      "0000100" when "01000111111100101", -- t[36837] = 4
      "0000100" when "01000111111100110", -- t[36838] = 4
      "0000100" when "01000111111100111", -- t[36839] = 4
      "0000100" when "01000111111101000", -- t[36840] = 4
      "0000100" when "01000111111101001", -- t[36841] = 4
      "0000100" when "01000111111101010", -- t[36842] = 4
      "0000100" when "01000111111101011", -- t[36843] = 4
      "0000100" when "01000111111101100", -- t[36844] = 4
      "0000100" when "01000111111101101", -- t[36845] = 4
      "0000100" when "01000111111101110", -- t[36846] = 4
      "0000100" when "01000111111101111", -- t[36847] = 4
      "0000100" when "01000111111110000", -- t[36848] = 4
      "0000100" when "01000111111110001", -- t[36849] = 4
      "0000100" when "01000111111110010", -- t[36850] = 4
      "0000100" when "01000111111110011", -- t[36851] = 4
      "0000100" when "01000111111110100", -- t[36852] = 4
      "0000100" when "01000111111110101", -- t[36853] = 4
      "0000100" when "01000111111110110", -- t[36854] = 4
      "0000100" when "01000111111110111", -- t[36855] = 4
      "0000100" when "01000111111111000", -- t[36856] = 4
      "0000100" when "01000111111111001", -- t[36857] = 4
      "0000100" when "01000111111111010", -- t[36858] = 4
      "0000100" when "01000111111111011", -- t[36859] = 4
      "0000100" when "01000111111111100", -- t[36860] = 4
      "0000100" when "01000111111111101", -- t[36861] = 4
      "0000100" when "01000111111111110", -- t[36862] = 4
      "0000100" when "01000111111111111", -- t[36863] = 4
      "0000100" when "01001000000000000", -- t[36864] = 4
      "0000100" when "01001000000000001", -- t[36865] = 4
      "0000100" when "01001000000000010", -- t[36866] = 4
      "0000100" when "01001000000000011", -- t[36867] = 4
      "0000100" when "01001000000000100", -- t[36868] = 4
      "0000100" when "01001000000000101", -- t[36869] = 4
      "0000100" when "01001000000000110", -- t[36870] = 4
      "0000100" when "01001000000000111", -- t[36871] = 4
      "0000100" when "01001000000001000", -- t[36872] = 4
      "0000100" when "01001000000001001", -- t[36873] = 4
      "0000100" when "01001000000001010", -- t[36874] = 4
      "0000100" when "01001000000001011", -- t[36875] = 4
      "0000100" when "01001000000001100", -- t[36876] = 4
      "0000100" when "01001000000001101", -- t[36877] = 4
      "0000100" when "01001000000001110", -- t[36878] = 4
      "0000100" when "01001000000001111", -- t[36879] = 4
      "0000100" when "01001000000010000", -- t[36880] = 4
      "0000100" when "01001000000010001", -- t[36881] = 4
      "0000100" when "01001000000010010", -- t[36882] = 4
      "0000100" when "01001000000010011", -- t[36883] = 4
      "0000100" when "01001000000010100", -- t[36884] = 4
      "0000100" when "01001000000010101", -- t[36885] = 4
      "0000100" when "01001000000010110", -- t[36886] = 4
      "0000100" when "01001000000010111", -- t[36887] = 4
      "0000100" when "01001000000011000", -- t[36888] = 4
      "0000100" when "01001000000011001", -- t[36889] = 4
      "0000100" when "01001000000011010", -- t[36890] = 4
      "0000100" when "01001000000011011", -- t[36891] = 4
      "0000100" when "01001000000011100", -- t[36892] = 4
      "0000100" when "01001000000011101", -- t[36893] = 4
      "0000100" when "01001000000011110", -- t[36894] = 4
      "0000100" when "01001000000011111", -- t[36895] = 4
      "0000100" when "01001000000100000", -- t[36896] = 4
      "0000100" when "01001000000100001", -- t[36897] = 4
      "0000100" when "01001000000100010", -- t[36898] = 4
      "0000100" when "01001000000100011", -- t[36899] = 4
      "0000100" when "01001000000100100", -- t[36900] = 4
      "0000100" when "01001000000100101", -- t[36901] = 4
      "0000100" when "01001000000100110", -- t[36902] = 4
      "0000100" when "01001000000100111", -- t[36903] = 4
      "0000100" when "01001000000101000", -- t[36904] = 4
      "0000100" when "01001000000101001", -- t[36905] = 4
      "0000100" when "01001000000101010", -- t[36906] = 4
      "0000100" when "01001000000101011", -- t[36907] = 4
      "0000100" when "01001000000101100", -- t[36908] = 4
      "0000100" when "01001000000101101", -- t[36909] = 4
      "0000100" when "01001000000101110", -- t[36910] = 4
      "0000100" when "01001000000101111", -- t[36911] = 4
      "0000100" when "01001000000110000", -- t[36912] = 4
      "0000100" when "01001000000110001", -- t[36913] = 4
      "0000100" when "01001000000110010", -- t[36914] = 4
      "0000100" when "01001000000110011", -- t[36915] = 4
      "0000100" when "01001000000110100", -- t[36916] = 4
      "0000100" when "01001000000110101", -- t[36917] = 4
      "0000100" when "01001000000110110", -- t[36918] = 4
      "0000100" when "01001000000110111", -- t[36919] = 4
      "0000100" when "01001000000111000", -- t[36920] = 4
      "0000100" when "01001000000111001", -- t[36921] = 4
      "0000100" when "01001000000111010", -- t[36922] = 4
      "0000100" when "01001000000111011", -- t[36923] = 4
      "0000100" when "01001000000111100", -- t[36924] = 4
      "0000100" when "01001000000111101", -- t[36925] = 4
      "0000100" when "01001000000111110", -- t[36926] = 4
      "0000100" when "01001000000111111", -- t[36927] = 4
      "0000100" when "01001000001000000", -- t[36928] = 4
      "0000100" when "01001000001000001", -- t[36929] = 4
      "0000100" when "01001000001000010", -- t[36930] = 4
      "0000100" when "01001000001000011", -- t[36931] = 4
      "0000100" when "01001000001000100", -- t[36932] = 4
      "0000100" when "01001000001000101", -- t[36933] = 4
      "0000100" when "01001000001000110", -- t[36934] = 4
      "0000100" when "01001000001000111", -- t[36935] = 4
      "0000100" when "01001000001001000", -- t[36936] = 4
      "0000100" when "01001000001001001", -- t[36937] = 4
      "0000100" when "01001000001001010", -- t[36938] = 4
      "0000100" when "01001000001001011", -- t[36939] = 4
      "0000100" when "01001000001001100", -- t[36940] = 4
      "0000100" when "01001000001001101", -- t[36941] = 4
      "0000100" when "01001000001001110", -- t[36942] = 4
      "0000100" when "01001000001001111", -- t[36943] = 4
      "0000100" when "01001000001010000", -- t[36944] = 4
      "0000100" when "01001000001010001", -- t[36945] = 4
      "0000100" when "01001000001010010", -- t[36946] = 4
      "0000100" when "01001000001010011", -- t[36947] = 4
      "0000100" when "01001000001010100", -- t[36948] = 4
      "0000100" when "01001000001010101", -- t[36949] = 4
      "0000100" when "01001000001010110", -- t[36950] = 4
      "0000100" when "01001000001010111", -- t[36951] = 4
      "0000100" when "01001000001011000", -- t[36952] = 4
      "0000100" when "01001000001011001", -- t[36953] = 4
      "0000100" when "01001000001011010", -- t[36954] = 4
      "0000100" when "01001000001011011", -- t[36955] = 4
      "0000100" when "01001000001011100", -- t[36956] = 4
      "0000100" when "01001000001011101", -- t[36957] = 4
      "0000100" when "01001000001011110", -- t[36958] = 4
      "0000100" when "01001000001011111", -- t[36959] = 4
      "0000100" when "01001000001100000", -- t[36960] = 4
      "0000100" when "01001000001100001", -- t[36961] = 4
      "0000100" when "01001000001100010", -- t[36962] = 4
      "0000100" when "01001000001100011", -- t[36963] = 4
      "0000100" when "01001000001100100", -- t[36964] = 4
      "0000100" when "01001000001100101", -- t[36965] = 4
      "0000100" when "01001000001100110", -- t[36966] = 4
      "0000100" when "01001000001100111", -- t[36967] = 4
      "0000100" when "01001000001101000", -- t[36968] = 4
      "0000100" when "01001000001101001", -- t[36969] = 4
      "0000100" when "01001000001101010", -- t[36970] = 4
      "0000100" when "01001000001101011", -- t[36971] = 4
      "0000100" when "01001000001101100", -- t[36972] = 4
      "0000100" when "01001000001101101", -- t[36973] = 4
      "0000100" when "01001000001101110", -- t[36974] = 4
      "0000100" when "01001000001101111", -- t[36975] = 4
      "0000100" when "01001000001110000", -- t[36976] = 4
      "0000100" when "01001000001110001", -- t[36977] = 4
      "0000100" when "01001000001110010", -- t[36978] = 4
      "0000100" when "01001000001110011", -- t[36979] = 4
      "0000100" when "01001000001110100", -- t[36980] = 4
      "0000100" when "01001000001110101", -- t[36981] = 4
      "0000100" when "01001000001110110", -- t[36982] = 4
      "0000100" when "01001000001110111", -- t[36983] = 4
      "0000100" when "01001000001111000", -- t[36984] = 4
      "0000100" when "01001000001111001", -- t[36985] = 4
      "0000100" when "01001000001111010", -- t[36986] = 4
      "0000100" when "01001000001111011", -- t[36987] = 4
      "0000100" when "01001000001111100", -- t[36988] = 4
      "0000100" when "01001000001111101", -- t[36989] = 4
      "0000100" when "01001000001111110", -- t[36990] = 4
      "0000100" when "01001000001111111", -- t[36991] = 4
      "0000100" when "01001000010000000", -- t[36992] = 4
      "0000100" when "01001000010000001", -- t[36993] = 4
      "0000100" when "01001000010000010", -- t[36994] = 4
      "0000100" when "01001000010000011", -- t[36995] = 4
      "0000100" when "01001000010000100", -- t[36996] = 4
      "0000100" when "01001000010000101", -- t[36997] = 4
      "0000100" when "01001000010000110", -- t[36998] = 4
      "0000100" when "01001000010000111", -- t[36999] = 4
      "0000100" when "01001000010001000", -- t[37000] = 4
      "0000100" when "01001000010001001", -- t[37001] = 4
      "0000100" when "01001000010001010", -- t[37002] = 4
      "0000100" when "01001000010001011", -- t[37003] = 4
      "0000100" when "01001000010001100", -- t[37004] = 4
      "0000100" when "01001000010001101", -- t[37005] = 4
      "0000100" when "01001000010001110", -- t[37006] = 4
      "0000100" when "01001000010001111", -- t[37007] = 4
      "0000100" when "01001000010010000", -- t[37008] = 4
      "0000100" when "01001000010010001", -- t[37009] = 4
      "0000100" when "01001000010010010", -- t[37010] = 4
      "0000100" when "01001000010010011", -- t[37011] = 4
      "0000100" when "01001000010010100", -- t[37012] = 4
      "0000100" when "01001000010010101", -- t[37013] = 4
      "0000100" when "01001000010010110", -- t[37014] = 4
      "0000100" when "01001000010010111", -- t[37015] = 4
      "0000100" when "01001000010011000", -- t[37016] = 4
      "0000100" when "01001000010011001", -- t[37017] = 4
      "0000100" when "01001000010011010", -- t[37018] = 4
      "0000100" when "01001000010011011", -- t[37019] = 4
      "0000100" when "01001000010011100", -- t[37020] = 4
      "0000100" when "01001000010011101", -- t[37021] = 4
      "0000100" when "01001000010011110", -- t[37022] = 4
      "0000100" when "01001000010011111", -- t[37023] = 4
      "0000100" when "01001000010100000", -- t[37024] = 4
      "0000100" when "01001000010100001", -- t[37025] = 4
      "0000100" when "01001000010100010", -- t[37026] = 4
      "0000100" when "01001000010100011", -- t[37027] = 4
      "0000100" when "01001000010100100", -- t[37028] = 4
      "0000100" when "01001000010100101", -- t[37029] = 4
      "0000100" when "01001000010100110", -- t[37030] = 4
      "0000100" when "01001000010100111", -- t[37031] = 4
      "0000100" when "01001000010101000", -- t[37032] = 4
      "0000100" when "01001000010101001", -- t[37033] = 4
      "0000100" when "01001000010101010", -- t[37034] = 4
      "0000100" when "01001000010101011", -- t[37035] = 4
      "0000100" when "01001000010101100", -- t[37036] = 4
      "0000100" when "01001000010101101", -- t[37037] = 4
      "0000100" when "01001000010101110", -- t[37038] = 4
      "0000100" when "01001000010101111", -- t[37039] = 4
      "0000100" when "01001000010110000", -- t[37040] = 4
      "0000100" when "01001000010110001", -- t[37041] = 4
      "0000100" when "01001000010110010", -- t[37042] = 4
      "0000100" when "01001000010110011", -- t[37043] = 4
      "0000100" when "01001000010110100", -- t[37044] = 4
      "0000100" when "01001000010110101", -- t[37045] = 4
      "0000100" when "01001000010110110", -- t[37046] = 4
      "0000100" when "01001000010110111", -- t[37047] = 4
      "0000100" when "01001000010111000", -- t[37048] = 4
      "0000100" when "01001000010111001", -- t[37049] = 4
      "0000100" when "01001000010111010", -- t[37050] = 4
      "0000100" when "01001000010111011", -- t[37051] = 4
      "0000100" when "01001000010111100", -- t[37052] = 4
      "0000100" when "01001000010111101", -- t[37053] = 4
      "0000100" when "01001000010111110", -- t[37054] = 4
      "0000100" when "01001000010111111", -- t[37055] = 4
      "0000100" when "01001000011000000", -- t[37056] = 4
      "0000100" when "01001000011000001", -- t[37057] = 4
      "0000100" when "01001000011000010", -- t[37058] = 4
      "0000100" when "01001000011000011", -- t[37059] = 4
      "0000100" when "01001000011000100", -- t[37060] = 4
      "0000100" when "01001000011000101", -- t[37061] = 4
      "0000100" when "01001000011000110", -- t[37062] = 4
      "0000100" when "01001000011000111", -- t[37063] = 4
      "0000100" when "01001000011001000", -- t[37064] = 4
      "0000100" when "01001000011001001", -- t[37065] = 4
      "0000100" when "01001000011001010", -- t[37066] = 4
      "0000100" when "01001000011001011", -- t[37067] = 4
      "0000100" when "01001000011001100", -- t[37068] = 4
      "0000100" when "01001000011001101", -- t[37069] = 4
      "0000100" when "01001000011001110", -- t[37070] = 4
      "0000100" when "01001000011001111", -- t[37071] = 4
      "0000100" when "01001000011010000", -- t[37072] = 4
      "0000100" when "01001000011010001", -- t[37073] = 4
      "0000100" when "01001000011010010", -- t[37074] = 4
      "0000100" when "01001000011010011", -- t[37075] = 4
      "0000100" when "01001000011010100", -- t[37076] = 4
      "0000100" when "01001000011010101", -- t[37077] = 4
      "0000100" when "01001000011010110", -- t[37078] = 4
      "0000100" when "01001000011010111", -- t[37079] = 4
      "0000100" when "01001000011011000", -- t[37080] = 4
      "0000100" when "01001000011011001", -- t[37081] = 4
      "0000100" when "01001000011011010", -- t[37082] = 4
      "0000100" when "01001000011011011", -- t[37083] = 4
      "0000100" when "01001000011011100", -- t[37084] = 4
      "0000100" when "01001000011011101", -- t[37085] = 4
      "0000100" when "01001000011011110", -- t[37086] = 4
      "0000100" when "01001000011011111", -- t[37087] = 4
      "0000100" when "01001000011100000", -- t[37088] = 4
      "0000100" when "01001000011100001", -- t[37089] = 4
      "0000100" when "01001000011100010", -- t[37090] = 4
      "0000100" when "01001000011100011", -- t[37091] = 4
      "0000100" when "01001000011100100", -- t[37092] = 4
      "0000100" when "01001000011100101", -- t[37093] = 4
      "0000100" when "01001000011100110", -- t[37094] = 4
      "0000100" when "01001000011100111", -- t[37095] = 4
      "0000100" when "01001000011101000", -- t[37096] = 4
      "0000100" when "01001000011101001", -- t[37097] = 4
      "0000100" when "01001000011101010", -- t[37098] = 4
      "0000100" when "01001000011101011", -- t[37099] = 4
      "0000100" when "01001000011101100", -- t[37100] = 4
      "0000100" when "01001000011101101", -- t[37101] = 4
      "0000100" when "01001000011101110", -- t[37102] = 4
      "0000100" when "01001000011101111", -- t[37103] = 4
      "0000100" when "01001000011110000", -- t[37104] = 4
      "0000100" when "01001000011110001", -- t[37105] = 4
      "0000100" when "01001000011110010", -- t[37106] = 4
      "0000100" when "01001000011110011", -- t[37107] = 4
      "0000100" when "01001000011110100", -- t[37108] = 4
      "0000100" when "01001000011110101", -- t[37109] = 4
      "0000100" when "01001000011110110", -- t[37110] = 4
      "0000100" when "01001000011110111", -- t[37111] = 4
      "0000100" when "01001000011111000", -- t[37112] = 4
      "0000100" when "01001000011111001", -- t[37113] = 4
      "0000100" when "01001000011111010", -- t[37114] = 4
      "0000100" when "01001000011111011", -- t[37115] = 4
      "0000100" when "01001000011111100", -- t[37116] = 4
      "0000100" when "01001000011111101", -- t[37117] = 4
      "0000100" when "01001000011111110", -- t[37118] = 4
      "0000100" when "01001000011111111", -- t[37119] = 4
      "0000100" when "01001000100000000", -- t[37120] = 4
      "0000100" when "01001000100000001", -- t[37121] = 4
      "0000100" when "01001000100000010", -- t[37122] = 4
      "0000100" when "01001000100000011", -- t[37123] = 4
      "0000100" when "01001000100000100", -- t[37124] = 4
      "0000100" when "01001000100000101", -- t[37125] = 4
      "0000100" when "01001000100000110", -- t[37126] = 4
      "0000100" when "01001000100000111", -- t[37127] = 4
      "0000100" when "01001000100001000", -- t[37128] = 4
      "0000100" when "01001000100001001", -- t[37129] = 4
      "0000100" when "01001000100001010", -- t[37130] = 4
      "0000100" when "01001000100001011", -- t[37131] = 4
      "0000100" when "01001000100001100", -- t[37132] = 4
      "0000100" when "01001000100001101", -- t[37133] = 4
      "0000100" when "01001000100001110", -- t[37134] = 4
      "0000100" when "01001000100001111", -- t[37135] = 4
      "0000100" when "01001000100010000", -- t[37136] = 4
      "0000100" when "01001000100010001", -- t[37137] = 4
      "0000100" when "01001000100010010", -- t[37138] = 4
      "0000100" when "01001000100010011", -- t[37139] = 4
      "0000100" when "01001000100010100", -- t[37140] = 4
      "0000100" when "01001000100010101", -- t[37141] = 4
      "0000100" when "01001000100010110", -- t[37142] = 4
      "0000100" when "01001000100010111", -- t[37143] = 4
      "0000100" when "01001000100011000", -- t[37144] = 4
      "0000100" when "01001000100011001", -- t[37145] = 4
      "0000100" when "01001000100011010", -- t[37146] = 4
      "0000100" when "01001000100011011", -- t[37147] = 4
      "0000100" when "01001000100011100", -- t[37148] = 4
      "0000100" when "01001000100011101", -- t[37149] = 4
      "0000100" when "01001000100011110", -- t[37150] = 4
      "0000100" when "01001000100011111", -- t[37151] = 4
      "0000100" when "01001000100100000", -- t[37152] = 4
      "0000100" when "01001000100100001", -- t[37153] = 4
      "0000100" when "01001000100100010", -- t[37154] = 4
      "0000100" when "01001000100100011", -- t[37155] = 4
      "0000100" when "01001000100100100", -- t[37156] = 4
      "0000100" when "01001000100100101", -- t[37157] = 4
      "0000100" when "01001000100100110", -- t[37158] = 4
      "0000100" when "01001000100100111", -- t[37159] = 4
      "0000100" when "01001000100101000", -- t[37160] = 4
      "0000100" when "01001000100101001", -- t[37161] = 4
      "0000100" when "01001000100101010", -- t[37162] = 4
      "0000100" when "01001000100101011", -- t[37163] = 4
      "0000100" when "01001000100101100", -- t[37164] = 4
      "0000100" when "01001000100101101", -- t[37165] = 4
      "0000100" when "01001000100101110", -- t[37166] = 4
      "0000100" when "01001000100101111", -- t[37167] = 4
      "0000100" when "01001000100110000", -- t[37168] = 4
      "0000100" when "01001000100110001", -- t[37169] = 4
      "0000100" when "01001000100110010", -- t[37170] = 4
      "0000100" when "01001000100110011", -- t[37171] = 4
      "0000100" when "01001000100110100", -- t[37172] = 4
      "0000100" when "01001000100110101", -- t[37173] = 4
      "0000100" when "01001000100110110", -- t[37174] = 4
      "0000100" when "01001000100110111", -- t[37175] = 4
      "0000100" when "01001000100111000", -- t[37176] = 4
      "0000100" when "01001000100111001", -- t[37177] = 4
      "0000100" when "01001000100111010", -- t[37178] = 4
      "0000100" when "01001000100111011", -- t[37179] = 4
      "0000100" when "01001000100111100", -- t[37180] = 4
      "0000100" when "01001000100111101", -- t[37181] = 4
      "0000100" when "01001000100111110", -- t[37182] = 4
      "0000100" when "01001000100111111", -- t[37183] = 4
      "0000100" when "01001000101000000", -- t[37184] = 4
      "0000100" when "01001000101000001", -- t[37185] = 4
      "0000100" when "01001000101000010", -- t[37186] = 4
      "0000100" when "01001000101000011", -- t[37187] = 4
      "0000100" when "01001000101000100", -- t[37188] = 4
      "0000100" when "01001000101000101", -- t[37189] = 4
      "0000100" when "01001000101000110", -- t[37190] = 4
      "0000100" when "01001000101000111", -- t[37191] = 4
      "0000100" when "01001000101001000", -- t[37192] = 4
      "0000100" when "01001000101001001", -- t[37193] = 4
      "0000100" when "01001000101001010", -- t[37194] = 4
      "0000100" when "01001000101001011", -- t[37195] = 4
      "0000100" when "01001000101001100", -- t[37196] = 4
      "0000100" when "01001000101001101", -- t[37197] = 4
      "0000100" when "01001000101001110", -- t[37198] = 4
      "0000100" when "01001000101001111", -- t[37199] = 4
      "0000100" when "01001000101010000", -- t[37200] = 4
      "0000100" when "01001000101010001", -- t[37201] = 4
      "0000100" when "01001000101010010", -- t[37202] = 4
      "0000100" when "01001000101010011", -- t[37203] = 4
      "0000100" when "01001000101010100", -- t[37204] = 4
      "0000100" when "01001000101010101", -- t[37205] = 4
      "0000100" when "01001000101010110", -- t[37206] = 4
      "0000100" when "01001000101010111", -- t[37207] = 4
      "0000100" when "01001000101011000", -- t[37208] = 4
      "0000100" when "01001000101011001", -- t[37209] = 4
      "0000100" when "01001000101011010", -- t[37210] = 4
      "0000100" when "01001000101011011", -- t[37211] = 4
      "0000100" when "01001000101011100", -- t[37212] = 4
      "0000100" when "01001000101011101", -- t[37213] = 4
      "0000100" when "01001000101011110", -- t[37214] = 4
      "0000100" when "01001000101011111", -- t[37215] = 4
      "0000100" when "01001000101100000", -- t[37216] = 4
      "0000100" when "01001000101100001", -- t[37217] = 4
      "0000100" when "01001000101100010", -- t[37218] = 4
      "0000100" when "01001000101100011", -- t[37219] = 4
      "0000100" when "01001000101100100", -- t[37220] = 4
      "0000100" when "01001000101100101", -- t[37221] = 4
      "0000100" when "01001000101100110", -- t[37222] = 4
      "0000100" when "01001000101100111", -- t[37223] = 4
      "0000100" when "01001000101101000", -- t[37224] = 4
      "0000100" when "01001000101101001", -- t[37225] = 4
      "0000100" when "01001000101101010", -- t[37226] = 4
      "0000100" when "01001000101101011", -- t[37227] = 4
      "0000100" when "01001000101101100", -- t[37228] = 4
      "0000100" when "01001000101101101", -- t[37229] = 4
      "0000100" when "01001000101101110", -- t[37230] = 4
      "0000100" when "01001000101101111", -- t[37231] = 4
      "0000100" when "01001000101110000", -- t[37232] = 4
      "0000100" when "01001000101110001", -- t[37233] = 4
      "0000100" when "01001000101110010", -- t[37234] = 4
      "0000100" when "01001000101110011", -- t[37235] = 4
      "0000100" when "01001000101110100", -- t[37236] = 4
      "0000100" when "01001000101110101", -- t[37237] = 4
      "0000100" when "01001000101110110", -- t[37238] = 4
      "0000100" when "01001000101110111", -- t[37239] = 4
      "0000100" when "01001000101111000", -- t[37240] = 4
      "0000100" when "01001000101111001", -- t[37241] = 4
      "0000100" when "01001000101111010", -- t[37242] = 4
      "0000100" when "01001000101111011", -- t[37243] = 4
      "0000100" when "01001000101111100", -- t[37244] = 4
      "0000100" when "01001000101111101", -- t[37245] = 4
      "0000100" when "01001000101111110", -- t[37246] = 4
      "0000100" when "01001000101111111", -- t[37247] = 4
      "0000100" when "01001000110000000", -- t[37248] = 4
      "0000100" when "01001000110000001", -- t[37249] = 4
      "0000100" when "01001000110000010", -- t[37250] = 4
      "0000100" when "01001000110000011", -- t[37251] = 4
      "0000100" when "01001000110000100", -- t[37252] = 4
      "0000100" when "01001000110000101", -- t[37253] = 4
      "0000100" when "01001000110000110", -- t[37254] = 4
      "0000100" when "01001000110000111", -- t[37255] = 4
      "0000100" when "01001000110001000", -- t[37256] = 4
      "0000100" when "01001000110001001", -- t[37257] = 4
      "0000100" when "01001000110001010", -- t[37258] = 4
      "0000100" when "01001000110001011", -- t[37259] = 4
      "0000100" when "01001000110001100", -- t[37260] = 4
      "0000100" when "01001000110001101", -- t[37261] = 4
      "0000100" when "01001000110001110", -- t[37262] = 4
      "0000100" when "01001000110001111", -- t[37263] = 4
      "0000100" when "01001000110010000", -- t[37264] = 4
      "0000100" when "01001000110010001", -- t[37265] = 4
      "0000100" when "01001000110010010", -- t[37266] = 4
      "0000100" when "01001000110010011", -- t[37267] = 4
      "0000100" when "01001000110010100", -- t[37268] = 4
      "0000100" when "01001000110010101", -- t[37269] = 4
      "0000100" when "01001000110010110", -- t[37270] = 4
      "0000100" when "01001000110010111", -- t[37271] = 4
      "0000100" when "01001000110011000", -- t[37272] = 4
      "0000100" when "01001000110011001", -- t[37273] = 4
      "0000100" when "01001000110011010", -- t[37274] = 4
      "0000100" when "01001000110011011", -- t[37275] = 4
      "0000100" when "01001000110011100", -- t[37276] = 4
      "0000100" when "01001000110011101", -- t[37277] = 4
      "0000100" when "01001000110011110", -- t[37278] = 4
      "0000100" when "01001000110011111", -- t[37279] = 4
      "0000100" when "01001000110100000", -- t[37280] = 4
      "0000100" when "01001000110100001", -- t[37281] = 4
      "0000100" when "01001000110100010", -- t[37282] = 4
      "0000100" when "01001000110100011", -- t[37283] = 4
      "0000100" when "01001000110100100", -- t[37284] = 4
      "0000100" when "01001000110100101", -- t[37285] = 4
      "0000100" when "01001000110100110", -- t[37286] = 4
      "0000100" when "01001000110100111", -- t[37287] = 4
      "0000100" when "01001000110101000", -- t[37288] = 4
      "0000100" when "01001000110101001", -- t[37289] = 4
      "0000100" when "01001000110101010", -- t[37290] = 4
      "0000100" when "01001000110101011", -- t[37291] = 4
      "0000100" when "01001000110101100", -- t[37292] = 4
      "0000100" when "01001000110101101", -- t[37293] = 4
      "0000100" when "01001000110101110", -- t[37294] = 4
      "0000100" when "01001000110101111", -- t[37295] = 4
      "0000100" when "01001000110110000", -- t[37296] = 4
      "0000100" when "01001000110110001", -- t[37297] = 4
      "0000100" when "01001000110110010", -- t[37298] = 4
      "0000100" when "01001000110110011", -- t[37299] = 4
      "0000100" when "01001000110110100", -- t[37300] = 4
      "0000100" when "01001000110110101", -- t[37301] = 4
      "0000100" when "01001000110110110", -- t[37302] = 4
      "0000100" when "01001000110110111", -- t[37303] = 4
      "0000100" when "01001000110111000", -- t[37304] = 4
      "0000100" when "01001000110111001", -- t[37305] = 4
      "0000100" when "01001000110111010", -- t[37306] = 4
      "0000100" when "01001000110111011", -- t[37307] = 4
      "0000100" when "01001000110111100", -- t[37308] = 4
      "0000100" when "01001000110111101", -- t[37309] = 4
      "0000100" when "01001000110111110", -- t[37310] = 4
      "0000100" when "01001000110111111", -- t[37311] = 4
      "0000100" when "01001000111000000", -- t[37312] = 4
      "0000100" when "01001000111000001", -- t[37313] = 4
      "0000100" when "01001000111000010", -- t[37314] = 4
      "0000100" when "01001000111000011", -- t[37315] = 4
      "0000100" when "01001000111000100", -- t[37316] = 4
      "0000100" when "01001000111000101", -- t[37317] = 4
      "0000100" when "01001000111000110", -- t[37318] = 4
      "0000100" when "01001000111000111", -- t[37319] = 4
      "0000100" when "01001000111001000", -- t[37320] = 4
      "0000100" when "01001000111001001", -- t[37321] = 4
      "0000100" when "01001000111001010", -- t[37322] = 4
      "0000100" when "01001000111001011", -- t[37323] = 4
      "0000100" when "01001000111001100", -- t[37324] = 4
      "0000100" when "01001000111001101", -- t[37325] = 4
      "0000100" when "01001000111001110", -- t[37326] = 4
      "0000100" when "01001000111001111", -- t[37327] = 4
      "0000100" when "01001000111010000", -- t[37328] = 4
      "0000100" when "01001000111010001", -- t[37329] = 4
      "0000100" when "01001000111010010", -- t[37330] = 4
      "0000100" when "01001000111010011", -- t[37331] = 4
      "0000100" when "01001000111010100", -- t[37332] = 4
      "0000100" when "01001000111010101", -- t[37333] = 4
      "0000100" when "01001000111010110", -- t[37334] = 4
      "0000100" when "01001000111010111", -- t[37335] = 4
      "0000100" when "01001000111011000", -- t[37336] = 4
      "0000100" when "01001000111011001", -- t[37337] = 4
      "0000100" when "01001000111011010", -- t[37338] = 4
      "0000100" when "01001000111011011", -- t[37339] = 4
      "0000100" when "01001000111011100", -- t[37340] = 4
      "0000100" when "01001000111011101", -- t[37341] = 4
      "0000100" when "01001000111011110", -- t[37342] = 4
      "0000100" when "01001000111011111", -- t[37343] = 4
      "0000100" when "01001000111100000", -- t[37344] = 4
      "0000100" when "01001000111100001", -- t[37345] = 4
      "0000100" when "01001000111100010", -- t[37346] = 4
      "0000100" when "01001000111100011", -- t[37347] = 4
      "0000100" when "01001000111100100", -- t[37348] = 4
      "0000100" when "01001000111100101", -- t[37349] = 4
      "0000100" when "01001000111100110", -- t[37350] = 4
      "0000100" when "01001000111100111", -- t[37351] = 4
      "0000100" when "01001000111101000", -- t[37352] = 4
      "0000100" when "01001000111101001", -- t[37353] = 4
      "0000100" when "01001000111101010", -- t[37354] = 4
      "0000100" when "01001000111101011", -- t[37355] = 4
      "0000100" when "01001000111101100", -- t[37356] = 4
      "0000100" when "01001000111101101", -- t[37357] = 4
      "0000100" when "01001000111101110", -- t[37358] = 4
      "0000100" when "01001000111101111", -- t[37359] = 4
      "0000100" when "01001000111110000", -- t[37360] = 4
      "0000100" when "01001000111110001", -- t[37361] = 4
      "0000100" when "01001000111110010", -- t[37362] = 4
      "0000100" when "01001000111110011", -- t[37363] = 4
      "0000100" when "01001000111110100", -- t[37364] = 4
      "0000100" when "01001000111110101", -- t[37365] = 4
      "0000100" when "01001000111110110", -- t[37366] = 4
      "0000100" when "01001000111110111", -- t[37367] = 4
      "0000100" when "01001000111111000", -- t[37368] = 4
      "0000100" when "01001000111111001", -- t[37369] = 4
      "0000100" when "01001000111111010", -- t[37370] = 4
      "0000100" when "01001000111111011", -- t[37371] = 4
      "0000100" when "01001000111111100", -- t[37372] = 4
      "0000100" when "01001000111111101", -- t[37373] = 4
      "0000100" when "01001000111111110", -- t[37374] = 4
      "0000100" when "01001000111111111", -- t[37375] = 4
      "0000100" when "01001001000000000", -- t[37376] = 4
      "0000100" when "01001001000000001", -- t[37377] = 4
      "0000100" when "01001001000000010", -- t[37378] = 4
      "0000100" when "01001001000000011", -- t[37379] = 4
      "0000100" when "01001001000000100", -- t[37380] = 4
      "0000100" when "01001001000000101", -- t[37381] = 4
      "0000100" when "01001001000000110", -- t[37382] = 4
      "0000100" when "01001001000000111", -- t[37383] = 4
      "0000100" when "01001001000001000", -- t[37384] = 4
      "0000100" when "01001001000001001", -- t[37385] = 4
      "0000100" when "01001001000001010", -- t[37386] = 4
      "0000100" when "01001001000001011", -- t[37387] = 4
      "0000100" when "01001001000001100", -- t[37388] = 4
      "0000100" when "01001001000001101", -- t[37389] = 4
      "0000100" when "01001001000001110", -- t[37390] = 4
      "0000100" when "01001001000001111", -- t[37391] = 4
      "0000100" when "01001001000010000", -- t[37392] = 4
      "0000100" when "01001001000010001", -- t[37393] = 4
      "0000100" when "01001001000010010", -- t[37394] = 4
      "0000100" when "01001001000010011", -- t[37395] = 4
      "0000100" when "01001001000010100", -- t[37396] = 4
      "0000100" when "01001001000010101", -- t[37397] = 4
      "0000100" when "01001001000010110", -- t[37398] = 4
      "0000100" when "01001001000010111", -- t[37399] = 4
      "0000100" when "01001001000011000", -- t[37400] = 4
      "0000100" when "01001001000011001", -- t[37401] = 4
      "0000100" when "01001001000011010", -- t[37402] = 4
      "0000100" when "01001001000011011", -- t[37403] = 4
      "0000100" when "01001001000011100", -- t[37404] = 4
      "0000100" when "01001001000011101", -- t[37405] = 4
      "0000100" when "01001001000011110", -- t[37406] = 4
      "0000100" when "01001001000011111", -- t[37407] = 4
      "0000100" when "01001001000100000", -- t[37408] = 4
      "0000100" when "01001001000100001", -- t[37409] = 4
      "0000100" when "01001001000100010", -- t[37410] = 4
      "0000100" when "01001001000100011", -- t[37411] = 4
      "0000100" when "01001001000100100", -- t[37412] = 4
      "0000100" when "01001001000100101", -- t[37413] = 4
      "0000100" when "01001001000100110", -- t[37414] = 4
      "0000100" when "01001001000100111", -- t[37415] = 4
      "0000100" when "01001001000101000", -- t[37416] = 4
      "0000100" when "01001001000101001", -- t[37417] = 4
      "0000100" when "01001001000101010", -- t[37418] = 4
      "0000100" when "01001001000101011", -- t[37419] = 4
      "0000100" when "01001001000101100", -- t[37420] = 4
      "0000100" when "01001001000101101", -- t[37421] = 4
      "0000100" when "01001001000101110", -- t[37422] = 4
      "0000100" when "01001001000101111", -- t[37423] = 4
      "0000100" when "01001001000110000", -- t[37424] = 4
      "0000100" when "01001001000110001", -- t[37425] = 4
      "0000100" when "01001001000110010", -- t[37426] = 4
      "0000100" when "01001001000110011", -- t[37427] = 4
      "0000100" when "01001001000110100", -- t[37428] = 4
      "0000100" when "01001001000110101", -- t[37429] = 4
      "0000100" when "01001001000110110", -- t[37430] = 4
      "0000100" when "01001001000110111", -- t[37431] = 4
      "0000100" when "01001001000111000", -- t[37432] = 4
      "0000100" when "01001001000111001", -- t[37433] = 4
      "0000100" when "01001001000111010", -- t[37434] = 4
      "0000100" when "01001001000111011", -- t[37435] = 4
      "0000100" when "01001001000111100", -- t[37436] = 4
      "0000100" when "01001001000111101", -- t[37437] = 4
      "0000100" when "01001001000111110", -- t[37438] = 4
      "0000100" when "01001001000111111", -- t[37439] = 4
      "0000100" when "01001001001000000", -- t[37440] = 4
      "0000100" when "01001001001000001", -- t[37441] = 4
      "0000100" when "01001001001000010", -- t[37442] = 4
      "0000100" when "01001001001000011", -- t[37443] = 4
      "0000100" when "01001001001000100", -- t[37444] = 4
      "0000100" when "01001001001000101", -- t[37445] = 4
      "0000100" when "01001001001000110", -- t[37446] = 4
      "0000100" when "01001001001000111", -- t[37447] = 4
      "0000100" when "01001001001001000", -- t[37448] = 4
      "0000100" when "01001001001001001", -- t[37449] = 4
      "0000100" when "01001001001001010", -- t[37450] = 4
      "0000100" when "01001001001001011", -- t[37451] = 4
      "0000100" when "01001001001001100", -- t[37452] = 4
      "0000100" when "01001001001001101", -- t[37453] = 4
      "0000100" when "01001001001001110", -- t[37454] = 4
      "0000100" when "01001001001001111", -- t[37455] = 4
      "0000100" when "01001001001010000", -- t[37456] = 4
      "0000100" when "01001001001010001", -- t[37457] = 4
      "0000100" when "01001001001010010", -- t[37458] = 4
      "0000100" when "01001001001010011", -- t[37459] = 4
      "0000100" when "01001001001010100", -- t[37460] = 4
      "0000100" when "01001001001010101", -- t[37461] = 4
      "0000100" when "01001001001010110", -- t[37462] = 4
      "0000100" when "01001001001010111", -- t[37463] = 4
      "0000100" when "01001001001011000", -- t[37464] = 4
      "0000100" when "01001001001011001", -- t[37465] = 4
      "0000100" when "01001001001011010", -- t[37466] = 4
      "0000100" when "01001001001011011", -- t[37467] = 4
      "0000100" when "01001001001011100", -- t[37468] = 4
      "0000100" when "01001001001011101", -- t[37469] = 4
      "0000100" when "01001001001011110", -- t[37470] = 4
      "0000100" when "01001001001011111", -- t[37471] = 4
      "0000100" when "01001001001100000", -- t[37472] = 4
      "0000100" when "01001001001100001", -- t[37473] = 4
      "0000100" when "01001001001100010", -- t[37474] = 4
      "0000100" when "01001001001100011", -- t[37475] = 4
      "0000100" when "01001001001100100", -- t[37476] = 4
      "0000100" when "01001001001100101", -- t[37477] = 4
      "0000100" when "01001001001100110", -- t[37478] = 4
      "0000100" when "01001001001100111", -- t[37479] = 4
      "0000100" when "01001001001101000", -- t[37480] = 4
      "0000100" when "01001001001101001", -- t[37481] = 4
      "0000100" when "01001001001101010", -- t[37482] = 4
      "0000100" when "01001001001101011", -- t[37483] = 4
      "0000100" when "01001001001101100", -- t[37484] = 4
      "0000100" when "01001001001101101", -- t[37485] = 4
      "0000100" when "01001001001101110", -- t[37486] = 4
      "0000100" when "01001001001101111", -- t[37487] = 4
      "0000100" when "01001001001110000", -- t[37488] = 4
      "0000100" when "01001001001110001", -- t[37489] = 4
      "0000100" when "01001001001110010", -- t[37490] = 4
      "0000100" when "01001001001110011", -- t[37491] = 4
      "0000100" when "01001001001110100", -- t[37492] = 4
      "0000100" when "01001001001110101", -- t[37493] = 4
      "0000100" when "01001001001110110", -- t[37494] = 4
      "0000100" when "01001001001110111", -- t[37495] = 4
      "0000100" when "01001001001111000", -- t[37496] = 4
      "0000100" when "01001001001111001", -- t[37497] = 4
      "0000100" when "01001001001111010", -- t[37498] = 4
      "0000100" when "01001001001111011", -- t[37499] = 4
      "0000100" when "01001001001111100", -- t[37500] = 4
      "0000100" when "01001001001111101", -- t[37501] = 4
      "0000100" when "01001001001111110", -- t[37502] = 4
      "0000100" when "01001001001111111", -- t[37503] = 4
      "0000100" when "01001001010000000", -- t[37504] = 4
      "0000100" when "01001001010000001", -- t[37505] = 4
      "0000100" when "01001001010000010", -- t[37506] = 4
      "0000100" when "01001001010000011", -- t[37507] = 4
      "0000100" when "01001001010000100", -- t[37508] = 4
      "0000100" when "01001001010000101", -- t[37509] = 4
      "0000100" when "01001001010000110", -- t[37510] = 4
      "0000100" when "01001001010000111", -- t[37511] = 4
      "0000100" when "01001001010001000", -- t[37512] = 4
      "0000100" when "01001001010001001", -- t[37513] = 4
      "0000100" when "01001001010001010", -- t[37514] = 4
      "0000100" when "01001001010001011", -- t[37515] = 4
      "0000100" when "01001001010001100", -- t[37516] = 4
      "0000100" when "01001001010001101", -- t[37517] = 4
      "0000100" when "01001001010001110", -- t[37518] = 4
      "0000100" when "01001001010001111", -- t[37519] = 4
      "0000100" when "01001001010010000", -- t[37520] = 4
      "0000100" when "01001001010010001", -- t[37521] = 4
      "0000100" when "01001001010010010", -- t[37522] = 4
      "0000100" when "01001001010010011", -- t[37523] = 4
      "0000100" when "01001001010010100", -- t[37524] = 4
      "0000100" when "01001001010010101", -- t[37525] = 4
      "0000100" when "01001001010010110", -- t[37526] = 4
      "0000100" when "01001001010010111", -- t[37527] = 4
      "0000100" when "01001001010011000", -- t[37528] = 4
      "0000100" when "01001001010011001", -- t[37529] = 4
      "0000100" when "01001001010011010", -- t[37530] = 4
      "0000100" when "01001001010011011", -- t[37531] = 4
      "0000100" when "01001001010011100", -- t[37532] = 4
      "0000100" when "01001001010011101", -- t[37533] = 4
      "0000100" when "01001001010011110", -- t[37534] = 4
      "0000100" when "01001001010011111", -- t[37535] = 4
      "0000100" when "01001001010100000", -- t[37536] = 4
      "0000100" when "01001001010100001", -- t[37537] = 4
      "0000100" when "01001001010100010", -- t[37538] = 4
      "0000100" when "01001001010100011", -- t[37539] = 4
      "0000100" when "01001001010100100", -- t[37540] = 4
      "0000100" when "01001001010100101", -- t[37541] = 4
      "0000100" when "01001001010100110", -- t[37542] = 4
      "0000100" when "01001001010100111", -- t[37543] = 4
      "0000100" when "01001001010101000", -- t[37544] = 4
      "0000100" when "01001001010101001", -- t[37545] = 4
      "0000100" when "01001001010101010", -- t[37546] = 4
      "0000100" when "01001001010101011", -- t[37547] = 4
      "0000100" when "01001001010101100", -- t[37548] = 4
      "0000100" when "01001001010101101", -- t[37549] = 4
      "0000100" when "01001001010101110", -- t[37550] = 4
      "0000100" when "01001001010101111", -- t[37551] = 4
      "0000100" when "01001001010110000", -- t[37552] = 4
      "0000100" when "01001001010110001", -- t[37553] = 4
      "0000100" when "01001001010110010", -- t[37554] = 4
      "0000100" when "01001001010110011", -- t[37555] = 4
      "0000100" when "01001001010110100", -- t[37556] = 4
      "0000100" when "01001001010110101", -- t[37557] = 4
      "0000100" when "01001001010110110", -- t[37558] = 4
      "0000100" when "01001001010110111", -- t[37559] = 4
      "0000100" when "01001001010111000", -- t[37560] = 4
      "0000100" when "01001001010111001", -- t[37561] = 4
      "0000100" when "01001001010111010", -- t[37562] = 4
      "0000100" when "01001001010111011", -- t[37563] = 4
      "0000100" when "01001001010111100", -- t[37564] = 4
      "0000100" when "01001001010111101", -- t[37565] = 4
      "0000100" when "01001001010111110", -- t[37566] = 4
      "0000100" when "01001001010111111", -- t[37567] = 4
      "0000100" when "01001001011000000", -- t[37568] = 4
      "0000100" when "01001001011000001", -- t[37569] = 4
      "0000100" when "01001001011000010", -- t[37570] = 4
      "0000100" when "01001001011000011", -- t[37571] = 4
      "0000100" when "01001001011000100", -- t[37572] = 4
      "0000100" when "01001001011000101", -- t[37573] = 4
      "0000100" when "01001001011000110", -- t[37574] = 4
      "0000100" when "01001001011000111", -- t[37575] = 4
      "0000100" when "01001001011001000", -- t[37576] = 4
      "0000100" when "01001001011001001", -- t[37577] = 4
      "0000100" when "01001001011001010", -- t[37578] = 4
      "0000100" when "01001001011001011", -- t[37579] = 4
      "0000100" when "01001001011001100", -- t[37580] = 4
      "0000100" when "01001001011001101", -- t[37581] = 4
      "0000100" when "01001001011001110", -- t[37582] = 4
      "0000100" when "01001001011001111", -- t[37583] = 4
      "0000100" when "01001001011010000", -- t[37584] = 4
      "0000100" when "01001001011010001", -- t[37585] = 4
      "0000100" when "01001001011010010", -- t[37586] = 4
      "0000100" when "01001001011010011", -- t[37587] = 4
      "0000100" when "01001001011010100", -- t[37588] = 4
      "0000100" when "01001001011010101", -- t[37589] = 4
      "0000100" when "01001001011010110", -- t[37590] = 4
      "0000100" when "01001001011010111", -- t[37591] = 4
      "0000100" when "01001001011011000", -- t[37592] = 4
      "0000100" when "01001001011011001", -- t[37593] = 4
      "0000100" when "01001001011011010", -- t[37594] = 4
      "0000100" when "01001001011011011", -- t[37595] = 4
      "0000100" when "01001001011011100", -- t[37596] = 4
      "0000100" when "01001001011011101", -- t[37597] = 4
      "0000100" when "01001001011011110", -- t[37598] = 4
      "0000100" when "01001001011011111", -- t[37599] = 4
      "0000100" when "01001001011100000", -- t[37600] = 4
      "0000100" when "01001001011100001", -- t[37601] = 4
      "0000100" when "01001001011100010", -- t[37602] = 4
      "0000100" when "01001001011100011", -- t[37603] = 4
      "0000100" when "01001001011100100", -- t[37604] = 4
      "0000100" when "01001001011100101", -- t[37605] = 4
      "0000100" when "01001001011100110", -- t[37606] = 4
      "0000100" when "01001001011100111", -- t[37607] = 4
      "0000100" when "01001001011101000", -- t[37608] = 4
      "0000100" when "01001001011101001", -- t[37609] = 4
      "0000100" when "01001001011101010", -- t[37610] = 4
      "0000100" when "01001001011101011", -- t[37611] = 4
      "0000100" when "01001001011101100", -- t[37612] = 4
      "0000100" when "01001001011101101", -- t[37613] = 4
      "0000100" when "01001001011101110", -- t[37614] = 4
      "0000100" when "01001001011101111", -- t[37615] = 4
      "0000100" when "01001001011110000", -- t[37616] = 4
      "0000100" when "01001001011110001", -- t[37617] = 4
      "0000100" when "01001001011110010", -- t[37618] = 4
      "0000100" when "01001001011110011", -- t[37619] = 4
      "0000100" when "01001001011110100", -- t[37620] = 4
      "0000100" when "01001001011110101", -- t[37621] = 4
      "0000100" when "01001001011110110", -- t[37622] = 4
      "0000100" when "01001001011110111", -- t[37623] = 4
      "0000100" when "01001001011111000", -- t[37624] = 4
      "0000100" when "01001001011111001", -- t[37625] = 4
      "0000100" when "01001001011111010", -- t[37626] = 4
      "0000100" when "01001001011111011", -- t[37627] = 4
      "0000100" when "01001001011111100", -- t[37628] = 4
      "0000100" when "01001001011111101", -- t[37629] = 4
      "0000100" when "01001001011111110", -- t[37630] = 4
      "0000100" when "01001001011111111", -- t[37631] = 4
      "0000100" when "01001001100000000", -- t[37632] = 4
      "0000100" when "01001001100000001", -- t[37633] = 4
      "0000100" when "01001001100000010", -- t[37634] = 4
      "0000100" when "01001001100000011", -- t[37635] = 4
      "0000100" when "01001001100000100", -- t[37636] = 4
      "0000100" when "01001001100000101", -- t[37637] = 4
      "0000100" when "01001001100000110", -- t[37638] = 4
      "0000100" when "01001001100000111", -- t[37639] = 4
      "0000100" when "01001001100001000", -- t[37640] = 4
      "0000100" when "01001001100001001", -- t[37641] = 4
      "0000100" when "01001001100001010", -- t[37642] = 4
      "0000100" when "01001001100001011", -- t[37643] = 4
      "0000100" when "01001001100001100", -- t[37644] = 4
      "0000100" when "01001001100001101", -- t[37645] = 4
      "0000100" when "01001001100001110", -- t[37646] = 4
      "0000100" when "01001001100001111", -- t[37647] = 4
      "0000100" when "01001001100010000", -- t[37648] = 4
      "0000100" when "01001001100010001", -- t[37649] = 4
      "0000100" when "01001001100010010", -- t[37650] = 4
      "0000100" when "01001001100010011", -- t[37651] = 4
      "0000100" when "01001001100010100", -- t[37652] = 4
      "0000100" when "01001001100010101", -- t[37653] = 4
      "0000100" when "01001001100010110", -- t[37654] = 4
      "0000100" when "01001001100010111", -- t[37655] = 4
      "0000100" when "01001001100011000", -- t[37656] = 4
      "0000100" when "01001001100011001", -- t[37657] = 4
      "0000100" when "01001001100011010", -- t[37658] = 4
      "0000100" when "01001001100011011", -- t[37659] = 4
      "0000100" when "01001001100011100", -- t[37660] = 4
      "0000100" when "01001001100011101", -- t[37661] = 4
      "0000100" when "01001001100011110", -- t[37662] = 4
      "0000100" when "01001001100011111", -- t[37663] = 4
      "0000100" when "01001001100100000", -- t[37664] = 4
      "0000100" when "01001001100100001", -- t[37665] = 4
      "0000100" when "01001001100100010", -- t[37666] = 4
      "0000100" when "01001001100100011", -- t[37667] = 4
      "0000100" when "01001001100100100", -- t[37668] = 4
      "0000100" when "01001001100100101", -- t[37669] = 4
      "0000100" when "01001001100100110", -- t[37670] = 4
      "0000100" when "01001001100100111", -- t[37671] = 4
      "0000100" when "01001001100101000", -- t[37672] = 4
      "0000100" when "01001001100101001", -- t[37673] = 4
      "0000100" when "01001001100101010", -- t[37674] = 4
      "0000100" when "01001001100101011", -- t[37675] = 4
      "0000100" when "01001001100101100", -- t[37676] = 4
      "0000100" when "01001001100101101", -- t[37677] = 4
      "0000100" when "01001001100101110", -- t[37678] = 4
      "0000100" when "01001001100101111", -- t[37679] = 4
      "0000100" when "01001001100110000", -- t[37680] = 4
      "0000100" when "01001001100110001", -- t[37681] = 4
      "0000100" when "01001001100110010", -- t[37682] = 4
      "0000100" when "01001001100110011", -- t[37683] = 4
      "0000100" when "01001001100110100", -- t[37684] = 4
      "0000100" when "01001001100110101", -- t[37685] = 4
      "0000100" when "01001001100110110", -- t[37686] = 4
      "0000100" when "01001001100110111", -- t[37687] = 4
      "0000100" when "01001001100111000", -- t[37688] = 4
      "0000100" when "01001001100111001", -- t[37689] = 4
      "0000100" when "01001001100111010", -- t[37690] = 4
      "0000100" when "01001001100111011", -- t[37691] = 4
      "0000100" when "01001001100111100", -- t[37692] = 4
      "0000100" when "01001001100111101", -- t[37693] = 4
      "0000100" when "01001001100111110", -- t[37694] = 4
      "0000100" when "01001001100111111", -- t[37695] = 4
      "0000100" when "01001001101000000", -- t[37696] = 4
      "0000100" when "01001001101000001", -- t[37697] = 4
      "0000100" when "01001001101000010", -- t[37698] = 4
      "0000100" when "01001001101000011", -- t[37699] = 4
      "0000100" when "01001001101000100", -- t[37700] = 4
      "0000100" when "01001001101000101", -- t[37701] = 4
      "0000100" when "01001001101000110", -- t[37702] = 4
      "0000100" when "01001001101000111", -- t[37703] = 4
      "0000100" when "01001001101001000", -- t[37704] = 4
      "0000100" when "01001001101001001", -- t[37705] = 4
      "0000100" when "01001001101001010", -- t[37706] = 4
      "0000100" when "01001001101001011", -- t[37707] = 4
      "0000100" when "01001001101001100", -- t[37708] = 4
      "0000100" when "01001001101001101", -- t[37709] = 4
      "0000100" when "01001001101001110", -- t[37710] = 4
      "0000100" when "01001001101001111", -- t[37711] = 4
      "0000100" when "01001001101010000", -- t[37712] = 4
      "0000100" when "01001001101010001", -- t[37713] = 4
      "0000100" when "01001001101010010", -- t[37714] = 4
      "0000100" when "01001001101010011", -- t[37715] = 4
      "0000100" when "01001001101010100", -- t[37716] = 4
      "0000100" when "01001001101010101", -- t[37717] = 4
      "0000100" when "01001001101010110", -- t[37718] = 4
      "0000100" when "01001001101010111", -- t[37719] = 4
      "0000100" when "01001001101011000", -- t[37720] = 4
      "0000100" when "01001001101011001", -- t[37721] = 4
      "0000100" when "01001001101011010", -- t[37722] = 4
      "0000100" when "01001001101011011", -- t[37723] = 4
      "0000100" when "01001001101011100", -- t[37724] = 4
      "0000100" when "01001001101011101", -- t[37725] = 4
      "0000100" when "01001001101011110", -- t[37726] = 4
      "0000100" when "01001001101011111", -- t[37727] = 4
      "0000100" when "01001001101100000", -- t[37728] = 4
      "0000100" when "01001001101100001", -- t[37729] = 4
      "0000100" when "01001001101100010", -- t[37730] = 4
      "0000100" when "01001001101100011", -- t[37731] = 4
      "0000100" when "01001001101100100", -- t[37732] = 4
      "0000100" when "01001001101100101", -- t[37733] = 4
      "0000100" when "01001001101100110", -- t[37734] = 4
      "0000100" when "01001001101100111", -- t[37735] = 4
      "0000100" when "01001001101101000", -- t[37736] = 4
      "0000100" when "01001001101101001", -- t[37737] = 4
      "0000100" when "01001001101101010", -- t[37738] = 4
      "0000100" when "01001001101101011", -- t[37739] = 4
      "0000100" when "01001001101101100", -- t[37740] = 4
      "0000100" when "01001001101101101", -- t[37741] = 4
      "0000100" when "01001001101101110", -- t[37742] = 4
      "0000100" when "01001001101101111", -- t[37743] = 4
      "0000100" when "01001001101110000", -- t[37744] = 4
      "0000100" when "01001001101110001", -- t[37745] = 4
      "0000100" when "01001001101110010", -- t[37746] = 4
      "0000100" when "01001001101110011", -- t[37747] = 4
      "0000100" when "01001001101110100", -- t[37748] = 4
      "0000100" when "01001001101110101", -- t[37749] = 4
      "0000100" when "01001001101110110", -- t[37750] = 4
      "0000100" when "01001001101110111", -- t[37751] = 4
      "0000100" when "01001001101111000", -- t[37752] = 4
      "0000100" when "01001001101111001", -- t[37753] = 4
      "0000100" when "01001001101111010", -- t[37754] = 4
      "0000100" when "01001001101111011", -- t[37755] = 4
      "0000100" when "01001001101111100", -- t[37756] = 4
      "0000100" when "01001001101111101", -- t[37757] = 4
      "0000100" when "01001001101111110", -- t[37758] = 4
      "0000100" when "01001001101111111", -- t[37759] = 4
      "0000100" when "01001001110000000", -- t[37760] = 4
      "0000100" when "01001001110000001", -- t[37761] = 4
      "0000100" when "01001001110000010", -- t[37762] = 4
      "0000100" when "01001001110000011", -- t[37763] = 4
      "0000100" when "01001001110000100", -- t[37764] = 4
      "0000100" when "01001001110000101", -- t[37765] = 4
      "0000100" when "01001001110000110", -- t[37766] = 4
      "0000100" when "01001001110000111", -- t[37767] = 4
      "0000100" when "01001001110001000", -- t[37768] = 4
      "0000100" when "01001001110001001", -- t[37769] = 4
      "0000100" when "01001001110001010", -- t[37770] = 4
      "0000100" when "01001001110001011", -- t[37771] = 4
      "0000100" when "01001001110001100", -- t[37772] = 4
      "0000100" when "01001001110001101", -- t[37773] = 4
      "0000100" when "01001001110001110", -- t[37774] = 4
      "0000100" when "01001001110001111", -- t[37775] = 4
      "0000100" when "01001001110010000", -- t[37776] = 4
      "0000100" when "01001001110010001", -- t[37777] = 4
      "0000100" when "01001001110010010", -- t[37778] = 4
      "0000100" when "01001001110010011", -- t[37779] = 4
      "0000100" when "01001001110010100", -- t[37780] = 4
      "0000100" when "01001001110010101", -- t[37781] = 4
      "0000100" when "01001001110010110", -- t[37782] = 4
      "0000100" when "01001001110010111", -- t[37783] = 4
      "0000100" when "01001001110011000", -- t[37784] = 4
      "0000100" when "01001001110011001", -- t[37785] = 4
      "0000100" when "01001001110011010", -- t[37786] = 4
      "0000100" when "01001001110011011", -- t[37787] = 4
      "0000100" when "01001001110011100", -- t[37788] = 4
      "0000100" when "01001001110011101", -- t[37789] = 4
      "0000100" when "01001001110011110", -- t[37790] = 4
      "0000100" when "01001001110011111", -- t[37791] = 4
      "0000100" when "01001001110100000", -- t[37792] = 4
      "0000100" when "01001001110100001", -- t[37793] = 4
      "0000100" when "01001001110100010", -- t[37794] = 4
      "0000100" when "01001001110100011", -- t[37795] = 4
      "0000100" when "01001001110100100", -- t[37796] = 4
      "0000100" when "01001001110100101", -- t[37797] = 4
      "0000100" when "01001001110100110", -- t[37798] = 4
      "0000100" when "01001001110100111", -- t[37799] = 4
      "0000100" when "01001001110101000", -- t[37800] = 4
      "0000100" when "01001001110101001", -- t[37801] = 4
      "0000100" when "01001001110101010", -- t[37802] = 4
      "0000100" when "01001001110101011", -- t[37803] = 4
      "0000100" when "01001001110101100", -- t[37804] = 4
      "0000100" when "01001001110101101", -- t[37805] = 4
      "0000100" when "01001001110101110", -- t[37806] = 4
      "0000100" when "01001001110101111", -- t[37807] = 4
      "0000100" when "01001001110110000", -- t[37808] = 4
      "0000100" when "01001001110110001", -- t[37809] = 4
      "0000100" when "01001001110110010", -- t[37810] = 4
      "0000100" when "01001001110110011", -- t[37811] = 4
      "0000100" when "01001001110110100", -- t[37812] = 4
      "0000100" when "01001001110110101", -- t[37813] = 4
      "0000100" when "01001001110110110", -- t[37814] = 4
      "0000100" when "01001001110110111", -- t[37815] = 4
      "0000100" when "01001001110111000", -- t[37816] = 4
      "0000100" when "01001001110111001", -- t[37817] = 4
      "0000100" when "01001001110111010", -- t[37818] = 4
      "0000100" when "01001001110111011", -- t[37819] = 4
      "0000100" when "01001001110111100", -- t[37820] = 4
      "0000100" when "01001001110111101", -- t[37821] = 4
      "0000100" when "01001001110111110", -- t[37822] = 4
      "0000100" when "01001001110111111", -- t[37823] = 4
      "0000100" when "01001001111000000", -- t[37824] = 4
      "0000100" when "01001001111000001", -- t[37825] = 4
      "0000100" when "01001001111000010", -- t[37826] = 4
      "0000100" when "01001001111000011", -- t[37827] = 4
      "0000100" when "01001001111000100", -- t[37828] = 4
      "0000100" when "01001001111000101", -- t[37829] = 4
      "0000100" when "01001001111000110", -- t[37830] = 4
      "0000100" when "01001001111000111", -- t[37831] = 4
      "0000100" when "01001001111001000", -- t[37832] = 4
      "0000100" when "01001001111001001", -- t[37833] = 4
      "0000100" when "01001001111001010", -- t[37834] = 4
      "0000100" when "01001001111001011", -- t[37835] = 4
      "0000100" when "01001001111001100", -- t[37836] = 4
      "0000100" when "01001001111001101", -- t[37837] = 4
      "0000100" when "01001001111001110", -- t[37838] = 4
      "0000100" when "01001001111001111", -- t[37839] = 4
      "0000100" when "01001001111010000", -- t[37840] = 4
      "0000100" when "01001001111010001", -- t[37841] = 4
      "0000100" when "01001001111010010", -- t[37842] = 4
      "0000100" when "01001001111010011", -- t[37843] = 4
      "0000100" when "01001001111010100", -- t[37844] = 4
      "0000100" when "01001001111010101", -- t[37845] = 4
      "0000100" when "01001001111010110", -- t[37846] = 4
      "0000100" when "01001001111010111", -- t[37847] = 4
      "0000100" when "01001001111011000", -- t[37848] = 4
      "0000100" when "01001001111011001", -- t[37849] = 4
      "0000100" when "01001001111011010", -- t[37850] = 4
      "0000100" when "01001001111011011", -- t[37851] = 4
      "0000100" when "01001001111011100", -- t[37852] = 4
      "0000100" when "01001001111011101", -- t[37853] = 4
      "0000100" when "01001001111011110", -- t[37854] = 4
      "0000100" when "01001001111011111", -- t[37855] = 4
      "0000100" when "01001001111100000", -- t[37856] = 4
      "0000100" when "01001001111100001", -- t[37857] = 4
      "0000100" when "01001001111100010", -- t[37858] = 4
      "0000100" when "01001001111100011", -- t[37859] = 4
      "0000100" when "01001001111100100", -- t[37860] = 4
      "0000100" when "01001001111100101", -- t[37861] = 4
      "0000100" when "01001001111100110", -- t[37862] = 4
      "0000100" when "01001001111100111", -- t[37863] = 4
      "0000100" when "01001001111101000", -- t[37864] = 4
      "0000100" when "01001001111101001", -- t[37865] = 4
      "0000100" when "01001001111101010", -- t[37866] = 4
      "0000100" when "01001001111101011", -- t[37867] = 4
      "0000100" when "01001001111101100", -- t[37868] = 4
      "0000100" when "01001001111101101", -- t[37869] = 4
      "0000100" when "01001001111101110", -- t[37870] = 4
      "0000100" when "01001001111101111", -- t[37871] = 4
      "0000100" when "01001001111110000", -- t[37872] = 4
      "0000100" when "01001001111110001", -- t[37873] = 4
      "0000100" when "01001001111110010", -- t[37874] = 4
      "0000100" when "01001001111110011", -- t[37875] = 4
      "0000100" when "01001001111110100", -- t[37876] = 4
      "0000100" when "01001001111110101", -- t[37877] = 4
      "0000100" when "01001001111110110", -- t[37878] = 4
      "0000100" when "01001001111110111", -- t[37879] = 4
      "0000100" when "01001001111111000", -- t[37880] = 4
      "0000100" when "01001001111111001", -- t[37881] = 4
      "0000100" when "01001001111111010", -- t[37882] = 4
      "0000100" when "01001001111111011", -- t[37883] = 4
      "0000100" when "01001001111111100", -- t[37884] = 4
      "0000100" when "01001001111111101", -- t[37885] = 4
      "0000100" when "01001001111111110", -- t[37886] = 4
      "0000100" when "01001001111111111", -- t[37887] = 4
      "0000100" when "01001010000000000", -- t[37888] = 4
      "0000100" when "01001010000000001", -- t[37889] = 4
      "0000100" when "01001010000000010", -- t[37890] = 4
      "0000100" when "01001010000000011", -- t[37891] = 4
      "0000100" when "01001010000000100", -- t[37892] = 4
      "0000100" when "01001010000000101", -- t[37893] = 4
      "0000100" when "01001010000000110", -- t[37894] = 4
      "0000100" when "01001010000000111", -- t[37895] = 4
      "0000100" when "01001010000001000", -- t[37896] = 4
      "0000100" when "01001010000001001", -- t[37897] = 4
      "0000100" when "01001010000001010", -- t[37898] = 4
      "0000100" when "01001010000001011", -- t[37899] = 4
      "0000100" when "01001010000001100", -- t[37900] = 4
      "0000100" when "01001010000001101", -- t[37901] = 4
      "0000100" when "01001010000001110", -- t[37902] = 4
      "0000100" when "01001010000001111", -- t[37903] = 4
      "0000100" when "01001010000010000", -- t[37904] = 4
      "0000100" when "01001010000010001", -- t[37905] = 4
      "0000100" when "01001010000010010", -- t[37906] = 4
      "0000100" when "01001010000010011", -- t[37907] = 4
      "0000100" when "01001010000010100", -- t[37908] = 4
      "0000100" when "01001010000010101", -- t[37909] = 4
      "0000100" when "01001010000010110", -- t[37910] = 4
      "0000100" when "01001010000010111", -- t[37911] = 4
      "0000100" when "01001010000011000", -- t[37912] = 4
      "0000100" when "01001010000011001", -- t[37913] = 4
      "0000100" when "01001010000011010", -- t[37914] = 4
      "0000100" when "01001010000011011", -- t[37915] = 4
      "0000100" when "01001010000011100", -- t[37916] = 4
      "0000100" when "01001010000011101", -- t[37917] = 4
      "0000100" when "01001010000011110", -- t[37918] = 4
      "0000100" when "01001010000011111", -- t[37919] = 4
      "0000100" when "01001010000100000", -- t[37920] = 4
      "0000100" when "01001010000100001", -- t[37921] = 4
      "0000100" when "01001010000100010", -- t[37922] = 4
      "0000100" when "01001010000100011", -- t[37923] = 4
      "0000100" when "01001010000100100", -- t[37924] = 4
      "0000100" when "01001010000100101", -- t[37925] = 4
      "0000100" when "01001010000100110", -- t[37926] = 4
      "0000100" when "01001010000100111", -- t[37927] = 4
      "0000100" when "01001010000101000", -- t[37928] = 4
      "0000100" when "01001010000101001", -- t[37929] = 4
      "0000100" when "01001010000101010", -- t[37930] = 4
      "0000100" when "01001010000101011", -- t[37931] = 4
      "0000100" when "01001010000101100", -- t[37932] = 4
      "0000100" when "01001010000101101", -- t[37933] = 4
      "0000100" when "01001010000101110", -- t[37934] = 4
      "0000100" when "01001010000101111", -- t[37935] = 4
      "0000100" when "01001010000110000", -- t[37936] = 4
      "0000100" when "01001010000110001", -- t[37937] = 4
      "0000100" when "01001010000110010", -- t[37938] = 4
      "0000100" when "01001010000110011", -- t[37939] = 4
      "0000100" when "01001010000110100", -- t[37940] = 4
      "0000100" when "01001010000110101", -- t[37941] = 4
      "0000100" when "01001010000110110", -- t[37942] = 4
      "0000100" when "01001010000110111", -- t[37943] = 4
      "0000100" when "01001010000111000", -- t[37944] = 4
      "0000100" when "01001010000111001", -- t[37945] = 4
      "0000100" when "01001010000111010", -- t[37946] = 4
      "0000100" when "01001010000111011", -- t[37947] = 4
      "0000100" when "01001010000111100", -- t[37948] = 4
      "0000100" when "01001010000111101", -- t[37949] = 4
      "0000100" when "01001010000111110", -- t[37950] = 4
      "0000100" when "01001010000111111", -- t[37951] = 4
      "0000100" when "01001010001000000", -- t[37952] = 4
      "0000100" when "01001010001000001", -- t[37953] = 4
      "0000100" when "01001010001000010", -- t[37954] = 4
      "0000100" when "01001010001000011", -- t[37955] = 4
      "0000100" when "01001010001000100", -- t[37956] = 4
      "0000100" when "01001010001000101", -- t[37957] = 4
      "0000100" when "01001010001000110", -- t[37958] = 4
      "0000100" when "01001010001000111", -- t[37959] = 4
      "0000100" when "01001010001001000", -- t[37960] = 4
      "0000100" when "01001010001001001", -- t[37961] = 4
      "0000100" when "01001010001001010", -- t[37962] = 4
      "0000100" when "01001010001001011", -- t[37963] = 4
      "0000100" when "01001010001001100", -- t[37964] = 4
      "0000100" when "01001010001001101", -- t[37965] = 4
      "0000100" when "01001010001001110", -- t[37966] = 4
      "0000100" when "01001010001001111", -- t[37967] = 4
      "0000100" when "01001010001010000", -- t[37968] = 4
      "0000100" when "01001010001010001", -- t[37969] = 4
      "0000100" when "01001010001010010", -- t[37970] = 4
      "0000100" when "01001010001010011", -- t[37971] = 4
      "0000100" when "01001010001010100", -- t[37972] = 4
      "0000100" when "01001010001010101", -- t[37973] = 4
      "0000100" when "01001010001010110", -- t[37974] = 4
      "0000100" when "01001010001010111", -- t[37975] = 4
      "0000100" when "01001010001011000", -- t[37976] = 4
      "0000100" when "01001010001011001", -- t[37977] = 4
      "0000100" when "01001010001011010", -- t[37978] = 4
      "0000100" when "01001010001011011", -- t[37979] = 4
      "0000100" when "01001010001011100", -- t[37980] = 4
      "0000100" when "01001010001011101", -- t[37981] = 4
      "0000100" when "01001010001011110", -- t[37982] = 4
      "0000100" when "01001010001011111", -- t[37983] = 4
      "0000100" when "01001010001100000", -- t[37984] = 4
      "0000100" when "01001010001100001", -- t[37985] = 4
      "0000100" when "01001010001100010", -- t[37986] = 4
      "0000100" when "01001010001100011", -- t[37987] = 4
      "0000100" when "01001010001100100", -- t[37988] = 4
      "0000100" when "01001010001100101", -- t[37989] = 4
      "0000100" when "01001010001100110", -- t[37990] = 4
      "0000100" when "01001010001100111", -- t[37991] = 4
      "0000100" when "01001010001101000", -- t[37992] = 4
      "0000100" when "01001010001101001", -- t[37993] = 4
      "0000100" when "01001010001101010", -- t[37994] = 4
      "0000100" when "01001010001101011", -- t[37995] = 4
      "0000100" when "01001010001101100", -- t[37996] = 4
      "0000100" when "01001010001101101", -- t[37997] = 4
      "0000100" when "01001010001101110", -- t[37998] = 4
      "0000100" when "01001010001101111", -- t[37999] = 4
      "0000100" when "01001010001110000", -- t[38000] = 4
      "0000100" when "01001010001110001", -- t[38001] = 4
      "0000100" when "01001010001110010", -- t[38002] = 4
      "0000100" when "01001010001110011", -- t[38003] = 4
      "0000100" when "01001010001110100", -- t[38004] = 4
      "0000100" when "01001010001110101", -- t[38005] = 4
      "0000100" when "01001010001110110", -- t[38006] = 4
      "0000100" when "01001010001110111", -- t[38007] = 4
      "0000100" when "01001010001111000", -- t[38008] = 4
      "0000100" when "01001010001111001", -- t[38009] = 4
      "0000100" when "01001010001111010", -- t[38010] = 4
      "0000100" when "01001010001111011", -- t[38011] = 4
      "0000100" when "01001010001111100", -- t[38012] = 4
      "0000100" when "01001010001111101", -- t[38013] = 4
      "0000100" when "01001010001111110", -- t[38014] = 4
      "0000100" when "01001010001111111", -- t[38015] = 4
      "0000100" when "01001010010000000", -- t[38016] = 4
      "0000100" when "01001010010000001", -- t[38017] = 4
      "0000100" when "01001010010000010", -- t[38018] = 4
      "0000101" when "01001010010000011", -- t[38019] = 5
      "0000101" when "01001010010000100", -- t[38020] = 5
      "0000101" when "01001010010000101", -- t[38021] = 5
      "0000101" when "01001010010000110", -- t[38022] = 5
      "0000101" when "01001010010000111", -- t[38023] = 5
      "0000101" when "01001010010001000", -- t[38024] = 5
      "0000101" when "01001010010001001", -- t[38025] = 5
      "0000101" when "01001010010001010", -- t[38026] = 5
      "0000101" when "01001010010001011", -- t[38027] = 5
      "0000101" when "01001010010001100", -- t[38028] = 5
      "0000101" when "01001010010001101", -- t[38029] = 5
      "0000101" when "01001010010001110", -- t[38030] = 5
      "0000101" when "01001010010001111", -- t[38031] = 5
      "0000101" when "01001010010010000", -- t[38032] = 5
      "0000101" when "01001010010010001", -- t[38033] = 5
      "0000101" when "01001010010010010", -- t[38034] = 5
      "0000101" when "01001010010010011", -- t[38035] = 5
      "0000101" when "01001010010010100", -- t[38036] = 5
      "0000101" when "01001010010010101", -- t[38037] = 5
      "0000101" when "01001010010010110", -- t[38038] = 5
      "0000101" when "01001010010010111", -- t[38039] = 5
      "0000101" when "01001010010011000", -- t[38040] = 5
      "0000101" when "01001010010011001", -- t[38041] = 5
      "0000101" when "01001010010011010", -- t[38042] = 5
      "0000101" when "01001010010011011", -- t[38043] = 5
      "0000101" when "01001010010011100", -- t[38044] = 5
      "0000101" when "01001010010011101", -- t[38045] = 5
      "0000101" when "01001010010011110", -- t[38046] = 5
      "0000101" when "01001010010011111", -- t[38047] = 5
      "0000101" when "01001010010100000", -- t[38048] = 5
      "0000101" when "01001010010100001", -- t[38049] = 5
      "0000101" when "01001010010100010", -- t[38050] = 5
      "0000101" when "01001010010100011", -- t[38051] = 5
      "0000101" when "01001010010100100", -- t[38052] = 5
      "0000101" when "01001010010100101", -- t[38053] = 5
      "0000101" when "01001010010100110", -- t[38054] = 5
      "0000101" when "01001010010100111", -- t[38055] = 5
      "0000101" when "01001010010101000", -- t[38056] = 5
      "0000101" when "01001010010101001", -- t[38057] = 5
      "0000101" when "01001010010101010", -- t[38058] = 5
      "0000101" when "01001010010101011", -- t[38059] = 5
      "0000101" when "01001010010101100", -- t[38060] = 5
      "0000101" when "01001010010101101", -- t[38061] = 5
      "0000101" when "01001010010101110", -- t[38062] = 5
      "0000101" when "01001010010101111", -- t[38063] = 5
      "0000101" when "01001010010110000", -- t[38064] = 5
      "0000101" when "01001010010110001", -- t[38065] = 5
      "0000101" when "01001010010110010", -- t[38066] = 5
      "0000101" when "01001010010110011", -- t[38067] = 5
      "0000101" when "01001010010110100", -- t[38068] = 5
      "0000101" when "01001010010110101", -- t[38069] = 5
      "0000101" when "01001010010110110", -- t[38070] = 5
      "0000101" when "01001010010110111", -- t[38071] = 5
      "0000101" when "01001010010111000", -- t[38072] = 5
      "0000101" when "01001010010111001", -- t[38073] = 5
      "0000101" when "01001010010111010", -- t[38074] = 5
      "0000101" when "01001010010111011", -- t[38075] = 5
      "0000101" when "01001010010111100", -- t[38076] = 5
      "0000101" when "01001010010111101", -- t[38077] = 5
      "0000101" when "01001010010111110", -- t[38078] = 5
      "0000101" when "01001010010111111", -- t[38079] = 5
      "0000101" when "01001010011000000", -- t[38080] = 5
      "0000101" when "01001010011000001", -- t[38081] = 5
      "0000101" when "01001010011000010", -- t[38082] = 5
      "0000101" when "01001010011000011", -- t[38083] = 5
      "0000101" when "01001010011000100", -- t[38084] = 5
      "0000101" when "01001010011000101", -- t[38085] = 5
      "0000101" when "01001010011000110", -- t[38086] = 5
      "0000101" when "01001010011000111", -- t[38087] = 5
      "0000101" when "01001010011001000", -- t[38088] = 5
      "0000101" when "01001010011001001", -- t[38089] = 5
      "0000101" when "01001010011001010", -- t[38090] = 5
      "0000101" when "01001010011001011", -- t[38091] = 5
      "0000101" when "01001010011001100", -- t[38092] = 5
      "0000101" when "01001010011001101", -- t[38093] = 5
      "0000101" when "01001010011001110", -- t[38094] = 5
      "0000101" when "01001010011001111", -- t[38095] = 5
      "0000101" when "01001010011010000", -- t[38096] = 5
      "0000101" when "01001010011010001", -- t[38097] = 5
      "0000101" when "01001010011010010", -- t[38098] = 5
      "0000101" when "01001010011010011", -- t[38099] = 5
      "0000101" when "01001010011010100", -- t[38100] = 5
      "0000101" when "01001010011010101", -- t[38101] = 5
      "0000101" when "01001010011010110", -- t[38102] = 5
      "0000101" when "01001010011010111", -- t[38103] = 5
      "0000101" when "01001010011011000", -- t[38104] = 5
      "0000101" when "01001010011011001", -- t[38105] = 5
      "0000101" when "01001010011011010", -- t[38106] = 5
      "0000101" when "01001010011011011", -- t[38107] = 5
      "0000101" when "01001010011011100", -- t[38108] = 5
      "0000101" when "01001010011011101", -- t[38109] = 5
      "0000101" when "01001010011011110", -- t[38110] = 5
      "0000101" when "01001010011011111", -- t[38111] = 5
      "0000101" when "01001010011100000", -- t[38112] = 5
      "0000101" when "01001010011100001", -- t[38113] = 5
      "0000101" when "01001010011100010", -- t[38114] = 5
      "0000101" when "01001010011100011", -- t[38115] = 5
      "0000101" when "01001010011100100", -- t[38116] = 5
      "0000101" when "01001010011100101", -- t[38117] = 5
      "0000101" when "01001010011100110", -- t[38118] = 5
      "0000101" when "01001010011100111", -- t[38119] = 5
      "0000101" when "01001010011101000", -- t[38120] = 5
      "0000101" when "01001010011101001", -- t[38121] = 5
      "0000101" when "01001010011101010", -- t[38122] = 5
      "0000101" when "01001010011101011", -- t[38123] = 5
      "0000101" when "01001010011101100", -- t[38124] = 5
      "0000101" when "01001010011101101", -- t[38125] = 5
      "0000101" when "01001010011101110", -- t[38126] = 5
      "0000101" when "01001010011101111", -- t[38127] = 5
      "0000101" when "01001010011110000", -- t[38128] = 5
      "0000101" when "01001010011110001", -- t[38129] = 5
      "0000101" when "01001010011110010", -- t[38130] = 5
      "0000101" when "01001010011110011", -- t[38131] = 5
      "0000101" when "01001010011110100", -- t[38132] = 5
      "0000101" when "01001010011110101", -- t[38133] = 5
      "0000101" when "01001010011110110", -- t[38134] = 5
      "0000101" when "01001010011110111", -- t[38135] = 5
      "0000101" when "01001010011111000", -- t[38136] = 5
      "0000101" when "01001010011111001", -- t[38137] = 5
      "0000101" when "01001010011111010", -- t[38138] = 5
      "0000101" when "01001010011111011", -- t[38139] = 5
      "0000101" when "01001010011111100", -- t[38140] = 5
      "0000101" when "01001010011111101", -- t[38141] = 5
      "0000101" when "01001010011111110", -- t[38142] = 5
      "0000101" when "01001010011111111", -- t[38143] = 5
      "0000101" when "01001010100000000", -- t[38144] = 5
      "0000101" when "01001010100000001", -- t[38145] = 5
      "0000101" when "01001010100000010", -- t[38146] = 5
      "0000101" when "01001010100000011", -- t[38147] = 5
      "0000101" when "01001010100000100", -- t[38148] = 5
      "0000101" when "01001010100000101", -- t[38149] = 5
      "0000101" when "01001010100000110", -- t[38150] = 5
      "0000101" when "01001010100000111", -- t[38151] = 5
      "0000101" when "01001010100001000", -- t[38152] = 5
      "0000101" when "01001010100001001", -- t[38153] = 5
      "0000101" when "01001010100001010", -- t[38154] = 5
      "0000101" when "01001010100001011", -- t[38155] = 5
      "0000101" when "01001010100001100", -- t[38156] = 5
      "0000101" when "01001010100001101", -- t[38157] = 5
      "0000101" when "01001010100001110", -- t[38158] = 5
      "0000101" when "01001010100001111", -- t[38159] = 5
      "0000101" when "01001010100010000", -- t[38160] = 5
      "0000101" when "01001010100010001", -- t[38161] = 5
      "0000101" when "01001010100010010", -- t[38162] = 5
      "0000101" when "01001010100010011", -- t[38163] = 5
      "0000101" when "01001010100010100", -- t[38164] = 5
      "0000101" when "01001010100010101", -- t[38165] = 5
      "0000101" when "01001010100010110", -- t[38166] = 5
      "0000101" when "01001010100010111", -- t[38167] = 5
      "0000101" when "01001010100011000", -- t[38168] = 5
      "0000101" when "01001010100011001", -- t[38169] = 5
      "0000101" when "01001010100011010", -- t[38170] = 5
      "0000101" when "01001010100011011", -- t[38171] = 5
      "0000101" when "01001010100011100", -- t[38172] = 5
      "0000101" when "01001010100011101", -- t[38173] = 5
      "0000101" when "01001010100011110", -- t[38174] = 5
      "0000101" when "01001010100011111", -- t[38175] = 5
      "0000101" when "01001010100100000", -- t[38176] = 5
      "0000101" when "01001010100100001", -- t[38177] = 5
      "0000101" when "01001010100100010", -- t[38178] = 5
      "0000101" when "01001010100100011", -- t[38179] = 5
      "0000101" when "01001010100100100", -- t[38180] = 5
      "0000101" when "01001010100100101", -- t[38181] = 5
      "0000101" when "01001010100100110", -- t[38182] = 5
      "0000101" when "01001010100100111", -- t[38183] = 5
      "0000101" when "01001010100101000", -- t[38184] = 5
      "0000101" when "01001010100101001", -- t[38185] = 5
      "0000101" when "01001010100101010", -- t[38186] = 5
      "0000101" when "01001010100101011", -- t[38187] = 5
      "0000101" when "01001010100101100", -- t[38188] = 5
      "0000101" when "01001010100101101", -- t[38189] = 5
      "0000101" when "01001010100101110", -- t[38190] = 5
      "0000101" when "01001010100101111", -- t[38191] = 5
      "0000101" when "01001010100110000", -- t[38192] = 5
      "0000101" when "01001010100110001", -- t[38193] = 5
      "0000101" when "01001010100110010", -- t[38194] = 5
      "0000101" when "01001010100110011", -- t[38195] = 5
      "0000101" when "01001010100110100", -- t[38196] = 5
      "0000101" when "01001010100110101", -- t[38197] = 5
      "0000101" when "01001010100110110", -- t[38198] = 5
      "0000101" when "01001010100110111", -- t[38199] = 5
      "0000101" when "01001010100111000", -- t[38200] = 5
      "0000101" when "01001010100111001", -- t[38201] = 5
      "0000101" when "01001010100111010", -- t[38202] = 5
      "0000101" when "01001010100111011", -- t[38203] = 5
      "0000101" when "01001010100111100", -- t[38204] = 5
      "0000101" when "01001010100111101", -- t[38205] = 5
      "0000101" when "01001010100111110", -- t[38206] = 5
      "0000101" when "01001010100111111", -- t[38207] = 5
      "0000101" when "01001010101000000", -- t[38208] = 5
      "0000101" when "01001010101000001", -- t[38209] = 5
      "0000101" when "01001010101000010", -- t[38210] = 5
      "0000101" when "01001010101000011", -- t[38211] = 5
      "0000101" when "01001010101000100", -- t[38212] = 5
      "0000101" when "01001010101000101", -- t[38213] = 5
      "0000101" when "01001010101000110", -- t[38214] = 5
      "0000101" when "01001010101000111", -- t[38215] = 5
      "0000101" when "01001010101001000", -- t[38216] = 5
      "0000101" when "01001010101001001", -- t[38217] = 5
      "0000101" when "01001010101001010", -- t[38218] = 5
      "0000101" when "01001010101001011", -- t[38219] = 5
      "0000101" when "01001010101001100", -- t[38220] = 5
      "0000101" when "01001010101001101", -- t[38221] = 5
      "0000101" when "01001010101001110", -- t[38222] = 5
      "0000101" when "01001010101001111", -- t[38223] = 5
      "0000101" when "01001010101010000", -- t[38224] = 5
      "0000101" when "01001010101010001", -- t[38225] = 5
      "0000101" when "01001010101010010", -- t[38226] = 5
      "0000101" when "01001010101010011", -- t[38227] = 5
      "0000101" when "01001010101010100", -- t[38228] = 5
      "0000101" when "01001010101010101", -- t[38229] = 5
      "0000101" when "01001010101010110", -- t[38230] = 5
      "0000101" when "01001010101010111", -- t[38231] = 5
      "0000101" when "01001010101011000", -- t[38232] = 5
      "0000101" when "01001010101011001", -- t[38233] = 5
      "0000101" when "01001010101011010", -- t[38234] = 5
      "0000101" when "01001010101011011", -- t[38235] = 5
      "0000101" when "01001010101011100", -- t[38236] = 5
      "0000101" when "01001010101011101", -- t[38237] = 5
      "0000101" when "01001010101011110", -- t[38238] = 5
      "0000101" when "01001010101011111", -- t[38239] = 5
      "0000101" when "01001010101100000", -- t[38240] = 5
      "0000101" when "01001010101100001", -- t[38241] = 5
      "0000101" when "01001010101100010", -- t[38242] = 5
      "0000101" when "01001010101100011", -- t[38243] = 5
      "0000101" when "01001010101100100", -- t[38244] = 5
      "0000101" when "01001010101100101", -- t[38245] = 5
      "0000101" when "01001010101100110", -- t[38246] = 5
      "0000101" when "01001010101100111", -- t[38247] = 5
      "0000101" when "01001010101101000", -- t[38248] = 5
      "0000101" when "01001010101101001", -- t[38249] = 5
      "0000101" when "01001010101101010", -- t[38250] = 5
      "0000101" when "01001010101101011", -- t[38251] = 5
      "0000101" when "01001010101101100", -- t[38252] = 5
      "0000101" when "01001010101101101", -- t[38253] = 5
      "0000101" when "01001010101101110", -- t[38254] = 5
      "0000101" when "01001010101101111", -- t[38255] = 5
      "0000101" when "01001010101110000", -- t[38256] = 5
      "0000101" when "01001010101110001", -- t[38257] = 5
      "0000101" when "01001010101110010", -- t[38258] = 5
      "0000101" when "01001010101110011", -- t[38259] = 5
      "0000101" when "01001010101110100", -- t[38260] = 5
      "0000101" when "01001010101110101", -- t[38261] = 5
      "0000101" when "01001010101110110", -- t[38262] = 5
      "0000101" when "01001010101110111", -- t[38263] = 5
      "0000101" when "01001010101111000", -- t[38264] = 5
      "0000101" when "01001010101111001", -- t[38265] = 5
      "0000101" when "01001010101111010", -- t[38266] = 5
      "0000101" when "01001010101111011", -- t[38267] = 5
      "0000101" when "01001010101111100", -- t[38268] = 5
      "0000101" when "01001010101111101", -- t[38269] = 5
      "0000101" when "01001010101111110", -- t[38270] = 5
      "0000101" when "01001010101111111", -- t[38271] = 5
      "0000101" when "01001010110000000", -- t[38272] = 5
      "0000101" when "01001010110000001", -- t[38273] = 5
      "0000101" when "01001010110000010", -- t[38274] = 5
      "0000101" when "01001010110000011", -- t[38275] = 5
      "0000101" when "01001010110000100", -- t[38276] = 5
      "0000101" when "01001010110000101", -- t[38277] = 5
      "0000101" when "01001010110000110", -- t[38278] = 5
      "0000101" when "01001010110000111", -- t[38279] = 5
      "0000101" when "01001010110001000", -- t[38280] = 5
      "0000101" when "01001010110001001", -- t[38281] = 5
      "0000101" when "01001010110001010", -- t[38282] = 5
      "0000101" when "01001010110001011", -- t[38283] = 5
      "0000101" when "01001010110001100", -- t[38284] = 5
      "0000101" when "01001010110001101", -- t[38285] = 5
      "0000101" when "01001010110001110", -- t[38286] = 5
      "0000101" when "01001010110001111", -- t[38287] = 5
      "0000101" when "01001010110010000", -- t[38288] = 5
      "0000101" when "01001010110010001", -- t[38289] = 5
      "0000101" when "01001010110010010", -- t[38290] = 5
      "0000101" when "01001010110010011", -- t[38291] = 5
      "0000101" when "01001010110010100", -- t[38292] = 5
      "0000101" when "01001010110010101", -- t[38293] = 5
      "0000101" when "01001010110010110", -- t[38294] = 5
      "0000101" when "01001010110010111", -- t[38295] = 5
      "0000101" when "01001010110011000", -- t[38296] = 5
      "0000101" when "01001010110011001", -- t[38297] = 5
      "0000101" when "01001010110011010", -- t[38298] = 5
      "0000101" when "01001010110011011", -- t[38299] = 5
      "0000101" when "01001010110011100", -- t[38300] = 5
      "0000101" when "01001010110011101", -- t[38301] = 5
      "0000101" when "01001010110011110", -- t[38302] = 5
      "0000101" when "01001010110011111", -- t[38303] = 5
      "0000101" when "01001010110100000", -- t[38304] = 5
      "0000101" when "01001010110100001", -- t[38305] = 5
      "0000101" when "01001010110100010", -- t[38306] = 5
      "0000101" when "01001010110100011", -- t[38307] = 5
      "0000101" when "01001010110100100", -- t[38308] = 5
      "0000101" when "01001010110100101", -- t[38309] = 5
      "0000101" when "01001010110100110", -- t[38310] = 5
      "0000101" when "01001010110100111", -- t[38311] = 5
      "0000101" when "01001010110101000", -- t[38312] = 5
      "0000101" when "01001010110101001", -- t[38313] = 5
      "0000101" when "01001010110101010", -- t[38314] = 5
      "0000101" when "01001010110101011", -- t[38315] = 5
      "0000101" when "01001010110101100", -- t[38316] = 5
      "0000101" when "01001010110101101", -- t[38317] = 5
      "0000101" when "01001010110101110", -- t[38318] = 5
      "0000101" when "01001010110101111", -- t[38319] = 5
      "0000101" when "01001010110110000", -- t[38320] = 5
      "0000101" when "01001010110110001", -- t[38321] = 5
      "0000101" when "01001010110110010", -- t[38322] = 5
      "0000101" when "01001010110110011", -- t[38323] = 5
      "0000101" when "01001010110110100", -- t[38324] = 5
      "0000101" when "01001010110110101", -- t[38325] = 5
      "0000101" when "01001010110110110", -- t[38326] = 5
      "0000101" when "01001010110110111", -- t[38327] = 5
      "0000101" when "01001010110111000", -- t[38328] = 5
      "0000101" when "01001010110111001", -- t[38329] = 5
      "0000101" when "01001010110111010", -- t[38330] = 5
      "0000101" when "01001010110111011", -- t[38331] = 5
      "0000101" when "01001010110111100", -- t[38332] = 5
      "0000101" when "01001010110111101", -- t[38333] = 5
      "0000101" when "01001010110111110", -- t[38334] = 5
      "0000101" when "01001010110111111", -- t[38335] = 5
      "0000101" when "01001010111000000", -- t[38336] = 5
      "0000101" when "01001010111000001", -- t[38337] = 5
      "0000101" when "01001010111000010", -- t[38338] = 5
      "0000101" when "01001010111000011", -- t[38339] = 5
      "0000101" when "01001010111000100", -- t[38340] = 5
      "0000101" when "01001010111000101", -- t[38341] = 5
      "0000101" when "01001010111000110", -- t[38342] = 5
      "0000101" when "01001010111000111", -- t[38343] = 5
      "0000101" when "01001010111001000", -- t[38344] = 5
      "0000101" when "01001010111001001", -- t[38345] = 5
      "0000101" when "01001010111001010", -- t[38346] = 5
      "0000101" when "01001010111001011", -- t[38347] = 5
      "0000101" when "01001010111001100", -- t[38348] = 5
      "0000101" when "01001010111001101", -- t[38349] = 5
      "0000101" when "01001010111001110", -- t[38350] = 5
      "0000101" when "01001010111001111", -- t[38351] = 5
      "0000101" when "01001010111010000", -- t[38352] = 5
      "0000101" when "01001010111010001", -- t[38353] = 5
      "0000101" when "01001010111010010", -- t[38354] = 5
      "0000101" when "01001010111010011", -- t[38355] = 5
      "0000101" when "01001010111010100", -- t[38356] = 5
      "0000101" when "01001010111010101", -- t[38357] = 5
      "0000101" when "01001010111010110", -- t[38358] = 5
      "0000101" when "01001010111010111", -- t[38359] = 5
      "0000101" when "01001010111011000", -- t[38360] = 5
      "0000101" when "01001010111011001", -- t[38361] = 5
      "0000101" when "01001010111011010", -- t[38362] = 5
      "0000101" when "01001010111011011", -- t[38363] = 5
      "0000101" when "01001010111011100", -- t[38364] = 5
      "0000101" when "01001010111011101", -- t[38365] = 5
      "0000101" when "01001010111011110", -- t[38366] = 5
      "0000101" when "01001010111011111", -- t[38367] = 5
      "0000101" when "01001010111100000", -- t[38368] = 5
      "0000101" when "01001010111100001", -- t[38369] = 5
      "0000101" when "01001010111100010", -- t[38370] = 5
      "0000101" when "01001010111100011", -- t[38371] = 5
      "0000101" when "01001010111100100", -- t[38372] = 5
      "0000101" when "01001010111100101", -- t[38373] = 5
      "0000101" when "01001010111100110", -- t[38374] = 5
      "0000101" when "01001010111100111", -- t[38375] = 5
      "0000101" when "01001010111101000", -- t[38376] = 5
      "0000101" when "01001010111101001", -- t[38377] = 5
      "0000101" when "01001010111101010", -- t[38378] = 5
      "0000101" when "01001010111101011", -- t[38379] = 5
      "0000101" when "01001010111101100", -- t[38380] = 5
      "0000101" when "01001010111101101", -- t[38381] = 5
      "0000101" when "01001010111101110", -- t[38382] = 5
      "0000101" when "01001010111101111", -- t[38383] = 5
      "0000101" when "01001010111110000", -- t[38384] = 5
      "0000101" when "01001010111110001", -- t[38385] = 5
      "0000101" when "01001010111110010", -- t[38386] = 5
      "0000101" when "01001010111110011", -- t[38387] = 5
      "0000101" when "01001010111110100", -- t[38388] = 5
      "0000101" when "01001010111110101", -- t[38389] = 5
      "0000101" when "01001010111110110", -- t[38390] = 5
      "0000101" when "01001010111110111", -- t[38391] = 5
      "0000101" when "01001010111111000", -- t[38392] = 5
      "0000101" when "01001010111111001", -- t[38393] = 5
      "0000101" when "01001010111111010", -- t[38394] = 5
      "0000101" when "01001010111111011", -- t[38395] = 5
      "0000101" when "01001010111111100", -- t[38396] = 5
      "0000101" when "01001010111111101", -- t[38397] = 5
      "0000101" when "01001010111111110", -- t[38398] = 5
      "0000101" when "01001010111111111", -- t[38399] = 5
      "0000101" when "01001011000000000", -- t[38400] = 5
      "0000101" when "01001011000000001", -- t[38401] = 5
      "0000101" when "01001011000000010", -- t[38402] = 5
      "0000101" when "01001011000000011", -- t[38403] = 5
      "0000101" when "01001011000000100", -- t[38404] = 5
      "0000101" when "01001011000000101", -- t[38405] = 5
      "0000101" when "01001011000000110", -- t[38406] = 5
      "0000101" when "01001011000000111", -- t[38407] = 5
      "0000101" when "01001011000001000", -- t[38408] = 5
      "0000101" when "01001011000001001", -- t[38409] = 5
      "0000101" when "01001011000001010", -- t[38410] = 5
      "0000101" when "01001011000001011", -- t[38411] = 5
      "0000101" when "01001011000001100", -- t[38412] = 5
      "0000101" when "01001011000001101", -- t[38413] = 5
      "0000101" when "01001011000001110", -- t[38414] = 5
      "0000101" when "01001011000001111", -- t[38415] = 5
      "0000101" when "01001011000010000", -- t[38416] = 5
      "0000101" when "01001011000010001", -- t[38417] = 5
      "0000101" when "01001011000010010", -- t[38418] = 5
      "0000101" when "01001011000010011", -- t[38419] = 5
      "0000101" when "01001011000010100", -- t[38420] = 5
      "0000101" when "01001011000010101", -- t[38421] = 5
      "0000101" when "01001011000010110", -- t[38422] = 5
      "0000101" when "01001011000010111", -- t[38423] = 5
      "0000101" when "01001011000011000", -- t[38424] = 5
      "0000101" when "01001011000011001", -- t[38425] = 5
      "0000101" when "01001011000011010", -- t[38426] = 5
      "0000101" when "01001011000011011", -- t[38427] = 5
      "0000101" when "01001011000011100", -- t[38428] = 5
      "0000101" when "01001011000011101", -- t[38429] = 5
      "0000101" when "01001011000011110", -- t[38430] = 5
      "0000101" when "01001011000011111", -- t[38431] = 5
      "0000101" when "01001011000100000", -- t[38432] = 5
      "0000101" when "01001011000100001", -- t[38433] = 5
      "0000101" when "01001011000100010", -- t[38434] = 5
      "0000101" when "01001011000100011", -- t[38435] = 5
      "0000101" when "01001011000100100", -- t[38436] = 5
      "0000101" when "01001011000100101", -- t[38437] = 5
      "0000101" when "01001011000100110", -- t[38438] = 5
      "0000101" when "01001011000100111", -- t[38439] = 5
      "0000101" when "01001011000101000", -- t[38440] = 5
      "0000101" when "01001011000101001", -- t[38441] = 5
      "0000101" when "01001011000101010", -- t[38442] = 5
      "0000101" when "01001011000101011", -- t[38443] = 5
      "0000101" when "01001011000101100", -- t[38444] = 5
      "0000101" when "01001011000101101", -- t[38445] = 5
      "0000101" when "01001011000101110", -- t[38446] = 5
      "0000101" when "01001011000101111", -- t[38447] = 5
      "0000101" when "01001011000110000", -- t[38448] = 5
      "0000101" when "01001011000110001", -- t[38449] = 5
      "0000101" when "01001011000110010", -- t[38450] = 5
      "0000101" when "01001011000110011", -- t[38451] = 5
      "0000101" when "01001011000110100", -- t[38452] = 5
      "0000101" when "01001011000110101", -- t[38453] = 5
      "0000101" when "01001011000110110", -- t[38454] = 5
      "0000101" when "01001011000110111", -- t[38455] = 5
      "0000101" when "01001011000111000", -- t[38456] = 5
      "0000101" when "01001011000111001", -- t[38457] = 5
      "0000101" when "01001011000111010", -- t[38458] = 5
      "0000101" when "01001011000111011", -- t[38459] = 5
      "0000101" when "01001011000111100", -- t[38460] = 5
      "0000101" when "01001011000111101", -- t[38461] = 5
      "0000101" when "01001011000111110", -- t[38462] = 5
      "0000101" when "01001011000111111", -- t[38463] = 5
      "0000101" when "01001011001000000", -- t[38464] = 5
      "0000101" when "01001011001000001", -- t[38465] = 5
      "0000101" when "01001011001000010", -- t[38466] = 5
      "0000101" when "01001011001000011", -- t[38467] = 5
      "0000101" when "01001011001000100", -- t[38468] = 5
      "0000101" when "01001011001000101", -- t[38469] = 5
      "0000101" when "01001011001000110", -- t[38470] = 5
      "0000101" when "01001011001000111", -- t[38471] = 5
      "0000101" when "01001011001001000", -- t[38472] = 5
      "0000101" when "01001011001001001", -- t[38473] = 5
      "0000101" when "01001011001001010", -- t[38474] = 5
      "0000101" when "01001011001001011", -- t[38475] = 5
      "0000101" when "01001011001001100", -- t[38476] = 5
      "0000101" when "01001011001001101", -- t[38477] = 5
      "0000101" when "01001011001001110", -- t[38478] = 5
      "0000101" when "01001011001001111", -- t[38479] = 5
      "0000101" when "01001011001010000", -- t[38480] = 5
      "0000101" when "01001011001010001", -- t[38481] = 5
      "0000101" when "01001011001010010", -- t[38482] = 5
      "0000101" when "01001011001010011", -- t[38483] = 5
      "0000101" when "01001011001010100", -- t[38484] = 5
      "0000101" when "01001011001010101", -- t[38485] = 5
      "0000101" when "01001011001010110", -- t[38486] = 5
      "0000101" when "01001011001010111", -- t[38487] = 5
      "0000101" when "01001011001011000", -- t[38488] = 5
      "0000101" when "01001011001011001", -- t[38489] = 5
      "0000101" when "01001011001011010", -- t[38490] = 5
      "0000101" when "01001011001011011", -- t[38491] = 5
      "0000101" when "01001011001011100", -- t[38492] = 5
      "0000101" when "01001011001011101", -- t[38493] = 5
      "0000101" when "01001011001011110", -- t[38494] = 5
      "0000101" when "01001011001011111", -- t[38495] = 5
      "0000101" when "01001011001100000", -- t[38496] = 5
      "0000101" when "01001011001100001", -- t[38497] = 5
      "0000101" when "01001011001100010", -- t[38498] = 5
      "0000101" when "01001011001100011", -- t[38499] = 5
      "0000101" when "01001011001100100", -- t[38500] = 5
      "0000101" when "01001011001100101", -- t[38501] = 5
      "0000101" when "01001011001100110", -- t[38502] = 5
      "0000101" when "01001011001100111", -- t[38503] = 5
      "0000101" when "01001011001101000", -- t[38504] = 5
      "0000101" when "01001011001101001", -- t[38505] = 5
      "0000101" when "01001011001101010", -- t[38506] = 5
      "0000101" when "01001011001101011", -- t[38507] = 5
      "0000101" when "01001011001101100", -- t[38508] = 5
      "0000101" when "01001011001101101", -- t[38509] = 5
      "0000101" when "01001011001101110", -- t[38510] = 5
      "0000101" when "01001011001101111", -- t[38511] = 5
      "0000101" when "01001011001110000", -- t[38512] = 5
      "0000101" when "01001011001110001", -- t[38513] = 5
      "0000101" when "01001011001110010", -- t[38514] = 5
      "0000101" when "01001011001110011", -- t[38515] = 5
      "0000101" when "01001011001110100", -- t[38516] = 5
      "0000101" when "01001011001110101", -- t[38517] = 5
      "0000101" when "01001011001110110", -- t[38518] = 5
      "0000101" when "01001011001110111", -- t[38519] = 5
      "0000101" when "01001011001111000", -- t[38520] = 5
      "0000101" when "01001011001111001", -- t[38521] = 5
      "0000101" when "01001011001111010", -- t[38522] = 5
      "0000101" when "01001011001111011", -- t[38523] = 5
      "0000101" when "01001011001111100", -- t[38524] = 5
      "0000101" when "01001011001111101", -- t[38525] = 5
      "0000101" when "01001011001111110", -- t[38526] = 5
      "0000101" when "01001011001111111", -- t[38527] = 5
      "0000101" when "01001011010000000", -- t[38528] = 5
      "0000101" when "01001011010000001", -- t[38529] = 5
      "0000101" when "01001011010000010", -- t[38530] = 5
      "0000101" when "01001011010000011", -- t[38531] = 5
      "0000101" when "01001011010000100", -- t[38532] = 5
      "0000101" when "01001011010000101", -- t[38533] = 5
      "0000101" when "01001011010000110", -- t[38534] = 5
      "0000101" when "01001011010000111", -- t[38535] = 5
      "0000101" when "01001011010001000", -- t[38536] = 5
      "0000101" when "01001011010001001", -- t[38537] = 5
      "0000101" when "01001011010001010", -- t[38538] = 5
      "0000101" when "01001011010001011", -- t[38539] = 5
      "0000101" when "01001011010001100", -- t[38540] = 5
      "0000101" when "01001011010001101", -- t[38541] = 5
      "0000101" when "01001011010001110", -- t[38542] = 5
      "0000101" when "01001011010001111", -- t[38543] = 5
      "0000101" when "01001011010010000", -- t[38544] = 5
      "0000101" when "01001011010010001", -- t[38545] = 5
      "0000101" when "01001011010010010", -- t[38546] = 5
      "0000101" when "01001011010010011", -- t[38547] = 5
      "0000101" when "01001011010010100", -- t[38548] = 5
      "0000101" when "01001011010010101", -- t[38549] = 5
      "0000101" when "01001011010010110", -- t[38550] = 5
      "0000101" when "01001011010010111", -- t[38551] = 5
      "0000101" when "01001011010011000", -- t[38552] = 5
      "0000101" when "01001011010011001", -- t[38553] = 5
      "0000101" when "01001011010011010", -- t[38554] = 5
      "0000101" when "01001011010011011", -- t[38555] = 5
      "0000101" when "01001011010011100", -- t[38556] = 5
      "0000101" when "01001011010011101", -- t[38557] = 5
      "0000101" when "01001011010011110", -- t[38558] = 5
      "0000101" when "01001011010011111", -- t[38559] = 5
      "0000101" when "01001011010100000", -- t[38560] = 5
      "0000101" when "01001011010100001", -- t[38561] = 5
      "0000101" when "01001011010100010", -- t[38562] = 5
      "0000101" when "01001011010100011", -- t[38563] = 5
      "0000101" when "01001011010100100", -- t[38564] = 5
      "0000101" when "01001011010100101", -- t[38565] = 5
      "0000101" when "01001011010100110", -- t[38566] = 5
      "0000101" when "01001011010100111", -- t[38567] = 5
      "0000101" when "01001011010101000", -- t[38568] = 5
      "0000101" when "01001011010101001", -- t[38569] = 5
      "0000101" when "01001011010101010", -- t[38570] = 5
      "0000101" when "01001011010101011", -- t[38571] = 5
      "0000101" when "01001011010101100", -- t[38572] = 5
      "0000101" when "01001011010101101", -- t[38573] = 5
      "0000101" when "01001011010101110", -- t[38574] = 5
      "0000101" when "01001011010101111", -- t[38575] = 5
      "0000101" when "01001011010110000", -- t[38576] = 5
      "0000101" when "01001011010110001", -- t[38577] = 5
      "0000101" when "01001011010110010", -- t[38578] = 5
      "0000101" when "01001011010110011", -- t[38579] = 5
      "0000101" when "01001011010110100", -- t[38580] = 5
      "0000101" when "01001011010110101", -- t[38581] = 5
      "0000101" when "01001011010110110", -- t[38582] = 5
      "0000101" when "01001011010110111", -- t[38583] = 5
      "0000101" when "01001011010111000", -- t[38584] = 5
      "0000101" when "01001011010111001", -- t[38585] = 5
      "0000101" when "01001011010111010", -- t[38586] = 5
      "0000101" when "01001011010111011", -- t[38587] = 5
      "0000101" when "01001011010111100", -- t[38588] = 5
      "0000101" when "01001011010111101", -- t[38589] = 5
      "0000101" when "01001011010111110", -- t[38590] = 5
      "0000101" when "01001011010111111", -- t[38591] = 5
      "0000101" when "01001011011000000", -- t[38592] = 5
      "0000101" when "01001011011000001", -- t[38593] = 5
      "0000101" when "01001011011000010", -- t[38594] = 5
      "0000101" when "01001011011000011", -- t[38595] = 5
      "0000101" when "01001011011000100", -- t[38596] = 5
      "0000101" when "01001011011000101", -- t[38597] = 5
      "0000101" when "01001011011000110", -- t[38598] = 5
      "0000101" when "01001011011000111", -- t[38599] = 5
      "0000101" when "01001011011001000", -- t[38600] = 5
      "0000101" when "01001011011001001", -- t[38601] = 5
      "0000101" when "01001011011001010", -- t[38602] = 5
      "0000101" when "01001011011001011", -- t[38603] = 5
      "0000101" when "01001011011001100", -- t[38604] = 5
      "0000101" when "01001011011001101", -- t[38605] = 5
      "0000101" when "01001011011001110", -- t[38606] = 5
      "0000101" when "01001011011001111", -- t[38607] = 5
      "0000101" when "01001011011010000", -- t[38608] = 5
      "0000101" when "01001011011010001", -- t[38609] = 5
      "0000101" when "01001011011010010", -- t[38610] = 5
      "0000101" when "01001011011010011", -- t[38611] = 5
      "0000101" when "01001011011010100", -- t[38612] = 5
      "0000101" when "01001011011010101", -- t[38613] = 5
      "0000101" when "01001011011010110", -- t[38614] = 5
      "0000101" when "01001011011010111", -- t[38615] = 5
      "0000101" when "01001011011011000", -- t[38616] = 5
      "0000101" when "01001011011011001", -- t[38617] = 5
      "0000101" when "01001011011011010", -- t[38618] = 5
      "0000101" when "01001011011011011", -- t[38619] = 5
      "0000101" when "01001011011011100", -- t[38620] = 5
      "0000101" when "01001011011011101", -- t[38621] = 5
      "0000101" when "01001011011011110", -- t[38622] = 5
      "0000101" when "01001011011011111", -- t[38623] = 5
      "0000101" when "01001011011100000", -- t[38624] = 5
      "0000101" when "01001011011100001", -- t[38625] = 5
      "0000101" when "01001011011100010", -- t[38626] = 5
      "0000101" when "01001011011100011", -- t[38627] = 5
      "0000101" when "01001011011100100", -- t[38628] = 5
      "0000101" when "01001011011100101", -- t[38629] = 5
      "0000101" when "01001011011100110", -- t[38630] = 5
      "0000101" when "01001011011100111", -- t[38631] = 5
      "0000101" when "01001011011101000", -- t[38632] = 5
      "0000101" when "01001011011101001", -- t[38633] = 5
      "0000101" when "01001011011101010", -- t[38634] = 5
      "0000101" when "01001011011101011", -- t[38635] = 5
      "0000101" when "01001011011101100", -- t[38636] = 5
      "0000101" when "01001011011101101", -- t[38637] = 5
      "0000101" when "01001011011101110", -- t[38638] = 5
      "0000101" when "01001011011101111", -- t[38639] = 5
      "0000101" when "01001011011110000", -- t[38640] = 5
      "0000101" when "01001011011110001", -- t[38641] = 5
      "0000101" when "01001011011110010", -- t[38642] = 5
      "0000101" when "01001011011110011", -- t[38643] = 5
      "0000101" when "01001011011110100", -- t[38644] = 5
      "0000101" when "01001011011110101", -- t[38645] = 5
      "0000101" when "01001011011110110", -- t[38646] = 5
      "0000101" when "01001011011110111", -- t[38647] = 5
      "0000101" when "01001011011111000", -- t[38648] = 5
      "0000101" when "01001011011111001", -- t[38649] = 5
      "0000101" when "01001011011111010", -- t[38650] = 5
      "0000101" when "01001011011111011", -- t[38651] = 5
      "0000101" when "01001011011111100", -- t[38652] = 5
      "0000101" when "01001011011111101", -- t[38653] = 5
      "0000101" when "01001011011111110", -- t[38654] = 5
      "0000101" when "01001011011111111", -- t[38655] = 5
      "0000101" when "01001011100000000", -- t[38656] = 5
      "0000101" when "01001011100000001", -- t[38657] = 5
      "0000101" when "01001011100000010", -- t[38658] = 5
      "0000101" when "01001011100000011", -- t[38659] = 5
      "0000101" when "01001011100000100", -- t[38660] = 5
      "0000101" when "01001011100000101", -- t[38661] = 5
      "0000101" when "01001011100000110", -- t[38662] = 5
      "0000101" when "01001011100000111", -- t[38663] = 5
      "0000101" when "01001011100001000", -- t[38664] = 5
      "0000101" when "01001011100001001", -- t[38665] = 5
      "0000101" when "01001011100001010", -- t[38666] = 5
      "0000101" when "01001011100001011", -- t[38667] = 5
      "0000101" when "01001011100001100", -- t[38668] = 5
      "0000101" when "01001011100001101", -- t[38669] = 5
      "0000101" when "01001011100001110", -- t[38670] = 5
      "0000101" when "01001011100001111", -- t[38671] = 5
      "0000101" when "01001011100010000", -- t[38672] = 5
      "0000101" when "01001011100010001", -- t[38673] = 5
      "0000101" when "01001011100010010", -- t[38674] = 5
      "0000101" when "01001011100010011", -- t[38675] = 5
      "0000101" when "01001011100010100", -- t[38676] = 5
      "0000101" when "01001011100010101", -- t[38677] = 5
      "0000101" when "01001011100010110", -- t[38678] = 5
      "0000101" when "01001011100010111", -- t[38679] = 5
      "0000101" when "01001011100011000", -- t[38680] = 5
      "0000101" when "01001011100011001", -- t[38681] = 5
      "0000101" when "01001011100011010", -- t[38682] = 5
      "0000101" when "01001011100011011", -- t[38683] = 5
      "0000101" when "01001011100011100", -- t[38684] = 5
      "0000101" when "01001011100011101", -- t[38685] = 5
      "0000101" when "01001011100011110", -- t[38686] = 5
      "0000101" when "01001011100011111", -- t[38687] = 5
      "0000101" when "01001011100100000", -- t[38688] = 5
      "0000101" when "01001011100100001", -- t[38689] = 5
      "0000101" when "01001011100100010", -- t[38690] = 5
      "0000101" when "01001011100100011", -- t[38691] = 5
      "0000101" when "01001011100100100", -- t[38692] = 5
      "0000101" when "01001011100100101", -- t[38693] = 5
      "0000101" when "01001011100100110", -- t[38694] = 5
      "0000101" when "01001011100100111", -- t[38695] = 5
      "0000101" when "01001011100101000", -- t[38696] = 5
      "0000101" when "01001011100101001", -- t[38697] = 5
      "0000101" when "01001011100101010", -- t[38698] = 5
      "0000101" when "01001011100101011", -- t[38699] = 5
      "0000101" when "01001011100101100", -- t[38700] = 5
      "0000101" when "01001011100101101", -- t[38701] = 5
      "0000101" when "01001011100101110", -- t[38702] = 5
      "0000101" when "01001011100101111", -- t[38703] = 5
      "0000101" when "01001011100110000", -- t[38704] = 5
      "0000101" when "01001011100110001", -- t[38705] = 5
      "0000101" when "01001011100110010", -- t[38706] = 5
      "0000101" when "01001011100110011", -- t[38707] = 5
      "0000101" when "01001011100110100", -- t[38708] = 5
      "0000101" when "01001011100110101", -- t[38709] = 5
      "0000101" when "01001011100110110", -- t[38710] = 5
      "0000101" when "01001011100110111", -- t[38711] = 5
      "0000101" when "01001011100111000", -- t[38712] = 5
      "0000101" when "01001011100111001", -- t[38713] = 5
      "0000101" when "01001011100111010", -- t[38714] = 5
      "0000101" when "01001011100111011", -- t[38715] = 5
      "0000101" when "01001011100111100", -- t[38716] = 5
      "0000101" when "01001011100111101", -- t[38717] = 5
      "0000101" when "01001011100111110", -- t[38718] = 5
      "0000101" when "01001011100111111", -- t[38719] = 5
      "0000101" when "01001011101000000", -- t[38720] = 5
      "0000101" when "01001011101000001", -- t[38721] = 5
      "0000101" when "01001011101000010", -- t[38722] = 5
      "0000101" when "01001011101000011", -- t[38723] = 5
      "0000101" when "01001011101000100", -- t[38724] = 5
      "0000101" when "01001011101000101", -- t[38725] = 5
      "0000101" when "01001011101000110", -- t[38726] = 5
      "0000101" when "01001011101000111", -- t[38727] = 5
      "0000101" when "01001011101001000", -- t[38728] = 5
      "0000101" when "01001011101001001", -- t[38729] = 5
      "0000101" when "01001011101001010", -- t[38730] = 5
      "0000101" when "01001011101001011", -- t[38731] = 5
      "0000101" when "01001011101001100", -- t[38732] = 5
      "0000101" when "01001011101001101", -- t[38733] = 5
      "0000101" when "01001011101001110", -- t[38734] = 5
      "0000101" when "01001011101001111", -- t[38735] = 5
      "0000101" when "01001011101010000", -- t[38736] = 5
      "0000101" when "01001011101010001", -- t[38737] = 5
      "0000101" when "01001011101010010", -- t[38738] = 5
      "0000101" when "01001011101010011", -- t[38739] = 5
      "0000101" when "01001011101010100", -- t[38740] = 5
      "0000101" when "01001011101010101", -- t[38741] = 5
      "0000101" when "01001011101010110", -- t[38742] = 5
      "0000101" when "01001011101010111", -- t[38743] = 5
      "0000101" when "01001011101011000", -- t[38744] = 5
      "0000101" when "01001011101011001", -- t[38745] = 5
      "0000101" when "01001011101011010", -- t[38746] = 5
      "0000101" when "01001011101011011", -- t[38747] = 5
      "0000101" when "01001011101011100", -- t[38748] = 5
      "0000101" when "01001011101011101", -- t[38749] = 5
      "0000101" when "01001011101011110", -- t[38750] = 5
      "0000101" when "01001011101011111", -- t[38751] = 5
      "0000101" when "01001011101100000", -- t[38752] = 5
      "0000101" when "01001011101100001", -- t[38753] = 5
      "0000101" when "01001011101100010", -- t[38754] = 5
      "0000101" when "01001011101100011", -- t[38755] = 5
      "0000101" when "01001011101100100", -- t[38756] = 5
      "0000101" when "01001011101100101", -- t[38757] = 5
      "0000101" when "01001011101100110", -- t[38758] = 5
      "0000101" when "01001011101100111", -- t[38759] = 5
      "0000101" when "01001011101101000", -- t[38760] = 5
      "0000101" when "01001011101101001", -- t[38761] = 5
      "0000101" when "01001011101101010", -- t[38762] = 5
      "0000101" when "01001011101101011", -- t[38763] = 5
      "0000101" when "01001011101101100", -- t[38764] = 5
      "0000101" when "01001011101101101", -- t[38765] = 5
      "0000101" when "01001011101101110", -- t[38766] = 5
      "0000101" when "01001011101101111", -- t[38767] = 5
      "0000101" when "01001011101110000", -- t[38768] = 5
      "0000101" when "01001011101110001", -- t[38769] = 5
      "0000101" when "01001011101110010", -- t[38770] = 5
      "0000101" when "01001011101110011", -- t[38771] = 5
      "0000101" when "01001011101110100", -- t[38772] = 5
      "0000101" when "01001011101110101", -- t[38773] = 5
      "0000101" when "01001011101110110", -- t[38774] = 5
      "0000101" when "01001011101110111", -- t[38775] = 5
      "0000101" when "01001011101111000", -- t[38776] = 5
      "0000101" when "01001011101111001", -- t[38777] = 5
      "0000101" when "01001011101111010", -- t[38778] = 5
      "0000101" when "01001011101111011", -- t[38779] = 5
      "0000101" when "01001011101111100", -- t[38780] = 5
      "0000101" when "01001011101111101", -- t[38781] = 5
      "0000101" when "01001011101111110", -- t[38782] = 5
      "0000101" when "01001011101111111", -- t[38783] = 5
      "0000101" when "01001011110000000", -- t[38784] = 5
      "0000101" when "01001011110000001", -- t[38785] = 5
      "0000101" when "01001011110000010", -- t[38786] = 5
      "0000101" when "01001011110000011", -- t[38787] = 5
      "0000101" when "01001011110000100", -- t[38788] = 5
      "0000101" when "01001011110000101", -- t[38789] = 5
      "0000101" when "01001011110000110", -- t[38790] = 5
      "0000101" when "01001011110000111", -- t[38791] = 5
      "0000101" when "01001011110001000", -- t[38792] = 5
      "0000101" when "01001011110001001", -- t[38793] = 5
      "0000101" when "01001011110001010", -- t[38794] = 5
      "0000101" when "01001011110001011", -- t[38795] = 5
      "0000101" when "01001011110001100", -- t[38796] = 5
      "0000101" when "01001011110001101", -- t[38797] = 5
      "0000101" when "01001011110001110", -- t[38798] = 5
      "0000101" when "01001011110001111", -- t[38799] = 5
      "0000101" when "01001011110010000", -- t[38800] = 5
      "0000101" when "01001011110010001", -- t[38801] = 5
      "0000101" when "01001011110010010", -- t[38802] = 5
      "0000101" when "01001011110010011", -- t[38803] = 5
      "0000101" when "01001011110010100", -- t[38804] = 5
      "0000101" when "01001011110010101", -- t[38805] = 5
      "0000101" when "01001011110010110", -- t[38806] = 5
      "0000101" when "01001011110010111", -- t[38807] = 5
      "0000101" when "01001011110011000", -- t[38808] = 5
      "0000101" when "01001011110011001", -- t[38809] = 5
      "0000101" when "01001011110011010", -- t[38810] = 5
      "0000101" when "01001011110011011", -- t[38811] = 5
      "0000101" when "01001011110011100", -- t[38812] = 5
      "0000101" when "01001011110011101", -- t[38813] = 5
      "0000101" when "01001011110011110", -- t[38814] = 5
      "0000101" when "01001011110011111", -- t[38815] = 5
      "0000101" when "01001011110100000", -- t[38816] = 5
      "0000101" when "01001011110100001", -- t[38817] = 5
      "0000101" when "01001011110100010", -- t[38818] = 5
      "0000101" when "01001011110100011", -- t[38819] = 5
      "0000101" when "01001011110100100", -- t[38820] = 5
      "0000101" when "01001011110100101", -- t[38821] = 5
      "0000101" when "01001011110100110", -- t[38822] = 5
      "0000101" when "01001011110100111", -- t[38823] = 5
      "0000101" when "01001011110101000", -- t[38824] = 5
      "0000101" when "01001011110101001", -- t[38825] = 5
      "0000101" when "01001011110101010", -- t[38826] = 5
      "0000101" when "01001011110101011", -- t[38827] = 5
      "0000101" when "01001011110101100", -- t[38828] = 5
      "0000101" when "01001011110101101", -- t[38829] = 5
      "0000101" when "01001011110101110", -- t[38830] = 5
      "0000101" when "01001011110101111", -- t[38831] = 5
      "0000101" when "01001011110110000", -- t[38832] = 5
      "0000101" when "01001011110110001", -- t[38833] = 5
      "0000101" when "01001011110110010", -- t[38834] = 5
      "0000101" when "01001011110110011", -- t[38835] = 5
      "0000101" when "01001011110110100", -- t[38836] = 5
      "0000101" when "01001011110110101", -- t[38837] = 5
      "0000101" when "01001011110110110", -- t[38838] = 5
      "0000101" when "01001011110110111", -- t[38839] = 5
      "0000101" when "01001011110111000", -- t[38840] = 5
      "0000101" when "01001011110111001", -- t[38841] = 5
      "0000101" when "01001011110111010", -- t[38842] = 5
      "0000101" when "01001011110111011", -- t[38843] = 5
      "0000101" when "01001011110111100", -- t[38844] = 5
      "0000101" when "01001011110111101", -- t[38845] = 5
      "0000101" when "01001011110111110", -- t[38846] = 5
      "0000101" when "01001011110111111", -- t[38847] = 5
      "0000101" when "01001011111000000", -- t[38848] = 5
      "0000101" when "01001011111000001", -- t[38849] = 5
      "0000101" when "01001011111000010", -- t[38850] = 5
      "0000101" when "01001011111000011", -- t[38851] = 5
      "0000101" when "01001011111000100", -- t[38852] = 5
      "0000101" when "01001011111000101", -- t[38853] = 5
      "0000101" when "01001011111000110", -- t[38854] = 5
      "0000101" when "01001011111000111", -- t[38855] = 5
      "0000101" when "01001011111001000", -- t[38856] = 5
      "0000101" when "01001011111001001", -- t[38857] = 5
      "0000101" when "01001011111001010", -- t[38858] = 5
      "0000101" when "01001011111001011", -- t[38859] = 5
      "0000101" when "01001011111001100", -- t[38860] = 5
      "0000101" when "01001011111001101", -- t[38861] = 5
      "0000101" when "01001011111001110", -- t[38862] = 5
      "0000101" when "01001011111001111", -- t[38863] = 5
      "0000101" when "01001011111010000", -- t[38864] = 5
      "0000101" when "01001011111010001", -- t[38865] = 5
      "0000101" when "01001011111010010", -- t[38866] = 5
      "0000101" when "01001011111010011", -- t[38867] = 5
      "0000101" when "01001011111010100", -- t[38868] = 5
      "0000101" when "01001011111010101", -- t[38869] = 5
      "0000101" when "01001011111010110", -- t[38870] = 5
      "0000101" when "01001011111010111", -- t[38871] = 5
      "0000101" when "01001011111011000", -- t[38872] = 5
      "0000101" when "01001011111011001", -- t[38873] = 5
      "0000101" when "01001011111011010", -- t[38874] = 5
      "0000101" when "01001011111011011", -- t[38875] = 5
      "0000101" when "01001011111011100", -- t[38876] = 5
      "0000101" when "01001011111011101", -- t[38877] = 5
      "0000101" when "01001011111011110", -- t[38878] = 5
      "0000101" when "01001011111011111", -- t[38879] = 5
      "0000101" when "01001011111100000", -- t[38880] = 5
      "0000101" when "01001011111100001", -- t[38881] = 5
      "0000101" when "01001011111100010", -- t[38882] = 5
      "0000101" when "01001011111100011", -- t[38883] = 5
      "0000101" when "01001011111100100", -- t[38884] = 5
      "0000101" when "01001011111100101", -- t[38885] = 5
      "0000101" when "01001011111100110", -- t[38886] = 5
      "0000101" when "01001011111100111", -- t[38887] = 5
      "0000101" when "01001011111101000", -- t[38888] = 5
      "0000101" when "01001011111101001", -- t[38889] = 5
      "0000101" when "01001011111101010", -- t[38890] = 5
      "0000101" when "01001011111101011", -- t[38891] = 5
      "0000101" when "01001011111101100", -- t[38892] = 5
      "0000101" when "01001011111101101", -- t[38893] = 5
      "0000101" when "01001011111101110", -- t[38894] = 5
      "0000101" when "01001011111101111", -- t[38895] = 5
      "0000101" when "01001011111110000", -- t[38896] = 5
      "0000101" when "01001011111110001", -- t[38897] = 5
      "0000101" when "01001011111110010", -- t[38898] = 5
      "0000101" when "01001011111110011", -- t[38899] = 5
      "0000101" when "01001011111110100", -- t[38900] = 5
      "0000101" when "01001011111110101", -- t[38901] = 5
      "0000101" when "01001011111110110", -- t[38902] = 5
      "0000101" when "01001011111110111", -- t[38903] = 5
      "0000101" when "01001011111111000", -- t[38904] = 5
      "0000101" when "01001011111111001", -- t[38905] = 5
      "0000101" when "01001011111111010", -- t[38906] = 5
      "0000101" when "01001011111111011", -- t[38907] = 5
      "0000101" when "01001011111111100", -- t[38908] = 5
      "0000101" when "01001011111111101", -- t[38909] = 5
      "0000101" when "01001011111111110", -- t[38910] = 5
      "0000101" when "01001011111111111", -- t[38911] = 5
      "0000101" when "01001100000000000", -- t[38912] = 5
      "0000101" when "01001100000000001", -- t[38913] = 5
      "0000101" when "01001100000000010", -- t[38914] = 5
      "0000101" when "01001100000000011", -- t[38915] = 5
      "0000101" when "01001100000000100", -- t[38916] = 5
      "0000101" when "01001100000000101", -- t[38917] = 5
      "0000101" when "01001100000000110", -- t[38918] = 5
      "0000101" when "01001100000000111", -- t[38919] = 5
      "0000101" when "01001100000001000", -- t[38920] = 5
      "0000101" when "01001100000001001", -- t[38921] = 5
      "0000101" when "01001100000001010", -- t[38922] = 5
      "0000101" when "01001100000001011", -- t[38923] = 5
      "0000101" when "01001100000001100", -- t[38924] = 5
      "0000101" when "01001100000001101", -- t[38925] = 5
      "0000101" when "01001100000001110", -- t[38926] = 5
      "0000101" when "01001100000001111", -- t[38927] = 5
      "0000101" when "01001100000010000", -- t[38928] = 5
      "0000101" when "01001100000010001", -- t[38929] = 5
      "0000101" when "01001100000010010", -- t[38930] = 5
      "0000101" when "01001100000010011", -- t[38931] = 5
      "0000101" when "01001100000010100", -- t[38932] = 5
      "0000101" when "01001100000010101", -- t[38933] = 5
      "0000101" when "01001100000010110", -- t[38934] = 5
      "0000101" when "01001100000010111", -- t[38935] = 5
      "0000101" when "01001100000011000", -- t[38936] = 5
      "0000101" when "01001100000011001", -- t[38937] = 5
      "0000101" when "01001100000011010", -- t[38938] = 5
      "0000101" when "01001100000011011", -- t[38939] = 5
      "0000101" when "01001100000011100", -- t[38940] = 5
      "0000101" when "01001100000011101", -- t[38941] = 5
      "0000101" when "01001100000011110", -- t[38942] = 5
      "0000101" when "01001100000011111", -- t[38943] = 5
      "0000101" when "01001100000100000", -- t[38944] = 5
      "0000101" when "01001100000100001", -- t[38945] = 5
      "0000101" when "01001100000100010", -- t[38946] = 5
      "0000101" when "01001100000100011", -- t[38947] = 5
      "0000101" when "01001100000100100", -- t[38948] = 5
      "0000101" when "01001100000100101", -- t[38949] = 5
      "0000101" when "01001100000100110", -- t[38950] = 5
      "0000101" when "01001100000100111", -- t[38951] = 5
      "0000101" when "01001100000101000", -- t[38952] = 5
      "0000101" when "01001100000101001", -- t[38953] = 5
      "0000101" when "01001100000101010", -- t[38954] = 5
      "0000101" when "01001100000101011", -- t[38955] = 5
      "0000101" when "01001100000101100", -- t[38956] = 5
      "0000101" when "01001100000101101", -- t[38957] = 5
      "0000101" when "01001100000101110", -- t[38958] = 5
      "0000101" when "01001100000101111", -- t[38959] = 5
      "0000101" when "01001100000110000", -- t[38960] = 5
      "0000101" when "01001100000110001", -- t[38961] = 5
      "0000101" when "01001100000110010", -- t[38962] = 5
      "0000101" when "01001100000110011", -- t[38963] = 5
      "0000101" when "01001100000110100", -- t[38964] = 5
      "0000101" when "01001100000110101", -- t[38965] = 5
      "0000101" when "01001100000110110", -- t[38966] = 5
      "0000101" when "01001100000110111", -- t[38967] = 5
      "0000101" when "01001100000111000", -- t[38968] = 5
      "0000101" when "01001100000111001", -- t[38969] = 5
      "0000101" when "01001100000111010", -- t[38970] = 5
      "0000101" when "01001100000111011", -- t[38971] = 5
      "0000101" when "01001100000111100", -- t[38972] = 5
      "0000101" when "01001100000111101", -- t[38973] = 5
      "0000101" when "01001100000111110", -- t[38974] = 5
      "0000101" when "01001100000111111", -- t[38975] = 5
      "0000101" when "01001100001000000", -- t[38976] = 5
      "0000101" when "01001100001000001", -- t[38977] = 5
      "0000101" when "01001100001000010", -- t[38978] = 5
      "0000101" when "01001100001000011", -- t[38979] = 5
      "0000101" when "01001100001000100", -- t[38980] = 5
      "0000101" when "01001100001000101", -- t[38981] = 5
      "0000101" when "01001100001000110", -- t[38982] = 5
      "0000101" when "01001100001000111", -- t[38983] = 5
      "0000101" when "01001100001001000", -- t[38984] = 5
      "0000101" when "01001100001001001", -- t[38985] = 5
      "0000101" when "01001100001001010", -- t[38986] = 5
      "0000101" when "01001100001001011", -- t[38987] = 5
      "0000101" when "01001100001001100", -- t[38988] = 5
      "0000101" when "01001100001001101", -- t[38989] = 5
      "0000101" when "01001100001001110", -- t[38990] = 5
      "0000101" when "01001100001001111", -- t[38991] = 5
      "0000101" when "01001100001010000", -- t[38992] = 5
      "0000101" when "01001100001010001", -- t[38993] = 5
      "0000101" when "01001100001010010", -- t[38994] = 5
      "0000101" when "01001100001010011", -- t[38995] = 5
      "0000101" when "01001100001010100", -- t[38996] = 5
      "0000101" when "01001100001010101", -- t[38997] = 5
      "0000101" when "01001100001010110", -- t[38998] = 5
      "0000101" when "01001100001010111", -- t[38999] = 5
      "0000101" when "01001100001011000", -- t[39000] = 5
      "0000101" when "01001100001011001", -- t[39001] = 5
      "0000101" when "01001100001011010", -- t[39002] = 5
      "0000101" when "01001100001011011", -- t[39003] = 5
      "0000101" when "01001100001011100", -- t[39004] = 5
      "0000101" when "01001100001011101", -- t[39005] = 5
      "0000101" when "01001100001011110", -- t[39006] = 5
      "0000101" when "01001100001011111", -- t[39007] = 5
      "0000101" when "01001100001100000", -- t[39008] = 5
      "0000101" when "01001100001100001", -- t[39009] = 5
      "0000101" when "01001100001100010", -- t[39010] = 5
      "0000101" when "01001100001100011", -- t[39011] = 5
      "0000101" when "01001100001100100", -- t[39012] = 5
      "0000101" when "01001100001100101", -- t[39013] = 5
      "0000101" when "01001100001100110", -- t[39014] = 5
      "0000101" when "01001100001100111", -- t[39015] = 5
      "0000101" when "01001100001101000", -- t[39016] = 5
      "0000101" when "01001100001101001", -- t[39017] = 5
      "0000101" when "01001100001101010", -- t[39018] = 5
      "0000101" when "01001100001101011", -- t[39019] = 5
      "0000101" when "01001100001101100", -- t[39020] = 5
      "0000101" when "01001100001101101", -- t[39021] = 5
      "0000101" when "01001100001101110", -- t[39022] = 5
      "0000101" when "01001100001101111", -- t[39023] = 5
      "0000101" when "01001100001110000", -- t[39024] = 5
      "0000101" when "01001100001110001", -- t[39025] = 5
      "0000101" when "01001100001110010", -- t[39026] = 5
      "0000101" when "01001100001110011", -- t[39027] = 5
      "0000101" when "01001100001110100", -- t[39028] = 5
      "0000101" when "01001100001110101", -- t[39029] = 5
      "0000101" when "01001100001110110", -- t[39030] = 5
      "0000101" when "01001100001110111", -- t[39031] = 5
      "0000101" when "01001100001111000", -- t[39032] = 5
      "0000101" when "01001100001111001", -- t[39033] = 5
      "0000101" when "01001100001111010", -- t[39034] = 5
      "0000101" when "01001100001111011", -- t[39035] = 5
      "0000101" when "01001100001111100", -- t[39036] = 5
      "0000101" when "01001100001111101", -- t[39037] = 5
      "0000101" when "01001100001111110", -- t[39038] = 5
      "0000101" when "01001100001111111", -- t[39039] = 5
      "0000101" when "01001100010000000", -- t[39040] = 5
      "0000101" when "01001100010000001", -- t[39041] = 5
      "0000101" when "01001100010000010", -- t[39042] = 5
      "0000101" when "01001100010000011", -- t[39043] = 5
      "0000101" when "01001100010000100", -- t[39044] = 5
      "0000101" when "01001100010000101", -- t[39045] = 5
      "0000101" when "01001100010000110", -- t[39046] = 5
      "0000101" when "01001100010000111", -- t[39047] = 5
      "0000101" when "01001100010001000", -- t[39048] = 5
      "0000101" when "01001100010001001", -- t[39049] = 5
      "0000101" when "01001100010001010", -- t[39050] = 5
      "0000101" when "01001100010001011", -- t[39051] = 5
      "0000101" when "01001100010001100", -- t[39052] = 5
      "0000101" when "01001100010001101", -- t[39053] = 5
      "0000101" when "01001100010001110", -- t[39054] = 5
      "0000101" when "01001100010001111", -- t[39055] = 5
      "0000101" when "01001100010010000", -- t[39056] = 5
      "0000101" when "01001100010010001", -- t[39057] = 5
      "0000101" when "01001100010010010", -- t[39058] = 5
      "0000101" when "01001100010010011", -- t[39059] = 5
      "0000101" when "01001100010010100", -- t[39060] = 5
      "0000101" when "01001100010010101", -- t[39061] = 5
      "0000101" when "01001100010010110", -- t[39062] = 5
      "0000101" when "01001100010010111", -- t[39063] = 5
      "0000101" when "01001100010011000", -- t[39064] = 5
      "0000101" when "01001100010011001", -- t[39065] = 5
      "0000101" when "01001100010011010", -- t[39066] = 5
      "0000101" when "01001100010011011", -- t[39067] = 5
      "0000101" when "01001100010011100", -- t[39068] = 5
      "0000101" when "01001100010011101", -- t[39069] = 5
      "0000101" when "01001100010011110", -- t[39070] = 5
      "0000101" when "01001100010011111", -- t[39071] = 5
      "0000101" when "01001100010100000", -- t[39072] = 5
      "0000101" when "01001100010100001", -- t[39073] = 5
      "0000101" when "01001100010100010", -- t[39074] = 5
      "0000101" when "01001100010100011", -- t[39075] = 5
      "0000101" when "01001100010100100", -- t[39076] = 5
      "0000101" when "01001100010100101", -- t[39077] = 5
      "0000101" when "01001100010100110", -- t[39078] = 5
      "0000101" when "01001100010100111", -- t[39079] = 5
      "0000101" when "01001100010101000", -- t[39080] = 5
      "0000101" when "01001100010101001", -- t[39081] = 5
      "0000101" when "01001100010101010", -- t[39082] = 5
      "0000101" when "01001100010101011", -- t[39083] = 5
      "0000101" when "01001100010101100", -- t[39084] = 5
      "0000101" when "01001100010101101", -- t[39085] = 5
      "0000101" when "01001100010101110", -- t[39086] = 5
      "0000101" when "01001100010101111", -- t[39087] = 5
      "0000101" when "01001100010110000", -- t[39088] = 5
      "0000101" when "01001100010110001", -- t[39089] = 5
      "0000101" when "01001100010110010", -- t[39090] = 5
      "0000101" when "01001100010110011", -- t[39091] = 5
      "0000101" when "01001100010110100", -- t[39092] = 5
      "0000101" when "01001100010110101", -- t[39093] = 5
      "0000101" when "01001100010110110", -- t[39094] = 5
      "0000101" when "01001100010110111", -- t[39095] = 5
      "0000101" when "01001100010111000", -- t[39096] = 5
      "0000101" when "01001100010111001", -- t[39097] = 5
      "0000101" when "01001100010111010", -- t[39098] = 5
      "0000101" when "01001100010111011", -- t[39099] = 5
      "0000101" when "01001100010111100", -- t[39100] = 5
      "0000101" when "01001100010111101", -- t[39101] = 5
      "0000101" when "01001100010111110", -- t[39102] = 5
      "0000101" when "01001100010111111", -- t[39103] = 5
      "0000101" when "01001100011000000", -- t[39104] = 5
      "0000101" when "01001100011000001", -- t[39105] = 5
      "0000101" when "01001100011000010", -- t[39106] = 5
      "0000101" when "01001100011000011", -- t[39107] = 5
      "0000101" when "01001100011000100", -- t[39108] = 5
      "0000101" when "01001100011000101", -- t[39109] = 5
      "0000101" when "01001100011000110", -- t[39110] = 5
      "0000101" when "01001100011000111", -- t[39111] = 5
      "0000101" when "01001100011001000", -- t[39112] = 5
      "0000101" when "01001100011001001", -- t[39113] = 5
      "0000101" when "01001100011001010", -- t[39114] = 5
      "0000101" when "01001100011001011", -- t[39115] = 5
      "0000101" when "01001100011001100", -- t[39116] = 5
      "0000101" when "01001100011001101", -- t[39117] = 5
      "0000101" when "01001100011001110", -- t[39118] = 5
      "0000101" when "01001100011001111", -- t[39119] = 5
      "0000101" when "01001100011010000", -- t[39120] = 5
      "0000101" when "01001100011010001", -- t[39121] = 5
      "0000101" when "01001100011010010", -- t[39122] = 5
      "0000101" when "01001100011010011", -- t[39123] = 5
      "0000101" when "01001100011010100", -- t[39124] = 5
      "0000101" when "01001100011010101", -- t[39125] = 5
      "0000101" when "01001100011010110", -- t[39126] = 5
      "0000101" when "01001100011010111", -- t[39127] = 5
      "0000101" when "01001100011011000", -- t[39128] = 5
      "0000101" when "01001100011011001", -- t[39129] = 5
      "0000101" when "01001100011011010", -- t[39130] = 5
      "0000101" when "01001100011011011", -- t[39131] = 5
      "0000101" when "01001100011011100", -- t[39132] = 5
      "0000101" when "01001100011011101", -- t[39133] = 5
      "0000101" when "01001100011011110", -- t[39134] = 5
      "0000101" when "01001100011011111", -- t[39135] = 5
      "0000101" when "01001100011100000", -- t[39136] = 5
      "0000101" when "01001100011100001", -- t[39137] = 5
      "0000101" when "01001100011100010", -- t[39138] = 5
      "0000101" when "01001100011100011", -- t[39139] = 5
      "0000101" when "01001100011100100", -- t[39140] = 5
      "0000101" when "01001100011100101", -- t[39141] = 5
      "0000101" when "01001100011100110", -- t[39142] = 5
      "0000101" when "01001100011100111", -- t[39143] = 5
      "0000101" when "01001100011101000", -- t[39144] = 5
      "0000101" when "01001100011101001", -- t[39145] = 5
      "0000101" when "01001100011101010", -- t[39146] = 5
      "0000101" when "01001100011101011", -- t[39147] = 5
      "0000101" when "01001100011101100", -- t[39148] = 5
      "0000101" when "01001100011101101", -- t[39149] = 5
      "0000101" when "01001100011101110", -- t[39150] = 5
      "0000101" when "01001100011101111", -- t[39151] = 5
      "0000101" when "01001100011110000", -- t[39152] = 5
      "0000101" when "01001100011110001", -- t[39153] = 5
      "0000101" when "01001100011110010", -- t[39154] = 5
      "0000101" when "01001100011110011", -- t[39155] = 5
      "0000101" when "01001100011110100", -- t[39156] = 5
      "0000101" when "01001100011110101", -- t[39157] = 5
      "0000101" when "01001100011110110", -- t[39158] = 5
      "0000101" when "01001100011110111", -- t[39159] = 5
      "0000101" when "01001100011111000", -- t[39160] = 5
      "0000101" when "01001100011111001", -- t[39161] = 5
      "0000101" when "01001100011111010", -- t[39162] = 5
      "0000101" when "01001100011111011", -- t[39163] = 5
      "0000101" when "01001100011111100", -- t[39164] = 5
      "0000101" when "01001100011111101", -- t[39165] = 5
      "0000101" when "01001100011111110", -- t[39166] = 5
      "0000101" when "01001100011111111", -- t[39167] = 5
      "0000101" when "01001100100000000", -- t[39168] = 5
      "0000101" when "01001100100000001", -- t[39169] = 5
      "0000101" when "01001100100000010", -- t[39170] = 5
      "0000101" when "01001100100000011", -- t[39171] = 5
      "0000101" when "01001100100000100", -- t[39172] = 5
      "0000101" when "01001100100000101", -- t[39173] = 5
      "0000101" when "01001100100000110", -- t[39174] = 5
      "0000101" when "01001100100000111", -- t[39175] = 5
      "0000101" when "01001100100001000", -- t[39176] = 5
      "0000101" when "01001100100001001", -- t[39177] = 5
      "0000101" when "01001100100001010", -- t[39178] = 5
      "0000101" when "01001100100001011", -- t[39179] = 5
      "0000101" when "01001100100001100", -- t[39180] = 5
      "0000101" when "01001100100001101", -- t[39181] = 5
      "0000101" when "01001100100001110", -- t[39182] = 5
      "0000101" when "01001100100001111", -- t[39183] = 5
      "0000101" when "01001100100010000", -- t[39184] = 5
      "0000101" when "01001100100010001", -- t[39185] = 5
      "0000101" when "01001100100010010", -- t[39186] = 5
      "0000101" when "01001100100010011", -- t[39187] = 5
      "0000101" when "01001100100010100", -- t[39188] = 5
      "0000101" when "01001100100010101", -- t[39189] = 5
      "0000101" when "01001100100010110", -- t[39190] = 5
      "0000101" when "01001100100010111", -- t[39191] = 5
      "0000101" when "01001100100011000", -- t[39192] = 5
      "0000101" when "01001100100011001", -- t[39193] = 5
      "0000101" when "01001100100011010", -- t[39194] = 5
      "0000101" when "01001100100011011", -- t[39195] = 5
      "0000101" when "01001100100011100", -- t[39196] = 5
      "0000101" when "01001100100011101", -- t[39197] = 5
      "0000101" when "01001100100011110", -- t[39198] = 5
      "0000101" when "01001100100011111", -- t[39199] = 5
      "0000101" when "01001100100100000", -- t[39200] = 5
      "0000101" when "01001100100100001", -- t[39201] = 5
      "0000101" when "01001100100100010", -- t[39202] = 5
      "0000101" when "01001100100100011", -- t[39203] = 5
      "0000101" when "01001100100100100", -- t[39204] = 5
      "0000101" when "01001100100100101", -- t[39205] = 5
      "0000101" when "01001100100100110", -- t[39206] = 5
      "0000101" when "01001100100100111", -- t[39207] = 5
      "0000101" when "01001100100101000", -- t[39208] = 5
      "0000101" when "01001100100101001", -- t[39209] = 5
      "0000101" when "01001100100101010", -- t[39210] = 5
      "0000101" when "01001100100101011", -- t[39211] = 5
      "0000101" when "01001100100101100", -- t[39212] = 5
      "0000101" when "01001100100101101", -- t[39213] = 5
      "0000101" when "01001100100101110", -- t[39214] = 5
      "0000101" when "01001100100101111", -- t[39215] = 5
      "0000101" when "01001100100110000", -- t[39216] = 5
      "0000101" when "01001100100110001", -- t[39217] = 5
      "0000101" when "01001100100110010", -- t[39218] = 5
      "0000101" when "01001100100110011", -- t[39219] = 5
      "0000101" when "01001100100110100", -- t[39220] = 5
      "0000101" when "01001100100110101", -- t[39221] = 5
      "0000101" when "01001100100110110", -- t[39222] = 5
      "0000101" when "01001100100110111", -- t[39223] = 5
      "0000101" when "01001100100111000", -- t[39224] = 5
      "0000101" when "01001100100111001", -- t[39225] = 5
      "0000101" when "01001100100111010", -- t[39226] = 5
      "0000101" when "01001100100111011", -- t[39227] = 5
      "0000101" when "01001100100111100", -- t[39228] = 5
      "0000101" when "01001100100111101", -- t[39229] = 5
      "0000101" when "01001100100111110", -- t[39230] = 5
      "0000101" when "01001100100111111", -- t[39231] = 5
      "0000101" when "01001100101000000", -- t[39232] = 5
      "0000101" when "01001100101000001", -- t[39233] = 5
      "0000101" when "01001100101000010", -- t[39234] = 5
      "0000101" when "01001100101000011", -- t[39235] = 5
      "0000101" when "01001100101000100", -- t[39236] = 5
      "0000101" when "01001100101000101", -- t[39237] = 5
      "0000101" when "01001100101000110", -- t[39238] = 5
      "0000101" when "01001100101000111", -- t[39239] = 5
      "0000101" when "01001100101001000", -- t[39240] = 5
      "0000101" when "01001100101001001", -- t[39241] = 5
      "0000101" when "01001100101001010", -- t[39242] = 5
      "0000101" when "01001100101001011", -- t[39243] = 5
      "0000101" when "01001100101001100", -- t[39244] = 5
      "0000101" when "01001100101001101", -- t[39245] = 5
      "0000101" when "01001100101001110", -- t[39246] = 5
      "0000101" when "01001100101001111", -- t[39247] = 5
      "0000101" when "01001100101010000", -- t[39248] = 5
      "0000101" when "01001100101010001", -- t[39249] = 5
      "0000101" when "01001100101010010", -- t[39250] = 5
      "0000101" when "01001100101010011", -- t[39251] = 5
      "0000101" when "01001100101010100", -- t[39252] = 5
      "0000101" when "01001100101010101", -- t[39253] = 5
      "0000101" when "01001100101010110", -- t[39254] = 5
      "0000101" when "01001100101010111", -- t[39255] = 5
      "0000101" when "01001100101011000", -- t[39256] = 5
      "0000101" when "01001100101011001", -- t[39257] = 5
      "0000101" when "01001100101011010", -- t[39258] = 5
      "0000101" when "01001100101011011", -- t[39259] = 5
      "0000101" when "01001100101011100", -- t[39260] = 5
      "0000101" when "01001100101011101", -- t[39261] = 5
      "0000101" when "01001100101011110", -- t[39262] = 5
      "0000101" when "01001100101011111", -- t[39263] = 5
      "0000101" when "01001100101100000", -- t[39264] = 5
      "0000101" when "01001100101100001", -- t[39265] = 5
      "0000101" when "01001100101100010", -- t[39266] = 5
      "0000101" when "01001100101100011", -- t[39267] = 5
      "0000101" when "01001100101100100", -- t[39268] = 5
      "0000101" when "01001100101100101", -- t[39269] = 5
      "0000101" when "01001100101100110", -- t[39270] = 5
      "0000101" when "01001100101100111", -- t[39271] = 5
      "0000101" when "01001100101101000", -- t[39272] = 5
      "0000101" when "01001100101101001", -- t[39273] = 5
      "0000101" when "01001100101101010", -- t[39274] = 5
      "0000101" when "01001100101101011", -- t[39275] = 5
      "0000101" when "01001100101101100", -- t[39276] = 5
      "0000101" when "01001100101101101", -- t[39277] = 5
      "0000101" when "01001100101101110", -- t[39278] = 5
      "0000101" when "01001100101101111", -- t[39279] = 5
      "0000101" when "01001100101110000", -- t[39280] = 5
      "0000101" when "01001100101110001", -- t[39281] = 5
      "0000101" when "01001100101110010", -- t[39282] = 5
      "0000101" when "01001100101110011", -- t[39283] = 5
      "0000101" when "01001100101110100", -- t[39284] = 5
      "0000101" when "01001100101110101", -- t[39285] = 5
      "0000101" when "01001100101110110", -- t[39286] = 5
      "0000101" when "01001100101110111", -- t[39287] = 5
      "0000101" when "01001100101111000", -- t[39288] = 5
      "0000101" when "01001100101111001", -- t[39289] = 5
      "0000101" when "01001100101111010", -- t[39290] = 5
      "0000101" when "01001100101111011", -- t[39291] = 5
      "0000101" when "01001100101111100", -- t[39292] = 5
      "0000101" when "01001100101111101", -- t[39293] = 5
      "0000101" when "01001100101111110", -- t[39294] = 5
      "0000101" when "01001100101111111", -- t[39295] = 5
      "0000101" when "01001100110000000", -- t[39296] = 5
      "0000101" when "01001100110000001", -- t[39297] = 5
      "0000101" when "01001100110000010", -- t[39298] = 5
      "0000101" when "01001100110000011", -- t[39299] = 5
      "0000101" when "01001100110000100", -- t[39300] = 5
      "0000101" when "01001100110000101", -- t[39301] = 5
      "0000101" when "01001100110000110", -- t[39302] = 5
      "0000101" when "01001100110000111", -- t[39303] = 5
      "0000101" when "01001100110001000", -- t[39304] = 5
      "0000101" when "01001100110001001", -- t[39305] = 5
      "0000101" when "01001100110001010", -- t[39306] = 5
      "0000101" when "01001100110001011", -- t[39307] = 5
      "0000101" when "01001100110001100", -- t[39308] = 5
      "0000101" when "01001100110001101", -- t[39309] = 5
      "0000101" when "01001100110001110", -- t[39310] = 5
      "0000101" when "01001100110001111", -- t[39311] = 5
      "0000101" when "01001100110010000", -- t[39312] = 5
      "0000101" when "01001100110010001", -- t[39313] = 5
      "0000101" when "01001100110010010", -- t[39314] = 5
      "0000101" when "01001100110010011", -- t[39315] = 5
      "0000101" when "01001100110010100", -- t[39316] = 5
      "0000101" when "01001100110010101", -- t[39317] = 5
      "0000101" when "01001100110010110", -- t[39318] = 5
      "0000101" when "01001100110010111", -- t[39319] = 5
      "0000101" when "01001100110011000", -- t[39320] = 5
      "0000101" when "01001100110011001", -- t[39321] = 5
      "0000101" when "01001100110011010", -- t[39322] = 5
      "0000101" when "01001100110011011", -- t[39323] = 5
      "0000101" when "01001100110011100", -- t[39324] = 5
      "0000101" when "01001100110011101", -- t[39325] = 5
      "0000101" when "01001100110011110", -- t[39326] = 5
      "0000101" when "01001100110011111", -- t[39327] = 5
      "0000101" when "01001100110100000", -- t[39328] = 5
      "0000101" when "01001100110100001", -- t[39329] = 5
      "0000101" when "01001100110100010", -- t[39330] = 5
      "0000101" when "01001100110100011", -- t[39331] = 5
      "0000101" when "01001100110100100", -- t[39332] = 5
      "0000101" when "01001100110100101", -- t[39333] = 5
      "0000101" when "01001100110100110", -- t[39334] = 5
      "0000101" when "01001100110100111", -- t[39335] = 5
      "0000101" when "01001100110101000", -- t[39336] = 5
      "0000101" when "01001100110101001", -- t[39337] = 5
      "0000101" when "01001100110101010", -- t[39338] = 5
      "0000101" when "01001100110101011", -- t[39339] = 5
      "0000101" when "01001100110101100", -- t[39340] = 5
      "0000101" when "01001100110101101", -- t[39341] = 5
      "0000101" when "01001100110101110", -- t[39342] = 5
      "0000101" when "01001100110101111", -- t[39343] = 5
      "0000101" when "01001100110110000", -- t[39344] = 5
      "0000101" when "01001100110110001", -- t[39345] = 5
      "0000101" when "01001100110110010", -- t[39346] = 5
      "0000101" when "01001100110110011", -- t[39347] = 5
      "0000101" when "01001100110110100", -- t[39348] = 5
      "0000101" when "01001100110110101", -- t[39349] = 5
      "0000101" when "01001100110110110", -- t[39350] = 5
      "0000101" when "01001100110110111", -- t[39351] = 5
      "0000101" when "01001100110111000", -- t[39352] = 5
      "0000101" when "01001100110111001", -- t[39353] = 5
      "0000101" when "01001100110111010", -- t[39354] = 5
      "0000101" when "01001100110111011", -- t[39355] = 5
      "0000101" when "01001100110111100", -- t[39356] = 5
      "0000101" when "01001100110111101", -- t[39357] = 5
      "0000101" when "01001100110111110", -- t[39358] = 5
      "0000101" when "01001100110111111", -- t[39359] = 5
      "0000101" when "01001100111000000", -- t[39360] = 5
      "0000101" when "01001100111000001", -- t[39361] = 5
      "0000101" when "01001100111000010", -- t[39362] = 5
      "0000101" when "01001100111000011", -- t[39363] = 5
      "0000101" when "01001100111000100", -- t[39364] = 5
      "0000101" when "01001100111000101", -- t[39365] = 5
      "0000101" when "01001100111000110", -- t[39366] = 5
      "0000101" when "01001100111000111", -- t[39367] = 5
      "0000101" when "01001100111001000", -- t[39368] = 5
      "0000101" when "01001100111001001", -- t[39369] = 5
      "0000101" when "01001100111001010", -- t[39370] = 5
      "0000101" when "01001100111001011", -- t[39371] = 5
      "0000101" when "01001100111001100", -- t[39372] = 5
      "0000101" when "01001100111001101", -- t[39373] = 5
      "0000101" when "01001100111001110", -- t[39374] = 5
      "0000101" when "01001100111001111", -- t[39375] = 5
      "0000101" when "01001100111010000", -- t[39376] = 5
      "0000101" when "01001100111010001", -- t[39377] = 5
      "0000101" when "01001100111010010", -- t[39378] = 5
      "0000101" when "01001100111010011", -- t[39379] = 5
      "0000101" when "01001100111010100", -- t[39380] = 5
      "0000101" when "01001100111010101", -- t[39381] = 5
      "0000101" when "01001100111010110", -- t[39382] = 5
      "0000101" when "01001100111010111", -- t[39383] = 5
      "0000101" when "01001100111011000", -- t[39384] = 5
      "0000101" when "01001100111011001", -- t[39385] = 5
      "0000101" when "01001100111011010", -- t[39386] = 5
      "0000101" when "01001100111011011", -- t[39387] = 5
      "0000101" when "01001100111011100", -- t[39388] = 5
      "0000101" when "01001100111011101", -- t[39389] = 5
      "0000101" when "01001100111011110", -- t[39390] = 5
      "0000101" when "01001100111011111", -- t[39391] = 5
      "0000101" when "01001100111100000", -- t[39392] = 5
      "0000101" when "01001100111100001", -- t[39393] = 5
      "0000101" when "01001100111100010", -- t[39394] = 5
      "0000101" when "01001100111100011", -- t[39395] = 5
      "0000101" when "01001100111100100", -- t[39396] = 5
      "0000101" when "01001100111100101", -- t[39397] = 5
      "0000101" when "01001100111100110", -- t[39398] = 5
      "0000101" when "01001100111100111", -- t[39399] = 5
      "0000101" when "01001100111101000", -- t[39400] = 5
      "0000101" when "01001100111101001", -- t[39401] = 5
      "0000101" when "01001100111101010", -- t[39402] = 5
      "0000101" when "01001100111101011", -- t[39403] = 5
      "0000101" when "01001100111101100", -- t[39404] = 5
      "0000101" when "01001100111101101", -- t[39405] = 5
      "0000101" when "01001100111101110", -- t[39406] = 5
      "0000101" when "01001100111101111", -- t[39407] = 5
      "0000101" when "01001100111110000", -- t[39408] = 5
      "0000101" when "01001100111110001", -- t[39409] = 5
      "0000101" when "01001100111110010", -- t[39410] = 5
      "0000101" when "01001100111110011", -- t[39411] = 5
      "0000101" when "01001100111110100", -- t[39412] = 5
      "0000101" when "01001100111110101", -- t[39413] = 5
      "0000101" when "01001100111110110", -- t[39414] = 5
      "0000101" when "01001100111110111", -- t[39415] = 5
      "0000101" when "01001100111111000", -- t[39416] = 5
      "0000101" when "01001100111111001", -- t[39417] = 5
      "0000101" when "01001100111111010", -- t[39418] = 5
      "0000101" when "01001100111111011", -- t[39419] = 5
      "0000101" when "01001100111111100", -- t[39420] = 5
      "0000101" when "01001100111111101", -- t[39421] = 5
      "0000101" when "01001100111111110", -- t[39422] = 5
      "0000101" when "01001100111111111", -- t[39423] = 5
      "0000101" when "01001101000000000", -- t[39424] = 5
      "0000101" when "01001101000000001", -- t[39425] = 5
      "0000101" when "01001101000000010", -- t[39426] = 5
      "0000101" when "01001101000000011", -- t[39427] = 5
      "0000101" when "01001101000000100", -- t[39428] = 5
      "0000101" when "01001101000000101", -- t[39429] = 5
      "0000101" when "01001101000000110", -- t[39430] = 5
      "0000101" when "01001101000000111", -- t[39431] = 5
      "0000101" when "01001101000001000", -- t[39432] = 5
      "0000101" when "01001101000001001", -- t[39433] = 5
      "0000101" when "01001101000001010", -- t[39434] = 5
      "0000101" when "01001101000001011", -- t[39435] = 5
      "0000101" when "01001101000001100", -- t[39436] = 5
      "0000101" when "01001101000001101", -- t[39437] = 5
      "0000101" when "01001101000001110", -- t[39438] = 5
      "0000101" when "01001101000001111", -- t[39439] = 5
      "0000101" when "01001101000010000", -- t[39440] = 5
      "0000101" when "01001101000010001", -- t[39441] = 5
      "0000101" when "01001101000010010", -- t[39442] = 5
      "0000101" when "01001101000010011", -- t[39443] = 5
      "0000101" when "01001101000010100", -- t[39444] = 5
      "0000101" when "01001101000010101", -- t[39445] = 5
      "0000101" when "01001101000010110", -- t[39446] = 5
      "0000101" when "01001101000010111", -- t[39447] = 5
      "0000101" when "01001101000011000", -- t[39448] = 5
      "0000101" when "01001101000011001", -- t[39449] = 5
      "0000101" when "01001101000011010", -- t[39450] = 5
      "0000101" when "01001101000011011", -- t[39451] = 5
      "0000101" when "01001101000011100", -- t[39452] = 5
      "0000101" when "01001101000011101", -- t[39453] = 5
      "0000101" when "01001101000011110", -- t[39454] = 5
      "0000101" when "01001101000011111", -- t[39455] = 5
      "0000101" when "01001101000100000", -- t[39456] = 5
      "0000101" when "01001101000100001", -- t[39457] = 5
      "0000101" when "01001101000100010", -- t[39458] = 5
      "0000101" when "01001101000100011", -- t[39459] = 5
      "0000101" when "01001101000100100", -- t[39460] = 5
      "0000101" when "01001101000100101", -- t[39461] = 5
      "0000101" when "01001101000100110", -- t[39462] = 5
      "0000101" when "01001101000100111", -- t[39463] = 5
      "0000101" when "01001101000101000", -- t[39464] = 5
      "0000101" when "01001101000101001", -- t[39465] = 5
      "0000101" when "01001101000101010", -- t[39466] = 5
      "0000101" when "01001101000101011", -- t[39467] = 5
      "0000101" when "01001101000101100", -- t[39468] = 5
      "0000101" when "01001101000101101", -- t[39469] = 5
      "0000101" when "01001101000101110", -- t[39470] = 5
      "0000101" when "01001101000101111", -- t[39471] = 5
      "0000101" when "01001101000110000", -- t[39472] = 5
      "0000101" when "01001101000110001", -- t[39473] = 5
      "0000101" when "01001101000110010", -- t[39474] = 5
      "0000101" when "01001101000110011", -- t[39475] = 5
      "0000101" when "01001101000110100", -- t[39476] = 5
      "0000101" when "01001101000110101", -- t[39477] = 5
      "0000101" when "01001101000110110", -- t[39478] = 5
      "0000101" when "01001101000110111", -- t[39479] = 5
      "0000101" when "01001101000111000", -- t[39480] = 5
      "0000101" when "01001101000111001", -- t[39481] = 5
      "0000101" when "01001101000111010", -- t[39482] = 5
      "0000101" when "01001101000111011", -- t[39483] = 5
      "0000101" when "01001101000111100", -- t[39484] = 5
      "0000101" when "01001101000111101", -- t[39485] = 5
      "0000101" when "01001101000111110", -- t[39486] = 5
      "0000101" when "01001101000111111", -- t[39487] = 5
      "0000101" when "01001101001000000", -- t[39488] = 5
      "0000101" when "01001101001000001", -- t[39489] = 5
      "0000101" when "01001101001000010", -- t[39490] = 5
      "0000101" when "01001101001000011", -- t[39491] = 5
      "0000101" when "01001101001000100", -- t[39492] = 5
      "0000101" when "01001101001000101", -- t[39493] = 5
      "0000101" when "01001101001000110", -- t[39494] = 5
      "0000101" when "01001101001000111", -- t[39495] = 5
      "0000101" when "01001101001001000", -- t[39496] = 5
      "0000101" when "01001101001001001", -- t[39497] = 5
      "0000101" when "01001101001001010", -- t[39498] = 5
      "0000101" when "01001101001001011", -- t[39499] = 5
      "0000101" when "01001101001001100", -- t[39500] = 5
      "0000101" when "01001101001001101", -- t[39501] = 5
      "0000101" when "01001101001001110", -- t[39502] = 5
      "0000101" when "01001101001001111", -- t[39503] = 5
      "0000101" when "01001101001010000", -- t[39504] = 5
      "0000101" when "01001101001010001", -- t[39505] = 5
      "0000101" when "01001101001010010", -- t[39506] = 5
      "0000101" when "01001101001010011", -- t[39507] = 5
      "0000101" when "01001101001010100", -- t[39508] = 5
      "0000101" when "01001101001010101", -- t[39509] = 5
      "0000101" when "01001101001010110", -- t[39510] = 5
      "0000101" when "01001101001010111", -- t[39511] = 5
      "0000101" when "01001101001011000", -- t[39512] = 5
      "0000101" when "01001101001011001", -- t[39513] = 5
      "0000101" when "01001101001011010", -- t[39514] = 5
      "0000101" when "01001101001011011", -- t[39515] = 5
      "0000101" when "01001101001011100", -- t[39516] = 5
      "0000101" when "01001101001011101", -- t[39517] = 5
      "0000101" when "01001101001011110", -- t[39518] = 5
      "0000101" when "01001101001011111", -- t[39519] = 5
      "0000101" when "01001101001100000", -- t[39520] = 5
      "0000101" when "01001101001100001", -- t[39521] = 5
      "0000101" when "01001101001100010", -- t[39522] = 5
      "0000101" when "01001101001100011", -- t[39523] = 5
      "0000101" when "01001101001100100", -- t[39524] = 5
      "0000101" when "01001101001100101", -- t[39525] = 5
      "0000101" when "01001101001100110", -- t[39526] = 5
      "0000101" when "01001101001100111", -- t[39527] = 5
      "0000101" when "01001101001101000", -- t[39528] = 5
      "0000101" when "01001101001101001", -- t[39529] = 5
      "0000101" when "01001101001101010", -- t[39530] = 5
      "0000101" when "01001101001101011", -- t[39531] = 5
      "0000101" when "01001101001101100", -- t[39532] = 5
      "0000101" when "01001101001101101", -- t[39533] = 5
      "0000101" when "01001101001101110", -- t[39534] = 5
      "0000101" when "01001101001101111", -- t[39535] = 5
      "0000101" when "01001101001110000", -- t[39536] = 5
      "0000101" when "01001101001110001", -- t[39537] = 5
      "0000101" when "01001101001110010", -- t[39538] = 5
      "0000101" when "01001101001110011", -- t[39539] = 5
      "0000101" when "01001101001110100", -- t[39540] = 5
      "0000101" when "01001101001110101", -- t[39541] = 5
      "0000101" when "01001101001110110", -- t[39542] = 5
      "0000101" when "01001101001110111", -- t[39543] = 5
      "0000101" when "01001101001111000", -- t[39544] = 5
      "0000101" when "01001101001111001", -- t[39545] = 5
      "0000101" when "01001101001111010", -- t[39546] = 5
      "0000101" when "01001101001111011", -- t[39547] = 5
      "0000101" when "01001101001111100", -- t[39548] = 5
      "0000101" when "01001101001111101", -- t[39549] = 5
      "0000101" when "01001101001111110", -- t[39550] = 5
      "0000101" when "01001101001111111", -- t[39551] = 5
      "0000101" when "01001101010000000", -- t[39552] = 5
      "0000101" when "01001101010000001", -- t[39553] = 5
      "0000101" when "01001101010000010", -- t[39554] = 5
      "0000101" when "01001101010000011", -- t[39555] = 5
      "0000101" when "01001101010000100", -- t[39556] = 5
      "0000101" when "01001101010000101", -- t[39557] = 5
      "0000101" when "01001101010000110", -- t[39558] = 5
      "0000101" when "01001101010000111", -- t[39559] = 5
      "0000101" when "01001101010001000", -- t[39560] = 5
      "0000101" when "01001101010001001", -- t[39561] = 5
      "0000101" when "01001101010001010", -- t[39562] = 5
      "0000101" when "01001101010001011", -- t[39563] = 5
      "0000101" when "01001101010001100", -- t[39564] = 5
      "0000101" when "01001101010001101", -- t[39565] = 5
      "0000101" when "01001101010001110", -- t[39566] = 5
      "0000101" when "01001101010001111", -- t[39567] = 5
      "0000101" when "01001101010010000", -- t[39568] = 5
      "0000101" when "01001101010010001", -- t[39569] = 5
      "0000101" when "01001101010010010", -- t[39570] = 5
      "0000101" when "01001101010010011", -- t[39571] = 5
      "0000101" when "01001101010010100", -- t[39572] = 5
      "0000101" when "01001101010010101", -- t[39573] = 5
      "0000101" when "01001101010010110", -- t[39574] = 5
      "0000101" when "01001101010010111", -- t[39575] = 5
      "0000101" when "01001101010011000", -- t[39576] = 5
      "0000101" when "01001101010011001", -- t[39577] = 5
      "0000101" when "01001101010011010", -- t[39578] = 5
      "0000101" when "01001101010011011", -- t[39579] = 5
      "0000101" when "01001101010011100", -- t[39580] = 5
      "0000101" when "01001101010011101", -- t[39581] = 5
      "0000101" when "01001101010011110", -- t[39582] = 5
      "0000101" when "01001101010011111", -- t[39583] = 5
      "0000101" when "01001101010100000", -- t[39584] = 5
      "0000101" when "01001101010100001", -- t[39585] = 5
      "0000101" when "01001101010100010", -- t[39586] = 5
      "0000101" when "01001101010100011", -- t[39587] = 5
      "0000101" when "01001101010100100", -- t[39588] = 5
      "0000101" when "01001101010100101", -- t[39589] = 5
      "0000101" when "01001101010100110", -- t[39590] = 5
      "0000101" when "01001101010100111", -- t[39591] = 5
      "0000101" when "01001101010101000", -- t[39592] = 5
      "0000101" when "01001101010101001", -- t[39593] = 5
      "0000101" when "01001101010101010", -- t[39594] = 5
      "0000101" when "01001101010101011", -- t[39595] = 5
      "0000101" when "01001101010101100", -- t[39596] = 5
      "0000101" when "01001101010101101", -- t[39597] = 5
      "0000101" when "01001101010101110", -- t[39598] = 5
      "0000101" when "01001101010101111", -- t[39599] = 5
      "0000101" when "01001101010110000", -- t[39600] = 5
      "0000101" when "01001101010110001", -- t[39601] = 5
      "0000101" when "01001101010110010", -- t[39602] = 5
      "0000101" when "01001101010110011", -- t[39603] = 5
      "0000101" when "01001101010110100", -- t[39604] = 5
      "0000101" when "01001101010110101", -- t[39605] = 5
      "0000101" when "01001101010110110", -- t[39606] = 5
      "0000101" when "01001101010110111", -- t[39607] = 5
      "0000101" when "01001101010111000", -- t[39608] = 5
      "0000101" when "01001101010111001", -- t[39609] = 5
      "0000101" when "01001101010111010", -- t[39610] = 5
      "0000101" when "01001101010111011", -- t[39611] = 5
      "0000101" when "01001101010111100", -- t[39612] = 5
      "0000101" when "01001101010111101", -- t[39613] = 5
      "0000101" when "01001101010111110", -- t[39614] = 5
      "0000101" when "01001101010111111", -- t[39615] = 5
      "0000101" when "01001101011000000", -- t[39616] = 5
      "0000101" when "01001101011000001", -- t[39617] = 5
      "0000101" when "01001101011000010", -- t[39618] = 5
      "0000101" when "01001101011000011", -- t[39619] = 5
      "0000101" when "01001101011000100", -- t[39620] = 5
      "0000101" when "01001101011000101", -- t[39621] = 5
      "0000101" when "01001101011000110", -- t[39622] = 5
      "0000101" when "01001101011000111", -- t[39623] = 5
      "0000101" when "01001101011001000", -- t[39624] = 5
      "0000101" when "01001101011001001", -- t[39625] = 5
      "0000101" when "01001101011001010", -- t[39626] = 5
      "0000101" when "01001101011001011", -- t[39627] = 5
      "0000101" when "01001101011001100", -- t[39628] = 5
      "0000101" when "01001101011001101", -- t[39629] = 5
      "0000101" when "01001101011001110", -- t[39630] = 5
      "0000101" when "01001101011001111", -- t[39631] = 5
      "0000101" when "01001101011010000", -- t[39632] = 5
      "0000101" when "01001101011010001", -- t[39633] = 5
      "0000101" when "01001101011010010", -- t[39634] = 5
      "0000101" when "01001101011010011", -- t[39635] = 5
      "0000101" when "01001101011010100", -- t[39636] = 5
      "0000101" when "01001101011010101", -- t[39637] = 5
      "0000101" when "01001101011010110", -- t[39638] = 5
      "0000101" when "01001101011010111", -- t[39639] = 5
      "0000101" when "01001101011011000", -- t[39640] = 5
      "0000101" when "01001101011011001", -- t[39641] = 5
      "0000101" when "01001101011011010", -- t[39642] = 5
      "0000101" when "01001101011011011", -- t[39643] = 5
      "0000101" when "01001101011011100", -- t[39644] = 5
      "0000101" when "01001101011011101", -- t[39645] = 5
      "0000101" when "01001101011011110", -- t[39646] = 5
      "0000101" when "01001101011011111", -- t[39647] = 5
      "0000101" when "01001101011100000", -- t[39648] = 5
      "0000101" when "01001101011100001", -- t[39649] = 5
      "0000101" when "01001101011100010", -- t[39650] = 5
      "0000101" when "01001101011100011", -- t[39651] = 5
      "0000101" when "01001101011100100", -- t[39652] = 5
      "0000101" when "01001101011100101", -- t[39653] = 5
      "0000101" when "01001101011100110", -- t[39654] = 5
      "0000101" when "01001101011100111", -- t[39655] = 5
      "0000101" when "01001101011101000", -- t[39656] = 5
      "0000101" when "01001101011101001", -- t[39657] = 5
      "0000101" when "01001101011101010", -- t[39658] = 5
      "0000101" when "01001101011101011", -- t[39659] = 5
      "0000101" when "01001101011101100", -- t[39660] = 5
      "0000101" when "01001101011101101", -- t[39661] = 5
      "0000101" when "01001101011101110", -- t[39662] = 5
      "0000101" when "01001101011101111", -- t[39663] = 5
      "0000101" when "01001101011110000", -- t[39664] = 5
      "0000101" when "01001101011110001", -- t[39665] = 5
      "0000101" when "01001101011110010", -- t[39666] = 5
      "0000101" when "01001101011110011", -- t[39667] = 5
      "0000101" when "01001101011110100", -- t[39668] = 5
      "0000101" when "01001101011110101", -- t[39669] = 5
      "0000101" when "01001101011110110", -- t[39670] = 5
      "0000101" when "01001101011110111", -- t[39671] = 5
      "0000101" when "01001101011111000", -- t[39672] = 5
      "0000101" when "01001101011111001", -- t[39673] = 5
      "0000101" when "01001101011111010", -- t[39674] = 5
      "0000101" when "01001101011111011", -- t[39675] = 5
      "0000101" when "01001101011111100", -- t[39676] = 5
      "0000101" when "01001101011111101", -- t[39677] = 5
      "0000101" when "01001101011111110", -- t[39678] = 5
      "0000101" when "01001101011111111", -- t[39679] = 5
      "0000101" when "01001101100000000", -- t[39680] = 5
      "0000101" when "01001101100000001", -- t[39681] = 5
      "0000101" when "01001101100000010", -- t[39682] = 5
      "0000101" when "01001101100000011", -- t[39683] = 5
      "0000101" when "01001101100000100", -- t[39684] = 5
      "0000101" when "01001101100000101", -- t[39685] = 5
      "0000101" when "01001101100000110", -- t[39686] = 5
      "0000101" when "01001101100000111", -- t[39687] = 5
      "0000101" when "01001101100001000", -- t[39688] = 5
      "0000101" when "01001101100001001", -- t[39689] = 5
      "0000101" when "01001101100001010", -- t[39690] = 5
      "0000101" when "01001101100001011", -- t[39691] = 5
      "0000101" when "01001101100001100", -- t[39692] = 5
      "0000101" when "01001101100001101", -- t[39693] = 5
      "0000101" when "01001101100001110", -- t[39694] = 5
      "0000101" when "01001101100001111", -- t[39695] = 5
      "0000101" when "01001101100010000", -- t[39696] = 5
      "0000101" when "01001101100010001", -- t[39697] = 5
      "0000101" when "01001101100010010", -- t[39698] = 5
      "0000101" when "01001101100010011", -- t[39699] = 5
      "0000101" when "01001101100010100", -- t[39700] = 5
      "0000101" when "01001101100010101", -- t[39701] = 5
      "0000101" when "01001101100010110", -- t[39702] = 5
      "0000101" when "01001101100010111", -- t[39703] = 5
      "0000101" when "01001101100011000", -- t[39704] = 5
      "0000101" when "01001101100011001", -- t[39705] = 5
      "0000101" when "01001101100011010", -- t[39706] = 5
      "0000101" when "01001101100011011", -- t[39707] = 5
      "0000101" when "01001101100011100", -- t[39708] = 5
      "0000101" when "01001101100011101", -- t[39709] = 5
      "0000101" when "01001101100011110", -- t[39710] = 5
      "0000101" when "01001101100011111", -- t[39711] = 5
      "0000101" when "01001101100100000", -- t[39712] = 5
      "0000101" when "01001101100100001", -- t[39713] = 5
      "0000101" when "01001101100100010", -- t[39714] = 5
      "0000101" when "01001101100100011", -- t[39715] = 5
      "0000101" when "01001101100100100", -- t[39716] = 5
      "0000101" when "01001101100100101", -- t[39717] = 5
      "0000101" when "01001101100100110", -- t[39718] = 5
      "0000101" when "01001101100100111", -- t[39719] = 5
      "0000101" when "01001101100101000", -- t[39720] = 5
      "0000101" when "01001101100101001", -- t[39721] = 5
      "0000101" when "01001101100101010", -- t[39722] = 5
      "0000101" when "01001101100101011", -- t[39723] = 5
      "0000101" when "01001101100101100", -- t[39724] = 5
      "0000101" when "01001101100101101", -- t[39725] = 5
      "0000101" when "01001101100101110", -- t[39726] = 5
      "0000101" when "01001101100101111", -- t[39727] = 5
      "0000101" when "01001101100110000", -- t[39728] = 5
      "0000101" when "01001101100110001", -- t[39729] = 5
      "0000101" when "01001101100110010", -- t[39730] = 5
      "0000101" when "01001101100110011", -- t[39731] = 5
      "0000101" when "01001101100110100", -- t[39732] = 5
      "0000101" when "01001101100110101", -- t[39733] = 5
      "0000101" when "01001101100110110", -- t[39734] = 5
      "0000101" when "01001101100110111", -- t[39735] = 5
      "0000101" when "01001101100111000", -- t[39736] = 5
      "0000101" when "01001101100111001", -- t[39737] = 5
      "0000101" when "01001101100111010", -- t[39738] = 5
      "0000101" when "01001101100111011", -- t[39739] = 5
      "0000101" when "01001101100111100", -- t[39740] = 5
      "0000101" when "01001101100111101", -- t[39741] = 5
      "0000101" when "01001101100111110", -- t[39742] = 5
      "0000101" when "01001101100111111", -- t[39743] = 5
      "0000101" when "01001101101000000", -- t[39744] = 5
      "0000101" when "01001101101000001", -- t[39745] = 5
      "0000101" when "01001101101000010", -- t[39746] = 5
      "0000101" when "01001101101000011", -- t[39747] = 5
      "0000101" when "01001101101000100", -- t[39748] = 5
      "0000101" when "01001101101000101", -- t[39749] = 5
      "0000101" when "01001101101000110", -- t[39750] = 5
      "0000101" when "01001101101000111", -- t[39751] = 5
      "0000101" when "01001101101001000", -- t[39752] = 5
      "0000101" when "01001101101001001", -- t[39753] = 5
      "0000101" when "01001101101001010", -- t[39754] = 5
      "0000101" when "01001101101001011", -- t[39755] = 5
      "0000101" when "01001101101001100", -- t[39756] = 5
      "0000101" when "01001101101001101", -- t[39757] = 5
      "0000101" when "01001101101001110", -- t[39758] = 5
      "0000101" when "01001101101001111", -- t[39759] = 5
      "0000101" when "01001101101010000", -- t[39760] = 5
      "0000101" when "01001101101010001", -- t[39761] = 5
      "0000101" when "01001101101010010", -- t[39762] = 5
      "0000101" when "01001101101010011", -- t[39763] = 5
      "0000101" when "01001101101010100", -- t[39764] = 5
      "0000101" when "01001101101010101", -- t[39765] = 5
      "0000101" when "01001101101010110", -- t[39766] = 5
      "0000101" when "01001101101010111", -- t[39767] = 5
      "0000101" when "01001101101011000", -- t[39768] = 5
      "0000101" when "01001101101011001", -- t[39769] = 5
      "0000101" when "01001101101011010", -- t[39770] = 5
      "0000101" when "01001101101011011", -- t[39771] = 5
      "0000101" when "01001101101011100", -- t[39772] = 5
      "0000101" when "01001101101011101", -- t[39773] = 5
      "0000101" when "01001101101011110", -- t[39774] = 5
      "0000101" when "01001101101011111", -- t[39775] = 5
      "0000101" when "01001101101100000", -- t[39776] = 5
      "0000101" when "01001101101100001", -- t[39777] = 5
      "0000101" when "01001101101100010", -- t[39778] = 5
      "0000101" when "01001101101100011", -- t[39779] = 5
      "0000101" when "01001101101100100", -- t[39780] = 5
      "0000101" when "01001101101100101", -- t[39781] = 5
      "0000101" when "01001101101100110", -- t[39782] = 5
      "0000101" when "01001101101100111", -- t[39783] = 5
      "0000101" when "01001101101101000", -- t[39784] = 5
      "0000101" when "01001101101101001", -- t[39785] = 5
      "0000101" when "01001101101101010", -- t[39786] = 5
      "0000101" when "01001101101101011", -- t[39787] = 5
      "0000101" when "01001101101101100", -- t[39788] = 5
      "0000101" when "01001101101101101", -- t[39789] = 5
      "0000101" when "01001101101101110", -- t[39790] = 5
      "0000101" when "01001101101101111", -- t[39791] = 5
      "0000101" when "01001101101110000", -- t[39792] = 5
      "0000101" when "01001101101110001", -- t[39793] = 5
      "0000101" when "01001101101110010", -- t[39794] = 5
      "0000101" when "01001101101110011", -- t[39795] = 5
      "0000101" when "01001101101110100", -- t[39796] = 5
      "0000101" when "01001101101110101", -- t[39797] = 5
      "0000101" when "01001101101110110", -- t[39798] = 5
      "0000101" when "01001101101110111", -- t[39799] = 5
      "0000101" when "01001101101111000", -- t[39800] = 5
      "0000101" when "01001101101111001", -- t[39801] = 5
      "0000101" when "01001101101111010", -- t[39802] = 5
      "0000101" when "01001101101111011", -- t[39803] = 5
      "0000101" when "01001101101111100", -- t[39804] = 5
      "0000101" when "01001101101111101", -- t[39805] = 5
      "0000101" when "01001101101111110", -- t[39806] = 5
      "0000101" when "01001101101111111", -- t[39807] = 5
      "0000101" when "01001101110000000", -- t[39808] = 5
      "0000101" when "01001101110000001", -- t[39809] = 5
      "0000101" when "01001101110000010", -- t[39810] = 5
      "0000101" when "01001101110000011", -- t[39811] = 5
      "0000101" when "01001101110000100", -- t[39812] = 5
      "0000101" when "01001101110000101", -- t[39813] = 5
      "0000101" when "01001101110000110", -- t[39814] = 5
      "0000101" when "01001101110000111", -- t[39815] = 5
      "0000101" when "01001101110001000", -- t[39816] = 5
      "0000101" when "01001101110001001", -- t[39817] = 5
      "0000101" when "01001101110001010", -- t[39818] = 5
      "0000101" when "01001101110001011", -- t[39819] = 5
      "0000101" when "01001101110001100", -- t[39820] = 5
      "0000101" when "01001101110001101", -- t[39821] = 5
      "0000101" when "01001101110001110", -- t[39822] = 5
      "0000101" when "01001101110001111", -- t[39823] = 5
      "0000101" when "01001101110010000", -- t[39824] = 5
      "0000101" when "01001101110010001", -- t[39825] = 5
      "0000101" when "01001101110010010", -- t[39826] = 5
      "0000101" when "01001101110010011", -- t[39827] = 5
      "0000101" when "01001101110010100", -- t[39828] = 5
      "0000101" when "01001101110010101", -- t[39829] = 5
      "0000101" when "01001101110010110", -- t[39830] = 5
      "0000101" when "01001101110010111", -- t[39831] = 5
      "0000101" when "01001101110011000", -- t[39832] = 5
      "0000101" when "01001101110011001", -- t[39833] = 5
      "0000101" when "01001101110011010", -- t[39834] = 5
      "0000101" when "01001101110011011", -- t[39835] = 5
      "0000101" when "01001101110011100", -- t[39836] = 5
      "0000101" when "01001101110011101", -- t[39837] = 5
      "0000101" when "01001101110011110", -- t[39838] = 5
      "0000101" when "01001101110011111", -- t[39839] = 5
      "0000101" when "01001101110100000", -- t[39840] = 5
      "0000101" when "01001101110100001", -- t[39841] = 5
      "0000101" when "01001101110100010", -- t[39842] = 5
      "0000101" when "01001101110100011", -- t[39843] = 5
      "0000101" when "01001101110100100", -- t[39844] = 5
      "0000101" when "01001101110100101", -- t[39845] = 5
      "0000101" when "01001101110100110", -- t[39846] = 5
      "0000101" when "01001101110100111", -- t[39847] = 5
      "0000101" when "01001101110101000", -- t[39848] = 5
      "0000101" when "01001101110101001", -- t[39849] = 5
      "0000101" when "01001101110101010", -- t[39850] = 5
      "0000101" when "01001101110101011", -- t[39851] = 5
      "0000101" when "01001101110101100", -- t[39852] = 5
      "0000101" when "01001101110101101", -- t[39853] = 5
      "0000101" when "01001101110101110", -- t[39854] = 5
      "0000101" when "01001101110101111", -- t[39855] = 5
      "0000101" when "01001101110110000", -- t[39856] = 5
      "0000101" when "01001101110110001", -- t[39857] = 5
      "0000101" when "01001101110110010", -- t[39858] = 5
      "0000101" when "01001101110110011", -- t[39859] = 5
      "0000101" when "01001101110110100", -- t[39860] = 5
      "0000101" when "01001101110110101", -- t[39861] = 5
      "0000101" when "01001101110110110", -- t[39862] = 5
      "0000101" when "01001101110110111", -- t[39863] = 5
      "0000101" when "01001101110111000", -- t[39864] = 5
      "0000101" when "01001101110111001", -- t[39865] = 5
      "0000101" when "01001101110111010", -- t[39866] = 5
      "0000101" when "01001101110111011", -- t[39867] = 5
      "0000101" when "01001101110111100", -- t[39868] = 5
      "0000101" when "01001101110111101", -- t[39869] = 5
      "0000101" when "01001101110111110", -- t[39870] = 5
      "0000101" when "01001101110111111", -- t[39871] = 5
      "0000101" when "01001101111000000", -- t[39872] = 5
      "0000101" when "01001101111000001", -- t[39873] = 5
      "0000101" when "01001101111000010", -- t[39874] = 5
      "0000101" when "01001101111000011", -- t[39875] = 5
      "0000101" when "01001101111000100", -- t[39876] = 5
      "0000101" when "01001101111000101", -- t[39877] = 5
      "0000101" when "01001101111000110", -- t[39878] = 5
      "0000101" when "01001101111000111", -- t[39879] = 5
      "0000101" when "01001101111001000", -- t[39880] = 5
      "0000101" when "01001101111001001", -- t[39881] = 5
      "0000101" when "01001101111001010", -- t[39882] = 5
      "0000101" when "01001101111001011", -- t[39883] = 5
      "0000101" when "01001101111001100", -- t[39884] = 5
      "0000101" when "01001101111001101", -- t[39885] = 5
      "0000101" when "01001101111001110", -- t[39886] = 5
      "0000101" when "01001101111001111", -- t[39887] = 5
      "0000101" when "01001101111010000", -- t[39888] = 5
      "0000101" when "01001101111010001", -- t[39889] = 5
      "0000101" when "01001101111010010", -- t[39890] = 5
      "0000101" when "01001101111010011", -- t[39891] = 5
      "0000101" when "01001101111010100", -- t[39892] = 5
      "0000101" when "01001101111010101", -- t[39893] = 5
      "0000101" when "01001101111010110", -- t[39894] = 5
      "0000101" when "01001101111010111", -- t[39895] = 5
      "0000101" when "01001101111011000", -- t[39896] = 5
      "0000101" when "01001101111011001", -- t[39897] = 5
      "0000101" when "01001101111011010", -- t[39898] = 5
      "0000101" when "01001101111011011", -- t[39899] = 5
      "0000101" when "01001101111011100", -- t[39900] = 5
      "0000101" when "01001101111011101", -- t[39901] = 5
      "0000101" when "01001101111011110", -- t[39902] = 5
      "0000101" when "01001101111011111", -- t[39903] = 5
      "0000101" when "01001101111100000", -- t[39904] = 5
      "0000101" when "01001101111100001", -- t[39905] = 5
      "0000101" when "01001101111100010", -- t[39906] = 5
      "0000101" when "01001101111100011", -- t[39907] = 5
      "0000101" when "01001101111100100", -- t[39908] = 5
      "0000101" when "01001101111100101", -- t[39909] = 5
      "0000101" when "01001101111100110", -- t[39910] = 5
      "0000101" when "01001101111100111", -- t[39911] = 5
      "0000101" when "01001101111101000", -- t[39912] = 5
      "0000101" when "01001101111101001", -- t[39913] = 5
      "0000101" when "01001101111101010", -- t[39914] = 5
      "0000101" when "01001101111101011", -- t[39915] = 5
      "0000101" when "01001101111101100", -- t[39916] = 5
      "0000101" when "01001101111101101", -- t[39917] = 5
      "0000101" when "01001101111101110", -- t[39918] = 5
      "0000101" when "01001101111101111", -- t[39919] = 5
      "0000101" when "01001101111110000", -- t[39920] = 5
      "0000101" when "01001101111110001", -- t[39921] = 5
      "0000101" when "01001101111110010", -- t[39922] = 5
      "0000101" when "01001101111110011", -- t[39923] = 5
      "0000101" when "01001101111110100", -- t[39924] = 5
      "0000101" when "01001101111110101", -- t[39925] = 5
      "0000101" when "01001101111110110", -- t[39926] = 5
      "0000101" when "01001101111110111", -- t[39927] = 5
      "0000101" when "01001101111111000", -- t[39928] = 5
      "0000101" when "01001101111111001", -- t[39929] = 5
      "0000101" when "01001101111111010", -- t[39930] = 5
      "0000101" when "01001101111111011", -- t[39931] = 5
      "0000101" when "01001101111111100", -- t[39932] = 5
      "0000101" when "01001101111111101", -- t[39933] = 5
      "0000101" when "01001101111111110", -- t[39934] = 5
      "0000101" when "01001101111111111", -- t[39935] = 5
      "0000101" when "01001110000000000", -- t[39936] = 5
      "0000101" when "01001110000000001", -- t[39937] = 5
      "0000101" when "01001110000000010", -- t[39938] = 5
      "0000101" when "01001110000000011", -- t[39939] = 5
      "0000101" when "01001110000000100", -- t[39940] = 5
      "0000101" when "01001110000000101", -- t[39941] = 5
      "0000101" when "01001110000000110", -- t[39942] = 5
      "0000101" when "01001110000000111", -- t[39943] = 5
      "0000101" when "01001110000001000", -- t[39944] = 5
      "0000101" when "01001110000001001", -- t[39945] = 5
      "0000101" when "01001110000001010", -- t[39946] = 5
      "0000101" when "01001110000001011", -- t[39947] = 5
      "0000101" when "01001110000001100", -- t[39948] = 5
      "0000101" when "01001110000001101", -- t[39949] = 5
      "0000101" when "01001110000001110", -- t[39950] = 5
      "0000101" when "01001110000001111", -- t[39951] = 5
      "0000101" when "01001110000010000", -- t[39952] = 5
      "0000101" when "01001110000010001", -- t[39953] = 5
      "0000101" when "01001110000010010", -- t[39954] = 5
      "0000101" when "01001110000010011", -- t[39955] = 5
      "0000101" when "01001110000010100", -- t[39956] = 5
      "0000101" when "01001110000010101", -- t[39957] = 5
      "0000101" when "01001110000010110", -- t[39958] = 5
      "0000101" when "01001110000010111", -- t[39959] = 5
      "0000101" when "01001110000011000", -- t[39960] = 5
      "0000101" when "01001110000011001", -- t[39961] = 5
      "0000101" when "01001110000011010", -- t[39962] = 5
      "0000101" when "01001110000011011", -- t[39963] = 5
      "0000101" when "01001110000011100", -- t[39964] = 5
      "0000101" when "01001110000011101", -- t[39965] = 5
      "0000101" when "01001110000011110", -- t[39966] = 5
      "0000101" when "01001110000011111", -- t[39967] = 5
      "0000101" when "01001110000100000", -- t[39968] = 5
      "0000101" when "01001110000100001", -- t[39969] = 5
      "0000101" when "01001110000100010", -- t[39970] = 5
      "0000101" when "01001110000100011", -- t[39971] = 5
      "0000101" when "01001110000100100", -- t[39972] = 5
      "0000101" when "01001110000100101", -- t[39973] = 5
      "0000101" when "01001110000100110", -- t[39974] = 5
      "0000101" when "01001110000100111", -- t[39975] = 5
      "0000101" when "01001110000101000", -- t[39976] = 5
      "0000101" when "01001110000101001", -- t[39977] = 5
      "0000101" when "01001110000101010", -- t[39978] = 5
      "0000101" when "01001110000101011", -- t[39979] = 5
      "0000101" when "01001110000101100", -- t[39980] = 5
      "0000101" when "01001110000101101", -- t[39981] = 5
      "0000101" when "01001110000101110", -- t[39982] = 5
      "0000101" when "01001110000101111", -- t[39983] = 5
      "0000101" when "01001110000110000", -- t[39984] = 5
      "0000101" when "01001110000110001", -- t[39985] = 5
      "0000101" when "01001110000110010", -- t[39986] = 5
      "0000101" when "01001110000110011", -- t[39987] = 5
      "0000101" when "01001110000110100", -- t[39988] = 5
      "0000101" when "01001110000110101", -- t[39989] = 5
      "0000101" when "01001110000110110", -- t[39990] = 5
      "0000101" when "01001110000110111", -- t[39991] = 5
      "0000101" when "01001110000111000", -- t[39992] = 5
      "0000101" when "01001110000111001", -- t[39993] = 5
      "0000101" when "01001110000111010", -- t[39994] = 5
      "0000101" when "01001110000111011", -- t[39995] = 5
      "0000101" when "01001110000111100", -- t[39996] = 5
      "0000101" when "01001110000111101", -- t[39997] = 5
      "0000101" when "01001110000111110", -- t[39998] = 5
      "0000101" when "01001110000111111", -- t[39999] = 5
      "0000101" when "01001110001000000", -- t[40000] = 5
      "0000101" when "01001110001000001", -- t[40001] = 5
      "0000101" when "01001110001000010", -- t[40002] = 5
      "0000101" when "01001110001000011", -- t[40003] = 5
      "0000101" when "01001110001000100", -- t[40004] = 5
      "0000101" when "01001110001000101", -- t[40005] = 5
      "0000101" when "01001110001000110", -- t[40006] = 5
      "0000101" when "01001110001000111", -- t[40007] = 5
      "0000101" when "01001110001001000", -- t[40008] = 5
      "0000101" when "01001110001001001", -- t[40009] = 5
      "0000101" when "01001110001001010", -- t[40010] = 5
      "0000101" when "01001110001001011", -- t[40011] = 5
      "0000101" when "01001110001001100", -- t[40012] = 5
      "0000101" when "01001110001001101", -- t[40013] = 5
      "0000101" when "01001110001001110", -- t[40014] = 5
      "0000101" when "01001110001001111", -- t[40015] = 5
      "0000101" when "01001110001010000", -- t[40016] = 5
      "0000101" when "01001110001010001", -- t[40017] = 5
      "0000101" when "01001110001010010", -- t[40018] = 5
      "0000101" when "01001110001010011", -- t[40019] = 5
      "0000101" when "01001110001010100", -- t[40020] = 5
      "0000101" when "01001110001010101", -- t[40021] = 5
      "0000101" when "01001110001010110", -- t[40022] = 5
      "0000101" when "01001110001010111", -- t[40023] = 5
      "0000101" when "01001110001011000", -- t[40024] = 5
      "0000101" when "01001110001011001", -- t[40025] = 5
      "0000101" when "01001110001011010", -- t[40026] = 5
      "0000101" when "01001110001011011", -- t[40027] = 5
      "0000101" when "01001110001011100", -- t[40028] = 5
      "0000101" when "01001110001011101", -- t[40029] = 5
      "0000101" when "01001110001011110", -- t[40030] = 5
      "0000101" when "01001110001011111", -- t[40031] = 5
      "0000101" when "01001110001100000", -- t[40032] = 5
      "0000101" when "01001110001100001", -- t[40033] = 5
      "0000101" when "01001110001100010", -- t[40034] = 5
      "0000101" when "01001110001100011", -- t[40035] = 5
      "0000101" when "01001110001100100", -- t[40036] = 5
      "0000101" when "01001110001100101", -- t[40037] = 5
      "0000101" when "01001110001100110", -- t[40038] = 5
      "0000101" when "01001110001100111", -- t[40039] = 5
      "0000101" when "01001110001101000", -- t[40040] = 5
      "0000101" when "01001110001101001", -- t[40041] = 5
      "0000101" when "01001110001101010", -- t[40042] = 5
      "0000101" when "01001110001101011", -- t[40043] = 5
      "0000101" when "01001110001101100", -- t[40044] = 5
      "0000101" when "01001110001101101", -- t[40045] = 5
      "0000101" when "01001110001101110", -- t[40046] = 5
      "0000101" when "01001110001101111", -- t[40047] = 5
      "0000101" when "01001110001110000", -- t[40048] = 5
      "0000101" when "01001110001110001", -- t[40049] = 5
      "0000101" when "01001110001110010", -- t[40050] = 5
      "0000101" when "01001110001110011", -- t[40051] = 5
      "0000101" when "01001110001110100", -- t[40052] = 5
      "0000101" when "01001110001110101", -- t[40053] = 5
      "0000101" when "01001110001110110", -- t[40054] = 5
      "0000101" when "01001110001110111", -- t[40055] = 5
      "0000101" when "01001110001111000", -- t[40056] = 5
      "0000101" when "01001110001111001", -- t[40057] = 5
      "0000101" when "01001110001111010", -- t[40058] = 5
      "0000101" when "01001110001111011", -- t[40059] = 5
      "0000101" when "01001110001111100", -- t[40060] = 5
      "0000101" when "01001110001111101", -- t[40061] = 5
      "0000101" when "01001110001111110", -- t[40062] = 5
      "0000101" when "01001110001111111", -- t[40063] = 5
      "0000101" when "01001110010000000", -- t[40064] = 5
      "0000101" when "01001110010000001", -- t[40065] = 5
      "0000101" when "01001110010000010", -- t[40066] = 5
      "0000101" when "01001110010000011", -- t[40067] = 5
      "0000101" when "01001110010000100", -- t[40068] = 5
      "0000101" when "01001110010000101", -- t[40069] = 5
      "0000101" when "01001110010000110", -- t[40070] = 5
      "0000101" when "01001110010000111", -- t[40071] = 5
      "0000101" when "01001110010001000", -- t[40072] = 5
      "0000101" when "01001110010001001", -- t[40073] = 5
      "0000101" when "01001110010001010", -- t[40074] = 5
      "0000101" when "01001110010001011", -- t[40075] = 5
      "0000101" when "01001110010001100", -- t[40076] = 5
      "0000101" when "01001110010001101", -- t[40077] = 5
      "0000101" when "01001110010001110", -- t[40078] = 5
      "0000101" when "01001110010001111", -- t[40079] = 5
      "0000101" when "01001110010010000", -- t[40080] = 5
      "0000101" when "01001110010010001", -- t[40081] = 5
      "0000101" when "01001110010010010", -- t[40082] = 5
      "0000101" when "01001110010010011", -- t[40083] = 5
      "0000101" when "01001110010010100", -- t[40084] = 5
      "0000101" when "01001110010010101", -- t[40085] = 5
      "0000101" when "01001110010010110", -- t[40086] = 5
      "0000101" when "01001110010010111", -- t[40087] = 5
      "0000101" when "01001110010011000", -- t[40088] = 5
      "0000101" when "01001110010011001", -- t[40089] = 5
      "0000101" when "01001110010011010", -- t[40090] = 5
      "0000101" when "01001110010011011", -- t[40091] = 5
      "0000101" when "01001110010011100", -- t[40092] = 5
      "0000101" when "01001110010011101", -- t[40093] = 5
      "0000101" when "01001110010011110", -- t[40094] = 5
      "0000101" when "01001110010011111", -- t[40095] = 5
      "0000101" when "01001110010100000", -- t[40096] = 5
      "0000101" when "01001110010100001", -- t[40097] = 5
      "0000101" when "01001110010100010", -- t[40098] = 5
      "0000101" when "01001110010100011", -- t[40099] = 5
      "0000101" when "01001110010100100", -- t[40100] = 5
      "0000101" when "01001110010100101", -- t[40101] = 5
      "0000101" when "01001110010100110", -- t[40102] = 5
      "0000101" when "01001110010100111", -- t[40103] = 5
      "0000101" when "01001110010101000", -- t[40104] = 5
      "0000101" when "01001110010101001", -- t[40105] = 5
      "0000101" when "01001110010101010", -- t[40106] = 5
      "0000101" when "01001110010101011", -- t[40107] = 5
      "0000101" when "01001110010101100", -- t[40108] = 5
      "0000101" when "01001110010101101", -- t[40109] = 5
      "0000101" when "01001110010101110", -- t[40110] = 5
      "0000101" when "01001110010101111", -- t[40111] = 5
      "0000101" when "01001110010110000", -- t[40112] = 5
      "0000101" when "01001110010110001", -- t[40113] = 5
      "0000101" when "01001110010110010", -- t[40114] = 5
      "0000101" when "01001110010110011", -- t[40115] = 5
      "0000101" when "01001110010110100", -- t[40116] = 5
      "0000101" when "01001110010110101", -- t[40117] = 5
      "0000101" when "01001110010110110", -- t[40118] = 5
      "0000101" when "01001110010110111", -- t[40119] = 5
      "0000101" when "01001110010111000", -- t[40120] = 5
      "0000101" when "01001110010111001", -- t[40121] = 5
      "0000101" when "01001110010111010", -- t[40122] = 5
      "0000101" when "01001110010111011", -- t[40123] = 5
      "0000101" when "01001110010111100", -- t[40124] = 5
      "0000101" when "01001110010111101", -- t[40125] = 5
      "0000101" when "01001110010111110", -- t[40126] = 5
      "0000101" when "01001110010111111", -- t[40127] = 5
      "0000101" when "01001110011000000", -- t[40128] = 5
      "0000101" when "01001110011000001", -- t[40129] = 5
      "0000101" when "01001110011000010", -- t[40130] = 5
      "0000101" when "01001110011000011", -- t[40131] = 5
      "0000101" when "01001110011000100", -- t[40132] = 5
      "0000101" when "01001110011000101", -- t[40133] = 5
      "0000101" when "01001110011000110", -- t[40134] = 5
      "0000101" when "01001110011000111", -- t[40135] = 5
      "0000101" when "01001110011001000", -- t[40136] = 5
      "0000101" when "01001110011001001", -- t[40137] = 5
      "0000101" when "01001110011001010", -- t[40138] = 5
      "0000101" when "01001110011001011", -- t[40139] = 5
      "0000101" when "01001110011001100", -- t[40140] = 5
      "0000101" when "01001110011001101", -- t[40141] = 5
      "0000101" when "01001110011001110", -- t[40142] = 5
      "0000101" when "01001110011001111", -- t[40143] = 5
      "0000101" when "01001110011010000", -- t[40144] = 5
      "0000101" when "01001110011010001", -- t[40145] = 5
      "0000101" when "01001110011010010", -- t[40146] = 5
      "0000101" when "01001110011010011", -- t[40147] = 5
      "0000101" when "01001110011010100", -- t[40148] = 5
      "0000101" when "01001110011010101", -- t[40149] = 5
      "0000101" when "01001110011010110", -- t[40150] = 5
      "0000101" when "01001110011010111", -- t[40151] = 5
      "0000101" when "01001110011011000", -- t[40152] = 5
      "0000101" when "01001110011011001", -- t[40153] = 5
      "0000101" when "01001110011011010", -- t[40154] = 5
      "0000101" when "01001110011011011", -- t[40155] = 5
      "0000101" when "01001110011011100", -- t[40156] = 5
      "0000101" when "01001110011011101", -- t[40157] = 5
      "0000101" when "01001110011011110", -- t[40158] = 5
      "0000101" when "01001110011011111", -- t[40159] = 5
      "0000101" when "01001110011100000", -- t[40160] = 5
      "0000101" when "01001110011100001", -- t[40161] = 5
      "0000101" when "01001110011100010", -- t[40162] = 5
      "0000101" when "01001110011100011", -- t[40163] = 5
      "0000101" when "01001110011100100", -- t[40164] = 5
      "0000101" when "01001110011100101", -- t[40165] = 5
      "0000101" when "01001110011100110", -- t[40166] = 5
      "0000101" when "01001110011100111", -- t[40167] = 5
      "0000101" when "01001110011101000", -- t[40168] = 5
      "0000101" when "01001110011101001", -- t[40169] = 5
      "0000101" when "01001110011101010", -- t[40170] = 5
      "0000101" when "01001110011101011", -- t[40171] = 5
      "0000101" when "01001110011101100", -- t[40172] = 5
      "0000101" when "01001110011101101", -- t[40173] = 5
      "0000101" when "01001110011101110", -- t[40174] = 5
      "0000101" when "01001110011101111", -- t[40175] = 5
      "0000101" when "01001110011110000", -- t[40176] = 5
      "0000101" when "01001110011110001", -- t[40177] = 5
      "0000101" when "01001110011110010", -- t[40178] = 5
      "0000101" when "01001110011110011", -- t[40179] = 5
      "0000101" when "01001110011110100", -- t[40180] = 5
      "0000101" when "01001110011110101", -- t[40181] = 5
      "0000101" when "01001110011110110", -- t[40182] = 5
      "0000101" when "01001110011110111", -- t[40183] = 5
      "0000101" when "01001110011111000", -- t[40184] = 5
      "0000101" when "01001110011111001", -- t[40185] = 5
      "0000101" when "01001110011111010", -- t[40186] = 5
      "0000101" when "01001110011111011", -- t[40187] = 5
      "0000101" when "01001110011111100", -- t[40188] = 5
      "0000101" when "01001110011111101", -- t[40189] = 5
      "0000101" when "01001110011111110", -- t[40190] = 5
      "0000101" when "01001110011111111", -- t[40191] = 5
      "0000101" when "01001110100000000", -- t[40192] = 5
      "0000101" when "01001110100000001", -- t[40193] = 5
      "0000101" when "01001110100000010", -- t[40194] = 5
      "0000101" when "01001110100000011", -- t[40195] = 5
      "0000101" when "01001110100000100", -- t[40196] = 5
      "0000101" when "01001110100000101", -- t[40197] = 5
      "0000101" when "01001110100000110", -- t[40198] = 5
      "0000101" when "01001110100000111", -- t[40199] = 5
      "0000101" when "01001110100001000", -- t[40200] = 5
      "0000101" when "01001110100001001", -- t[40201] = 5
      "0000101" when "01001110100001010", -- t[40202] = 5
      "0000101" when "01001110100001011", -- t[40203] = 5
      "0000101" when "01001110100001100", -- t[40204] = 5
      "0000101" when "01001110100001101", -- t[40205] = 5
      "0000101" when "01001110100001110", -- t[40206] = 5
      "0000101" when "01001110100001111", -- t[40207] = 5
      "0000101" when "01001110100010000", -- t[40208] = 5
      "0000101" when "01001110100010001", -- t[40209] = 5
      "0000101" when "01001110100010010", -- t[40210] = 5
      "0000101" when "01001110100010011", -- t[40211] = 5
      "0000101" when "01001110100010100", -- t[40212] = 5
      "0000101" when "01001110100010101", -- t[40213] = 5
      "0000101" when "01001110100010110", -- t[40214] = 5
      "0000101" when "01001110100010111", -- t[40215] = 5
      "0000101" when "01001110100011000", -- t[40216] = 5
      "0000101" when "01001110100011001", -- t[40217] = 5
      "0000101" when "01001110100011010", -- t[40218] = 5
      "0000101" when "01001110100011011", -- t[40219] = 5
      "0000101" when "01001110100011100", -- t[40220] = 5
      "0000101" when "01001110100011101", -- t[40221] = 5
      "0000101" when "01001110100011110", -- t[40222] = 5
      "0000101" when "01001110100011111", -- t[40223] = 5
      "0000101" when "01001110100100000", -- t[40224] = 5
      "0000101" when "01001110100100001", -- t[40225] = 5
      "0000101" when "01001110100100010", -- t[40226] = 5
      "0000101" when "01001110100100011", -- t[40227] = 5
      "0000101" when "01001110100100100", -- t[40228] = 5
      "0000101" when "01001110100100101", -- t[40229] = 5
      "0000101" when "01001110100100110", -- t[40230] = 5
      "0000101" when "01001110100100111", -- t[40231] = 5
      "0000101" when "01001110100101000", -- t[40232] = 5
      "0000101" when "01001110100101001", -- t[40233] = 5
      "0000101" when "01001110100101010", -- t[40234] = 5
      "0000101" when "01001110100101011", -- t[40235] = 5
      "0000101" when "01001110100101100", -- t[40236] = 5
      "0000101" when "01001110100101101", -- t[40237] = 5
      "0000101" when "01001110100101110", -- t[40238] = 5
      "0000101" when "01001110100101111", -- t[40239] = 5
      "0000101" when "01001110100110000", -- t[40240] = 5
      "0000101" when "01001110100110001", -- t[40241] = 5
      "0000101" when "01001110100110010", -- t[40242] = 5
      "0000101" when "01001110100110011", -- t[40243] = 5
      "0000101" when "01001110100110100", -- t[40244] = 5
      "0000101" when "01001110100110101", -- t[40245] = 5
      "0000101" when "01001110100110110", -- t[40246] = 5
      "0000101" when "01001110100110111", -- t[40247] = 5
      "0000101" when "01001110100111000", -- t[40248] = 5
      "0000101" when "01001110100111001", -- t[40249] = 5
      "0000101" when "01001110100111010", -- t[40250] = 5
      "0000101" when "01001110100111011", -- t[40251] = 5
      "0000101" when "01001110100111100", -- t[40252] = 5
      "0000101" when "01001110100111101", -- t[40253] = 5
      "0000101" when "01001110100111110", -- t[40254] = 5
      "0000101" when "01001110100111111", -- t[40255] = 5
      "0000101" when "01001110101000000", -- t[40256] = 5
      "0000101" when "01001110101000001", -- t[40257] = 5
      "0000101" when "01001110101000010", -- t[40258] = 5
      "0000101" when "01001110101000011", -- t[40259] = 5
      "0000101" when "01001110101000100", -- t[40260] = 5
      "0000101" when "01001110101000101", -- t[40261] = 5
      "0000101" when "01001110101000110", -- t[40262] = 5
      "0000101" when "01001110101000111", -- t[40263] = 5
      "0000101" when "01001110101001000", -- t[40264] = 5
      "0000101" when "01001110101001001", -- t[40265] = 5
      "0000101" when "01001110101001010", -- t[40266] = 5
      "0000101" when "01001110101001011", -- t[40267] = 5
      "0000101" when "01001110101001100", -- t[40268] = 5
      "0000101" when "01001110101001101", -- t[40269] = 5
      "0000101" when "01001110101001110", -- t[40270] = 5
      "0000101" when "01001110101001111", -- t[40271] = 5
      "0000101" when "01001110101010000", -- t[40272] = 5
      "0000101" when "01001110101010001", -- t[40273] = 5
      "0000101" when "01001110101010010", -- t[40274] = 5
      "0000101" when "01001110101010011", -- t[40275] = 5
      "0000101" when "01001110101010100", -- t[40276] = 5
      "0000101" when "01001110101010101", -- t[40277] = 5
      "0000101" when "01001110101010110", -- t[40278] = 5
      "0000101" when "01001110101010111", -- t[40279] = 5
      "0000101" when "01001110101011000", -- t[40280] = 5
      "0000101" when "01001110101011001", -- t[40281] = 5
      "0000101" when "01001110101011010", -- t[40282] = 5
      "0000101" when "01001110101011011", -- t[40283] = 5
      "0000101" when "01001110101011100", -- t[40284] = 5
      "0000101" when "01001110101011101", -- t[40285] = 5
      "0000101" when "01001110101011110", -- t[40286] = 5
      "0000101" when "01001110101011111", -- t[40287] = 5
      "0000101" when "01001110101100000", -- t[40288] = 5
      "0000101" when "01001110101100001", -- t[40289] = 5
      "0000101" when "01001110101100010", -- t[40290] = 5
      "0000101" when "01001110101100011", -- t[40291] = 5
      "0000101" when "01001110101100100", -- t[40292] = 5
      "0000101" when "01001110101100101", -- t[40293] = 5
      "0000101" when "01001110101100110", -- t[40294] = 5
      "0000101" when "01001110101100111", -- t[40295] = 5
      "0000101" when "01001110101101000", -- t[40296] = 5
      "0000101" when "01001110101101001", -- t[40297] = 5
      "0000101" when "01001110101101010", -- t[40298] = 5
      "0000101" when "01001110101101011", -- t[40299] = 5
      "0000101" when "01001110101101100", -- t[40300] = 5
      "0000101" when "01001110101101101", -- t[40301] = 5
      "0000101" when "01001110101101110", -- t[40302] = 5
      "0000101" when "01001110101101111", -- t[40303] = 5
      "0000101" when "01001110101110000", -- t[40304] = 5
      "0000101" when "01001110101110001", -- t[40305] = 5
      "0000101" when "01001110101110010", -- t[40306] = 5
      "0000101" when "01001110101110011", -- t[40307] = 5
      "0000101" when "01001110101110100", -- t[40308] = 5
      "0000101" when "01001110101110101", -- t[40309] = 5
      "0000101" when "01001110101110110", -- t[40310] = 5
      "0000101" when "01001110101110111", -- t[40311] = 5
      "0000101" when "01001110101111000", -- t[40312] = 5
      "0000101" when "01001110101111001", -- t[40313] = 5
      "0000101" when "01001110101111010", -- t[40314] = 5
      "0000101" when "01001110101111011", -- t[40315] = 5
      "0000101" when "01001110101111100", -- t[40316] = 5
      "0000101" when "01001110101111101", -- t[40317] = 5
      "0000101" when "01001110101111110", -- t[40318] = 5
      "0000101" when "01001110101111111", -- t[40319] = 5
      "0000101" when "01001110110000000", -- t[40320] = 5
      "0000101" when "01001110110000001", -- t[40321] = 5
      "0000101" when "01001110110000010", -- t[40322] = 5
      "0000101" when "01001110110000011", -- t[40323] = 5
      "0000101" when "01001110110000100", -- t[40324] = 5
      "0000101" when "01001110110000101", -- t[40325] = 5
      "0000101" when "01001110110000110", -- t[40326] = 5
      "0000101" when "01001110110000111", -- t[40327] = 5
      "0000101" when "01001110110001000", -- t[40328] = 5
      "0000101" when "01001110110001001", -- t[40329] = 5
      "0000101" when "01001110110001010", -- t[40330] = 5
      "0000101" when "01001110110001011", -- t[40331] = 5
      "0000101" when "01001110110001100", -- t[40332] = 5
      "0000101" when "01001110110001101", -- t[40333] = 5
      "0000101" when "01001110110001110", -- t[40334] = 5
      "0000101" when "01001110110001111", -- t[40335] = 5
      "0000101" when "01001110110010000", -- t[40336] = 5
      "0000101" when "01001110110010001", -- t[40337] = 5
      "0000101" when "01001110110010010", -- t[40338] = 5
      "0000101" when "01001110110010011", -- t[40339] = 5
      "0000101" when "01001110110010100", -- t[40340] = 5
      "0000101" when "01001110110010101", -- t[40341] = 5
      "0000101" when "01001110110010110", -- t[40342] = 5
      "0000101" when "01001110110010111", -- t[40343] = 5
      "0000101" when "01001110110011000", -- t[40344] = 5
      "0000101" when "01001110110011001", -- t[40345] = 5
      "0000101" when "01001110110011010", -- t[40346] = 5
      "0000101" when "01001110110011011", -- t[40347] = 5
      "0000101" when "01001110110011100", -- t[40348] = 5
      "0000101" when "01001110110011101", -- t[40349] = 5
      "0000101" when "01001110110011110", -- t[40350] = 5
      "0000101" when "01001110110011111", -- t[40351] = 5
      "0000101" when "01001110110100000", -- t[40352] = 5
      "0000101" when "01001110110100001", -- t[40353] = 5
      "0000101" when "01001110110100010", -- t[40354] = 5
      "0000101" when "01001110110100011", -- t[40355] = 5
      "0000101" when "01001110110100100", -- t[40356] = 5
      "0000101" when "01001110110100101", -- t[40357] = 5
      "0000101" when "01001110110100110", -- t[40358] = 5
      "0000101" when "01001110110100111", -- t[40359] = 5
      "0000101" when "01001110110101000", -- t[40360] = 5
      "0000101" when "01001110110101001", -- t[40361] = 5
      "0000101" when "01001110110101010", -- t[40362] = 5
      "0000101" when "01001110110101011", -- t[40363] = 5
      "0000101" when "01001110110101100", -- t[40364] = 5
      "0000101" when "01001110110101101", -- t[40365] = 5
      "0000101" when "01001110110101110", -- t[40366] = 5
      "0000101" when "01001110110101111", -- t[40367] = 5
      "0000101" when "01001110110110000", -- t[40368] = 5
      "0000101" when "01001110110110001", -- t[40369] = 5
      "0000101" when "01001110110110010", -- t[40370] = 5
      "0000101" when "01001110110110011", -- t[40371] = 5
      "0000101" when "01001110110110100", -- t[40372] = 5
      "0000101" when "01001110110110101", -- t[40373] = 5
      "0000101" when "01001110110110110", -- t[40374] = 5
      "0000101" when "01001110110110111", -- t[40375] = 5
      "0000101" when "01001110110111000", -- t[40376] = 5
      "0000101" when "01001110110111001", -- t[40377] = 5
      "0000101" when "01001110110111010", -- t[40378] = 5
      "0000101" when "01001110110111011", -- t[40379] = 5
      "0000101" when "01001110110111100", -- t[40380] = 5
      "0000101" when "01001110110111101", -- t[40381] = 5
      "0000101" when "01001110110111110", -- t[40382] = 5
      "0000101" when "01001110110111111", -- t[40383] = 5
      "0000101" when "01001110111000000", -- t[40384] = 5
      "0000101" when "01001110111000001", -- t[40385] = 5
      "0000101" when "01001110111000010", -- t[40386] = 5
      "0000101" when "01001110111000011", -- t[40387] = 5
      "0000101" when "01001110111000100", -- t[40388] = 5
      "0000101" when "01001110111000101", -- t[40389] = 5
      "0000110" when "01001110111000110", -- t[40390] = 6
      "0000110" when "01001110111000111", -- t[40391] = 6
      "0000110" when "01001110111001000", -- t[40392] = 6
      "0000110" when "01001110111001001", -- t[40393] = 6
      "0000110" when "01001110111001010", -- t[40394] = 6
      "0000110" when "01001110111001011", -- t[40395] = 6
      "0000110" when "01001110111001100", -- t[40396] = 6
      "0000110" when "01001110111001101", -- t[40397] = 6
      "0000110" when "01001110111001110", -- t[40398] = 6
      "0000110" when "01001110111001111", -- t[40399] = 6
      "0000110" when "01001110111010000", -- t[40400] = 6
      "0000110" when "01001110111010001", -- t[40401] = 6
      "0000110" when "01001110111010010", -- t[40402] = 6
      "0000110" when "01001110111010011", -- t[40403] = 6
      "0000110" when "01001110111010100", -- t[40404] = 6
      "0000110" when "01001110111010101", -- t[40405] = 6
      "0000110" when "01001110111010110", -- t[40406] = 6
      "0000110" when "01001110111010111", -- t[40407] = 6
      "0000110" when "01001110111011000", -- t[40408] = 6
      "0000110" when "01001110111011001", -- t[40409] = 6
      "0000110" when "01001110111011010", -- t[40410] = 6
      "0000110" when "01001110111011011", -- t[40411] = 6
      "0000110" when "01001110111011100", -- t[40412] = 6
      "0000110" when "01001110111011101", -- t[40413] = 6
      "0000110" when "01001110111011110", -- t[40414] = 6
      "0000110" when "01001110111011111", -- t[40415] = 6
      "0000110" when "01001110111100000", -- t[40416] = 6
      "0000110" when "01001110111100001", -- t[40417] = 6
      "0000110" when "01001110111100010", -- t[40418] = 6
      "0000110" when "01001110111100011", -- t[40419] = 6
      "0000110" when "01001110111100100", -- t[40420] = 6
      "0000110" when "01001110111100101", -- t[40421] = 6
      "0000110" when "01001110111100110", -- t[40422] = 6
      "0000110" when "01001110111100111", -- t[40423] = 6
      "0000110" when "01001110111101000", -- t[40424] = 6
      "0000110" when "01001110111101001", -- t[40425] = 6
      "0000110" when "01001110111101010", -- t[40426] = 6
      "0000110" when "01001110111101011", -- t[40427] = 6
      "0000110" when "01001110111101100", -- t[40428] = 6
      "0000110" when "01001110111101101", -- t[40429] = 6
      "0000110" when "01001110111101110", -- t[40430] = 6
      "0000110" when "01001110111101111", -- t[40431] = 6
      "0000110" when "01001110111110000", -- t[40432] = 6
      "0000110" when "01001110111110001", -- t[40433] = 6
      "0000110" when "01001110111110010", -- t[40434] = 6
      "0000110" when "01001110111110011", -- t[40435] = 6
      "0000110" when "01001110111110100", -- t[40436] = 6
      "0000110" when "01001110111110101", -- t[40437] = 6
      "0000110" when "01001110111110110", -- t[40438] = 6
      "0000110" when "01001110111110111", -- t[40439] = 6
      "0000110" when "01001110111111000", -- t[40440] = 6
      "0000110" when "01001110111111001", -- t[40441] = 6
      "0000110" when "01001110111111010", -- t[40442] = 6
      "0000110" when "01001110111111011", -- t[40443] = 6
      "0000110" when "01001110111111100", -- t[40444] = 6
      "0000110" when "01001110111111101", -- t[40445] = 6
      "0000110" when "01001110111111110", -- t[40446] = 6
      "0000110" when "01001110111111111", -- t[40447] = 6
      "0000110" when "01001111000000000", -- t[40448] = 6
      "0000110" when "01001111000000001", -- t[40449] = 6
      "0000110" when "01001111000000010", -- t[40450] = 6
      "0000110" when "01001111000000011", -- t[40451] = 6
      "0000110" when "01001111000000100", -- t[40452] = 6
      "0000110" when "01001111000000101", -- t[40453] = 6
      "0000110" when "01001111000000110", -- t[40454] = 6
      "0000110" when "01001111000000111", -- t[40455] = 6
      "0000110" when "01001111000001000", -- t[40456] = 6
      "0000110" when "01001111000001001", -- t[40457] = 6
      "0000110" when "01001111000001010", -- t[40458] = 6
      "0000110" when "01001111000001011", -- t[40459] = 6
      "0000110" when "01001111000001100", -- t[40460] = 6
      "0000110" when "01001111000001101", -- t[40461] = 6
      "0000110" when "01001111000001110", -- t[40462] = 6
      "0000110" when "01001111000001111", -- t[40463] = 6
      "0000110" when "01001111000010000", -- t[40464] = 6
      "0000110" when "01001111000010001", -- t[40465] = 6
      "0000110" when "01001111000010010", -- t[40466] = 6
      "0000110" when "01001111000010011", -- t[40467] = 6
      "0000110" when "01001111000010100", -- t[40468] = 6
      "0000110" when "01001111000010101", -- t[40469] = 6
      "0000110" when "01001111000010110", -- t[40470] = 6
      "0000110" when "01001111000010111", -- t[40471] = 6
      "0000110" when "01001111000011000", -- t[40472] = 6
      "0000110" when "01001111000011001", -- t[40473] = 6
      "0000110" when "01001111000011010", -- t[40474] = 6
      "0000110" when "01001111000011011", -- t[40475] = 6
      "0000110" when "01001111000011100", -- t[40476] = 6
      "0000110" when "01001111000011101", -- t[40477] = 6
      "0000110" when "01001111000011110", -- t[40478] = 6
      "0000110" when "01001111000011111", -- t[40479] = 6
      "0000110" when "01001111000100000", -- t[40480] = 6
      "0000110" when "01001111000100001", -- t[40481] = 6
      "0000110" when "01001111000100010", -- t[40482] = 6
      "0000110" when "01001111000100011", -- t[40483] = 6
      "0000110" when "01001111000100100", -- t[40484] = 6
      "0000110" when "01001111000100101", -- t[40485] = 6
      "0000110" when "01001111000100110", -- t[40486] = 6
      "0000110" when "01001111000100111", -- t[40487] = 6
      "0000110" when "01001111000101000", -- t[40488] = 6
      "0000110" when "01001111000101001", -- t[40489] = 6
      "0000110" when "01001111000101010", -- t[40490] = 6
      "0000110" when "01001111000101011", -- t[40491] = 6
      "0000110" when "01001111000101100", -- t[40492] = 6
      "0000110" when "01001111000101101", -- t[40493] = 6
      "0000110" when "01001111000101110", -- t[40494] = 6
      "0000110" when "01001111000101111", -- t[40495] = 6
      "0000110" when "01001111000110000", -- t[40496] = 6
      "0000110" when "01001111000110001", -- t[40497] = 6
      "0000110" when "01001111000110010", -- t[40498] = 6
      "0000110" when "01001111000110011", -- t[40499] = 6
      "0000110" when "01001111000110100", -- t[40500] = 6
      "0000110" when "01001111000110101", -- t[40501] = 6
      "0000110" when "01001111000110110", -- t[40502] = 6
      "0000110" when "01001111000110111", -- t[40503] = 6
      "0000110" when "01001111000111000", -- t[40504] = 6
      "0000110" when "01001111000111001", -- t[40505] = 6
      "0000110" when "01001111000111010", -- t[40506] = 6
      "0000110" when "01001111000111011", -- t[40507] = 6
      "0000110" when "01001111000111100", -- t[40508] = 6
      "0000110" when "01001111000111101", -- t[40509] = 6
      "0000110" when "01001111000111110", -- t[40510] = 6
      "0000110" when "01001111000111111", -- t[40511] = 6
      "0000110" when "01001111001000000", -- t[40512] = 6
      "0000110" when "01001111001000001", -- t[40513] = 6
      "0000110" when "01001111001000010", -- t[40514] = 6
      "0000110" when "01001111001000011", -- t[40515] = 6
      "0000110" when "01001111001000100", -- t[40516] = 6
      "0000110" when "01001111001000101", -- t[40517] = 6
      "0000110" when "01001111001000110", -- t[40518] = 6
      "0000110" when "01001111001000111", -- t[40519] = 6
      "0000110" when "01001111001001000", -- t[40520] = 6
      "0000110" when "01001111001001001", -- t[40521] = 6
      "0000110" when "01001111001001010", -- t[40522] = 6
      "0000110" when "01001111001001011", -- t[40523] = 6
      "0000110" when "01001111001001100", -- t[40524] = 6
      "0000110" when "01001111001001101", -- t[40525] = 6
      "0000110" when "01001111001001110", -- t[40526] = 6
      "0000110" when "01001111001001111", -- t[40527] = 6
      "0000110" when "01001111001010000", -- t[40528] = 6
      "0000110" when "01001111001010001", -- t[40529] = 6
      "0000110" when "01001111001010010", -- t[40530] = 6
      "0000110" when "01001111001010011", -- t[40531] = 6
      "0000110" when "01001111001010100", -- t[40532] = 6
      "0000110" when "01001111001010101", -- t[40533] = 6
      "0000110" when "01001111001010110", -- t[40534] = 6
      "0000110" when "01001111001010111", -- t[40535] = 6
      "0000110" when "01001111001011000", -- t[40536] = 6
      "0000110" when "01001111001011001", -- t[40537] = 6
      "0000110" when "01001111001011010", -- t[40538] = 6
      "0000110" when "01001111001011011", -- t[40539] = 6
      "0000110" when "01001111001011100", -- t[40540] = 6
      "0000110" when "01001111001011101", -- t[40541] = 6
      "0000110" when "01001111001011110", -- t[40542] = 6
      "0000110" when "01001111001011111", -- t[40543] = 6
      "0000110" when "01001111001100000", -- t[40544] = 6
      "0000110" when "01001111001100001", -- t[40545] = 6
      "0000110" when "01001111001100010", -- t[40546] = 6
      "0000110" when "01001111001100011", -- t[40547] = 6
      "0000110" when "01001111001100100", -- t[40548] = 6
      "0000110" when "01001111001100101", -- t[40549] = 6
      "0000110" when "01001111001100110", -- t[40550] = 6
      "0000110" when "01001111001100111", -- t[40551] = 6
      "0000110" when "01001111001101000", -- t[40552] = 6
      "0000110" when "01001111001101001", -- t[40553] = 6
      "0000110" when "01001111001101010", -- t[40554] = 6
      "0000110" when "01001111001101011", -- t[40555] = 6
      "0000110" when "01001111001101100", -- t[40556] = 6
      "0000110" when "01001111001101101", -- t[40557] = 6
      "0000110" when "01001111001101110", -- t[40558] = 6
      "0000110" when "01001111001101111", -- t[40559] = 6
      "0000110" when "01001111001110000", -- t[40560] = 6
      "0000110" when "01001111001110001", -- t[40561] = 6
      "0000110" when "01001111001110010", -- t[40562] = 6
      "0000110" when "01001111001110011", -- t[40563] = 6
      "0000110" when "01001111001110100", -- t[40564] = 6
      "0000110" when "01001111001110101", -- t[40565] = 6
      "0000110" when "01001111001110110", -- t[40566] = 6
      "0000110" when "01001111001110111", -- t[40567] = 6
      "0000110" when "01001111001111000", -- t[40568] = 6
      "0000110" when "01001111001111001", -- t[40569] = 6
      "0000110" when "01001111001111010", -- t[40570] = 6
      "0000110" when "01001111001111011", -- t[40571] = 6
      "0000110" when "01001111001111100", -- t[40572] = 6
      "0000110" when "01001111001111101", -- t[40573] = 6
      "0000110" when "01001111001111110", -- t[40574] = 6
      "0000110" when "01001111001111111", -- t[40575] = 6
      "0000110" when "01001111010000000", -- t[40576] = 6
      "0000110" when "01001111010000001", -- t[40577] = 6
      "0000110" when "01001111010000010", -- t[40578] = 6
      "0000110" when "01001111010000011", -- t[40579] = 6
      "0000110" when "01001111010000100", -- t[40580] = 6
      "0000110" when "01001111010000101", -- t[40581] = 6
      "0000110" when "01001111010000110", -- t[40582] = 6
      "0000110" when "01001111010000111", -- t[40583] = 6
      "0000110" when "01001111010001000", -- t[40584] = 6
      "0000110" when "01001111010001001", -- t[40585] = 6
      "0000110" when "01001111010001010", -- t[40586] = 6
      "0000110" when "01001111010001011", -- t[40587] = 6
      "0000110" when "01001111010001100", -- t[40588] = 6
      "0000110" when "01001111010001101", -- t[40589] = 6
      "0000110" when "01001111010001110", -- t[40590] = 6
      "0000110" when "01001111010001111", -- t[40591] = 6
      "0000110" when "01001111010010000", -- t[40592] = 6
      "0000110" when "01001111010010001", -- t[40593] = 6
      "0000110" when "01001111010010010", -- t[40594] = 6
      "0000110" when "01001111010010011", -- t[40595] = 6
      "0000110" when "01001111010010100", -- t[40596] = 6
      "0000110" when "01001111010010101", -- t[40597] = 6
      "0000110" when "01001111010010110", -- t[40598] = 6
      "0000110" when "01001111010010111", -- t[40599] = 6
      "0000110" when "01001111010011000", -- t[40600] = 6
      "0000110" when "01001111010011001", -- t[40601] = 6
      "0000110" when "01001111010011010", -- t[40602] = 6
      "0000110" when "01001111010011011", -- t[40603] = 6
      "0000110" when "01001111010011100", -- t[40604] = 6
      "0000110" when "01001111010011101", -- t[40605] = 6
      "0000110" when "01001111010011110", -- t[40606] = 6
      "0000110" when "01001111010011111", -- t[40607] = 6
      "0000110" when "01001111010100000", -- t[40608] = 6
      "0000110" when "01001111010100001", -- t[40609] = 6
      "0000110" when "01001111010100010", -- t[40610] = 6
      "0000110" when "01001111010100011", -- t[40611] = 6
      "0000110" when "01001111010100100", -- t[40612] = 6
      "0000110" when "01001111010100101", -- t[40613] = 6
      "0000110" when "01001111010100110", -- t[40614] = 6
      "0000110" when "01001111010100111", -- t[40615] = 6
      "0000110" when "01001111010101000", -- t[40616] = 6
      "0000110" when "01001111010101001", -- t[40617] = 6
      "0000110" when "01001111010101010", -- t[40618] = 6
      "0000110" when "01001111010101011", -- t[40619] = 6
      "0000110" when "01001111010101100", -- t[40620] = 6
      "0000110" when "01001111010101101", -- t[40621] = 6
      "0000110" when "01001111010101110", -- t[40622] = 6
      "0000110" when "01001111010101111", -- t[40623] = 6
      "0000110" when "01001111010110000", -- t[40624] = 6
      "0000110" when "01001111010110001", -- t[40625] = 6
      "0000110" when "01001111010110010", -- t[40626] = 6
      "0000110" when "01001111010110011", -- t[40627] = 6
      "0000110" when "01001111010110100", -- t[40628] = 6
      "0000110" when "01001111010110101", -- t[40629] = 6
      "0000110" when "01001111010110110", -- t[40630] = 6
      "0000110" when "01001111010110111", -- t[40631] = 6
      "0000110" when "01001111010111000", -- t[40632] = 6
      "0000110" when "01001111010111001", -- t[40633] = 6
      "0000110" when "01001111010111010", -- t[40634] = 6
      "0000110" when "01001111010111011", -- t[40635] = 6
      "0000110" when "01001111010111100", -- t[40636] = 6
      "0000110" when "01001111010111101", -- t[40637] = 6
      "0000110" when "01001111010111110", -- t[40638] = 6
      "0000110" when "01001111010111111", -- t[40639] = 6
      "0000110" when "01001111011000000", -- t[40640] = 6
      "0000110" when "01001111011000001", -- t[40641] = 6
      "0000110" when "01001111011000010", -- t[40642] = 6
      "0000110" when "01001111011000011", -- t[40643] = 6
      "0000110" when "01001111011000100", -- t[40644] = 6
      "0000110" when "01001111011000101", -- t[40645] = 6
      "0000110" when "01001111011000110", -- t[40646] = 6
      "0000110" when "01001111011000111", -- t[40647] = 6
      "0000110" when "01001111011001000", -- t[40648] = 6
      "0000110" when "01001111011001001", -- t[40649] = 6
      "0000110" when "01001111011001010", -- t[40650] = 6
      "0000110" when "01001111011001011", -- t[40651] = 6
      "0000110" when "01001111011001100", -- t[40652] = 6
      "0000110" when "01001111011001101", -- t[40653] = 6
      "0000110" when "01001111011001110", -- t[40654] = 6
      "0000110" when "01001111011001111", -- t[40655] = 6
      "0000110" when "01001111011010000", -- t[40656] = 6
      "0000110" when "01001111011010001", -- t[40657] = 6
      "0000110" when "01001111011010010", -- t[40658] = 6
      "0000110" when "01001111011010011", -- t[40659] = 6
      "0000110" when "01001111011010100", -- t[40660] = 6
      "0000110" when "01001111011010101", -- t[40661] = 6
      "0000110" when "01001111011010110", -- t[40662] = 6
      "0000110" when "01001111011010111", -- t[40663] = 6
      "0000110" when "01001111011011000", -- t[40664] = 6
      "0000110" when "01001111011011001", -- t[40665] = 6
      "0000110" when "01001111011011010", -- t[40666] = 6
      "0000110" when "01001111011011011", -- t[40667] = 6
      "0000110" when "01001111011011100", -- t[40668] = 6
      "0000110" when "01001111011011101", -- t[40669] = 6
      "0000110" when "01001111011011110", -- t[40670] = 6
      "0000110" when "01001111011011111", -- t[40671] = 6
      "0000110" when "01001111011100000", -- t[40672] = 6
      "0000110" when "01001111011100001", -- t[40673] = 6
      "0000110" when "01001111011100010", -- t[40674] = 6
      "0000110" when "01001111011100011", -- t[40675] = 6
      "0000110" when "01001111011100100", -- t[40676] = 6
      "0000110" when "01001111011100101", -- t[40677] = 6
      "0000110" when "01001111011100110", -- t[40678] = 6
      "0000110" when "01001111011100111", -- t[40679] = 6
      "0000110" when "01001111011101000", -- t[40680] = 6
      "0000110" when "01001111011101001", -- t[40681] = 6
      "0000110" when "01001111011101010", -- t[40682] = 6
      "0000110" when "01001111011101011", -- t[40683] = 6
      "0000110" when "01001111011101100", -- t[40684] = 6
      "0000110" when "01001111011101101", -- t[40685] = 6
      "0000110" when "01001111011101110", -- t[40686] = 6
      "0000110" when "01001111011101111", -- t[40687] = 6
      "0000110" when "01001111011110000", -- t[40688] = 6
      "0000110" when "01001111011110001", -- t[40689] = 6
      "0000110" when "01001111011110010", -- t[40690] = 6
      "0000110" when "01001111011110011", -- t[40691] = 6
      "0000110" when "01001111011110100", -- t[40692] = 6
      "0000110" when "01001111011110101", -- t[40693] = 6
      "0000110" when "01001111011110110", -- t[40694] = 6
      "0000110" when "01001111011110111", -- t[40695] = 6
      "0000110" when "01001111011111000", -- t[40696] = 6
      "0000110" when "01001111011111001", -- t[40697] = 6
      "0000110" when "01001111011111010", -- t[40698] = 6
      "0000110" when "01001111011111011", -- t[40699] = 6
      "0000110" when "01001111011111100", -- t[40700] = 6
      "0000110" when "01001111011111101", -- t[40701] = 6
      "0000110" when "01001111011111110", -- t[40702] = 6
      "0000110" when "01001111011111111", -- t[40703] = 6
      "0000110" when "01001111100000000", -- t[40704] = 6
      "0000110" when "01001111100000001", -- t[40705] = 6
      "0000110" when "01001111100000010", -- t[40706] = 6
      "0000110" when "01001111100000011", -- t[40707] = 6
      "0000110" when "01001111100000100", -- t[40708] = 6
      "0000110" when "01001111100000101", -- t[40709] = 6
      "0000110" when "01001111100000110", -- t[40710] = 6
      "0000110" when "01001111100000111", -- t[40711] = 6
      "0000110" when "01001111100001000", -- t[40712] = 6
      "0000110" when "01001111100001001", -- t[40713] = 6
      "0000110" when "01001111100001010", -- t[40714] = 6
      "0000110" when "01001111100001011", -- t[40715] = 6
      "0000110" when "01001111100001100", -- t[40716] = 6
      "0000110" when "01001111100001101", -- t[40717] = 6
      "0000110" when "01001111100001110", -- t[40718] = 6
      "0000110" when "01001111100001111", -- t[40719] = 6
      "0000110" when "01001111100010000", -- t[40720] = 6
      "0000110" when "01001111100010001", -- t[40721] = 6
      "0000110" when "01001111100010010", -- t[40722] = 6
      "0000110" when "01001111100010011", -- t[40723] = 6
      "0000110" when "01001111100010100", -- t[40724] = 6
      "0000110" when "01001111100010101", -- t[40725] = 6
      "0000110" when "01001111100010110", -- t[40726] = 6
      "0000110" when "01001111100010111", -- t[40727] = 6
      "0000110" when "01001111100011000", -- t[40728] = 6
      "0000110" when "01001111100011001", -- t[40729] = 6
      "0000110" when "01001111100011010", -- t[40730] = 6
      "0000110" when "01001111100011011", -- t[40731] = 6
      "0000110" when "01001111100011100", -- t[40732] = 6
      "0000110" when "01001111100011101", -- t[40733] = 6
      "0000110" when "01001111100011110", -- t[40734] = 6
      "0000110" when "01001111100011111", -- t[40735] = 6
      "0000110" when "01001111100100000", -- t[40736] = 6
      "0000110" when "01001111100100001", -- t[40737] = 6
      "0000110" when "01001111100100010", -- t[40738] = 6
      "0000110" when "01001111100100011", -- t[40739] = 6
      "0000110" when "01001111100100100", -- t[40740] = 6
      "0000110" when "01001111100100101", -- t[40741] = 6
      "0000110" when "01001111100100110", -- t[40742] = 6
      "0000110" when "01001111100100111", -- t[40743] = 6
      "0000110" when "01001111100101000", -- t[40744] = 6
      "0000110" when "01001111100101001", -- t[40745] = 6
      "0000110" when "01001111100101010", -- t[40746] = 6
      "0000110" when "01001111100101011", -- t[40747] = 6
      "0000110" when "01001111100101100", -- t[40748] = 6
      "0000110" when "01001111100101101", -- t[40749] = 6
      "0000110" when "01001111100101110", -- t[40750] = 6
      "0000110" when "01001111100101111", -- t[40751] = 6
      "0000110" when "01001111100110000", -- t[40752] = 6
      "0000110" when "01001111100110001", -- t[40753] = 6
      "0000110" when "01001111100110010", -- t[40754] = 6
      "0000110" when "01001111100110011", -- t[40755] = 6
      "0000110" when "01001111100110100", -- t[40756] = 6
      "0000110" when "01001111100110101", -- t[40757] = 6
      "0000110" when "01001111100110110", -- t[40758] = 6
      "0000110" when "01001111100110111", -- t[40759] = 6
      "0000110" when "01001111100111000", -- t[40760] = 6
      "0000110" when "01001111100111001", -- t[40761] = 6
      "0000110" when "01001111100111010", -- t[40762] = 6
      "0000110" when "01001111100111011", -- t[40763] = 6
      "0000110" when "01001111100111100", -- t[40764] = 6
      "0000110" when "01001111100111101", -- t[40765] = 6
      "0000110" when "01001111100111110", -- t[40766] = 6
      "0000110" when "01001111100111111", -- t[40767] = 6
      "0000110" when "01001111101000000", -- t[40768] = 6
      "0000110" when "01001111101000001", -- t[40769] = 6
      "0000110" when "01001111101000010", -- t[40770] = 6
      "0000110" when "01001111101000011", -- t[40771] = 6
      "0000110" when "01001111101000100", -- t[40772] = 6
      "0000110" when "01001111101000101", -- t[40773] = 6
      "0000110" when "01001111101000110", -- t[40774] = 6
      "0000110" when "01001111101000111", -- t[40775] = 6
      "0000110" when "01001111101001000", -- t[40776] = 6
      "0000110" when "01001111101001001", -- t[40777] = 6
      "0000110" when "01001111101001010", -- t[40778] = 6
      "0000110" when "01001111101001011", -- t[40779] = 6
      "0000110" when "01001111101001100", -- t[40780] = 6
      "0000110" when "01001111101001101", -- t[40781] = 6
      "0000110" when "01001111101001110", -- t[40782] = 6
      "0000110" when "01001111101001111", -- t[40783] = 6
      "0000110" when "01001111101010000", -- t[40784] = 6
      "0000110" when "01001111101010001", -- t[40785] = 6
      "0000110" when "01001111101010010", -- t[40786] = 6
      "0000110" when "01001111101010011", -- t[40787] = 6
      "0000110" when "01001111101010100", -- t[40788] = 6
      "0000110" when "01001111101010101", -- t[40789] = 6
      "0000110" when "01001111101010110", -- t[40790] = 6
      "0000110" when "01001111101010111", -- t[40791] = 6
      "0000110" when "01001111101011000", -- t[40792] = 6
      "0000110" when "01001111101011001", -- t[40793] = 6
      "0000110" when "01001111101011010", -- t[40794] = 6
      "0000110" when "01001111101011011", -- t[40795] = 6
      "0000110" when "01001111101011100", -- t[40796] = 6
      "0000110" when "01001111101011101", -- t[40797] = 6
      "0000110" when "01001111101011110", -- t[40798] = 6
      "0000110" when "01001111101011111", -- t[40799] = 6
      "0000110" when "01001111101100000", -- t[40800] = 6
      "0000110" when "01001111101100001", -- t[40801] = 6
      "0000110" when "01001111101100010", -- t[40802] = 6
      "0000110" when "01001111101100011", -- t[40803] = 6
      "0000110" when "01001111101100100", -- t[40804] = 6
      "0000110" when "01001111101100101", -- t[40805] = 6
      "0000110" when "01001111101100110", -- t[40806] = 6
      "0000110" when "01001111101100111", -- t[40807] = 6
      "0000110" when "01001111101101000", -- t[40808] = 6
      "0000110" when "01001111101101001", -- t[40809] = 6
      "0000110" when "01001111101101010", -- t[40810] = 6
      "0000110" when "01001111101101011", -- t[40811] = 6
      "0000110" when "01001111101101100", -- t[40812] = 6
      "0000110" when "01001111101101101", -- t[40813] = 6
      "0000110" when "01001111101101110", -- t[40814] = 6
      "0000110" when "01001111101101111", -- t[40815] = 6
      "0000110" when "01001111101110000", -- t[40816] = 6
      "0000110" when "01001111101110001", -- t[40817] = 6
      "0000110" when "01001111101110010", -- t[40818] = 6
      "0000110" when "01001111101110011", -- t[40819] = 6
      "0000110" when "01001111101110100", -- t[40820] = 6
      "0000110" when "01001111101110101", -- t[40821] = 6
      "0000110" when "01001111101110110", -- t[40822] = 6
      "0000110" when "01001111101110111", -- t[40823] = 6
      "0000110" when "01001111101111000", -- t[40824] = 6
      "0000110" when "01001111101111001", -- t[40825] = 6
      "0000110" when "01001111101111010", -- t[40826] = 6
      "0000110" when "01001111101111011", -- t[40827] = 6
      "0000110" when "01001111101111100", -- t[40828] = 6
      "0000110" when "01001111101111101", -- t[40829] = 6
      "0000110" when "01001111101111110", -- t[40830] = 6
      "0000110" when "01001111101111111", -- t[40831] = 6
      "0000110" when "01001111110000000", -- t[40832] = 6
      "0000110" when "01001111110000001", -- t[40833] = 6
      "0000110" when "01001111110000010", -- t[40834] = 6
      "0000110" when "01001111110000011", -- t[40835] = 6
      "0000110" when "01001111110000100", -- t[40836] = 6
      "0000110" when "01001111110000101", -- t[40837] = 6
      "0000110" when "01001111110000110", -- t[40838] = 6
      "0000110" when "01001111110000111", -- t[40839] = 6
      "0000110" when "01001111110001000", -- t[40840] = 6
      "0000110" when "01001111110001001", -- t[40841] = 6
      "0000110" when "01001111110001010", -- t[40842] = 6
      "0000110" when "01001111110001011", -- t[40843] = 6
      "0000110" when "01001111110001100", -- t[40844] = 6
      "0000110" when "01001111110001101", -- t[40845] = 6
      "0000110" when "01001111110001110", -- t[40846] = 6
      "0000110" when "01001111110001111", -- t[40847] = 6
      "0000110" when "01001111110010000", -- t[40848] = 6
      "0000110" when "01001111110010001", -- t[40849] = 6
      "0000110" when "01001111110010010", -- t[40850] = 6
      "0000110" when "01001111110010011", -- t[40851] = 6
      "0000110" when "01001111110010100", -- t[40852] = 6
      "0000110" when "01001111110010101", -- t[40853] = 6
      "0000110" when "01001111110010110", -- t[40854] = 6
      "0000110" when "01001111110010111", -- t[40855] = 6
      "0000110" when "01001111110011000", -- t[40856] = 6
      "0000110" when "01001111110011001", -- t[40857] = 6
      "0000110" when "01001111110011010", -- t[40858] = 6
      "0000110" when "01001111110011011", -- t[40859] = 6
      "0000110" when "01001111110011100", -- t[40860] = 6
      "0000110" when "01001111110011101", -- t[40861] = 6
      "0000110" when "01001111110011110", -- t[40862] = 6
      "0000110" when "01001111110011111", -- t[40863] = 6
      "0000110" when "01001111110100000", -- t[40864] = 6
      "0000110" when "01001111110100001", -- t[40865] = 6
      "0000110" when "01001111110100010", -- t[40866] = 6
      "0000110" when "01001111110100011", -- t[40867] = 6
      "0000110" when "01001111110100100", -- t[40868] = 6
      "0000110" when "01001111110100101", -- t[40869] = 6
      "0000110" when "01001111110100110", -- t[40870] = 6
      "0000110" when "01001111110100111", -- t[40871] = 6
      "0000110" when "01001111110101000", -- t[40872] = 6
      "0000110" when "01001111110101001", -- t[40873] = 6
      "0000110" when "01001111110101010", -- t[40874] = 6
      "0000110" when "01001111110101011", -- t[40875] = 6
      "0000110" when "01001111110101100", -- t[40876] = 6
      "0000110" when "01001111110101101", -- t[40877] = 6
      "0000110" when "01001111110101110", -- t[40878] = 6
      "0000110" when "01001111110101111", -- t[40879] = 6
      "0000110" when "01001111110110000", -- t[40880] = 6
      "0000110" when "01001111110110001", -- t[40881] = 6
      "0000110" when "01001111110110010", -- t[40882] = 6
      "0000110" when "01001111110110011", -- t[40883] = 6
      "0000110" when "01001111110110100", -- t[40884] = 6
      "0000110" when "01001111110110101", -- t[40885] = 6
      "0000110" when "01001111110110110", -- t[40886] = 6
      "0000110" when "01001111110110111", -- t[40887] = 6
      "0000110" when "01001111110111000", -- t[40888] = 6
      "0000110" when "01001111110111001", -- t[40889] = 6
      "0000110" when "01001111110111010", -- t[40890] = 6
      "0000110" when "01001111110111011", -- t[40891] = 6
      "0000110" when "01001111110111100", -- t[40892] = 6
      "0000110" when "01001111110111101", -- t[40893] = 6
      "0000110" when "01001111110111110", -- t[40894] = 6
      "0000110" when "01001111110111111", -- t[40895] = 6
      "0000110" when "01001111111000000", -- t[40896] = 6
      "0000110" when "01001111111000001", -- t[40897] = 6
      "0000110" when "01001111111000010", -- t[40898] = 6
      "0000110" when "01001111111000011", -- t[40899] = 6
      "0000110" when "01001111111000100", -- t[40900] = 6
      "0000110" when "01001111111000101", -- t[40901] = 6
      "0000110" when "01001111111000110", -- t[40902] = 6
      "0000110" when "01001111111000111", -- t[40903] = 6
      "0000110" when "01001111111001000", -- t[40904] = 6
      "0000110" when "01001111111001001", -- t[40905] = 6
      "0000110" when "01001111111001010", -- t[40906] = 6
      "0000110" when "01001111111001011", -- t[40907] = 6
      "0000110" when "01001111111001100", -- t[40908] = 6
      "0000110" when "01001111111001101", -- t[40909] = 6
      "0000110" when "01001111111001110", -- t[40910] = 6
      "0000110" when "01001111111001111", -- t[40911] = 6
      "0000110" when "01001111111010000", -- t[40912] = 6
      "0000110" when "01001111111010001", -- t[40913] = 6
      "0000110" when "01001111111010010", -- t[40914] = 6
      "0000110" when "01001111111010011", -- t[40915] = 6
      "0000110" when "01001111111010100", -- t[40916] = 6
      "0000110" when "01001111111010101", -- t[40917] = 6
      "0000110" when "01001111111010110", -- t[40918] = 6
      "0000110" when "01001111111010111", -- t[40919] = 6
      "0000110" when "01001111111011000", -- t[40920] = 6
      "0000110" when "01001111111011001", -- t[40921] = 6
      "0000110" when "01001111111011010", -- t[40922] = 6
      "0000110" when "01001111111011011", -- t[40923] = 6
      "0000110" when "01001111111011100", -- t[40924] = 6
      "0000110" when "01001111111011101", -- t[40925] = 6
      "0000110" when "01001111111011110", -- t[40926] = 6
      "0000110" when "01001111111011111", -- t[40927] = 6
      "0000110" when "01001111111100000", -- t[40928] = 6
      "0000110" when "01001111111100001", -- t[40929] = 6
      "0000110" when "01001111111100010", -- t[40930] = 6
      "0000110" when "01001111111100011", -- t[40931] = 6
      "0000110" when "01001111111100100", -- t[40932] = 6
      "0000110" when "01001111111100101", -- t[40933] = 6
      "0000110" when "01001111111100110", -- t[40934] = 6
      "0000110" when "01001111111100111", -- t[40935] = 6
      "0000110" when "01001111111101000", -- t[40936] = 6
      "0000110" when "01001111111101001", -- t[40937] = 6
      "0000110" when "01001111111101010", -- t[40938] = 6
      "0000110" when "01001111111101011", -- t[40939] = 6
      "0000110" when "01001111111101100", -- t[40940] = 6
      "0000110" when "01001111111101101", -- t[40941] = 6
      "0000110" when "01001111111101110", -- t[40942] = 6
      "0000110" when "01001111111101111", -- t[40943] = 6
      "0000110" when "01001111111110000", -- t[40944] = 6
      "0000110" when "01001111111110001", -- t[40945] = 6
      "0000110" when "01001111111110010", -- t[40946] = 6
      "0000110" when "01001111111110011", -- t[40947] = 6
      "0000110" when "01001111111110100", -- t[40948] = 6
      "0000110" when "01001111111110101", -- t[40949] = 6
      "0000110" when "01001111111110110", -- t[40950] = 6
      "0000110" when "01001111111110111", -- t[40951] = 6
      "0000110" when "01001111111111000", -- t[40952] = 6
      "0000110" when "01001111111111001", -- t[40953] = 6
      "0000110" when "01001111111111010", -- t[40954] = 6
      "0000110" when "01001111111111011", -- t[40955] = 6
      "0000110" when "01001111111111100", -- t[40956] = 6
      "0000110" when "01001111111111101", -- t[40957] = 6
      "0000110" when "01001111111111110", -- t[40958] = 6
      "0000110" when "01001111111111111", -- t[40959] = 6
      "0000110" when "01010000000000000", -- t[40960] = 6
      "0000110" when "01010000000000001", -- t[40961] = 6
      "0000110" when "01010000000000010", -- t[40962] = 6
      "0000110" when "01010000000000011", -- t[40963] = 6
      "0000110" when "01010000000000100", -- t[40964] = 6
      "0000110" when "01010000000000101", -- t[40965] = 6
      "0000110" when "01010000000000110", -- t[40966] = 6
      "0000110" when "01010000000000111", -- t[40967] = 6
      "0000110" when "01010000000001000", -- t[40968] = 6
      "0000110" when "01010000000001001", -- t[40969] = 6
      "0000110" when "01010000000001010", -- t[40970] = 6
      "0000110" when "01010000000001011", -- t[40971] = 6
      "0000110" when "01010000000001100", -- t[40972] = 6
      "0000110" when "01010000000001101", -- t[40973] = 6
      "0000110" when "01010000000001110", -- t[40974] = 6
      "0000110" when "01010000000001111", -- t[40975] = 6
      "0000110" when "01010000000010000", -- t[40976] = 6
      "0000110" when "01010000000010001", -- t[40977] = 6
      "0000110" when "01010000000010010", -- t[40978] = 6
      "0000110" when "01010000000010011", -- t[40979] = 6
      "0000110" when "01010000000010100", -- t[40980] = 6
      "0000110" when "01010000000010101", -- t[40981] = 6
      "0000110" when "01010000000010110", -- t[40982] = 6
      "0000110" when "01010000000010111", -- t[40983] = 6
      "0000110" when "01010000000011000", -- t[40984] = 6
      "0000110" when "01010000000011001", -- t[40985] = 6
      "0000110" when "01010000000011010", -- t[40986] = 6
      "0000110" when "01010000000011011", -- t[40987] = 6
      "0000110" when "01010000000011100", -- t[40988] = 6
      "0000110" when "01010000000011101", -- t[40989] = 6
      "0000110" when "01010000000011110", -- t[40990] = 6
      "0000110" when "01010000000011111", -- t[40991] = 6
      "0000110" when "01010000000100000", -- t[40992] = 6
      "0000110" when "01010000000100001", -- t[40993] = 6
      "0000110" when "01010000000100010", -- t[40994] = 6
      "0000110" when "01010000000100011", -- t[40995] = 6
      "0000110" when "01010000000100100", -- t[40996] = 6
      "0000110" when "01010000000100101", -- t[40997] = 6
      "0000110" when "01010000000100110", -- t[40998] = 6
      "0000110" when "01010000000100111", -- t[40999] = 6
      "0000110" when "01010000000101000", -- t[41000] = 6
      "0000110" when "01010000000101001", -- t[41001] = 6
      "0000110" when "01010000000101010", -- t[41002] = 6
      "0000110" when "01010000000101011", -- t[41003] = 6
      "0000110" when "01010000000101100", -- t[41004] = 6
      "0000110" when "01010000000101101", -- t[41005] = 6
      "0000110" when "01010000000101110", -- t[41006] = 6
      "0000110" when "01010000000101111", -- t[41007] = 6
      "0000110" when "01010000000110000", -- t[41008] = 6
      "0000110" when "01010000000110001", -- t[41009] = 6
      "0000110" when "01010000000110010", -- t[41010] = 6
      "0000110" when "01010000000110011", -- t[41011] = 6
      "0000110" when "01010000000110100", -- t[41012] = 6
      "0000110" when "01010000000110101", -- t[41013] = 6
      "0000110" when "01010000000110110", -- t[41014] = 6
      "0000110" when "01010000000110111", -- t[41015] = 6
      "0000110" when "01010000000111000", -- t[41016] = 6
      "0000110" when "01010000000111001", -- t[41017] = 6
      "0000110" when "01010000000111010", -- t[41018] = 6
      "0000110" when "01010000000111011", -- t[41019] = 6
      "0000110" when "01010000000111100", -- t[41020] = 6
      "0000110" when "01010000000111101", -- t[41021] = 6
      "0000110" when "01010000000111110", -- t[41022] = 6
      "0000110" when "01010000000111111", -- t[41023] = 6
      "0000110" when "01010000001000000", -- t[41024] = 6
      "0000110" when "01010000001000001", -- t[41025] = 6
      "0000110" when "01010000001000010", -- t[41026] = 6
      "0000110" when "01010000001000011", -- t[41027] = 6
      "0000110" when "01010000001000100", -- t[41028] = 6
      "0000110" when "01010000001000101", -- t[41029] = 6
      "0000110" when "01010000001000110", -- t[41030] = 6
      "0000110" when "01010000001000111", -- t[41031] = 6
      "0000110" when "01010000001001000", -- t[41032] = 6
      "0000110" when "01010000001001001", -- t[41033] = 6
      "0000110" when "01010000001001010", -- t[41034] = 6
      "0000110" when "01010000001001011", -- t[41035] = 6
      "0000110" when "01010000001001100", -- t[41036] = 6
      "0000110" when "01010000001001101", -- t[41037] = 6
      "0000110" when "01010000001001110", -- t[41038] = 6
      "0000110" when "01010000001001111", -- t[41039] = 6
      "0000110" when "01010000001010000", -- t[41040] = 6
      "0000110" when "01010000001010001", -- t[41041] = 6
      "0000110" when "01010000001010010", -- t[41042] = 6
      "0000110" when "01010000001010011", -- t[41043] = 6
      "0000110" when "01010000001010100", -- t[41044] = 6
      "0000110" when "01010000001010101", -- t[41045] = 6
      "0000110" when "01010000001010110", -- t[41046] = 6
      "0000110" when "01010000001010111", -- t[41047] = 6
      "0000110" when "01010000001011000", -- t[41048] = 6
      "0000110" when "01010000001011001", -- t[41049] = 6
      "0000110" when "01010000001011010", -- t[41050] = 6
      "0000110" when "01010000001011011", -- t[41051] = 6
      "0000110" when "01010000001011100", -- t[41052] = 6
      "0000110" when "01010000001011101", -- t[41053] = 6
      "0000110" when "01010000001011110", -- t[41054] = 6
      "0000110" when "01010000001011111", -- t[41055] = 6
      "0000110" when "01010000001100000", -- t[41056] = 6
      "0000110" when "01010000001100001", -- t[41057] = 6
      "0000110" when "01010000001100010", -- t[41058] = 6
      "0000110" when "01010000001100011", -- t[41059] = 6
      "0000110" when "01010000001100100", -- t[41060] = 6
      "0000110" when "01010000001100101", -- t[41061] = 6
      "0000110" when "01010000001100110", -- t[41062] = 6
      "0000110" when "01010000001100111", -- t[41063] = 6
      "0000110" when "01010000001101000", -- t[41064] = 6
      "0000110" when "01010000001101001", -- t[41065] = 6
      "0000110" when "01010000001101010", -- t[41066] = 6
      "0000110" when "01010000001101011", -- t[41067] = 6
      "0000110" when "01010000001101100", -- t[41068] = 6
      "0000110" when "01010000001101101", -- t[41069] = 6
      "0000110" when "01010000001101110", -- t[41070] = 6
      "0000110" when "01010000001101111", -- t[41071] = 6
      "0000110" when "01010000001110000", -- t[41072] = 6
      "0000110" when "01010000001110001", -- t[41073] = 6
      "0000110" when "01010000001110010", -- t[41074] = 6
      "0000110" when "01010000001110011", -- t[41075] = 6
      "0000110" when "01010000001110100", -- t[41076] = 6
      "0000110" when "01010000001110101", -- t[41077] = 6
      "0000110" when "01010000001110110", -- t[41078] = 6
      "0000110" when "01010000001110111", -- t[41079] = 6
      "0000110" when "01010000001111000", -- t[41080] = 6
      "0000110" when "01010000001111001", -- t[41081] = 6
      "0000110" when "01010000001111010", -- t[41082] = 6
      "0000110" when "01010000001111011", -- t[41083] = 6
      "0000110" when "01010000001111100", -- t[41084] = 6
      "0000110" when "01010000001111101", -- t[41085] = 6
      "0000110" when "01010000001111110", -- t[41086] = 6
      "0000110" when "01010000001111111", -- t[41087] = 6
      "0000110" when "01010000010000000", -- t[41088] = 6
      "0000110" when "01010000010000001", -- t[41089] = 6
      "0000110" when "01010000010000010", -- t[41090] = 6
      "0000110" when "01010000010000011", -- t[41091] = 6
      "0000110" when "01010000010000100", -- t[41092] = 6
      "0000110" when "01010000010000101", -- t[41093] = 6
      "0000110" when "01010000010000110", -- t[41094] = 6
      "0000110" when "01010000010000111", -- t[41095] = 6
      "0000110" when "01010000010001000", -- t[41096] = 6
      "0000110" when "01010000010001001", -- t[41097] = 6
      "0000110" when "01010000010001010", -- t[41098] = 6
      "0000110" when "01010000010001011", -- t[41099] = 6
      "0000110" when "01010000010001100", -- t[41100] = 6
      "0000110" when "01010000010001101", -- t[41101] = 6
      "0000110" when "01010000010001110", -- t[41102] = 6
      "0000110" when "01010000010001111", -- t[41103] = 6
      "0000110" when "01010000010010000", -- t[41104] = 6
      "0000110" when "01010000010010001", -- t[41105] = 6
      "0000110" when "01010000010010010", -- t[41106] = 6
      "0000110" when "01010000010010011", -- t[41107] = 6
      "0000110" when "01010000010010100", -- t[41108] = 6
      "0000110" when "01010000010010101", -- t[41109] = 6
      "0000110" when "01010000010010110", -- t[41110] = 6
      "0000110" when "01010000010010111", -- t[41111] = 6
      "0000110" when "01010000010011000", -- t[41112] = 6
      "0000110" when "01010000010011001", -- t[41113] = 6
      "0000110" when "01010000010011010", -- t[41114] = 6
      "0000110" when "01010000010011011", -- t[41115] = 6
      "0000110" when "01010000010011100", -- t[41116] = 6
      "0000110" when "01010000010011101", -- t[41117] = 6
      "0000110" when "01010000010011110", -- t[41118] = 6
      "0000110" when "01010000010011111", -- t[41119] = 6
      "0000110" when "01010000010100000", -- t[41120] = 6
      "0000110" when "01010000010100001", -- t[41121] = 6
      "0000110" when "01010000010100010", -- t[41122] = 6
      "0000110" when "01010000010100011", -- t[41123] = 6
      "0000110" when "01010000010100100", -- t[41124] = 6
      "0000110" when "01010000010100101", -- t[41125] = 6
      "0000110" when "01010000010100110", -- t[41126] = 6
      "0000110" when "01010000010100111", -- t[41127] = 6
      "0000110" when "01010000010101000", -- t[41128] = 6
      "0000110" when "01010000010101001", -- t[41129] = 6
      "0000110" when "01010000010101010", -- t[41130] = 6
      "0000110" when "01010000010101011", -- t[41131] = 6
      "0000110" when "01010000010101100", -- t[41132] = 6
      "0000110" when "01010000010101101", -- t[41133] = 6
      "0000110" when "01010000010101110", -- t[41134] = 6
      "0000110" when "01010000010101111", -- t[41135] = 6
      "0000110" when "01010000010110000", -- t[41136] = 6
      "0000110" when "01010000010110001", -- t[41137] = 6
      "0000110" when "01010000010110010", -- t[41138] = 6
      "0000110" when "01010000010110011", -- t[41139] = 6
      "0000110" when "01010000010110100", -- t[41140] = 6
      "0000110" when "01010000010110101", -- t[41141] = 6
      "0000110" when "01010000010110110", -- t[41142] = 6
      "0000110" when "01010000010110111", -- t[41143] = 6
      "0000110" when "01010000010111000", -- t[41144] = 6
      "0000110" when "01010000010111001", -- t[41145] = 6
      "0000110" when "01010000010111010", -- t[41146] = 6
      "0000110" when "01010000010111011", -- t[41147] = 6
      "0000110" when "01010000010111100", -- t[41148] = 6
      "0000110" when "01010000010111101", -- t[41149] = 6
      "0000110" when "01010000010111110", -- t[41150] = 6
      "0000110" when "01010000010111111", -- t[41151] = 6
      "0000110" when "01010000011000000", -- t[41152] = 6
      "0000110" when "01010000011000001", -- t[41153] = 6
      "0000110" when "01010000011000010", -- t[41154] = 6
      "0000110" when "01010000011000011", -- t[41155] = 6
      "0000110" when "01010000011000100", -- t[41156] = 6
      "0000110" when "01010000011000101", -- t[41157] = 6
      "0000110" when "01010000011000110", -- t[41158] = 6
      "0000110" when "01010000011000111", -- t[41159] = 6
      "0000110" when "01010000011001000", -- t[41160] = 6
      "0000110" when "01010000011001001", -- t[41161] = 6
      "0000110" when "01010000011001010", -- t[41162] = 6
      "0000110" when "01010000011001011", -- t[41163] = 6
      "0000110" when "01010000011001100", -- t[41164] = 6
      "0000110" when "01010000011001101", -- t[41165] = 6
      "0000110" when "01010000011001110", -- t[41166] = 6
      "0000110" when "01010000011001111", -- t[41167] = 6
      "0000110" when "01010000011010000", -- t[41168] = 6
      "0000110" when "01010000011010001", -- t[41169] = 6
      "0000110" when "01010000011010010", -- t[41170] = 6
      "0000110" when "01010000011010011", -- t[41171] = 6
      "0000110" when "01010000011010100", -- t[41172] = 6
      "0000110" when "01010000011010101", -- t[41173] = 6
      "0000110" when "01010000011010110", -- t[41174] = 6
      "0000110" when "01010000011010111", -- t[41175] = 6
      "0000110" when "01010000011011000", -- t[41176] = 6
      "0000110" when "01010000011011001", -- t[41177] = 6
      "0000110" when "01010000011011010", -- t[41178] = 6
      "0000110" when "01010000011011011", -- t[41179] = 6
      "0000110" when "01010000011011100", -- t[41180] = 6
      "0000110" when "01010000011011101", -- t[41181] = 6
      "0000110" when "01010000011011110", -- t[41182] = 6
      "0000110" when "01010000011011111", -- t[41183] = 6
      "0000110" when "01010000011100000", -- t[41184] = 6
      "0000110" when "01010000011100001", -- t[41185] = 6
      "0000110" when "01010000011100010", -- t[41186] = 6
      "0000110" when "01010000011100011", -- t[41187] = 6
      "0000110" when "01010000011100100", -- t[41188] = 6
      "0000110" when "01010000011100101", -- t[41189] = 6
      "0000110" when "01010000011100110", -- t[41190] = 6
      "0000110" when "01010000011100111", -- t[41191] = 6
      "0000110" when "01010000011101000", -- t[41192] = 6
      "0000110" when "01010000011101001", -- t[41193] = 6
      "0000110" when "01010000011101010", -- t[41194] = 6
      "0000110" when "01010000011101011", -- t[41195] = 6
      "0000110" when "01010000011101100", -- t[41196] = 6
      "0000110" when "01010000011101101", -- t[41197] = 6
      "0000110" when "01010000011101110", -- t[41198] = 6
      "0000110" when "01010000011101111", -- t[41199] = 6
      "0000110" when "01010000011110000", -- t[41200] = 6
      "0000110" when "01010000011110001", -- t[41201] = 6
      "0000110" when "01010000011110010", -- t[41202] = 6
      "0000110" when "01010000011110011", -- t[41203] = 6
      "0000110" when "01010000011110100", -- t[41204] = 6
      "0000110" when "01010000011110101", -- t[41205] = 6
      "0000110" when "01010000011110110", -- t[41206] = 6
      "0000110" when "01010000011110111", -- t[41207] = 6
      "0000110" when "01010000011111000", -- t[41208] = 6
      "0000110" when "01010000011111001", -- t[41209] = 6
      "0000110" when "01010000011111010", -- t[41210] = 6
      "0000110" when "01010000011111011", -- t[41211] = 6
      "0000110" when "01010000011111100", -- t[41212] = 6
      "0000110" when "01010000011111101", -- t[41213] = 6
      "0000110" when "01010000011111110", -- t[41214] = 6
      "0000110" when "01010000011111111", -- t[41215] = 6
      "0000110" when "01010000100000000", -- t[41216] = 6
      "0000110" when "01010000100000001", -- t[41217] = 6
      "0000110" when "01010000100000010", -- t[41218] = 6
      "0000110" when "01010000100000011", -- t[41219] = 6
      "0000110" when "01010000100000100", -- t[41220] = 6
      "0000110" when "01010000100000101", -- t[41221] = 6
      "0000110" when "01010000100000110", -- t[41222] = 6
      "0000110" when "01010000100000111", -- t[41223] = 6
      "0000110" when "01010000100001000", -- t[41224] = 6
      "0000110" when "01010000100001001", -- t[41225] = 6
      "0000110" when "01010000100001010", -- t[41226] = 6
      "0000110" when "01010000100001011", -- t[41227] = 6
      "0000110" when "01010000100001100", -- t[41228] = 6
      "0000110" when "01010000100001101", -- t[41229] = 6
      "0000110" when "01010000100001110", -- t[41230] = 6
      "0000110" when "01010000100001111", -- t[41231] = 6
      "0000110" when "01010000100010000", -- t[41232] = 6
      "0000110" when "01010000100010001", -- t[41233] = 6
      "0000110" when "01010000100010010", -- t[41234] = 6
      "0000110" when "01010000100010011", -- t[41235] = 6
      "0000110" when "01010000100010100", -- t[41236] = 6
      "0000110" when "01010000100010101", -- t[41237] = 6
      "0000110" when "01010000100010110", -- t[41238] = 6
      "0000110" when "01010000100010111", -- t[41239] = 6
      "0000110" when "01010000100011000", -- t[41240] = 6
      "0000110" when "01010000100011001", -- t[41241] = 6
      "0000110" when "01010000100011010", -- t[41242] = 6
      "0000110" when "01010000100011011", -- t[41243] = 6
      "0000110" when "01010000100011100", -- t[41244] = 6
      "0000110" when "01010000100011101", -- t[41245] = 6
      "0000110" when "01010000100011110", -- t[41246] = 6
      "0000110" when "01010000100011111", -- t[41247] = 6
      "0000110" when "01010000100100000", -- t[41248] = 6
      "0000110" when "01010000100100001", -- t[41249] = 6
      "0000110" when "01010000100100010", -- t[41250] = 6
      "0000110" when "01010000100100011", -- t[41251] = 6
      "0000110" when "01010000100100100", -- t[41252] = 6
      "0000110" when "01010000100100101", -- t[41253] = 6
      "0000110" when "01010000100100110", -- t[41254] = 6
      "0000110" when "01010000100100111", -- t[41255] = 6
      "0000110" when "01010000100101000", -- t[41256] = 6
      "0000110" when "01010000100101001", -- t[41257] = 6
      "0000110" when "01010000100101010", -- t[41258] = 6
      "0000110" when "01010000100101011", -- t[41259] = 6
      "0000110" when "01010000100101100", -- t[41260] = 6
      "0000110" when "01010000100101101", -- t[41261] = 6
      "0000110" when "01010000100101110", -- t[41262] = 6
      "0000110" when "01010000100101111", -- t[41263] = 6
      "0000110" when "01010000100110000", -- t[41264] = 6
      "0000110" when "01010000100110001", -- t[41265] = 6
      "0000110" when "01010000100110010", -- t[41266] = 6
      "0000110" when "01010000100110011", -- t[41267] = 6
      "0000110" when "01010000100110100", -- t[41268] = 6
      "0000110" when "01010000100110101", -- t[41269] = 6
      "0000110" when "01010000100110110", -- t[41270] = 6
      "0000110" when "01010000100110111", -- t[41271] = 6
      "0000110" when "01010000100111000", -- t[41272] = 6
      "0000110" when "01010000100111001", -- t[41273] = 6
      "0000110" when "01010000100111010", -- t[41274] = 6
      "0000110" when "01010000100111011", -- t[41275] = 6
      "0000110" when "01010000100111100", -- t[41276] = 6
      "0000110" when "01010000100111101", -- t[41277] = 6
      "0000110" when "01010000100111110", -- t[41278] = 6
      "0000110" when "01010000100111111", -- t[41279] = 6
      "0000110" when "01010000101000000", -- t[41280] = 6
      "0000110" when "01010000101000001", -- t[41281] = 6
      "0000110" when "01010000101000010", -- t[41282] = 6
      "0000110" when "01010000101000011", -- t[41283] = 6
      "0000110" when "01010000101000100", -- t[41284] = 6
      "0000110" when "01010000101000101", -- t[41285] = 6
      "0000110" when "01010000101000110", -- t[41286] = 6
      "0000110" when "01010000101000111", -- t[41287] = 6
      "0000110" when "01010000101001000", -- t[41288] = 6
      "0000110" when "01010000101001001", -- t[41289] = 6
      "0000110" when "01010000101001010", -- t[41290] = 6
      "0000110" when "01010000101001011", -- t[41291] = 6
      "0000110" when "01010000101001100", -- t[41292] = 6
      "0000110" when "01010000101001101", -- t[41293] = 6
      "0000110" when "01010000101001110", -- t[41294] = 6
      "0000110" when "01010000101001111", -- t[41295] = 6
      "0000110" when "01010000101010000", -- t[41296] = 6
      "0000110" when "01010000101010001", -- t[41297] = 6
      "0000110" when "01010000101010010", -- t[41298] = 6
      "0000110" when "01010000101010011", -- t[41299] = 6
      "0000110" when "01010000101010100", -- t[41300] = 6
      "0000110" when "01010000101010101", -- t[41301] = 6
      "0000110" when "01010000101010110", -- t[41302] = 6
      "0000110" when "01010000101010111", -- t[41303] = 6
      "0000110" when "01010000101011000", -- t[41304] = 6
      "0000110" when "01010000101011001", -- t[41305] = 6
      "0000110" when "01010000101011010", -- t[41306] = 6
      "0000110" when "01010000101011011", -- t[41307] = 6
      "0000110" when "01010000101011100", -- t[41308] = 6
      "0000110" when "01010000101011101", -- t[41309] = 6
      "0000110" when "01010000101011110", -- t[41310] = 6
      "0000110" when "01010000101011111", -- t[41311] = 6
      "0000110" when "01010000101100000", -- t[41312] = 6
      "0000110" when "01010000101100001", -- t[41313] = 6
      "0000110" when "01010000101100010", -- t[41314] = 6
      "0000110" when "01010000101100011", -- t[41315] = 6
      "0000110" when "01010000101100100", -- t[41316] = 6
      "0000110" when "01010000101100101", -- t[41317] = 6
      "0000110" when "01010000101100110", -- t[41318] = 6
      "0000110" when "01010000101100111", -- t[41319] = 6
      "0000110" when "01010000101101000", -- t[41320] = 6
      "0000110" when "01010000101101001", -- t[41321] = 6
      "0000110" when "01010000101101010", -- t[41322] = 6
      "0000110" when "01010000101101011", -- t[41323] = 6
      "0000110" when "01010000101101100", -- t[41324] = 6
      "0000110" when "01010000101101101", -- t[41325] = 6
      "0000110" when "01010000101101110", -- t[41326] = 6
      "0000110" when "01010000101101111", -- t[41327] = 6
      "0000110" when "01010000101110000", -- t[41328] = 6
      "0000110" when "01010000101110001", -- t[41329] = 6
      "0000110" when "01010000101110010", -- t[41330] = 6
      "0000110" when "01010000101110011", -- t[41331] = 6
      "0000110" when "01010000101110100", -- t[41332] = 6
      "0000110" when "01010000101110101", -- t[41333] = 6
      "0000110" when "01010000101110110", -- t[41334] = 6
      "0000110" when "01010000101110111", -- t[41335] = 6
      "0000110" when "01010000101111000", -- t[41336] = 6
      "0000110" when "01010000101111001", -- t[41337] = 6
      "0000110" when "01010000101111010", -- t[41338] = 6
      "0000110" when "01010000101111011", -- t[41339] = 6
      "0000110" when "01010000101111100", -- t[41340] = 6
      "0000110" when "01010000101111101", -- t[41341] = 6
      "0000110" when "01010000101111110", -- t[41342] = 6
      "0000110" when "01010000101111111", -- t[41343] = 6
      "0000110" when "01010000110000000", -- t[41344] = 6
      "0000110" when "01010000110000001", -- t[41345] = 6
      "0000110" when "01010000110000010", -- t[41346] = 6
      "0000110" when "01010000110000011", -- t[41347] = 6
      "0000110" when "01010000110000100", -- t[41348] = 6
      "0000110" when "01010000110000101", -- t[41349] = 6
      "0000110" when "01010000110000110", -- t[41350] = 6
      "0000110" when "01010000110000111", -- t[41351] = 6
      "0000110" when "01010000110001000", -- t[41352] = 6
      "0000110" when "01010000110001001", -- t[41353] = 6
      "0000110" when "01010000110001010", -- t[41354] = 6
      "0000110" when "01010000110001011", -- t[41355] = 6
      "0000110" when "01010000110001100", -- t[41356] = 6
      "0000110" when "01010000110001101", -- t[41357] = 6
      "0000110" when "01010000110001110", -- t[41358] = 6
      "0000110" when "01010000110001111", -- t[41359] = 6
      "0000110" when "01010000110010000", -- t[41360] = 6
      "0000110" when "01010000110010001", -- t[41361] = 6
      "0000110" when "01010000110010010", -- t[41362] = 6
      "0000110" when "01010000110010011", -- t[41363] = 6
      "0000110" when "01010000110010100", -- t[41364] = 6
      "0000110" when "01010000110010101", -- t[41365] = 6
      "0000110" when "01010000110010110", -- t[41366] = 6
      "0000110" when "01010000110010111", -- t[41367] = 6
      "0000110" when "01010000110011000", -- t[41368] = 6
      "0000110" when "01010000110011001", -- t[41369] = 6
      "0000110" when "01010000110011010", -- t[41370] = 6
      "0000110" when "01010000110011011", -- t[41371] = 6
      "0000110" when "01010000110011100", -- t[41372] = 6
      "0000110" when "01010000110011101", -- t[41373] = 6
      "0000110" when "01010000110011110", -- t[41374] = 6
      "0000110" when "01010000110011111", -- t[41375] = 6
      "0000110" when "01010000110100000", -- t[41376] = 6
      "0000110" when "01010000110100001", -- t[41377] = 6
      "0000110" when "01010000110100010", -- t[41378] = 6
      "0000110" when "01010000110100011", -- t[41379] = 6
      "0000110" when "01010000110100100", -- t[41380] = 6
      "0000110" when "01010000110100101", -- t[41381] = 6
      "0000110" when "01010000110100110", -- t[41382] = 6
      "0000110" when "01010000110100111", -- t[41383] = 6
      "0000110" when "01010000110101000", -- t[41384] = 6
      "0000110" when "01010000110101001", -- t[41385] = 6
      "0000110" when "01010000110101010", -- t[41386] = 6
      "0000110" when "01010000110101011", -- t[41387] = 6
      "0000110" when "01010000110101100", -- t[41388] = 6
      "0000110" when "01010000110101101", -- t[41389] = 6
      "0000110" when "01010000110101110", -- t[41390] = 6
      "0000110" when "01010000110101111", -- t[41391] = 6
      "0000110" when "01010000110110000", -- t[41392] = 6
      "0000110" when "01010000110110001", -- t[41393] = 6
      "0000110" when "01010000110110010", -- t[41394] = 6
      "0000110" when "01010000110110011", -- t[41395] = 6
      "0000110" when "01010000110110100", -- t[41396] = 6
      "0000110" when "01010000110110101", -- t[41397] = 6
      "0000110" when "01010000110110110", -- t[41398] = 6
      "0000110" when "01010000110110111", -- t[41399] = 6
      "0000110" when "01010000110111000", -- t[41400] = 6
      "0000110" when "01010000110111001", -- t[41401] = 6
      "0000110" when "01010000110111010", -- t[41402] = 6
      "0000110" when "01010000110111011", -- t[41403] = 6
      "0000110" when "01010000110111100", -- t[41404] = 6
      "0000110" when "01010000110111101", -- t[41405] = 6
      "0000110" when "01010000110111110", -- t[41406] = 6
      "0000110" when "01010000110111111", -- t[41407] = 6
      "0000110" when "01010000111000000", -- t[41408] = 6
      "0000110" when "01010000111000001", -- t[41409] = 6
      "0000110" when "01010000111000010", -- t[41410] = 6
      "0000110" when "01010000111000011", -- t[41411] = 6
      "0000110" when "01010000111000100", -- t[41412] = 6
      "0000110" when "01010000111000101", -- t[41413] = 6
      "0000110" when "01010000111000110", -- t[41414] = 6
      "0000110" when "01010000111000111", -- t[41415] = 6
      "0000110" when "01010000111001000", -- t[41416] = 6
      "0000110" when "01010000111001001", -- t[41417] = 6
      "0000110" when "01010000111001010", -- t[41418] = 6
      "0000110" when "01010000111001011", -- t[41419] = 6
      "0000110" when "01010000111001100", -- t[41420] = 6
      "0000110" when "01010000111001101", -- t[41421] = 6
      "0000110" when "01010000111001110", -- t[41422] = 6
      "0000110" when "01010000111001111", -- t[41423] = 6
      "0000110" when "01010000111010000", -- t[41424] = 6
      "0000110" when "01010000111010001", -- t[41425] = 6
      "0000110" when "01010000111010010", -- t[41426] = 6
      "0000110" when "01010000111010011", -- t[41427] = 6
      "0000110" when "01010000111010100", -- t[41428] = 6
      "0000110" when "01010000111010101", -- t[41429] = 6
      "0000110" when "01010000111010110", -- t[41430] = 6
      "0000110" when "01010000111010111", -- t[41431] = 6
      "0000110" when "01010000111011000", -- t[41432] = 6
      "0000110" when "01010000111011001", -- t[41433] = 6
      "0000110" when "01010000111011010", -- t[41434] = 6
      "0000110" when "01010000111011011", -- t[41435] = 6
      "0000110" when "01010000111011100", -- t[41436] = 6
      "0000110" when "01010000111011101", -- t[41437] = 6
      "0000110" when "01010000111011110", -- t[41438] = 6
      "0000110" when "01010000111011111", -- t[41439] = 6
      "0000110" when "01010000111100000", -- t[41440] = 6
      "0000110" when "01010000111100001", -- t[41441] = 6
      "0000110" when "01010000111100010", -- t[41442] = 6
      "0000110" when "01010000111100011", -- t[41443] = 6
      "0000110" when "01010000111100100", -- t[41444] = 6
      "0000110" when "01010000111100101", -- t[41445] = 6
      "0000110" when "01010000111100110", -- t[41446] = 6
      "0000110" when "01010000111100111", -- t[41447] = 6
      "0000110" when "01010000111101000", -- t[41448] = 6
      "0000110" when "01010000111101001", -- t[41449] = 6
      "0000110" when "01010000111101010", -- t[41450] = 6
      "0000110" when "01010000111101011", -- t[41451] = 6
      "0000110" when "01010000111101100", -- t[41452] = 6
      "0000110" when "01010000111101101", -- t[41453] = 6
      "0000110" when "01010000111101110", -- t[41454] = 6
      "0000110" when "01010000111101111", -- t[41455] = 6
      "0000110" when "01010000111110000", -- t[41456] = 6
      "0000110" when "01010000111110001", -- t[41457] = 6
      "0000110" when "01010000111110010", -- t[41458] = 6
      "0000110" when "01010000111110011", -- t[41459] = 6
      "0000110" when "01010000111110100", -- t[41460] = 6
      "0000110" when "01010000111110101", -- t[41461] = 6
      "0000110" when "01010000111110110", -- t[41462] = 6
      "0000110" when "01010000111110111", -- t[41463] = 6
      "0000110" when "01010000111111000", -- t[41464] = 6
      "0000110" when "01010000111111001", -- t[41465] = 6
      "0000110" when "01010000111111010", -- t[41466] = 6
      "0000110" when "01010000111111011", -- t[41467] = 6
      "0000110" when "01010000111111100", -- t[41468] = 6
      "0000110" when "01010000111111101", -- t[41469] = 6
      "0000110" when "01010000111111110", -- t[41470] = 6
      "0000110" when "01010000111111111", -- t[41471] = 6
      "0000110" when "01010001000000000", -- t[41472] = 6
      "0000110" when "01010001000000001", -- t[41473] = 6
      "0000110" when "01010001000000010", -- t[41474] = 6
      "0000110" when "01010001000000011", -- t[41475] = 6
      "0000110" when "01010001000000100", -- t[41476] = 6
      "0000110" when "01010001000000101", -- t[41477] = 6
      "0000110" when "01010001000000110", -- t[41478] = 6
      "0000110" when "01010001000000111", -- t[41479] = 6
      "0000110" when "01010001000001000", -- t[41480] = 6
      "0000110" when "01010001000001001", -- t[41481] = 6
      "0000110" when "01010001000001010", -- t[41482] = 6
      "0000110" when "01010001000001011", -- t[41483] = 6
      "0000110" when "01010001000001100", -- t[41484] = 6
      "0000110" when "01010001000001101", -- t[41485] = 6
      "0000110" when "01010001000001110", -- t[41486] = 6
      "0000110" when "01010001000001111", -- t[41487] = 6
      "0000110" when "01010001000010000", -- t[41488] = 6
      "0000110" when "01010001000010001", -- t[41489] = 6
      "0000110" when "01010001000010010", -- t[41490] = 6
      "0000110" when "01010001000010011", -- t[41491] = 6
      "0000110" when "01010001000010100", -- t[41492] = 6
      "0000110" when "01010001000010101", -- t[41493] = 6
      "0000110" when "01010001000010110", -- t[41494] = 6
      "0000110" when "01010001000010111", -- t[41495] = 6
      "0000110" when "01010001000011000", -- t[41496] = 6
      "0000110" when "01010001000011001", -- t[41497] = 6
      "0000110" when "01010001000011010", -- t[41498] = 6
      "0000110" when "01010001000011011", -- t[41499] = 6
      "0000110" when "01010001000011100", -- t[41500] = 6
      "0000110" when "01010001000011101", -- t[41501] = 6
      "0000110" when "01010001000011110", -- t[41502] = 6
      "0000110" when "01010001000011111", -- t[41503] = 6
      "0000110" when "01010001000100000", -- t[41504] = 6
      "0000110" when "01010001000100001", -- t[41505] = 6
      "0000110" when "01010001000100010", -- t[41506] = 6
      "0000110" when "01010001000100011", -- t[41507] = 6
      "0000110" when "01010001000100100", -- t[41508] = 6
      "0000110" when "01010001000100101", -- t[41509] = 6
      "0000110" when "01010001000100110", -- t[41510] = 6
      "0000110" when "01010001000100111", -- t[41511] = 6
      "0000110" when "01010001000101000", -- t[41512] = 6
      "0000110" when "01010001000101001", -- t[41513] = 6
      "0000110" when "01010001000101010", -- t[41514] = 6
      "0000110" when "01010001000101011", -- t[41515] = 6
      "0000110" when "01010001000101100", -- t[41516] = 6
      "0000110" when "01010001000101101", -- t[41517] = 6
      "0000110" when "01010001000101110", -- t[41518] = 6
      "0000110" when "01010001000101111", -- t[41519] = 6
      "0000110" when "01010001000110000", -- t[41520] = 6
      "0000110" when "01010001000110001", -- t[41521] = 6
      "0000110" when "01010001000110010", -- t[41522] = 6
      "0000110" when "01010001000110011", -- t[41523] = 6
      "0000110" when "01010001000110100", -- t[41524] = 6
      "0000110" when "01010001000110101", -- t[41525] = 6
      "0000110" when "01010001000110110", -- t[41526] = 6
      "0000110" when "01010001000110111", -- t[41527] = 6
      "0000110" when "01010001000111000", -- t[41528] = 6
      "0000110" when "01010001000111001", -- t[41529] = 6
      "0000110" when "01010001000111010", -- t[41530] = 6
      "0000110" when "01010001000111011", -- t[41531] = 6
      "0000110" when "01010001000111100", -- t[41532] = 6
      "0000110" when "01010001000111101", -- t[41533] = 6
      "0000110" when "01010001000111110", -- t[41534] = 6
      "0000110" when "01010001000111111", -- t[41535] = 6
      "0000110" when "01010001001000000", -- t[41536] = 6
      "0000110" when "01010001001000001", -- t[41537] = 6
      "0000110" when "01010001001000010", -- t[41538] = 6
      "0000110" when "01010001001000011", -- t[41539] = 6
      "0000110" when "01010001001000100", -- t[41540] = 6
      "0000110" when "01010001001000101", -- t[41541] = 6
      "0000110" when "01010001001000110", -- t[41542] = 6
      "0000110" when "01010001001000111", -- t[41543] = 6
      "0000110" when "01010001001001000", -- t[41544] = 6
      "0000110" when "01010001001001001", -- t[41545] = 6
      "0000110" when "01010001001001010", -- t[41546] = 6
      "0000110" when "01010001001001011", -- t[41547] = 6
      "0000110" when "01010001001001100", -- t[41548] = 6
      "0000110" when "01010001001001101", -- t[41549] = 6
      "0000110" when "01010001001001110", -- t[41550] = 6
      "0000110" when "01010001001001111", -- t[41551] = 6
      "0000110" when "01010001001010000", -- t[41552] = 6
      "0000110" when "01010001001010001", -- t[41553] = 6
      "0000110" when "01010001001010010", -- t[41554] = 6
      "0000110" when "01010001001010011", -- t[41555] = 6
      "0000110" when "01010001001010100", -- t[41556] = 6
      "0000110" when "01010001001010101", -- t[41557] = 6
      "0000110" when "01010001001010110", -- t[41558] = 6
      "0000110" when "01010001001010111", -- t[41559] = 6
      "0000110" when "01010001001011000", -- t[41560] = 6
      "0000110" when "01010001001011001", -- t[41561] = 6
      "0000110" when "01010001001011010", -- t[41562] = 6
      "0000110" when "01010001001011011", -- t[41563] = 6
      "0000110" when "01010001001011100", -- t[41564] = 6
      "0000110" when "01010001001011101", -- t[41565] = 6
      "0000110" when "01010001001011110", -- t[41566] = 6
      "0000110" when "01010001001011111", -- t[41567] = 6
      "0000110" when "01010001001100000", -- t[41568] = 6
      "0000110" when "01010001001100001", -- t[41569] = 6
      "0000110" when "01010001001100010", -- t[41570] = 6
      "0000110" when "01010001001100011", -- t[41571] = 6
      "0000110" when "01010001001100100", -- t[41572] = 6
      "0000110" when "01010001001100101", -- t[41573] = 6
      "0000110" when "01010001001100110", -- t[41574] = 6
      "0000110" when "01010001001100111", -- t[41575] = 6
      "0000110" when "01010001001101000", -- t[41576] = 6
      "0000110" when "01010001001101001", -- t[41577] = 6
      "0000110" when "01010001001101010", -- t[41578] = 6
      "0000110" when "01010001001101011", -- t[41579] = 6
      "0000110" when "01010001001101100", -- t[41580] = 6
      "0000110" when "01010001001101101", -- t[41581] = 6
      "0000110" when "01010001001101110", -- t[41582] = 6
      "0000110" when "01010001001101111", -- t[41583] = 6
      "0000110" when "01010001001110000", -- t[41584] = 6
      "0000110" when "01010001001110001", -- t[41585] = 6
      "0000110" when "01010001001110010", -- t[41586] = 6
      "0000110" when "01010001001110011", -- t[41587] = 6
      "0000110" when "01010001001110100", -- t[41588] = 6
      "0000110" when "01010001001110101", -- t[41589] = 6
      "0000110" when "01010001001110110", -- t[41590] = 6
      "0000110" when "01010001001110111", -- t[41591] = 6
      "0000110" when "01010001001111000", -- t[41592] = 6
      "0000110" when "01010001001111001", -- t[41593] = 6
      "0000110" when "01010001001111010", -- t[41594] = 6
      "0000110" when "01010001001111011", -- t[41595] = 6
      "0000110" when "01010001001111100", -- t[41596] = 6
      "0000110" when "01010001001111101", -- t[41597] = 6
      "0000110" when "01010001001111110", -- t[41598] = 6
      "0000110" when "01010001001111111", -- t[41599] = 6
      "0000110" when "01010001010000000", -- t[41600] = 6
      "0000110" when "01010001010000001", -- t[41601] = 6
      "0000110" when "01010001010000010", -- t[41602] = 6
      "0000110" when "01010001010000011", -- t[41603] = 6
      "0000110" when "01010001010000100", -- t[41604] = 6
      "0000110" when "01010001010000101", -- t[41605] = 6
      "0000110" when "01010001010000110", -- t[41606] = 6
      "0000110" when "01010001010000111", -- t[41607] = 6
      "0000110" when "01010001010001000", -- t[41608] = 6
      "0000110" when "01010001010001001", -- t[41609] = 6
      "0000110" when "01010001010001010", -- t[41610] = 6
      "0000110" when "01010001010001011", -- t[41611] = 6
      "0000110" when "01010001010001100", -- t[41612] = 6
      "0000110" when "01010001010001101", -- t[41613] = 6
      "0000110" when "01010001010001110", -- t[41614] = 6
      "0000110" when "01010001010001111", -- t[41615] = 6
      "0000110" when "01010001010010000", -- t[41616] = 6
      "0000110" when "01010001010010001", -- t[41617] = 6
      "0000110" when "01010001010010010", -- t[41618] = 6
      "0000110" when "01010001010010011", -- t[41619] = 6
      "0000110" when "01010001010010100", -- t[41620] = 6
      "0000110" when "01010001010010101", -- t[41621] = 6
      "0000110" when "01010001010010110", -- t[41622] = 6
      "0000110" when "01010001010010111", -- t[41623] = 6
      "0000110" when "01010001010011000", -- t[41624] = 6
      "0000110" when "01010001010011001", -- t[41625] = 6
      "0000110" when "01010001010011010", -- t[41626] = 6
      "0000110" when "01010001010011011", -- t[41627] = 6
      "0000110" when "01010001010011100", -- t[41628] = 6
      "0000110" when "01010001010011101", -- t[41629] = 6
      "0000110" when "01010001010011110", -- t[41630] = 6
      "0000110" when "01010001010011111", -- t[41631] = 6
      "0000110" when "01010001010100000", -- t[41632] = 6
      "0000110" when "01010001010100001", -- t[41633] = 6
      "0000110" when "01010001010100010", -- t[41634] = 6
      "0000110" when "01010001010100011", -- t[41635] = 6
      "0000110" when "01010001010100100", -- t[41636] = 6
      "0000110" when "01010001010100101", -- t[41637] = 6
      "0000110" when "01010001010100110", -- t[41638] = 6
      "0000110" when "01010001010100111", -- t[41639] = 6
      "0000110" when "01010001010101000", -- t[41640] = 6
      "0000110" when "01010001010101001", -- t[41641] = 6
      "0000110" when "01010001010101010", -- t[41642] = 6
      "0000110" when "01010001010101011", -- t[41643] = 6
      "0000110" when "01010001010101100", -- t[41644] = 6
      "0000110" when "01010001010101101", -- t[41645] = 6
      "0000110" when "01010001010101110", -- t[41646] = 6
      "0000110" when "01010001010101111", -- t[41647] = 6
      "0000110" when "01010001010110000", -- t[41648] = 6
      "0000110" when "01010001010110001", -- t[41649] = 6
      "0000110" when "01010001010110010", -- t[41650] = 6
      "0000110" when "01010001010110011", -- t[41651] = 6
      "0000110" when "01010001010110100", -- t[41652] = 6
      "0000110" when "01010001010110101", -- t[41653] = 6
      "0000110" when "01010001010110110", -- t[41654] = 6
      "0000110" when "01010001010110111", -- t[41655] = 6
      "0000110" when "01010001010111000", -- t[41656] = 6
      "0000110" when "01010001010111001", -- t[41657] = 6
      "0000110" when "01010001010111010", -- t[41658] = 6
      "0000110" when "01010001010111011", -- t[41659] = 6
      "0000110" when "01010001010111100", -- t[41660] = 6
      "0000110" when "01010001010111101", -- t[41661] = 6
      "0000110" when "01010001010111110", -- t[41662] = 6
      "0000110" when "01010001010111111", -- t[41663] = 6
      "0000110" when "01010001011000000", -- t[41664] = 6
      "0000110" when "01010001011000001", -- t[41665] = 6
      "0000110" when "01010001011000010", -- t[41666] = 6
      "0000110" when "01010001011000011", -- t[41667] = 6
      "0000110" when "01010001011000100", -- t[41668] = 6
      "0000110" when "01010001011000101", -- t[41669] = 6
      "0000110" when "01010001011000110", -- t[41670] = 6
      "0000110" when "01010001011000111", -- t[41671] = 6
      "0000110" when "01010001011001000", -- t[41672] = 6
      "0000110" when "01010001011001001", -- t[41673] = 6
      "0000110" when "01010001011001010", -- t[41674] = 6
      "0000110" when "01010001011001011", -- t[41675] = 6
      "0000110" when "01010001011001100", -- t[41676] = 6
      "0000110" when "01010001011001101", -- t[41677] = 6
      "0000110" when "01010001011001110", -- t[41678] = 6
      "0000110" when "01010001011001111", -- t[41679] = 6
      "0000110" when "01010001011010000", -- t[41680] = 6
      "0000110" when "01010001011010001", -- t[41681] = 6
      "0000110" when "01010001011010010", -- t[41682] = 6
      "0000110" when "01010001011010011", -- t[41683] = 6
      "0000110" when "01010001011010100", -- t[41684] = 6
      "0000110" when "01010001011010101", -- t[41685] = 6
      "0000110" when "01010001011010110", -- t[41686] = 6
      "0000110" when "01010001011010111", -- t[41687] = 6
      "0000110" when "01010001011011000", -- t[41688] = 6
      "0000110" when "01010001011011001", -- t[41689] = 6
      "0000110" when "01010001011011010", -- t[41690] = 6
      "0000110" when "01010001011011011", -- t[41691] = 6
      "0000110" when "01010001011011100", -- t[41692] = 6
      "0000110" when "01010001011011101", -- t[41693] = 6
      "0000110" when "01010001011011110", -- t[41694] = 6
      "0000110" when "01010001011011111", -- t[41695] = 6
      "0000110" when "01010001011100000", -- t[41696] = 6
      "0000110" when "01010001011100001", -- t[41697] = 6
      "0000110" when "01010001011100010", -- t[41698] = 6
      "0000110" when "01010001011100011", -- t[41699] = 6
      "0000110" when "01010001011100100", -- t[41700] = 6
      "0000110" when "01010001011100101", -- t[41701] = 6
      "0000110" when "01010001011100110", -- t[41702] = 6
      "0000110" when "01010001011100111", -- t[41703] = 6
      "0000110" when "01010001011101000", -- t[41704] = 6
      "0000110" when "01010001011101001", -- t[41705] = 6
      "0000110" when "01010001011101010", -- t[41706] = 6
      "0000110" when "01010001011101011", -- t[41707] = 6
      "0000110" when "01010001011101100", -- t[41708] = 6
      "0000110" when "01010001011101101", -- t[41709] = 6
      "0000110" when "01010001011101110", -- t[41710] = 6
      "0000110" when "01010001011101111", -- t[41711] = 6
      "0000110" when "01010001011110000", -- t[41712] = 6
      "0000110" when "01010001011110001", -- t[41713] = 6
      "0000110" when "01010001011110010", -- t[41714] = 6
      "0000110" when "01010001011110011", -- t[41715] = 6
      "0000110" when "01010001011110100", -- t[41716] = 6
      "0000110" when "01010001011110101", -- t[41717] = 6
      "0000110" when "01010001011110110", -- t[41718] = 6
      "0000110" when "01010001011110111", -- t[41719] = 6
      "0000110" when "01010001011111000", -- t[41720] = 6
      "0000110" when "01010001011111001", -- t[41721] = 6
      "0000110" when "01010001011111010", -- t[41722] = 6
      "0000110" when "01010001011111011", -- t[41723] = 6
      "0000110" when "01010001011111100", -- t[41724] = 6
      "0000110" when "01010001011111101", -- t[41725] = 6
      "0000110" when "01010001011111110", -- t[41726] = 6
      "0000110" when "01010001011111111", -- t[41727] = 6
      "0000110" when "01010001100000000", -- t[41728] = 6
      "0000110" when "01010001100000001", -- t[41729] = 6
      "0000110" when "01010001100000010", -- t[41730] = 6
      "0000110" when "01010001100000011", -- t[41731] = 6
      "0000110" when "01010001100000100", -- t[41732] = 6
      "0000110" when "01010001100000101", -- t[41733] = 6
      "0000110" when "01010001100000110", -- t[41734] = 6
      "0000110" when "01010001100000111", -- t[41735] = 6
      "0000110" when "01010001100001000", -- t[41736] = 6
      "0000110" when "01010001100001001", -- t[41737] = 6
      "0000110" when "01010001100001010", -- t[41738] = 6
      "0000110" when "01010001100001011", -- t[41739] = 6
      "0000110" when "01010001100001100", -- t[41740] = 6
      "0000110" when "01010001100001101", -- t[41741] = 6
      "0000110" when "01010001100001110", -- t[41742] = 6
      "0000110" when "01010001100001111", -- t[41743] = 6
      "0000110" when "01010001100010000", -- t[41744] = 6
      "0000110" when "01010001100010001", -- t[41745] = 6
      "0000110" when "01010001100010010", -- t[41746] = 6
      "0000110" when "01010001100010011", -- t[41747] = 6
      "0000110" when "01010001100010100", -- t[41748] = 6
      "0000110" when "01010001100010101", -- t[41749] = 6
      "0000110" when "01010001100010110", -- t[41750] = 6
      "0000110" when "01010001100010111", -- t[41751] = 6
      "0000110" when "01010001100011000", -- t[41752] = 6
      "0000110" when "01010001100011001", -- t[41753] = 6
      "0000110" when "01010001100011010", -- t[41754] = 6
      "0000110" when "01010001100011011", -- t[41755] = 6
      "0000110" when "01010001100011100", -- t[41756] = 6
      "0000110" when "01010001100011101", -- t[41757] = 6
      "0000110" when "01010001100011110", -- t[41758] = 6
      "0000110" when "01010001100011111", -- t[41759] = 6
      "0000110" when "01010001100100000", -- t[41760] = 6
      "0000110" when "01010001100100001", -- t[41761] = 6
      "0000110" when "01010001100100010", -- t[41762] = 6
      "0000110" when "01010001100100011", -- t[41763] = 6
      "0000110" when "01010001100100100", -- t[41764] = 6
      "0000110" when "01010001100100101", -- t[41765] = 6
      "0000110" when "01010001100100110", -- t[41766] = 6
      "0000110" when "01010001100100111", -- t[41767] = 6
      "0000110" when "01010001100101000", -- t[41768] = 6
      "0000110" when "01010001100101001", -- t[41769] = 6
      "0000110" when "01010001100101010", -- t[41770] = 6
      "0000110" when "01010001100101011", -- t[41771] = 6
      "0000110" when "01010001100101100", -- t[41772] = 6
      "0000110" when "01010001100101101", -- t[41773] = 6
      "0000110" when "01010001100101110", -- t[41774] = 6
      "0000110" when "01010001100101111", -- t[41775] = 6
      "0000110" when "01010001100110000", -- t[41776] = 6
      "0000110" when "01010001100110001", -- t[41777] = 6
      "0000110" when "01010001100110010", -- t[41778] = 6
      "0000110" when "01010001100110011", -- t[41779] = 6
      "0000110" when "01010001100110100", -- t[41780] = 6
      "0000110" when "01010001100110101", -- t[41781] = 6
      "0000110" when "01010001100110110", -- t[41782] = 6
      "0000110" when "01010001100110111", -- t[41783] = 6
      "0000110" when "01010001100111000", -- t[41784] = 6
      "0000110" when "01010001100111001", -- t[41785] = 6
      "0000110" when "01010001100111010", -- t[41786] = 6
      "0000110" when "01010001100111011", -- t[41787] = 6
      "0000110" when "01010001100111100", -- t[41788] = 6
      "0000110" when "01010001100111101", -- t[41789] = 6
      "0000110" when "01010001100111110", -- t[41790] = 6
      "0000110" when "01010001100111111", -- t[41791] = 6
      "0000110" when "01010001101000000", -- t[41792] = 6
      "0000110" when "01010001101000001", -- t[41793] = 6
      "0000110" when "01010001101000010", -- t[41794] = 6
      "0000110" when "01010001101000011", -- t[41795] = 6
      "0000110" when "01010001101000100", -- t[41796] = 6
      "0000110" when "01010001101000101", -- t[41797] = 6
      "0000110" when "01010001101000110", -- t[41798] = 6
      "0000110" when "01010001101000111", -- t[41799] = 6
      "0000110" when "01010001101001000", -- t[41800] = 6
      "0000110" when "01010001101001001", -- t[41801] = 6
      "0000110" when "01010001101001010", -- t[41802] = 6
      "0000110" when "01010001101001011", -- t[41803] = 6
      "0000110" when "01010001101001100", -- t[41804] = 6
      "0000110" when "01010001101001101", -- t[41805] = 6
      "0000110" when "01010001101001110", -- t[41806] = 6
      "0000110" when "01010001101001111", -- t[41807] = 6
      "0000110" when "01010001101010000", -- t[41808] = 6
      "0000110" when "01010001101010001", -- t[41809] = 6
      "0000110" when "01010001101010010", -- t[41810] = 6
      "0000110" when "01010001101010011", -- t[41811] = 6
      "0000110" when "01010001101010100", -- t[41812] = 6
      "0000110" when "01010001101010101", -- t[41813] = 6
      "0000110" when "01010001101010110", -- t[41814] = 6
      "0000110" when "01010001101010111", -- t[41815] = 6
      "0000110" when "01010001101011000", -- t[41816] = 6
      "0000110" when "01010001101011001", -- t[41817] = 6
      "0000110" when "01010001101011010", -- t[41818] = 6
      "0000110" when "01010001101011011", -- t[41819] = 6
      "0000110" when "01010001101011100", -- t[41820] = 6
      "0000110" when "01010001101011101", -- t[41821] = 6
      "0000110" when "01010001101011110", -- t[41822] = 6
      "0000110" when "01010001101011111", -- t[41823] = 6
      "0000110" when "01010001101100000", -- t[41824] = 6
      "0000110" when "01010001101100001", -- t[41825] = 6
      "0000110" when "01010001101100010", -- t[41826] = 6
      "0000110" when "01010001101100011", -- t[41827] = 6
      "0000110" when "01010001101100100", -- t[41828] = 6
      "0000110" when "01010001101100101", -- t[41829] = 6
      "0000110" when "01010001101100110", -- t[41830] = 6
      "0000110" when "01010001101100111", -- t[41831] = 6
      "0000110" when "01010001101101000", -- t[41832] = 6
      "0000110" when "01010001101101001", -- t[41833] = 6
      "0000110" when "01010001101101010", -- t[41834] = 6
      "0000110" when "01010001101101011", -- t[41835] = 6
      "0000110" when "01010001101101100", -- t[41836] = 6
      "0000110" when "01010001101101101", -- t[41837] = 6
      "0000110" when "01010001101101110", -- t[41838] = 6
      "0000110" when "01010001101101111", -- t[41839] = 6
      "0000110" when "01010001101110000", -- t[41840] = 6
      "0000110" when "01010001101110001", -- t[41841] = 6
      "0000110" when "01010001101110010", -- t[41842] = 6
      "0000110" when "01010001101110011", -- t[41843] = 6
      "0000110" when "01010001101110100", -- t[41844] = 6
      "0000110" when "01010001101110101", -- t[41845] = 6
      "0000110" when "01010001101110110", -- t[41846] = 6
      "0000110" when "01010001101110111", -- t[41847] = 6
      "0000110" when "01010001101111000", -- t[41848] = 6
      "0000110" when "01010001101111001", -- t[41849] = 6
      "0000110" when "01010001101111010", -- t[41850] = 6
      "0000110" when "01010001101111011", -- t[41851] = 6
      "0000110" when "01010001101111100", -- t[41852] = 6
      "0000110" when "01010001101111101", -- t[41853] = 6
      "0000110" when "01010001101111110", -- t[41854] = 6
      "0000110" when "01010001101111111", -- t[41855] = 6
      "0000110" when "01010001110000000", -- t[41856] = 6
      "0000110" when "01010001110000001", -- t[41857] = 6
      "0000110" when "01010001110000010", -- t[41858] = 6
      "0000110" when "01010001110000011", -- t[41859] = 6
      "0000110" when "01010001110000100", -- t[41860] = 6
      "0000110" when "01010001110000101", -- t[41861] = 6
      "0000110" when "01010001110000110", -- t[41862] = 6
      "0000110" when "01010001110000111", -- t[41863] = 6
      "0000110" when "01010001110001000", -- t[41864] = 6
      "0000110" when "01010001110001001", -- t[41865] = 6
      "0000110" when "01010001110001010", -- t[41866] = 6
      "0000110" when "01010001110001011", -- t[41867] = 6
      "0000110" when "01010001110001100", -- t[41868] = 6
      "0000110" when "01010001110001101", -- t[41869] = 6
      "0000110" when "01010001110001110", -- t[41870] = 6
      "0000110" when "01010001110001111", -- t[41871] = 6
      "0000110" when "01010001110010000", -- t[41872] = 6
      "0000110" when "01010001110010001", -- t[41873] = 6
      "0000110" when "01010001110010010", -- t[41874] = 6
      "0000110" when "01010001110010011", -- t[41875] = 6
      "0000110" when "01010001110010100", -- t[41876] = 6
      "0000110" when "01010001110010101", -- t[41877] = 6
      "0000110" when "01010001110010110", -- t[41878] = 6
      "0000110" when "01010001110010111", -- t[41879] = 6
      "0000110" when "01010001110011000", -- t[41880] = 6
      "0000110" when "01010001110011001", -- t[41881] = 6
      "0000110" when "01010001110011010", -- t[41882] = 6
      "0000110" when "01010001110011011", -- t[41883] = 6
      "0000110" when "01010001110011100", -- t[41884] = 6
      "0000110" when "01010001110011101", -- t[41885] = 6
      "0000110" when "01010001110011110", -- t[41886] = 6
      "0000110" when "01010001110011111", -- t[41887] = 6
      "0000110" when "01010001110100000", -- t[41888] = 6
      "0000110" when "01010001110100001", -- t[41889] = 6
      "0000110" when "01010001110100010", -- t[41890] = 6
      "0000110" when "01010001110100011", -- t[41891] = 6
      "0000110" when "01010001110100100", -- t[41892] = 6
      "0000110" when "01010001110100101", -- t[41893] = 6
      "0000110" when "01010001110100110", -- t[41894] = 6
      "0000110" when "01010001110100111", -- t[41895] = 6
      "0000110" when "01010001110101000", -- t[41896] = 6
      "0000110" when "01010001110101001", -- t[41897] = 6
      "0000110" when "01010001110101010", -- t[41898] = 6
      "0000110" when "01010001110101011", -- t[41899] = 6
      "0000110" when "01010001110101100", -- t[41900] = 6
      "0000110" when "01010001110101101", -- t[41901] = 6
      "0000110" when "01010001110101110", -- t[41902] = 6
      "0000110" when "01010001110101111", -- t[41903] = 6
      "0000110" when "01010001110110000", -- t[41904] = 6
      "0000110" when "01010001110110001", -- t[41905] = 6
      "0000110" when "01010001110110010", -- t[41906] = 6
      "0000110" when "01010001110110011", -- t[41907] = 6
      "0000110" when "01010001110110100", -- t[41908] = 6
      "0000110" when "01010001110110101", -- t[41909] = 6
      "0000110" when "01010001110110110", -- t[41910] = 6
      "0000110" when "01010001110110111", -- t[41911] = 6
      "0000110" when "01010001110111000", -- t[41912] = 6
      "0000110" when "01010001110111001", -- t[41913] = 6
      "0000110" when "01010001110111010", -- t[41914] = 6
      "0000110" when "01010001110111011", -- t[41915] = 6
      "0000110" when "01010001110111100", -- t[41916] = 6
      "0000110" when "01010001110111101", -- t[41917] = 6
      "0000110" when "01010001110111110", -- t[41918] = 6
      "0000110" when "01010001110111111", -- t[41919] = 6
      "0000110" when "01010001111000000", -- t[41920] = 6
      "0000110" when "01010001111000001", -- t[41921] = 6
      "0000110" when "01010001111000010", -- t[41922] = 6
      "0000110" when "01010001111000011", -- t[41923] = 6
      "0000110" when "01010001111000100", -- t[41924] = 6
      "0000110" when "01010001111000101", -- t[41925] = 6
      "0000110" when "01010001111000110", -- t[41926] = 6
      "0000110" when "01010001111000111", -- t[41927] = 6
      "0000110" when "01010001111001000", -- t[41928] = 6
      "0000110" when "01010001111001001", -- t[41929] = 6
      "0000110" when "01010001111001010", -- t[41930] = 6
      "0000110" when "01010001111001011", -- t[41931] = 6
      "0000110" when "01010001111001100", -- t[41932] = 6
      "0000110" when "01010001111001101", -- t[41933] = 6
      "0000110" when "01010001111001110", -- t[41934] = 6
      "0000110" when "01010001111001111", -- t[41935] = 6
      "0000110" when "01010001111010000", -- t[41936] = 6
      "0000110" when "01010001111010001", -- t[41937] = 6
      "0000110" when "01010001111010010", -- t[41938] = 6
      "0000110" when "01010001111010011", -- t[41939] = 6
      "0000110" when "01010001111010100", -- t[41940] = 6
      "0000110" when "01010001111010101", -- t[41941] = 6
      "0000110" when "01010001111010110", -- t[41942] = 6
      "0000110" when "01010001111010111", -- t[41943] = 6
      "0000110" when "01010001111011000", -- t[41944] = 6
      "0000110" when "01010001111011001", -- t[41945] = 6
      "0000110" when "01010001111011010", -- t[41946] = 6
      "0000110" when "01010001111011011", -- t[41947] = 6
      "0000110" when "01010001111011100", -- t[41948] = 6
      "0000110" when "01010001111011101", -- t[41949] = 6
      "0000110" when "01010001111011110", -- t[41950] = 6
      "0000110" when "01010001111011111", -- t[41951] = 6
      "0000110" when "01010001111100000", -- t[41952] = 6
      "0000110" when "01010001111100001", -- t[41953] = 6
      "0000110" when "01010001111100010", -- t[41954] = 6
      "0000110" when "01010001111100011", -- t[41955] = 6
      "0000110" when "01010001111100100", -- t[41956] = 6
      "0000110" when "01010001111100101", -- t[41957] = 6
      "0000110" when "01010001111100110", -- t[41958] = 6
      "0000110" when "01010001111100111", -- t[41959] = 6
      "0000110" when "01010001111101000", -- t[41960] = 6
      "0000110" when "01010001111101001", -- t[41961] = 6
      "0000110" when "01010001111101010", -- t[41962] = 6
      "0000110" when "01010001111101011", -- t[41963] = 6
      "0000110" when "01010001111101100", -- t[41964] = 6
      "0000110" when "01010001111101101", -- t[41965] = 6
      "0000110" when "01010001111101110", -- t[41966] = 6
      "0000110" when "01010001111101111", -- t[41967] = 6
      "0000110" when "01010001111110000", -- t[41968] = 6
      "0000110" when "01010001111110001", -- t[41969] = 6
      "0000110" when "01010001111110010", -- t[41970] = 6
      "0000110" when "01010001111110011", -- t[41971] = 6
      "0000110" when "01010001111110100", -- t[41972] = 6
      "0000110" when "01010001111110101", -- t[41973] = 6
      "0000110" when "01010001111110110", -- t[41974] = 6
      "0000110" when "01010001111110111", -- t[41975] = 6
      "0000110" when "01010001111111000", -- t[41976] = 6
      "0000110" when "01010001111111001", -- t[41977] = 6
      "0000110" when "01010001111111010", -- t[41978] = 6
      "0000110" when "01010001111111011", -- t[41979] = 6
      "0000110" when "01010001111111100", -- t[41980] = 6
      "0000110" when "01010001111111101", -- t[41981] = 6
      "0000110" when "01010001111111110", -- t[41982] = 6
      "0000110" when "01010001111111111", -- t[41983] = 6
      "0000110" when "01010010000000000", -- t[41984] = 6
      "0000110" when "01010010000000001", -- t[41985] = 6
      "0000110" when "01010010000000010", -- t[41986] = 6
      "0000110" when "01010010000000011", -- t[41987] = 6
      "0000110" when "01010010000000100", -- t[41988] = 6
      "0000110" when "01010010000000101", -- t[41989] = 6
      "0000110" when "01010010000000110", -- t[41990] = 6
      "0000110" when "01010010000000111", -- t[41991] = 6
      "0000110" when "01010010000001000", -- t[41992] = 6
      "0000110" when "01010010000001001", -- t[41993] = 6
      "0000110" when "01010010000001010", -- t[41994] = 6
      "0000110" when "01010010000001011", -- t[41995] = 6
      "0000110" when "01010010000001100", -- t[41996] = 6
      "0000110" when "01010010000001101", -- t[41997] = 6
      "0000110" when "01010010000001110", -- t[41998] = 6
      "0000110" when "01010010000001111", -- t[41999] = 6
      "0000110" when "01010010000010000", -- t[42000] = 6
      "0000110" when "01010010000010001", -- t[42001] = 6
      "0000110" when "01010010000010010", -- t[42002] = 6
      "0000110" when "01010010000010011", -- t[42003] = 6
      "0000110" when "01010010000010100", -- t[42004] = 6
      "0000110" when "01010010000010101", -- t[42005] = 6
      "0000110" when "01010010000010110", -- t[42006] = 6
      "0000110" when "01010010000010111", -- t[42007] = 6
      "0000110" when "01010010000011000", -- t[42008] = 6
      "0000110" when "01010010000011001", -- t[42009] = 6
      "0000110" when "01010010000011010", -- t[42010] = 6
      "0000110" when "01010010000011011", -- t[42011] = 6
      "0000110" when "01010010000011100", -- t[42012] = 6
      "0000110" when "01010010000011101", -- t[42013] = 6
      "0000110" when "01010010000011110", -- t[42014] = 6
      "0000110" when "01010010000011111", -- t[42015] = 6
      "0000110" when "01010010000100000", -- t[42016] = 6
      "0000110" when "01010010000100001", -- t[42017] = 6
      "0000110" when "01010010000100010", -- t[42018] = 6
      "0000110" when "01010010000100011", -- t[42019] = 6
      "0000110" when "01010010000100100", -- t[42020] = 6
      "0000110" when "01010010000100101", -- t[42021] = 6
      "0000110" when "01010010000100110", -- t[42022] = 6
      "0000110" when "01010010000100111", -- t[42023] = 6
      "0000110" when "01010010000101000", -- t[42024] = 6
      "0000110" when "01010010000101001", -- t[42025] = 6
      "0000110" when "01010010000101010", -- t[42026] = 6
      "0000110" when "01010010000101011", -- t[42027] = 6
      "0000110" when "01010010000101100", -- t[42028] = 6
      "0000110" when "01010010000101101", -- t[42029] = 6
      "0000110" when "01010010000101110", -- t[42030] = 6
      "0000110" when "01010010000101111", -- t[42031] = 6
      "0000110" when "01010010000110000", -- t[42032] = 6
      "0000110" when "01010010000110001", -- t[42033] = 6
      "0000110" when "01010010000110010", -- t[42034] = 6
      "0000110" when "01010010000110011", -- t[42035] = 6
      "0000110" when "01010010000110100", -- t[42036] = 6
      "0000110" when "01010010000110101", -- t[42037] = 6
      "0000110" when "01010010000110110", -- t[42038] = 6
      "0000110" when "01010010000110111", -- t[42039] = 6
      "0000110" when "01010010000111000", -- t[42040] = 6
      "0000110" when "01010010000111001", -- t[42041] = 6
      "0000110" when "01010010000111010", -- t[42042] = 6
      "0000110" when "01010010000111011", -- t[42043] = 6
      "0000110" when "01010010000111100", -- t[42044] = 6
      "0000110" when "01010010000111101", -- t[42045] = 6
      "0000110" when "01010010000111110", -- t[42046] = 6
      "0000110" when "01010010000111111", -- t[42047] = 6
      "0000110" when "01010010001000000", -- t[42048] = 6
      "0000110" when "01010010001000001", -- t[42049] = 6
      "0000110" when "01010010001000010", -- t[42050] = 6
      "0000110" when "01010010001000011", -- t[42051] = 6
      "0000110" when "01010010001000100", -- t[42052] = 6
      "0000110" when "01010010001000101", -- t[42053] = 6
      "0000110" when "01010010001000110", -- t[42054] = 6
      "0000110" when "01010010001000111", -- t[42055] = 6
      "0000110" when "01010010001001000", -- t[42056] = 6
      "0000110" when "01010010001001001", -- t[42057] = 6
      "0000110" when "01010010001001010", -- t[42058] = 6
      "0000110" when "01010010001001011", -- t[42059] = 6
      "0000110" when "01010010001001100", -- t[42060] = 6
      "0000110" when "01010010001001101", -- t[42061] = 6
      "0000110" when "01010010001001110", -- t[42062] = 6
      "0000110" when "01010010001001111", -- t[42063] = 6
      "0000110" when "01010010001010000", -- t[42064] = 6
      "0000110" when "01010010001010001", -- t[42065] = 6
      "0000110" when "01010010001010010", -- t[42066] = 6
      "0000110" when "01010010001010011", -- t[42067] = 6
      "0000110" when "01010010001010100", -- t[42068] = 6
      "0000110" when "01010010001010101", -- t[42069] = 6
      "0000110" when "01010010001010110", -- t[42070] = 6
      "0000110" when "01010010001010111", -- t[42071] = 6
      "0000110" when "01010010001011000", -- t[42072] = 6
      "0000110" when "01010010001011001", -- t[42073] = 6
      "0000110" when "01010010001011010", -- t[42074] = 6
      "0000110" when "01010010001011011", -- t[42075] = 6
      "0000110" when "01010010001011100", -- t[42076] = 6
      "0000110" when "01010010001011101", -- t[42077] = 6
      "0000110" when "01010010001011110", -- t[42078] = 6
      "0000110" when "01010010001011111", -- t[42079] = 6
      "0000110" when "01010010001100000", -- t[42080] = 6
      "0000110" when "01010010001100001", -- t[42081] = 6
      "0000110" when "01010010001100010", -- t[42082] = 6
      "0000110" when "01010010001100011", -- t[42083] = 6
      "0000110" when "01010010001100100", -- t[42084] = 6
      "0000110" when "01010010001100101", -- t[42085] = 6
      "0000110" when "01010010001100110", -- t[42086] = 6
      "0000110" when "01010010001100111", -- t[42087] = 6
      "0000110" when "01010010001101000", -- t[42088] = 6
      "0000110" when "01010010001101001", -- t[42089] = 6
      "0000110" when "01010010001101010", -- t[42090] = 6
      "0000110" when "01010010001101011", -- t[42091] = 6
      "0000110" when "01010010001101100", -- t[42092] = 6
      "0000110" when "01010010001101101", -- t[42093] = 6
      "0000110" when "01010010001101110", -- t[42094] = 6
      "0000110" when "01010010001101111", -- t[42095] = 6
      "0000110" when "01010010001110000", -- t[42096] = 6
      "0000110" when "01010010001110001", -- t[42097] = 6
      "0000110" when "01010010001110010", -- t[42098] = 6
      "0000110" when "01010010001110011", -- t[42099] = 6
      "0000110" when "01010010001110100", -- t[42100] = 6
      "0000110" when "01010010001110101", -- t[42101] = 6
      "0000110" when "01010010001110110", -- t[42102] = 6
      "0000110" when "01010010001110111", -- t[42103] = 6
      "0000110" when "01010010001111000", -- t[42104] = 6
      "0000110" when "01010010001111001", -- t[42105] = 6
      "0000110" when "01010010001111010", -- t[42106] = 6
      "0000110" when "01010010001111011", -- t[42107] = 6
      "0000110" when "01010010001111100", -- t[42108] = 6
      "0000110" when "01010010001111101", -- t[42109] = 6
      "0000110" when "01010010001111110", -- t[42110] = 6
      "0000110" when "01010010001111111", -- t[42111] = 6
      "0000110" when "01010010010000000", -- t[42112] = 6
      "0000110" when "01010010010000001", -- t[42113] = 6
      "0000110" when "01010010010000010", -- t[42114] = 6
      "0000110" when "01010010010000011", -- t[42115] = 6
      "0000110" when "01010010010000100", -- t[42116] = 6
      "0000110" when "01010010010000101", -- t[42117] = 6
      "0000110" when "01010010010000110", -- t[42118] = 6
      "0000110" when "01010010010000111", -- t[42119] = 6
      "0000110" when "01010010010001000", -- t[42120] = 6
      "0000110" when "01010010010001001", -- t[42121] = 6
      "0000110" when "01010010010001010", -- t[42122] = 6
      "0000110" when "01010010010001011", -- t[42123] = 6
      "0000110" when "01010010010001100", -- t[42124] = 6
      "0000110" when "01010010010001101", -- t[42125] = 6
      "0000110" when "01010010010001110", -- t[42126] = 6
      "0000110" when "01010010010001111", -- t[42127] = 6
      "0000110" when "01010010010010000", -- t[42128] = 6
      "0000110" when "01010010010010001", -- t[42129] = 6
      "0000110" when "01010010010010010", -- t[42130] = 6
      "0000110" when "01010010010010011", -- t[42131] = 6
      "0000110" when "01010010010010100", -- t[42132] = 6
      "0000110" when "01010010010010101", -- t[42133] = 6
      "0000110" when "01010010010010110", -- t[42134] = 6
      "0000110" when "01010010010010111", -- t[42135] = 6
      "0000110" when "01010010010011000", -- t[42136] = 6
      "0000110" when "01010010010011001", -- t[42137] = 6
      "0000110" when "01010010010011010", -- t[42138] = 6
      "0000110" when "01010010010011011", -- t[42139] = 6
      "0000110" when "01010010010011100", -- t[42140] = 6
      "0000110" when "01010010010011101", -- t[42141] = 6
      "0000110" when "01010010010011110", -- t[42142] = 6
      "0000110" when "01010010010011111", -- t[42143] = 6
      "0000110" when "01010010010100000", -- t[42144] = 6
      "0000110" when "01010010010100001", -- t[42145] = 6
      "0000110" when "01010010010100010", -- t[42146] = 6
      "0000110" when "01010010010100011", -- t[42147] = 6
      "0000110" when "01010010010100100", -- t[42148] = 6
      "0000110" when "01010010010100101", -- t[42149] = 6
      "0000110" when "01010010010100110", -- t[42150] = 6
      "0000110" when "01010010010100111", -- t[42151] = 6
      "0000110" when "01010010010101000", -- t[42152] = 6
      "0000110" when "01010010010101001", -- t[42153] = 6
      "0000110" when "01010010010101010", -- t[42154] = 6
      "0000110" when "01010010010101011", -- t[42155] = 6
      "0000110" when "01010010010101100", -- t[42156] = 6
      "0000110" when "01010010010101101", -- t[42157] = 6
      "0000110" when "01010010010101110", -- t[42158] = 6
      "0000110" when "01010010010101111", -- t[42159] = 6
      "0000110" when "01010010010110000", -- t[42160] = 6
      "0000110" when "01010010010110001", -- t[42161] = 6
      "0000110" when "01010010010110010", -- t[42162] = 6
      "0000110" when "01010010010110011", -- t[42163] = 6
      "0000110" when "01010010010110100", -- t[42164] = 6
      "0000110" when "01010010010110101", -- t[42165] = 6
      "0000110" when "01010010010110110", -- t[42166] = 6
      "0000110" when "01010010010110111", -- t[42167] = 6
      "0000110" when "01010010010111000", -- t[42168] = 6
      "0000110" when "01010010010111001", -- t[42169] = 6
      "0000110" when "01010010010111010", -- t[42170] = 6
      "0000110" when "01010010010111011", -- t[42171] = 6
      "0000110" when "01010010010111100", -- t[42172] = 6
      "0000110" when "01010010010111101", -- t[42173] = 6
      "0000110" when "01010010010111110", -- t[42174] = 6
      "0000110" when "01010010010111111", -- t[42175] = 6
      "0000110" when "01010010011000000", -- t[42176] = 6
      "0000110" when "01010010011000001", -- t[42177] = 6
      "0000110" when "01010010011000010", -- t[42178] = 6
      "0000110" when "01010010011000011", -- t[42179] = 6
      "0000110" when "01010010011000100", -- t[42180] = 6
      "0000110" when "01010010011000101", -- t[42181] = 6
      "0000110" when "01010010011000110", -- t[42182] = 6
      "0000110" when "01010010011000111", -- t[42183] = 6
      "0000110" when "01010010011001000", -- t[42184] = 6
      "0000110" when "01010010011001001", -- t[42185] = 6
      "0000110" when "01010010011001010", -- t[42186] = 6
      "0000110" when "01010010011001011", -- t[42187] = 6
      "0000110" when "01010010011001100", -- t[42188] = 6
      "0000110" when "01010010011001101", -- t[42189] = 6
      "0000110" when "01010010011001110", -- t[42190] = 6
      "0000110" when "01010010011001111", -- t[42191] = 6
      "0000110" when "01010010011010000", -- t[42192] = 6
      "0000110" when "01010010011010001", -- t[42193] = 6
      "0000110" when "01010010011010010", -- t[42194] = 6
      "0000110" when "01010010011010011", -- t[42195] = 6
      "0000110" when "01010010011010100", -- t[42196] = 6
      "0000110" when "01010010011010101", -- t[42197] = 6
      "0000110" when "01010010011010110", -- t[42198] = 6
      "0000110" when "01010010011010111", -- t[42199] = 6
      "0000110" when "01010010011011000", -- t[42200] = 6
      "0000110" when "01010010011011001", -- t[42201] = 6
      "0000110" when "01010010011011010", -- t[42202] = 6
      "0000110" when "01010010011011011", -- t[42203] = 6
      "0000110" when "01010010011011100", -- t[42204] = 6
      "0000110" when "01010010011011101", -- t[42205] = 6
      "0000110" when "01010010011011110", -- t[42206] = 6
      "0000110" when "01010010011011111", -- t[42207] = 6
      "0000110" when "01010010011100000", -- t[42208] = 6
      "0000110" when "01010010011100001", -- t[42209] = 6
      "0000110" when "01010010011100010", -- t[42210] = 6
      "0000110" when "01010010011100011", -- t[42211] = 6
      "0000110" when "01010010011100100", -- t[42212] = 6
      "0000110" when "01010010011100101", -- t[42213] = 6
      "0000110" when "01010010011100110", -- t[42214] = 6
      "0000110" when "01010010011100111", -- t[42215] = 6
      "0000110" when "01010010011101000", -- t[42216] = 6
      "0000110" when "01010010011101001", -- t[42217] = 6
      "0000110" when "01010010011101010", -- t[42218] = 6
      "0000110" when "01010010011101011", -- t[42219] = 6
      "0000110" when "01010010011101100", -- t[42220] = 6
      "0000110" when "01010010011101101", -- t[42221] = 6
      "0000110" when "01010010011101110", -- t[42222] = 6
      "0000110" when "01010010011101111", -- t[42223] = 6
      "0000110" when "01010010011110000", -- t[42224] = 6
      "0000110" when "01010010011110001", -- t[42225] = 6
      "0000110" when "01010010011110010", -- t[42226] = 6
      "0000110" when "01010010011110011", -- t[42227] = 6
      "0000110" when "01010010011110100", -- t[42228] = 6
      "0000110" when "01010010011110101", -- t[42229] = 6
      "0000110" when "01010010011110110", -- t[42230] = 6
      "0000110" when "01010010011110111", -- t[42231] = 6
      "0000110" when "01010010011111000", -- t[42232] = 6
      "0000110" when "01010010011111001", -- t[42233] = 6
      "0000110" when "01010010011111010", -- t[42234] = 6
      "0000110" when "01010010011111011", -- t[42235] = 6
      "0000110" when "01010010011111100", -- t[42236] = 6
      "0000110" when "01010010011111101", -- t[42237] = 6
      "0000110" when "01010010011111110", -- t[42238] = 6
      "0000110" when "01010010011111111", -- t[42239] = 6
      "0000110" when "01010010100000000", -- t[42240] = 6
      "0000110" when "01010010100000001", -- t[42241] = 6
      "0000110" when "01010010100000010", -- t[42242] = 6
      "0000110" when "01010010100000011", -- t[42243] = 6
      "0000110" when "01010010100000100", -- t[42244] = 6
      "0000110" when "01010010100000101", -- t[42245] = 6
      "0000110" when "01010010100000110", -- t[42246] = 6
      "0000110" when "01010010100000111", -- t[42247] = 6
      "0000110" when "01010010100001000", -- t[42248] = 6
      "0000110" when "01010010100001001", -- t[42249] = 6
      "0000110" when "01010010100001010", -- t[42250] = 6
      "0000110" when "01010010100001011", -- t[42251] = 6
      "0000110" when "01010010100001100", -- t[42252] = 6
      "0000110" when "01010010100001101", -- t[42253] = 6
      "0000110" when "01010010100001110", -- t[42254] = 6
      "0000110" when "01010010100001111", -- t[42255] = 6
      "0000110" when "01010010100010000", -- t[42256] = 6
      "0000110" when "01010010100010001", -- t[42257] = 6
      "0000110" when "01010010100010010", -- t[42258] = 6
      "0000110" when "01010010100010011", -- t[42259] = 6
      "0000110" when "01010010100010100", -- t[42260] = 6
      "0000110" when "01010010100010101", -- t[42261] = 6
      "0000110" when "01010010100010110", -- t[42262] = 6
      "0000110" when "01010010100010111", -- t[42263] = 6
      "0000110" when "01010010100011000", -- t[42264] = 6
      "0000110" when "01010010100011001", -- t[42265] = 6
      "0000110" when "01010010100011010", -- t[42266] = 6
      "0000110" when "01010010100011011", -- t[42267] = 6
      "0000110" when "01010010100011100", -- t[42268] = 6
      "0000110" when "01010010100011101", -- t[42269] = 6
      "0000110" when "01010010100011110", -- t[42270] = 6
      "0000110" when "01010010100011111", -- t[42271] = 6
      "0000110" when "01010010100100000", -- t[42272] = 6
      "0000110" when "01010010100100001", -- t[42273] = 6
      "0000110" when "01010010100100010", -- t[42274] = 6
      "0000110" when "01010010100100011", -- t[42275] = 6
      "0000110" when "01010010100100100", -- t[42276] = 6
      "0000110" when "01010010100100101", -- t[42277] = 6
      "0000110" when "01010010100100110", -- t[42278] = 6
      "0000110" when "01010010100100111", -- t[42279] = 6
      "0000110" when "01010010100101000", -- t[42280] = 6
      "0000110" when "01010010100101001", -- t[42281] = 6
      "0000110" when "01010010100101010", -- t[42282] = 6
      "0000110" when "01010010100101011", -- t[42283] = 6
      "0000110" when "01010010100101100", -- t[42284] = 6
      "0000110" when "01010010100101101", -- t[42285] = 6
      "0000110" when "01010010100101110", -- t[42286] = 6
      "0000110" when "01010010100101111", -- t[42287] = 6
      "0000110" when "01010010100110000", -- t[42288] = 6
      "0000110" when "01010010100110001", -- t[42289] = 6
      "0000110" when "01010010100110010", -- t[42290] = 6
      "0000110" when "01010010100110011", -- t[42291] = 6
      "0000110" when "01010010100110100", -- t[42292] = 6
      "0000110" when "01010010100110101", -- t[42293] = 6
      "0000110" when "01010010100110110", -- t[42294] = 6
      "0000110" when "01010010100110111", -- t[42295] = 6
      "0000110" when "01010010100111000", -- t[42296] = 6
      "0000110" when "01010010100111001", -- t[42297] = 6
      "0000110" when "01010010100111010", -- t[42298] = 6
      "0000110" when "01010010100111011", -- t[42299] = 6
      "0000110" when "01010010100111100", -- t[42300] = 6
      "0000110" when "01010010100111101", -- t[42301] = 6
      "0000110" when "01010010100111110", -- t[42302] = 6
      "0000110" when "01010010100111111", -- t[42303] = 6
      "0000110" when "01010010101000000", -- t[42304] = 6
      "0000110" when "01010010101000001", -- t[42305] = 6
      "0000110" when "01010010101000010", -- t[42306] = 6
      "0000110" when "01010010101000011", -- t[42307] = 6
      "0000110" when "01010010101000100", -- t[42308] = 6
      "0000110" when "01010010101000101", -- t[42309] = 6
      "0000110" when "01010010101000110", -- t[42310] = 6
      "0000110" when "01010010101000111", -- t[42311] = 6
      "0000110" when "01010010101001000", -- t[42312] = 6
      "0000110" when "01010010101001001", -- t[42313] = 6
      "0000110" when "01010010101001010", -- t[42314] = 6
      "0000110" when "01010010101001011", -- t[42315] = 6
      "0000110" when "01010010101001100", -- t[42316] = 6
      "0000110" when "01010010101001101", -- t[42317] = 6
      "0000110" when "01010010101001110", -- t[42318] = 6
      "0000110" when "01010010101001111", -- t[42319] = 6
      "0000110" when "01010010101010000", -- t[42320] = 6
      "0000110" when "01010010101010001", -- t[42321] = 6
      "0000110" when "01010010101010010", -- t[42322] = 6
      "0000110" when "01010010101010011", -- t[42323] = 6
      "0000110" when "01010010101010100", -- t[42324] = 6
      "0000110" when "01010010101010101", -- t[42325] = 6
      "0000110" when "01010010101010110", -- t[42326] = 6
      "0000110" when "01010010101010111", -- t[42327] = 6
      "0000110" when "01010010101011000", -- t[42328] = 6
      "0000110" when "01010010101011001", -- t[42329] = 6
      "0000110" when "01010010101011010", -- t[42330] = 6
      "0000110" when "01010010101011011", -- t[42331] = 6
      "0000110" when "01010010101011100", -- t[42332] = 6
      "0000110" when "01010010101011101", -- t[42333] = 6
      "0000110" when "01010010101011110", -- t[42334] = 6
      "0000110" when "01010010101011111", -- t[42335] = 6
      "0000110" when "01010010101100000", -- t[42336] = 6
      "0000110" when "01010010101100001", -- t[42337] = 6
      "0000110" when "01010010101100010", -- t[42338] = 6
      "0000110" when "01010010101100011", -- t[42339] = 6
      "0000110" when "01010010101100100", -- t[42340] = 6
      "0000110" when "01010010101100101", -- t[42341] = 6
      "0000110" when "01010010101100110", -- t[42342] = 6
      "0000110" when "01010010101100111", -- t[42343] = 6
      "0000110" when "01010010101101000", -- t[42344] = 6
      "0000110" when "01010010101101001", -- t[42345] = 6
      "0000110" when "01010010101101010", -- t[42346] = 6
      "0000110" when "01010010101101011", -- t[42347] = 6
      "0000110" when "01010010101101100", -- t[42348] = 6
      "0000110" when "01010010101101101", -- t[42349] = 6
      "0000110" when "01010010101101110", -- t[42350] = 6
      "0000110" when "01010010101101111", -- t[42351] = 6
      "0000110" when "01010010101110000", -- t[42352] = 6
      "0000110" when "01010010101110001", -- t[42353] = 6
      "0000110" when "01010010101110010", -- t[42354] = 6
      "0000110" when "01010010101110011", -- t[42355] = 6
      "0000110" when "01010010101110100", -- t[42356] = 6
      "0000110" when "01010010101110101", -- t[42357] = 6
      "0000110" when "01010010101110110", -- t[42358] = 6
      "0000110" when "01010010101110111", -- t[42359] = 6
      "0000110" when "01010010101111000", -- t[42360] = 6
      "0000110" when "01010010101111001", -- t[42361] = 6
      "0000110" when "01010010101111010", -- t[42362] = 6
      "0000110" when "01010010101111011", -- t[42363] = 6
      "0000111" when "01010010101111100", -- t[42364] = 7
      "0000111" when "01010010101111101", -- t[42365] = 7
      "0000111" when "01010010101111110", -- t[42366] = 7
      "0000111" when "01010010101111111", -- t[42367] = 7
      "0000111" when "01010010110000000", -- t[42368] = 7
      "0000111" when "01010010110000001", -- t[42369] = 7
      "0000111" when "01010010110000010", -- t[42370] = 7
      "0000111" when "01010010110000011", -- t[42371] = 7
      "0000111" when "01010010110000100", -- t[42372] = 7
      "0000111" when "01010010110000101", -- t[42373] = 7
      "0000111" when "01010010110000110", -- t[42374] = 7
      "0000111" when "01010010110000111", -- t[42375] = 7
      "0000111" when "01010010110001000", -- t[42376] = 7
      "0000111" when "01010010110001001", -- t[42377] = 7
      "0000111" when "01010010110001010", -- t[42378] = 7
      "0000111" when "01010010110001011", -- t[42379] = 7
      "0000111" when "01010010110001100", -- t[42380] = 7
      "0000111" when "01010010110001101", -- t[42381] = 7
      "0000111" when "01010010110001110", -- t[42382] = 7
      "0000111" when "01010010110001111", -- t[42383] = 7
      "0000111" when "01010010110010000", -- t[42384] = 7
      "0000111" when "01010010110010001", -- t[42385] = 7
      "0000111" when "01010010110010010", -- t[42386] = 7
      "0000111" when "01010010110010011", -- t[42387] = 7
      "0000111" when "01010010110010100", -- t[42388] = 7
      "0000111" when "01010010110010101", -- t[42389] = 7
      "0000111" when "01010010110010110", -- t[42390] = 7
      "0000111" when "01010010110010111", -- t[42391] = 7
      "0000111" when "01010010110011000", -- t[42392] = 7
      "0000111" when "01010010110011001", -- t[42393] = 7
      "0000111" when "01010010110011010", -- t[42394] = 7
      "0000111" when "01010010110011011", -- t[42395] = 7
      "0000111" when "01010010110011100", -- t[42396] = 7
      "0000111" when "01010010110011101", -- t[42397] = 7
      "0000111" when "01010010110011110", -- t[42398] = 7
      "0000111" when "01010010110011111", -- t[42399] = 7
      "0000111" when "01010010110100000", -- t[42400] = 7
      "0000111" when "01010010110100001", -- t[42401] = 7
      "0000111" when "01010010110100010", -- t[42402] = 7
      "0000111" when "01010010110100011", -- t[42403] = 7
      "0000111" when "01010010110100100", -- t[42404] = 7
      "0000111" when "01010010110100101", -- t[42405] = 7
      "0000111" when "01010010110100110", -- t[42406] = 7
      "0000111" when "01010010110100111", -- t[42407] = 7
      "0000111" when "01010010110101000", -- t[42408] = 7
      "0000111" when "01010010110101001", -- t[42409] = 7
      "0000111" when "01010010110101010", -- t[42410] = 7
      "0000111" when "01010010110101011", -- t[42411] = 7
      "0000111" when "01010010110101100", -- t[42412] = 7
      "0000111" when "01010010110101101", -- t[42413] = 7
      "0000111" when "01010010110101110", -- t[42414] = 7
      "0000111" when "01010010110101111", -- t[42415] = 7
      "0000111" when "01010010110110000", -- t[42416] = 7
      "0000111" when "01010010110110001", -- t[42417] = 7
      "0000111" when "01010010110110010", -- t[42418] = 7
      "0000111" when "01010010110110011", -- t[42419] = 7
      "0000111" when "01010010110110100", -- t[42420] = 7
      "0000111" when "01010010110110101", -- t[42421] = 7
      "0000111" when "01010010110110110", -- t[42422] = 7
      "0000111" when "01010010110110111", -- t[42423] = 7
      "0000111" when "01010010110111000", -- t[42424] = 7
      "0000111" when "01010010110111001", -- t[42425] = 7
      "0000111" when "01010010110111010", -- t[42426] = 7
      "0000111" when "01010010110111011", -- t[42427] = 7
      "0000111" when "01010010110111100", -- t[42428] = 7
      "0000111" when "01010010110111101", -- t[42429] = 7
      "0000111" when "01010010110111110", -- t[42430] = 7
      "0000111" when "01010010110111111", -- t[42431] = 7
      "0000111" when "01010010111000000", -- t[42432] = 7
      "0000111" when "01010010111000001", -- t[42433] = 7
      "0000111" when "01010010111000010", -- t[42434] = 7
      "0000111" when "01010010111000011", -- t[42435] = 7
      "0000111" when "01010010111000100", -- t[42436] = 7
      "0000111" when "01010010111000101", -- t[42437] = 7
      "0000111" when "01010010111000110", -- t[42438] = 7
      "0000111" when "01010010111000111", -- t[42439] = 7
      "0000111" when "01010010111001000", -- t[42440] = 7
      "0000111" when "01010010111001001", -- t[42441] = 7
      "0000111" when "01010010111001010", -- t[42442] = 7
      "0000111" when "01010010111001011", -- t[42443] = 7
      "0000111" when "01010010111001100", -- t[42444] = 7
      "0000111" when "01010010111001101", -- t[42445] = 7
      "0000111" when "01010010111001110", -- t[42446] = 7
      "0000111" when "01010010111001111", -- t[42447] = 7
      "0000111" when "01010010111010000", -- t[42448] = 7
      "0000111" when "01010010111010001", -- t[42449] = 7
      "0000111" when "01010010111010010", -- t[42450] = 7
      "0000111" when "01010010111010011", -- t[42451] = 7
      "0000111" when "01010010111010100", -- t[42452] = 7
      "0000111" when "01010010111010101", -- t[42453] = 7
      "0000111" when "01010010111010110", -- t[42454] = 7
      "0000111" when "01010010111010111", -- t[42455] = 7
      "0000111" when "01010010111011000", -- t[42456] = 7
      "0000111" when "01010010111011001", -- t[42457] = 7
      "0000111" when "01010010111011010", -- t[42458] = 7
      "0000111" when "01010010111011011", -- t[42459] = 7
      "0000111" when "01010010111011100", -- t[42460] = 7
      "0000111" when "01010010111011101", -- t[42461] = 7
      "0000111" when "01010010111011110", -- t[42462] = 7
      "0000111" when "01010010111011111", -- t[42463] = 7
      "0000111" when "01010010111100000", -- t[42464] = 7
      "0000111" when "01010010111100001", -- t[42465] = 7
      "0000111" when "01010010111100010", -- t[42466] = 7
      "0000111" when "01010010111100011", -- t[42467] = 7
      "0000111" when "01010010111100100", -- t[42468] = 7
      "0000111" when "01010010111100101", -- t[42469] = 7
      "0000111" when "01010010111100110", -- t[42470] = 7
      "0000111" when "01010010111100111", -- t[42471] = 7
      "0000111" when "01010010111101000", -- t[42472] = 7
      "0000111" when "01010010111101001", -- t[42473] = 7
      "0000111" when "01010010111101010", -- t[42474] = 7
      "0000111" when "01010010111101011", -- t[42475] = 7
      "0000111" when "01010010111101100", -- t[42476] = 7
      "0000111" when "01010010111101101", -- t[42477] = 7
      "0000111" when "01010010111101110", -- t[42478] = 7
      "0000111" when "01010010111101111", -- t[42479] = 7
      "0000111" when "01010010111110000", -- t[42480] = 7
      "0000111" when "01010010111110001", -- t[42481] = 7
      "0000111" when "01010010111110010", -- t[42482] = 7
      "0000111" when "01010010111110011", -- t[42483] = 7
      "0000111" when "01010010111110100", -- t[42484] = 7
      "0000111" when "01010010111110101", -- t[42485] = 7
      "0000111" when "01010010111110110", -- t[42486] = 7
      "0000111" when "01010010111110111", -- t[42487] = 7
      "0000111" when "01010010111111000", -- t[42488] = 7
      "0000111" when "01010010111111001", -- t[42489] = 7
      "0000111" when "01010010111111010", -- t[42490] = 7
      "0000111" when "01010010111111011", -- t[42491] = 7
      "0000111" when "01010010111111100", -- t[42492] = 7
      "0000111" when "01010010111111101", -- t[42493] = 7
      "0000111" when "01010010111111110", -- t[42494] = 7
      "0000111" when "01010010111111111", -- t[42495] = 7
      "0000111" when "01010011000000000", -- t[42496] = 7
      "0000111" when "01010011000000001", -- t[42497] = 7
      "0000111" when "01010011000000010", -- t[42498] = 7
      "0000111" when "01010011000000011", -- t[42499] = 7
      "0000111" when "01010011000000100", -- t[42500] = 7
      "0000111" when "01010011000000101", -- t[42501] = 7
      "0000111" when "01010011000000110", -- t[42502] = 7
      "0000111" when "01010011000000111", -- t[42503] = 7
      "0000111" when "01010011000001000", -- t[42504] = 7
      "0000111" when "01010011000001001", -- t[42505] = 7
      "0000111" when "01010011000001010", -- t[42506] = 7
      "0000111" when "01010011000001011", -- t[42507] = 7
      "0000111" when "01010011000001100", -- t[42508] = 7
      "0000111" when "01010011000001101", -- t[42509] = 7
      "0000111" when "01010011000001110", -- t[42510] = 7
      "0000111" when "01010011000001111", -- t[42511] = 7
      "0000111" when "01010011000010000", -- t[42512] = 7
      "0000111" when "01010011000010001", -- t[42513] = 7
      "0000111" when "01010011000010010", -- t[42514] = 7
      "0000111" when "01010011000010011", -- t[42515] = 7
      "0000111" when "01010011000010100", -- t[42516] = 7
      "0000111" when "01010011000010101", -- t[42517] = 7
      "0000111" when "01010011000010110", -- t[42518] = 7
      "0000111" when "01010011000010111", -- t[42519] = 7
      "0000111" when "01010011000011000", -- t[42520] = 7
      "0000111" when "01010011000011001", -- t[42521] = 7
      "0000111" when "01010011000011010", -- t[42522] = 7
      "0000111" when "01010011000011011", -- t[42523] = 7
      "0000111" when "01010011000011100", -- t[42524] = 7
      "0000111" when "01010011000011101", -- t[42525] = 7
      "0000111" when "01010011000011110", -- t[42526] = 7
      "0000111" when "01010011000011111", -- t[42527] = 7
      "0000111" when "01010011000100000", -- t[42528] = 7
      "0000111" when "01010011000100001", -- t[42529] = 7
      "0000111" when "01010011000100010", -- t[42530] = 7
      "0000111" when "01010011000100011", -- t[42531] = 7
      "0000111" when "01010011000100100", -- t[42532] = 7
      "0000111" when "01010011000100101", -- t[42533] = 7
      "0000111" when "01010011000100110", -- t[42534] = 7
      "0000111" when "01010011000100111", -- t[42535] = 7
      "0000111" when "01010011000101000", -- t[42536] = 7
      "0000111" when "01010011000101001", -- t[42537] = 7
      "0000111" when "01010011000101010", -- t[42538] = 7
      "0000111" when "01010011000101011", -- t[42539] = 7
      "0000111" when "01010011000101100", -- t[42540] = 7
      "0000111" when "01010011000101101", -- t[42541] = 7
      "0000111" when "01010011000101110", -- t[42542] = 7
      "0000111" when "01010011000101111", -- t[42543] = 7
      "0000111" when "01010011000110000", -- t[42544] = 7
      "0000111" when "01010011000110001", -- t[42545] = 7
      "0000111" when "01010011000110010", -- t[42546] = 7
      "0000111" when "01010011000110011", -- t[42547] = 7
      "0000111" when "01010011000110100", -- t[42548] = 7
      "0000111" when "01010011000110101", -- t[42549] = 7
      "0000111" when "01010011000110110", -- t[42550] = 7
      "0000111" when "01010011000110111", -- t[42551] = 7
      "0000111" when "01010011000111000", -- t[42552] = 7
      "0000111" when "01010011000111001", -- t[42553] = 7
      "0000111" when "01010011000111010", -- t[42554] = 7
      "0000111" when "01010011000111011", -- t[42555] = 7
      "0000111" when "01010011000111100", -- t[42556] = 7
      "0000111" when "01010011000111101", -- t[42557] = 7
      "0000111" when "01010011000111110", -- t[42558] = 7
      "0000111" when "01010011000111111", -- t[42559] = 7
      "0000111" when "01010011001000000", -- t[42560] = 7
      "0000111" when "01010011001000001", -- t[42561] = 7
      "0000111" when "01010011001000010", -- t[42562] = 7
      "0000111" when "01010011001000011", -- t[42563] = 7
      "0000111" when "01010011001000100", -- t[42564] = 7
      "0000111" when "01010011001000101", -- t[42565] = 7
      "0000111" when "01010011001000110", -- t[42566] = 7
      "0000111" when "01010011001000111", -- t[42567] = 7
      "0000111" when "01010011001001000", -- t[42568] = 7
      "0000111" when "01010011001001001", -- t[42569] = 7
      "0000111" when "01010011001001010", -- t[42570] = 7
      "0000111" when "01010011001001011", -- t[42571] = 7
      "0000111" when "01010011001001100", -- t[42572] = 7
      "0000111" when "01010011001001101", -- t[42573] = 7
      "0000111" when "01010011001001110", -- t[42574] = 7
      "0000111" when "01010011001001111", -- t[42575] = 7
      "0000111" when "01010011001010000", -- t[42576] = 7
      "0000111" when "01010011001010001", -- t[42577] = 7
      "0000111" when "01010011001010010", -- t[42578] = 7
      "0000111" when "01010011001010011", -- t[42579] = 7
      "0000111" when "01010011001010100", -- t[42580] = 7
      "0000111" when "01010011001010101", -- t[42581] = 7
      "0000111" when "01010011001010110", -- t[42582] = 7
      "0000111" when "01010011001010111", -- t[42583] = 7
      "0000111" when "01010011001011000", -- t[42584] = 7
      "0000111" when "01010011001011001", -- t[42585] = 7
      "0000111" when "01010011001011010", -- t[42586] = 7
      "0000111" when "01010011001011011", -- t[42587] = 7
      "0000111" when "01010011001011100", -- t[42588] = 7
      "0000111" when "01010011001011101", -- t[42589] = 7
      "0000111" when "01010011001011110", -- t[42590] = 7
      "0000111" when "01010011001011111", -- t[42591] = 7
      "0000111" when "01010011001100000", -- t[42592] = 7
      "0000111" when "01010011001100001", -- t[42593] = 7
      "0000111" when "01010011001100010", -- t[42594] = 7
      "0000111" when "01010011001100011", -- t[42595] = 7
      "0000111" when "01010011001100100", -- t[42596] = 7
      "0000111" when "01010011001100101", -- t[42597] = 7
      "0000111" when "01010011001100110", -- t[42598] = 7
      "0000111" when "01010011001100111", -- t[42599] = 7
      "0000111" when "01010011001101000", -- t[42600] = 7
      "0000111" when "01010011001101001", -- t[42601] = 7
      "0000111" when "01010011001101010", -- t[42602] = 7
      "0000111" when "01010011001101011", -- t[42603] = 7
      "0000111" when "01010011001101100", -- t[42604] = 7
      "0000111" when "01010011001101101", -- t[42605] = 7
      "0000111" when "01010011001101110", -- t[42606] = 7
      "0000111" when "01010011001101111", -- t[42607] = 7
      "0000111" when "01010011001110000", -- t[42608] = 7
      "0000111" when "01010011001110001", -- t[42609] = 7
      "0000111" when "01010011001110010", -- t[42610] = 7
      "0000111" when "01010011001110011", -- t[42611] = 7
      "0000111" when "01010011001110100", -- t[42612] = 7
      "0000111" when "01010011001110101", -- t[42613] = 7
      "0000111" when "01010011001110110", -- t[42614] = 7
      "0000111" when "01010011001110111", -- t[42615] = 7
      "0000111" when "01010011001111000", -- t[42616] = 7
      "0000111" when "01010011001111001", -- t[42617] = 7
      "0000111" when "01010011001111010", -- t[42618] = 7
      "0000111" when "01010011001111011", -- t[42619] = 7
      "0000111" when "01010011001111100", -- t[42620] = 7
      "0000111" when "01010011001111101", -- t[42621] = 7
      "0000111" when "01010011001111110", -- t[42622] = 7
      "0000111" when "01010011001111111", -- t[42623] = 7
      "0000111" when "01010011010000000", -- t[42624] = 7
      "0000111" when "01010011010000001", -- t[42625] = 7
      "0000111" when "01010011010000010", -- t[42626] = 7
      "0000111" when "01010011010000011", -- t[42627] = 7
      "0000111" when "01010011010000100", -- t[42628] = 7
      "0000111" when "01010011010000101", -- t[42629] = 7
      "0000111" when "01010011010000110", -- t[42630] = 7
      "0000111" when "01010011010000111", -- t[42631] = 7
      "0000111" when "01010011010001000", -- t[42632] = 7
      "0000111" when "01010011010001001", -- t[42633] = 7
      "0000111" when "01010011010001010", -- t[42634] = 7
      "0000111" when "01010011010001011", -- t[42635] = 7
      "0000111" when "01010011010001100", -- t[42636] = 7
      "0000111" when "01010011010001101", -- t[42637] = 7
      "0000111" when "01010011010001110", -- t[42638] = 7
      "0000111" when "01010011010001111", -- t[42639] = 7
      "0000111" when "01010011010010000", -- t[42640] = 7
      "0000111" when "01010011010010001", -- t[42641] = 7
      "0000111" when "01010011010010010", -- t[42642] = 7
      "0000111" when "01010011010010011", -- t[42643] = 7
      "0000111" when "01010011010010100", -- t[42644] = 7
      "0000111" when "01010011010010101", -- t[42645] = 7
      "0000111" when "01010011010010110", -- t[42646] = 7
      "0000111" when "01010011010010111", -- t[42647] = 7
      "0000111" when "01010011010011000", -- t[42648] = 7
      "0000111" when "01010011010011001", -- t[42649] = 7
      "0000111" when "01010011010011010", -- t[42650] = 7
      "0000111" when "01010011010011011", -- t[42651] = 7
      "0000111" when "01010011010011100", -- t[42652] = 7
      "0000111" when "01010011010011101", -- t[42653] = 7
      "0000111" when "01010011010011110", -- t[42654] = 7
      "0000111" when "01010011010011111", -- t[42655] = 7
      "0000111" when "01010011010100000", -- t[42656] = 7
      "0000111" when "01010011010100001", -- t[42657] = 7
      "0000111" when "01010011010100010", -- t[42658] = 7
      "0000111" when "01010011010100011", -- t[42659] = 7
      "0000111" when "01010011010100100", -- t[42660] = 7
      "0000111" when "01010011010100101", -- t[42661] = 7
      "0000111" when "01010011010100110", -- t[42662] = 7
      "0000111" when "01010011010100111", -- t[42663] = 7
      "0000111" when "01010011010101000", -- t[42664] = 7
      "0000111" when "01010011010101001", -- t[42665] = 7
      "0000111" when "01010011010101010", -- t[42666] = 7
      "0000111" when "01010011010101011", -- t[42667] = 7
      "0000111" when "01010011010101100", -- t[42668] = 7
      "0000111" when "01010011010101101", -- t[42669] = 7
      "0000111" when "01010011010101110", -- t[42670] = 7
      "0000111" when "01010011010101111", -- t[42671] = 7
      "0000111" when "01010011010110000", -- t[42672] = 7
      "0000111" when "01010011010110001", -- t[42673] = 7
      "0000111" when "01010011010110010", -- t[42674] = 7
      "0000111" when "01010011010110011", -- t[42675] = 7
      "0000111" when "01010011010110100", -- t[42676] = 7
      "0000111" when "01010011010110101", -- t[42677] = 7
      "0000111" when "01010011010110110", -- t[42678] = 7
      "0000111" when "01010011010110111", -- t[42679] = 7
      "0000111" when "01010011010111000", -- t[42680] = 7
      "0000111" when "01010011010111001", -- t[42681] = 7
      "0000111" when "01010011010111010", -- t[42682] = 7
      "0000111" when "01010011010111011", -- t[42683] = 7
      "0000111" when "01010011010111100", -- t[42684] = 7
      "0000111" when "01010011010111101", -- t[42685] = 7
      "0000111" when "01010011010111110", -- t[42686] = 7
      "0000111" when "01010011010111111", -- t[42687] = 7
      "0000111" when "01010011011000000", -- t[42688] = 7
      "0000111" when "01010011011000001", -- t[42689] = 7
      "0000111" when "01010011011000010", -- t[42690] = 7
      "0000111" when "01010011011000011", -- t[42691] = 7
      "0000111" when "01010011011000100", -- t[42692] = 7
      "0000111" when "01010011011000101", -- t[42693] = 7
      "0000111" when "01010011011000110", -- t[42694] = 7
      "0000111" when "01010011011000111", -- t[42695] = 7
      "0000111" when "01010011011001000", -- t[42696] = 7
      "0000111" when "01010011011001001", -- t[42697] = 7
      "0000111" when "01010011011001010", -- t[42698] = 7
      "0000111" when "01010011011001011", -- t[42699] = 7
      "0000111" when "01010011011001100", -- t[42700] = 7
      "0000111" when "01010011011001101", -- t[42701] = 7
      "0000111" when "01010011011001110", -- t[42702] = 7
      "0000111" when "01010011011001111", -- t[42703] = 7
      "0000111" when "01010011011010000", -- t[42704] = 7
      "0000111" when "01010011011010001", -- t[42705] = 7
      "0000111" when "01010011011010010", -- t[42706] = 7
      "0000111" when "01010011011010011", -- t[42707] = 7
      "0000111" when "01010011011010100", -- t[42708] = 7
      "0000111" when "01010011011010101", -- t[42709] = 7
      "0000111" when "01010011011010110", -- t[42710] = 7
      "0000111" when "01010011011010111", -- t[42711] = 7
      "0000111" when "01010011011011000", -- t[42712] = 7
      "0000111" when "01010011011011001", -- t[42713] = 7
      "0000111" when "01010011011011010", -- t[42714] = 7
      "0000111" when "01010011011011011", -- t[42715] = 7
      "0000111" when "01010011011011100", -- t[42716] = 7
      "0000111" when "01010011011011101", -- t[42717] = 7
      "0000111" when "01010011011011110", -- t[42718] = 7
      "0000111" when "01010011011011111", -- t[42719] = 7
      "0000111" when "01010011011100000", -- t[42720] = 7
      "0000111" when "01010011011100001", -- t[42721] = 7
      "0000111" when "01010011011100010", -- t[42722] = 7
      "0000111" when "01010011011100011", -- t[42723] = 7
      "0000111" when "01010011011100100", -- t[42724] = 7
      "0000111" when "01010011011100101", -- t[42725] = 7
      "0000111" when "01010011011100110", -- t[42726] = 7
      "0000111" when "01010011011100111", -- t[42727] = 7
      "0000111" when "01010011011101000", -- t[42728] = 7
      "0000111" when "01010011011101001", -- t[42729] = 7
      "0000111" when "01010011011101010", -- t[42730] = 7
      "0000111" when "01010011011101011", -- t[42731] = 7
      "0000111" when "01010011011101100", -- t[42732] = 7
      "0000111" when "01010011011101101", -- t[42733] = 7
      "0000111" when "01010011011101110", -- t[42734] = 7
      "0000111" when "01010011011101111", -- t[42735] = 7
      "0000111" when "01010011011110000", -- t[42736] = 7
      "0000111" when "01010011011110001", -- t[42737] = 7
      "0000111" when "01010011011110010", -- t[42738] = 7
      "0000111" when "01010011011110011", -- t[42739] = 7
      "0000111" when "01010011011110100", -- t[42740] = 7
      "0000111" when "01010011011110101", -- t[42741] = 7
      "0000111" when "01010011011110110", -- t[42742] = 7
      "0000111" when "01010011011110111", -- t[42743] = 7
      "0000111" when "01010011011111000", -- t[42744] = 7
      "0000111" when "01010011011111001", -- t[42745] = 7
      "0000111" when "01010011011111010", -- t[42746] = 7
      "0000111" when "01010011011111011", -- t[42747] = 7
      "0000111" when "01010011011111100", -- t[42748] = 7
      "0000111" when "01010011011111101", -- t[42749] = 7
      "0000111" when "01010011011111110", -- t[42750] = 7
      "0000111" when "01010011011111111", -- t[42751] = 7
      "0000111" when "01010011100000000", -- t[42752] = 7
      "0000111" when "01010011100000001", -- t[42753] = 7
      "0000111" when "01010011100000010", -- t[42754] = 7
      "0000111" when "01010011100000011", -- t[42755] = 7
      "0000111" when "01010011100000100", -- t[42756] = 7
      "0000111" when "01010011100000101", -- t[42757] = 7
      "0000111" when "01010011100000110", -- t[42758] = 7
      "0000111" when "01010011100000111", -- t[42759] = 7
      "0000111" when "01010011100001000", -- t[42760] = 7
      "0000111" when "01010011100001001", -- t[42761] = 7
      "0000111" when "01010011100001010", -- t[42762] = 7
      "0000111" when "01010011100001011", -- t[42763] = 7
      "0000111" when "01010011100001100", -- t[42764] = 7
      "0000111" when "01010011100001101", -- t[42765] = 7
      "0000111" when "01010011100001110", -- t[42766] = 7
      "0000111" when "01010011100001111", -- t[42767] = 7
      "0000111" when "01010011100010000", -- t[42768] = 7
      "0000111" when "01010011100010001", -- t[42769] = 7
      "0000111" when "01010011100010010", -- t[42770] = 7
      "0000111" when "01010011100010011", -- t[42771] = 7
      "0000111" when "01010011100010100", -- t[42772] = 7
      "0000111" when "01010011100010101", -- t[42773] = 7
      "0000111" when "01010011100010110", -- t[42774] = 7
      "0000111" when "01010011100010111", -- t[42775] = 7
      "0000111" when "01010011100011000", -- t[42776] = 7
      "0000111" when "01010011100011001", -- t[42777] = 7
      "0000111" when "01010011100011010", -- t[42778] = 7
      "0000111" when "01010011100011011", -- t[42779] = 7
      "0000111" when "01010011100011100", -- t[42780] = 7
      "0000111" when "01010011100011101", -- t[42781] = 7
      "0000111" when "01010011100011110", -- t[42782] = 7
      "0000111" when "01010011100011111", -- t[42783] = 7
      "0000111" when "01010011100100000", -- t[42784] = 7
      "0000111" when "01010011100100001", -- t[42785] = 7
      "0000111" when "01010011100100010", -- t[42786] = 7
      "0000111" when "01010011100100011", -- t[42787] = 7
      "0000111" when "01010011100100100", -- t[42788] = 7
      "0000111" when "01010011100100101", -- t[42789] = 7
      "0000111" when "01010011100100110", -- t[42790] = 7
      "0000111" when "01010011100100111", -- t[42791] = 7
      "0000111" when "01010011100101000", -- t[42792] = 7
      "0000111" when "01010011100101001", -- t[42793] = 7
      "0000111" when "01010011100101010", -- t[42794] = 7
      "0000111" when "01010011100101011", -- t[42795] = 7
      "0000111" when "01010011100101100", -- t[42796] = 7
      "0000111" when "01010011100101101", -- t[42797] = 7
      "0000111" when "01010011100101110", -- t[42798] = 7
      "0000111" when "01010011100101111", -- t[42799] = 7
      "0000111" when "01010011100110000", -- t[42800] = 7
      "0000111" when "01010011100110001", -- t[42801] = 7
      "0000111" when "01010011100110010", -- t[42802] = 7
      "0000111" when "01010011100110011", -- t[42803] = 7
      "0000111" when "01010011100110100", -- t[42804] = 7
      "0000111" when "01010011100110101", -- t[42805] = 7
      "0000111" when "01010011100110110", -- t[42806] = 7
      "0000111" when "01010011100110111", -- t[42807] = 7
      "0000111" when "01010011100111000", -- t[42808] = 7
      "0000111" when "01010011100111001", -- t[42809] = 7
      "0000111" when "01010011100111010", -- t[42810] = 7
      "0000111" when "01010011100111011", -- t[42811] = 7
      "0000111" when "01010011100111100", -- t[42812] = 7
      "0000111" when "01010011100111101", -- t[42813] = 7
      "0000111" when "01010011100111110", -- t[42814] = 7
      "0000111" when "01010011100111111", -- t[42815] = 7
      "0000111" when "01010011101000000", -- t[42816] = 7
      "0000111" when "01010011101000001", -- t[42817] = 7
      "0000111" when "01010011101000010", -- t[42818] = 7
      "0000111" when "01010011101000011", -- t[42819] = 7
      "0000111" when "01010011101000100", -- t[42820] = 7
      "0000111" when "01010011101000101", -- t[42821] = 7
      "0000111" when "01010011101000110", -- t[42822] = 7
      "0000111" when "01010011101000111", -- t[42823] = 7
      "0000111" when "01010011101001000", -- t[42824] = 7
      "0000111" when "01010011101001001", -- t[42825] = 7
      "0000111" when "01010011101001010", -- t[42826] = 7
      "0000111" when "01010011101001011", -- t[42827] = 7
      "0000111" when "01010011101001100", -- t[42828] = 7
      "0000111" when "01010011101001101", -- t[42829] = 7
      "0000111" when "01010011101001110", -- t[42830] = 7
      "0000111" when "01010011101001111", -- t[42831] = 7
      "0000111" when "01010011101010000", -- t[42832] = 7
      "0000111" when "01010011101010001", -- t[42833] = 7
      "0000111" when "01010011101010010", -- t[42834] = 7
      "0000111" when "01010011101010011", -- t[42835] = 7
      "0000111" when "01010011101010100", -- t[42836] = 7
      "0000111" when "01010011101010101", -- t[42837] = 7
      "0000111" when "01010011101010110", -- t[42838] = 7
      "0000111" when "01010011101010111", -- t[42839] = 7
      "0000111" when "01010011101011000", -- t[42840] = 7
      "0000111" when "01010011101011001", -- t[42841] = 7
      "0000111" when "01010011101011010", -- t[42842] = 7
      "0000111" when "01010011101011011", -- t[42843] = 7
      "0000111" when "01010011101011100", -- t[42844] = 7
      "0000111" when "01010011101011101", -- t[42845] = 7
      "0000111" when "01010011101011110", -- t[42846] = 7
      "0000111" when "01010011101011111", -- t[42847] = 7
      "0000111" when "01010011101100000", -- t[42848] = 7
      "0000111" when "01010011101100001", -- t[42849] = 7
      "0000111" when "01010011101100010", -- t[42850] = 7
      "0000111" when "01010011101100011", -- t[42851] = 7
      "0000111" when "01010011101100100", -- t[42852] = 7
      "0000111" when "01010011101100101", -- t[42853] = 7
      "0000111" when "01010011101100110", -- t[42854] = 7
      "0000111" when "01010011101100111", -- t[42855] = 7
      "0000111" when "01010011101101000", -- t[42856] = 7
      "0000111" when "01010011101101001", -- t[42857] = 7
      "0000111" when "01010011101101010", -- t[42858] = 7
      "0000111" when "01010011101101011", -- t[42859] = 7
      "0000111" when "01010011101101100", -- t[42860] = 7
      "0000111" when "01010011101101101", -- t[42861] = 7
      "0000111" when "01010011101101110", -- t[42862] = 7
      "0000111" when "01010011101101111", -- t[42863] = 7
      "0000111" when "01010011101110000", -- t[42864] = 7
      "0000111" when "01010011101110001", -- t[42865] = 7
      "0000111" when "01010011101110010", -- t[42866] = 7
      "0000111" when "01010011101110011", -- t[42867] = 7
      "0000111" when "01010011101110100", -- t[42868] = 7
      "0000111" when "01010011101110101", -- t[42869] = 7
      "0000111" when "01010011101110110", -- t[42870] = 7
      "0000111" when "01010011101110111", -- t[42871] = 7
      "0000111" when "01010011101111000", -- t[42872] = 7
      "0000111" when "01010011101111001", -- t[42873] = 7
      "0000111" when "01010011101111010", -- t[42874] = 7
      "0000111" when "01010011101111011", -- t[42875] = 7
      "0000111" when "01010011101111100", -- t[42876] = 7
      "0000111" when "01010011101111101", -- t[42877] = 7
      "0000111" when "01010011101111110", -- t[42878] = 7
      "0000111" when "01010011101111111", -- t[42879] = 7
      "0000111" when "01010011110000000", -- t[42880] = 7
      "0000111" when "01010011110000001", -- t[42881] = 7
      "0000111" when "01010011110000010", -- t[42882] = 7
      "0000111" when "01010011110000011", -- t[42883] = 7
      "0000111" when "01010011110000100", -- t[42884] = 7
      "0000111" when "01010011110000101", -- t[42885] = 7
      "0000111" when "01010011110000110", -- t[42886] = 7
      "0000111" when "01010011110000111", -- t[42887] = 7
      "0000111" when "01010011110001000", -- t[42888] = 7
      "0000111" when "01010011110001001", -- t[42889] = 7
      "0000111" when "01010011110001010", -- t[42890] = 7
      "0000111" when "01010011110001011", -- t[42891] = 7
      "0000111" when "01010011110001100", -- t[42892] = 7
      "0000111" when "01010011110001101", -- t[42893] = 7
      "0000111" when "01010011110001110", -- t[42894] = 7
      "0000111" when "01010011110001111", -- t[42895] = 7
      "0000111" when "01010011110010000", -- t[42896] = 7
      "0000111" when "01010011110010001", -- t[42897] = 7
      "0000111" when "01010011110010010", -- t[42898] = 7
      "0000111" when "01010011110010011", -- t[42899] = 7
      "0000111" when "01010011110010100", -- t[42900] = 7
      "0000111" when "01010011110010101", -- t[42901] = 7
      "0000111" when "01010011110010110", -- t[42902] = 7
      "0000111" when "01010011110010111", -- t[42903] = 7
      "0000111" when "01010011110011000", -- t[42904] = 7
      "0000111" when "01010011110011001", -- t[42905] = 7
      "0000111" when "01010011110011010", -- t[42906] = 7
      "0000111" when "01010011110011011", -- t[42907] = 7
      "0000111" when "01010011110011100", -- t[42908] = 7
      "0000111" when "01010011110011101", -- t[42909] = 7
      "0000111" when "01010011110011110", -- t[42910] = 7
      "0000111" when "01010011110011111", -- t[42911] = 7
      "0000111" when "01010011110100000", -- t[42912] = 7
      "0000111" when "01010011110100001", -- t[42913] = 7
      "0000111" when "01010011110100010", -- t[42914] = 7
      "0000111" when "01010011110100011", -- t[42915] = 7
      "0000111" when "01010011110100100", -- t[42916] = 7
      "0000111" when "01010011110100101", -- t[42917] = 7
      "0000111" when "01010011110100110", -- t[42918] = 7
      "0000111" when "01010011110100111", -- t[42919] = 7
      "0000111" when "01010011110101000", -- t[42920] = 7
      "0000111" when "01010011110101001", -- t[42921] = 7
      "0000111" when "01010011110101010", -- t[42922] = 7
      "0000111" when "01010011110101011", -- t[42923] = 7
      "0000111" when "01010011110101100", -- t[42924] = 7
      "0000111" when "01010011110101101", -- t[42925] = 7
      "0000111" when "01010011110101110", -- t[42926] = 7
      "0000111" when "01010011110101111", -- t[42927] = 7
      "0000111" when "01010011110110000", -- t[42928] = 7
      "0000111" when "01010011110110001", -- t[42929] = 7
      "0000111" when "01010011110110010", -- t[42930] = 7
      "0000111" when "01010011110110011", -- t[42931] = 7
      "0000111" when "01010011110110100", -- t[42932] = 7
      "0000111" when "01010011110110101", -- t[42933] = 7
      "0000111" when "01010011110110110", -- t[42934] = 7
      "0000111" when "01010011110110111", -- t[42935] = 7
      "0000111" when "01010011110111000", -- t[42936] = 7
      "0000111" when "01010011110111001", -- t[42937] = 7
      "0000111" when "01010011110111010", -- t[42938] = 7
      "0000111" when "01010011110111011", -- t[42939] = 7
      "0000111" when "01010011110111100", -- t[42940] = 7
      "0000111" when "01010011110111101", -- t[42941] = 7
      "0000111" when "01010011110111110", -- t[42942] = 7
      "0000111" when "01010011110111111", -- t[42943] = 7
      "0000111" when "01010011111000000", -- t[42944] = 7
      "0000111" when "01010011111000001", -- t[42945] = 7
      "0000111" when "01010011111000010", -- t[42946] = 7
      "0000111" when "01010011111000011", -- t[42947] = 7
      "0000111" when "01010011111000100", -- t[42948] = 7
      "0000111" when "01010011111000101", -- t[42949] = 7
      "0000111" when "01010011111000110", -- t[42950] = 7
      "0000111" when "01010011111000111", -- t[42951] = 7
      "0000111" when "01010011111001000", -- t[42952] = 7
      "0000111" when "01010011111001001", -- t[42953] = 7
      "0000111" when "01010011111001010", -- t[42954] = 7
      "0000111" when "01010011111001011", -- t[42955] = 7
      "0000111" when "01010011111001100", -- t[42956] = 7
      "0000111" when "01010011111001101", -- t[42957] = 7
      "0000111" when "01010011111001110", -- t[42958] = 7
      "0000111" when "01010011111001111", -- t[42959] = 7
      "0000111" when "01010011111010000", -- t[42960] = 7
      "0000111" when "01010011111010001", -- t[42961] = 7
      "0000111" when "01010011111010010", -- t[42962] = 7
      "0000111" when "01010011111010011", -- t[42963] = 7
      "0000111" when "01010011111010100", -- t[42964] = 7
      "0000111" when "01010011111010101", -- t[42965] = 7
      "0000111" when "01010011111010110", -- t[42966] = 7
      "0000111" when "01010011111010111", -- t[42967] = 7
      "0000111" when "01010011111011000", -- t[42968] = 7
      "0000111" when "01010011111011001", -- t[42969] = 7
      "0000111" when "01010011111011010", -- t[42970] = 7
      "0000111" when "01010011111011011", -- t[42971] = 7
      "0000111" when "01010011111011100", -- t[42972] = 7
      "0000111" when "01010011111011101", -- t[42973] = 7
      "0000111" when "01010011111011110", -- t[42974] = 7
      "0000111" when "01010011111011111", -- t[42975] = 7
      "0000111" when "01010011111100000", -- t[42976] = 7
      "0000111" when "01010011111100001", -- t[42977] = 7
      "0000111" when "01010011111100010", -- t[42978] = 7
      "0000111" when "01010011111100011", -- t[42979] = 7
      "0000111" when "01010011111100100", -- t[42980] = 7
      "0000111" when "01010011111100101", -- t[42981] = 7
      "0000111" when "01010011111100110", -- t[42982] = 7
      "0000111" when "01010011111100111", -- t[42983] = 7
      "0000111" when "01010011111101000", -- t[42984] = 7
      "0000111" when "01010011111101001", -- t[42985] = 7
      "0000111" when "01010011111101010", -- t[42986] = 7
      "0000111" when "01010011111101011", -- t[42987] = 7
      "0000111" when "01010011111101100", -- t[42988] = 7
      "0000111" when "01010011111101101", -- t[42989] = 7
      "0000111" when "01010011111101110", -- t[42990] = 7
      "0000111" when "01010011111101111", -- t[42991] = 7
      "0000111" when "01010011111110000", -- t[42992] = 7
      "0000111" when "01010011111110001", -- t[42993] = 7
      "0000111" when "01010011111110010", -- t[42994] = 7
      "0000111" when "01010011111110011", -- t[42995] = 7
      "0000111" when "01010011111110100", -- t[42996] = 7
      "0000111" when "01010011111110101", -- t[42997] = 7
      "0000111" when "01010011111110110", -- t[42998] = 7
      "0000111" when "01010011111110111", -- t[42999] = 7
      "0000111" when "01010011111111000", -- t[43000] = 7
      "0000111" when "01010011111111001", -- t[43001] = 7
      "0000111" when "01010011111111010", -- t[43002] = 7
      "0000111" when "01010011111111011", -- t[43003] = 7
      "0000111" when "01010011111111100", -- t[43004] = 7
      "0000111" when "01010011111111101", -- t[43005] = 7
      "0000111" when "01010011111111110", -- t[43006] = 7
      "0000111" when "01010011111111111", -- t[43007] = 7
      "0000111" when "01010100000000000", -- t[43008] = 7
      "0000111" when "01010100000000001", -- t[43009] = 7
      "0000111" when "01010100000000010", -- t[43010] = 7
      "0000111" when "01010100000000011", -- t[43011] = 7
      "0000111" when "01010100000000100", -- t[43012] = 7
      "0000111" when "01010100000000101", -- t[43013] = 7
      "0000111" when "01010100000000110", -- t[43014] = 7
      "0000111" when "01010100000000111", -- t[43015] = 7
      "0000111" when "01010100000001000", -- t[43016] = 7
      "0000111" when "01010100000001001", -- t[43017] = 7
      "0000111" when "01010100000001010", -- t[43018] = 7
      "0000111" when "01010100000001011", -- t[43019] = 7
      "0000111" when "01010100000001100", -- t[43020] = 7
      "0000111" when "01010100000001101", -- t[43021] = 7
      "0000111" when "01010100000001110", -- t[43022] = 7
      "0000111" when "01010100000001111", -- t[43023] = 7
      "0000111" when "01010100000010000", -- t[43024] = 7
      "0000111" when "01010100000010001", -- t[43025] = 7
      "0000111" when "01010100000010010", -- t[43026] = 7
      "0000111" when "01010100000010011", -- t[43027] = 7
      "0000111" when "01010100000010100", -- t[43028] = 7
      "0000111" when "01010100000010101", -- t[43029] = 7
      "0000111" when "01010100000010110", -- t[43030] = 7
      "0000111" when "01010100000010111", -- t[43031] = 7
      "0000111" when "01010100000011000", -- t[43032] = 7
      "0000111" when "01010100000011001", -- t[43033] = 7
      "0000111" when "01010100000011010", -- t[43034] = 7
      "0000111" when "01010100000011011", -- t[43035] = 7
      "0000111" when "01010100000011100", -- t[43036] = 7
      "0000111" when "01010100000011101", -- t[43037] = 7
      "0000111" when "01010100000011110", -- t[43038] = 7
      "0000111" when "01010100000011111", -- t[43039] = 7
      "0000111" when "01010100000100000", -- t[43040] = 7
      "0000111" when "01010100000100001", -- t[43041] = 7
      "0000111" when "01010100000100010", -- t[43042] = 7
      "0000111" when "01010100000100011", -- t[43043] = 7
      "0000111" when "01010100000100100", -- t[43044] = 7
      "0000111" when "01010100000100101", -- t[43045] = 7
      "0000111" when "01010100000100110", -- t[43046] = 7
      "0000111" when "01010100000100111", -- t[43047] = 7
      "0000111" when "01010100000101000", -- t[43048] = 7
      "0000111" when "01010100000101001", -- t[43049] = 7
      "0000111" when "01010100000101010", -- t[43050] = 7
      "0000111" when "01010100000101011", -- t[43051] = 7
      "0000111" when "01010100000101100", -- t[43052] = 7
      "0000111" when "01010100000101101", -- t[43053] = 7
      "0000111" when "01010100000101110", -- t[43054] = 7
      "0000111" when "01010100000101111", -- t[43055] = 7
      "0000111" when "01010100000110000", -- t[43056] = 7
      "0000111" when "01010100000110001", -- t[43057] = 7
      "0000111" when "01010100000110010", -- t[43058] = 7
      "0000111" when "01010100000110011", -- t[43059] = 7
      "0000111" when "01010100000110100", -- t[43060] = 7
      "0000111" when "01010100000110101", -- t[43061] = 7
      "0000111" when "01010100000110110", -- t[43062] = 7
      "0000111" when "01010100000110111", -- t[43063] = 7
      "0000111" when "01010100000111000", -- t[43064] = 7
      "0000111" when "01010100000111001", -- t[43065] = 7
      "0000111" when "01010100000111010", -- t[43066] = 7
      "0000111" when "01010100000111011", -- t[43067] = 7
      "0000111" when "01010100000111100", -- t[43068] = 7
      "0000111" when "01010100000111101", -- t[43069] = 7
      "0000111" when "01010100000111110", -- t[43070] = 7
      "0000111" when "01010100000111111", -- t[43071] = 7
      "0000111" when "01010100001000000", -- t[43072] = 7
      "0000111" when "01010100001000001", -- t[43073] = 7
      "0000111" when "01010100001000010", -- t[43074] = 7
      "0000111" when "01010100001000011", -- t[43075] = 7
      "0000111" when "01010100001000100", -- t[43076] = 7
      "0000111" when "01010100001000101", -- t[43077] = 7
      "0000111" when "01010100001000110", -- t[43078] = 7
      "0000111" when "01010100001000111", -- t[43079] = 7
      "0000111" when "01010100001001000", -- t[43080] = 7
      "0000111" when "01010100001001001", -- t[43081] = 7
      "0000111" when "01010100001001010", -- t[43082] = 7
      "0000111" when "01010100001001011", -- t[43083] = 7
      "0000111" when "01010100001001100", -- t[43084] = 7
      "0000111" when "01010100001001101", -- t[43085] = 7
      "0000111" when "01010100001001110", -- t[43086] = 7
      "0000111" when "01010100001001111", -- t[43087] = 7
      "0000111" when "01010100001010000", -- t[43088] = 7
      "0000111" when "01010100001010001", -- t[43089] = 7
      "0000111" when "01010100001010010", -- t[43090] = 7
      "0000111" when "01010100001010011", -- t[43091] = 7
      "0000111" when "01010100001010100", -- t[43092] = 7
      "0000111" when "01010100001010101", -- t[43093] = 7
      "0000111" when "01010100001010110", -- t[43094] = 7
      "0000111" when "01010100001010111", -- t[43095] = 7
      "0000111" when "01010100001011000", -- t[43096] = 7
      "0000111" when "01010100001011001", -- t[43097] = 7
      "0000111" when "01010100001011010", -- t[43098] = 7
      "0000111" when "01010100001011011", -- t[43099] = 7
      "0000111" when "01010100001011100", -- t[43100] = 7
      "0000111" when "01010100001011101", -- t[43101] = 7
      "0000111" when "01010100001011110", -- t[43102] = 7
      "0000111" when "01010100001011111", -- t[43103] = 7
      "0000111" when "01010100001100000", -- t[43104] = 7
      "0000111" when "01010100001100001", -- t[43105] = 7
      "0000111" when "01010100001100010", -- t[43106] = 7
      "0000111" when "01010100001100011", -- t[43107] = 7
      "0000111" when "01010100001100100", -- t[43108] = 7
      "0000111" when "01010100001100101", -- t[43109] = 7
      "0000111" when "01010100001100110", -- t[43110] = 7
      "0000111" when "01010100001100111", -- t[43111] = 7
      "0000111" when "01010100001101000", -- t[43112] = 7
      "0000111" when "01010100001101001", -- t[43113] = 7
      "0000111" when "01010100001101010", -- t[43114] = 7
      "0000111" when "01010100001101011", -- t[43115] = 7
      "0000111" when "01010100001101100", -- t[43116] = 7
      "0000111" when "01010100001101101", -- t[43117] = 7
      "0000111" when "01010100001101110", -- t[43118] = 7
      "0000111" when "01010100001101111", -- t[43119] = 7
      "0000111" when "01010100001110000", -- t[43120] = 7
      "0000111" when "01010100001110001", -- t[43121] = 7
      "0000111" when "01010100001110010", -- t[43122] = 7
      "0000111" when "01010100001110011", -- t[43123] = 7
      "0000111" when "01010100001110100", -- t[43124] = 7
      "0000111" when "01010100001110101", -- t[43125] = 7
      "0000111" when "01010100001110110", -- t[43126] = 7
      "0000111" when "01010100001110111", -- t[43127] = 7
      "0000111" when "01010100001111000", -- t[43128] = 7
      "0000111" when "01010100001111001", -- t[43129] = 7
      "0000111" when "01010100001111010", -- t[43130] = 7
      "0000111" when "01010100001111011", -- t[43131] = 7
      "0000111" when "01010100001111100", -- t[43132] = 7
      "0000111" when "01010100001111101", -- t[43133] = 7
      "0000111" when "01010100001111110", -- t[43134] = 7
      "0000111" when "01010100001111111", -- t[43135] = 7
      "0000111" when "01010100010000000", -- t[43136] = 7
      "0000111" when "01010100010000001", -- t[43137] = 7
      "0000111" when "01010100010000010", -- t[43138] = 7
      "0000111" when "01010100010000011", -- t[43139] = 7
      "0000111" when "01010100010000100", -- t[43140] = 7
      "0000111" when "01010100010000101", -- t[43141] = 7
      "0000111" when "01010100010000110", -- t[43142] = 7
      "0000111" when "01010100010000111", -- t[43143] = 7
      "0000111" when "01010100010001000", -- t[43144] = 7
      "0000111" when "01010100010001001", -- t[43145] = 7
      "0000111" when "01010100010001010", -- t[43146] = 7
      "0000111" when "01010100010001011", -- t[43147] = 7
      "0000111" when "01010100010001100", -- t[43148] = 7
      "0000111" when "01010100010001101", -- t[43149] = 7
      "0000111" when "01010100010001110", -- t[43150] = 7
      "0000111" when "01010100010001111", -- t[43151] = 7
      "0000111" when "01010100010010000", -- t[43152] = 7
      "0000111" when "01010100010010001", -- t[43153] = 7
      "0000111" when "01010100010010010", -- t[43154] = 7
      "0000111" when "01010100010010011", -- t[43155] = 7
      "0000111" when "01010100010010100", -- t[43156] = 7
      "0000111" when "01010100010010101", -- t[43157] = 7
      "0000111" when "01010100010010110", -- t[43158] = 7
      "0000111" when "01010100010010111", -- t[43159] = 7
      "0000111" when "01010100010011000", -- t[43160] = 7
      "0000111" when "01010100010011001", -- t[43161] = 7
      "0000111" when "01010100010011010", -- t[43162] = 7
      "0000111" when "01010100010011011", -- t[43163] = 7
      "0000111" when "01010100010011100", -- t[43164] = 7
      "0000111" when "01010100010011101", -- t[43165] = 7
      "0000111" when "01010100010011110", -- t[43166] = 7
      "0000111" when "01010100010011111", -- t[43167] = 7
      "0000111" when "01010100010100000", -- t[43168] = 7
      "0000111" when "01010100010100001", -- t[43169] = 7
      "0000111" when "01010100010100010", -- t[43170] = 7
      "0000111" when "01010100010100011", -- t[43171] = 7
      "0000111" when "01010100010100100", -- t[43172] = 7
      "0000111" when "01010100010100101", -- t[43173] = 7
      "0000111" when "01010100010100110", -- t[43174] = 7
      "0000111" when "01010100010100111", -- t[43175] = 7
      "0000111" when "01010100010101000", -- t[43176] = 7
      "0000111" when "01010100010101001", -- t[43177] = 7
      "0000111" when "01010100010101010", -- t[43178] = 7
      "0000111" when "01010100010101011", -- t[43179] = 7
      "0000111" when "01010100010101100", -- t[43180] = 7
      "0000111" when "01010100010101101", -- t[43181] = 7
      "0000111" when "01010100010101110", -- t[43182] = 7
      "0000111" when "01010100010101111", -- t[43183] = 7
      "0000111" when "01010100010110000", -- t[43184] = 7
      "0000111" when "01010100010110001", -- t[43185] = 7
      "0000111" when "01010100010110010", -- t[43186] = 7
      "0000111" when "01010100010110011", -- t[43187] = 7
      "0000111" when "01010100010110100", -- t[43188] = 7
      "0000111" when "01010100010110101", -- t[43189] = 7
      "0000111" when "01010100010110110", -- t[43190] = 7
      "0000111" when "01010100010110111", -- t[43191] = 7
      "0000111" when "01010100010111000", -- t[43192] = 7
      "0000111" when "01010100010111001", -- t[43193] = 7
      "0000111" when "01010100010111010", -- t[43194] = 7
      "0000111" when "01010100010111011", -- t[43195] = 7
      "0000111" when "01010100010111100", -- t[43196] = 7
      "0000111" when "01010100010111101", -- t[43197] = 7
      "0000111" when "01010100010111110", -- t[43198] = 7
      "0000111" when "01010100010111111", -- t[43199] = 7
      "0000111" when "01010100011000000", -- t[43200] = 7
      "0000111" when "01010100011000001", -- t[43201] = 7
      "0000111" when "01010100011000010", -- t[43202] = 7
      "0000111" when "01010100011000011", -- t[43203] = 7
      "0000111" when "01010100011000100", -- t[43204] = 7
      "0000111" when "01010100011000101", -- t[43205] = 7
      "0000111" when "01010100011000110", -- t[43206] = 7
      "0000111" when "01010100011000111", -- t[43207] = 7
      "0000111" when "01010100011001000", -- t[43208] = 7
      "0000111" when "01010100011001001", -- t[43209] = 7
      "0000111" when "01010100011001010", -- t[43210] = 7
      "0000111" when "01010100011001011", -- t[43211] = 7
      "0000111" when "01010100011001100", -- t[43212] = 7
      "0000111" when "01010100011001101", -- t[43213] = 7
      "0000111" when "01010100011001110", -- t[43214] = 7
      "0000111" when "01010100011001111", -- t[43215] = 7
      "0000111" when "01010100011010000", -- t[43216] = 7
      "0000111" when "01010100011010001", -- t[43217] = 7
      "0000111" when "01010100011010010", -- t[43218] = 7
      "0000111" when "01010100011010011", -- t[43219] = 7
      "0000111" when "01010100011010100", -- t[43220] = 7
      "0000111" when "01010100011010101", -- t[43221] = 7
      "0000111" when "01010100011010110", -- t[43222] = 7
      "0000111" when "01010100011010111", -- t[43223] = 7
      "0000111" when "01010100011011000", -- t[43224] = 7
      "0000111" when "01010100011011001", -- t[43225] = 7
      "0000111" when "01010100011011010", -- t[43226] = 7
      "0000111" when "01010100011011011", -- t[43227] = 7
      "0000111" when "01010100011011100", -- t[43228] = 7
      "0000111" when "01010100011011101", -- t[43229] = 7
      "0000111" when "01010100011011110", -- t[43230] = 7
      "0000111" when "01010100011011111", -- t[43231] = 7
      "0000111" when "01010100011100000", -- t[43232] = 7
      "0000111" when "01010100011100001", -- t[43233] = 7
      "0000111" when "01010100011100010", -- t[43234] = 7
      "0000111" when "01010100011100011", -- t[43235] = 7
      "0000111" when "01010100011100100", -- t[43236] = 7
      "0000111" when "01010100011100101", -- t[43237] = 7
      "0000111" when "01010100011100110", -- t[43238] = 7
      "0000111" when "01010100011100111", -- t[43239] = 7
      "0000111" when "01010100011101000", -- t[43240] = 7
      "0000111" when "01010100011101001", -- t[43241] = 7
      "0000111" when "01010100011101010", -- t[43242] = 7
      "0000111" when "01010100011101011", -- t[43243] = 7
      "0000111" when "01010100011101100", -- t[43244] = 7
      "0000111" when "01010100011101101", -- t[43245] = 7
      "0000111" when "01010100011101110", -- t[43246] = 7
      "0000111" when "01010100011101111", -- t[43247] = 7
      "0000111" when "01010100011110000", -- t[43248] = 7
      "0000111" when "01010100011110001", -- t[43249] = 7
      "0000111" when "01010100011110010", -- t[43250] = 7
      "0000111" when "01010100011110011", -- t[43251] = 7
      "0000111" when "01010100011110100", -- t[43252] = 7
      "0000111" when "01010100011110101", -- t[43253] = 7
      "0000111" when "01010100011110110", -- t[43254] = 7
      "0000111" when "01010100011110111", -- t[43255] = 7
      "0000111" when "01010100011111000", -- t[43256] = 7
      "0000111" when "01010100011111001", -- t[43257] = 7
      "0000111" when "01010100011111010", -- t[43258] = 7
      "0000111" when "01010100011111011", -- t[43259] = 7
      "0000111" when "01010100011111100", -- t[43260] = 7
      "0000111" when "01010100011111101", -- t[43261] = 7
      "0000111" when "01010100011111110", -- t[43262] = 7
      "0000111" when "01010100011111111", -- t[43263] = 7
      "0000111" when "01010100100000000", -- t[43264] = 7
      "0000111" when "01010100100000001", -- t[43265] = 7
      "0000111" when "01010100100000010", -- t[43266] = 7
      "0000111" when "01010100100000011", -- t[43267] = 7
      "0000111" when "01010100100000100", -- t[43268] = 7
      "0000111" when "01010100100000101", -- t[43269] = 7
      "0000111" when "01010100100000110", -- t[43270] = 7
      "0000111" when "01010100100000111", -- t[43271] = 7
      "0000111" when "01010100100001000", -- t[43272] = 7
      "0000111" when "01010100100001001", -- t[43273] = 7
      "0000111" when "01010100100001010", -- t[43274] = 7
      "0000111" when "01010100100001011", -- t[43275] = 7
      "0000111" when "01010100100001100", -- t[43276] = 7
      "0000111" when "01010100100001101", -- t[43277] = 7
      "0000111" when "01010100100001110", -- t[43278] = 7
      "0000111" when "01010100100001111", -- t[43279] = 7
      "0000111" when "01010100100010000", -- t[43280] = 7
      "0000111" when "01010100100010001", -- t[43281] = 7
      "0000111" when "01010100100010010", -- t[43282] = 7
      "0000111" when "01010100100010011", -- t[43283] = 7
      "0000111" when "01010100100010100", -- t[43284] = 7
      "0000111" when "01010100100010101", -- t[43285] = 7
      "0000111" when "01010100100010110", -- t[43286] = 7
      "0000111" when "01010100100010111", -- t[43287] = 7
      "0000111" when "01010100100011000", -- t[43288] = 7
      "0000111" when "01010100100011001", -- t[43289] = 7
      "0000111" when "01010100100011010", -- t[43290] = 7
      "0000111" when "01010100100011011", -- t[43291] = 7
      "0000111" when "01010100100011100", -- t[43292] = 7
      "0000111" when "01010100100011101", -- t[43293] = 7
      "0000111" when "01010100100011110", -- t[43294] = 7
      "0000111" when "01010100100011111", -- t[43295] = 7
      "0000111" when "01010100100100000", -- t[43296] = 7
      "0000111" when "01010100100100001", -- t[43297] = 7
      "0000111" when "01010100100100010", -- t[43298] = 7
      "0000111" when "01010100100100011", -- t[43299] = 7
      "0000111" when "01010100100100100", -- t[43300] = 7
      "0000111" when "01010100100100101", -- t[43301] = 7
      "0000111" when "01010100100100110", -- t[43302] = 7
      "0000111" when "01010100100100111", -- t[43303] = 7
      "0000111" when "01010100100101000", -- t[43304] = 7
      "0000111" when "01010100100101001", -- t[43305] = 7
      "0000111" when "01010100100101010", -- t[43306] = 7
      "0000111" when "01010100100101011", -- t[43307] = 7
      "0000111" when "01010100100101100", -- t[43308] = 7
      "0000111" when "01010100100101101", -- t[43309] = 7
      "0000111" when "01010100100101110", -- t[43310] = 7
      "0000111" when "01010100100101111", -- t[43311] = 7
      "0000111" when "01010100100110000", -- t[43312] = 7
      "0000111" when "01010100100110001", -- t[43313] = 7
      "0000111" when "01010100100110010", -- t[43314] = 7
      "0000111" when "01010100100110011", -- t[43315] = 7
      "0000111" when "01010100100110100", -- t[43316] = 7
      "0000111" when "01010100100110101", -- t[43317] = 7
      "0000111" when "01010100100110110", -- t[43318] = 7
      "0000111" when "01010100100110111", -- t[43319] = 7
      "0000111" when "01010100100111000", -- t[43320] = 7
      "0000111" when "01010100100111001", -- t[43321] = 7
      "0000111" when "01010100100111010", -- t[43322] = 7
      "0000111" when "01010100100111011", -- t[43323] = 7
      "0000111" when "01010100100111100", -- t[43324] = 7
      "0000111" when "01010100100111101", -- t[43325] = 7
      "0000111" when "01010100100111110", -- t[43326] = 7
      "0000111" when "01010100100111111", -- t[43327] = 7
      "0000111" when "01010100101000000", -- t[43328] = 7
      "0000111" when "01010100101000001", -- t[43329] = 7
      "0000111" when "01010100101000010", -- t[43330] = 7
      "0000111" when "01010100101000011", -- t[43331] = 7
      "0000111" when "01010100101000100", -- t[43332] = 7
      "0000111" when "01010100101000101", -- t[43333] = 7
      "0000111" when "01010100101000110", -- t[43334] = 7
      "0000111" when "01010100101000111", -- t[43335] = 7
      "0000111" when "01010100101001000", -- t[43336] = 7
      "0000111" when "01010100101001001", -- t[43337] = 7
      "0000111" when "01010100101001010", -- t[43338] = 7
      "0000111" when "01010100101001011", -- t[43339] = 7
      "0000111" when "01010100101001100", -- t[43340] = 7
      "0000111" when "01010100101001101", -- t[43341] = 7
      "0000111" when "01010100101001110", -- t[43342] = 7
      "0000111" when "01010100101001111", -- t[43343] = 7
      "0000111" when "01010100101010000", -- t[43344] = 7
      "0000111" when "01010100101010001", -- t[43345] = 7
      "0000111" when "01010100101010010", -- t[43346] = 7
      "0000111" when "01010100101010011", -- t[43347] = 7
      "0000111" when "01010100101010100", -- t[43348] = 7
      "0000111" when "01010100101010101", -- t[43349] = 7
      "0000111" when "01010100101010110", -- t[43350] = 7
      "0000111" when "01010100101010111", -- t[43351] = 7
      "0000111" when "01010100101011000", -- t[43352] = 7
      "0000111" when "01010100101011001", -- t[43353] = 7
      "0000111" when "01010100101011010", -- t[43354] = 7
      "0000111" when "01010100101011011", -- t[43355] = 7
      "0000111" when "01010100101011100", -- t[43356] = 7
      "0000111" when "01010100101011101", -- t[43357] = 7
      "0000111" when "01010100101011110", -- t[43358] = 7
      "0000111" when "01010100101011111", -- t[43359] = 7
      "0000111" when "01010100101100000", -- t[43360] = 7
      "0000111" when "01010100101100001", -- t[43361] = 7
      "0000111" when "01010100101100010", -- t[43362] = 7
      "0000111" when "01010100101100011", -- t[43363] = 7
      "0000111" when "01010100101100100", -- t[43364] = 7
      "0000111" when "01010100101100101", -- t[43365] = 7
      "0000111" when "01010100101100110", -- t[43366] = 7
      "0000111" when "01010100101100111", -- t[43367] = 7
      "0000111" when "01010100101101000", -- t[43368] = 7
      "0000111" when "01010100101101001", -- t[43369] = 7
      "0000111" when "01010100101101010", -- t[43370] = 7
      "0000111" when "01010100101101011", -- t[43371] = 7
      "0000111" when "01010100101101100", -- t[43372] = 7
      "0000111" when "01010100101101101", -- t[43373] = 7
      "0000111" when "01010100101101110", -- t[43374] = 7
      "0000111" when "01010100101101111", -- t[43375] = 7
      "0000111" when "01010100101110000", -- t[43376] = 7
      "0000111" when "01010100101110001", -- t[43377] = 7
      "0000111" when "01010100101110010", -- t[43378] = 7
      "0000111" when "01010100101110011", -- t[43379] = 7
      "0000111" when "01010100101110100", -- t[43380] = 7
      "0000111" when "01010100101110101", -- t[43381] = 7
      "0000111" when "01010100101110110", -- t[43382] = 7
      "0000111" when "01010100101110111", -- t[43383] = 7
      "0000111" when "01010100101111000", -- t[43384] = 7
      "0000111" when "01010100101111001", -- t[43385] = 7
      "0000111" when "01010100101111010", -- t[43386] = 7
      "0000111" when "01010100101111011", -- t[43387] = 7
      "0000111" when "01010100101111100", -- t[43388] = 7
      "0000111" when "01010100101111101", -- t[43389] = 7
      "0000111" when "01010100101111110", -- t[43390] = 7
      "0000111" when "01010100101111111", -- t[43391] = 7
      "0000111" when "01010100110000000", -- t[43392] = 7
      "0000111" when "01010100110000001", -- t[43393] = 7
      "0000111" when "01010100110000010", -- t[43394] = 7
      "0000111" when "01010100110000011", -- t[43395] = 7
      "0000111" when "01010100110000100", -- t[43396] = 7
      "0000111" when "01010100110000101", -- t[43397] = 7
      "0000111" when "01010100110000110", -- t[43398] = 7
      "0000111" when "01010100110000111", -- t[43399] = 7
      "0000111" when "01010100110001000", -- t[43400] = 7
      "0000111" when "01010100110001001", -- t[43401] = 7
      "0000111" when "01010100110001010", -- t[43402] = 7
      "0000111" when "01010100110001011", -- t[43403] = 7
      "0000111" when "01010100110001100", -- t[43404] = 7
      "0000111" when "01010100110001101", -- t[43405] = 7
      "0000111" when "01010100110001110", -- t[43406] = 7
      "0000111" when "01010100110001111", -- t[43407] = 7
      "0000111" when "01010100110010000", -- t[43408] = 7
      "0000111" when "01010100110010001", -- t[43409] = 7
      "0000111" when "01010100110010010", -- t[43410] = 7
      "0000111" when "01010100110010011", -- t[43411] = 7
      "0000111" when "01010100110010100", -- t[43412] = 7
      "0000111" when "01010100110010101", -- t[43413] = 7
      "0000111" when "01010100110010110", -- t[43414] = 7
      "0000111" when "01010100110010111", -- t[43415] = 7
      "0000111" when "01010100110011000", -- t[43416] = 7
      "0000111" when "01010100110011001", -- t[43417] = 7
      "0000111" when "01010100110011010", -- t[43418] = 7
      "0000111" when "01010100110011011", -- t[43419] = 7
      "0000111" when "01010100110011100", -- t[43420] = 7
      "0000111" when "01010100110011101", -- t[43421] = 7
      "0000111" when "01010100110011110", -- t[43422] = 7
      "0000111" when "01010100110011111", -- t[43423] = 7
      "0000111" when "01010100110100000", -- t[43424] = 7
      "0000111" when "01010100110100001", -- t[43425] = 7
      "0000111" when "01010100110100010", -- t[43426] = 7
      "0000111" when "01010100110100011", -- t[43427] = 7
      "0000111" when "01010100110100100", -- t[43428] = 7
      "0000111" when "01010100110100101", -- t[43429] = 7
      "0000111" when "01010100110100110", -- t[43430] = 7
      "0000111" when "01010100110100111", -- t[43431] = 7
      "0000111" when "01010100110101000", -- t[43432] = 7
      "0000111" when "01010100110101001", -- t[43433] = 7
      "0000111" when "01010100110101010", -- t[43434] = 7
      "0000111" when "01010100110101011", -- t[43435] = 7
      "0000111" when "01010100110101100", -- t[43436] = 7
      "0000111" when "01010100110101101", -- t[43437] = 7
      "0000111" when "01010100110101110", -- t[43438] = 7
      "0000111" when "01010100110101111", -- t[43439] = 7
      "0000111" when "01010100110110000", -- t[43440] = 7
      "0000111" when "01010100110110001", -- t[43441] = 7
      "0000111" when "01010100110110010", -- t[43442] = 7
      "0000111" when "01010100110110011", -- t[43443] = 7
      "0000111" when "01010100110110100", -- t[43444] = 7
      "0000111" when "01010100110110101", -- t[43445] = 7
      "0000111" when "01010100110110110", -- t[43446] = 7
      "0000111" when "01010100110110111", -- t[43447] = 7
      "0000111" when "01010100110111000", -- t[43448] = 7
      "0000111" when "01010100110111001", -- t[43449] = 7
      "0000111" when "01010100110111010", -- t[43450] = 7
      "0000111" when "01010100110111011", -- t[43451] = 7
      "0000111" when "01010100110111100", -- t[43452] = 7
      "0000111" when "01010100110111101", -- t[43453] = 7
      "0000111" when "01010100110111110", -- t[43454] = 7
      "0000111" when "01010100110111111", -- t[43455] = 7
      "0000111" when "01010100111000000", -- t[43456] = 7
      "0000111" when "01010100111000001", -- t[43457] = 7
      "0000111" when "01010100111000010", -- t[43458] = 7
      "0000111" when "01010100111000011", -- t[43459] = 7
      "0000111" when "01010100111000100", -- t[43460] = 7
      "0000111" when "01010100111000101", -- t[43461] = 7
      "0000111" when "01010100111000110", -- t[43462] = 7
      "0000111" when "01010100111000111", -- t[43463] = 7
      "0000111" when "01010100111001000", -- t[43464] = 7
      "0000111" when "01010100111001001", -- t[43465] = 7
      "0000111" when "01010100111001010", -- t[43466] = 7
      "0000111" when "01010100111001011", -- t[43467] = 7
      "0000111" when "01010100111001100", -- t[43468] = 7
      "0000111" when "01010100111001101", -- t[43469] = 7
      "0000111" when "01010100111001110", -- t[43470] = 7
      "0000111" when "01010100111001111", -- t[43471] = 7
      "0000111" when "01010100111010000", -- t[43472] = 7
      "0000111" when "01010100111010001", -- t[43473] = 7
      "0000111" when "01010100111010010", -- t[43474] = 7
      "0000111" when "01010100111010011", -- t[43475] = 7
      "0000111" when "01010100111010100", -- t[43476] = 7
      "0000111" when "01010100111010101", -- t[43477] = 7
      "0000111" when "01010100111010110", -- t[43478] = 7
      "0000111" when "01010100111010111", -- t[43479] = 7
      "0000111" when "01010100111011000", -- t[43480] = 7
      "0000111" when "01010100111011001", -- t[43481] = 7
      "0000111" when "01010100111011010", -- t[43482] = 7
      "0000111" when "01010100111011011", -- t[43483] = 7
      "0000111" when "01010100111011100", -- t[43484] = 7
      "0000111" when "01010100111011101", -- t[43485] = 7
      "0000111" when "01010100111011110", -- t[43486] = 7
      "0000111" when "01010100111011111", -- t[43487] = 7
      "0000111" when "01010100111100000", -- t[43488] = 7
      "0000111" when "01010100111100001", -- t[43489] = 7
      "0000111" when "01010100111100010", -- t[43490] = 7
      "0000111" when "01010100111100011", -- t[43491] = 7
      "0000111" when "01010100111100100", -- t[43492] = 7
      "0000111" when "01010100111100101", -- t[43493] = 7
      "0000111" when "01010100111100110", -- t[43494] = 7
      "0000111" when "01010100111100111", -- t[43495] = 7
      "0000111" when "01010100111101000", -- t[43496] = 7
      "0000111" when "01010100111101001", -- t[43497] = 7
      "0000111" when "01010100111101010", -- t[43498] = 7
      "0000111" when "01010100111101011", -- t[43499] = 7
      "0000111" when "01010100111101100", -- t[43500] = 7
      "0000111" when "01010100111101101", -- t[43501] = 7
      "0000111" when "01010100111101110", -- t[43502] = 7
      "0000111" when "01010100111101111", -- t[43503] = 7
      "0000111" when "01010100111110000", -- t[43504] = 7
      "0000111" when "01010100111110001", -- t[43505] = 7
      "0000111" when "01010100111110010", -- t[43506] = 7
      "0000111" when "01010100111110011", -- t[43507] = 7
      "0000111" when "01010100111110100", -- t[43508] = 7
      "0000111" when "01010100111110101", -- t[43509] = 7
      "0000111" when "01010100111110110", -- t[43510] = 7
      "0000111" when "01010100111110111", -- t[43511] = 7
      "0000111" when "01010100111111000", -- t[43512] = 7
      "0000111" when "01010100111111001", -- t[43513] = 7
      "0000111" when "01010100111111010", -- t[43514] = 7
      "0000111" when "01010100111111011", -- t[43515] = 7
      "0000111" when "01010100111111100", -- t[43516] = 7
      "0000111" when "01010100111111101", -- t[43517] = 7
      "0000111" when "01010100111111110", -- t[43518] = 7
      "0000111" when "01010100111111111", -- t[43519] = 7
      "0000111" when "01010101000000000", -- t[43520] = 7
      "0000111" when "01010101000000001", -- t[43521] = 7
      "0000111" when "01010101000000010", -- t[43522] = 7
      "0000111" when "01010101000000011", -- t[43523] = 7
      "0000111" when "01010101000000100", -- t[43524] = 7
      "0000111" when "01010101000000101", -- t[43525] = 7
      "0000111" when "01010101000000110", -- t[43526] = 7
      "0000111" when "01010101000000111", -- t[43527] = 7
      "0000111" when "01010101000001000", -- t[43528] = 7
      "0000111" when "01010101000001001", -- t[43529] = 7
      "0000111" when "01010101000001010", -- t[43530] = 7
      "0000111" when "01010101000001011", -- t[43531] = 7
      "0000111" when "01010101000001100", -- t[43532] = 7
      "0000111" when "01010101000001101", -- t[43533] = 7
      "0000111" when "01010101000001110", -- t[43534] = 7
      "0000111" when "01010101000001111", -- t[43535] = 7
      "0000111" when "01010101000010000", -- t[43536] = 7
      "0000111" when "01010101000010001", -- t[43537] = 7
      "0000111" when "01010101000010010", -- t[43538] = 7
      "0000111" when "01010101000010011", -- t[43539] = 7
      "0000111" when "01010101000010100", -- t[43540] = 7
      "0000111" when "01010101000010101", -- t[43541] = 7
      "0000111" when "01010101000010110", -- t[43542] = 7
      "0000111" when "01010101000010111", -- t[43543] = 7
      "0000111" when "01010101000011000", -- t[43544] = 7
      "0000111" when "01010101000011001", -- t[43545] = 7
      "0000111" when "01010101000011010", -- t[43546] = 7
      "0000111" when "01010101000011011", -- t[43547] = 7
      "0000111" when "01010101000011100", -- t[43548] = 7
      "0000111" when "01010101000011101", -- t[43549] = 7
      "0000111" when "01010101000011110", -- t[43550] = 7
      "0000111" when "01010101000011111", -- t[43551] = 7
      "0000111" when "01010101000100000", -- t[43552] = 7
      "0000111" when "01010101000100001", -- t[43553] = 7
      "0000111" when "01010101000100010", -- t[43554] = 7
      "0000111" when "01010101000100011", -- t[43555] = 7
      "0000111" when "01010101000100100", -- t[43556] = 7
      "0000111" when "01010101000100101", -- t[43557] = 7
      "0000111" when "01010101000100110", -- t[43558] = 7
      "0000111" when "01010101000100111", -- t[43559] = 7
      "0000111" when "01010101000101000", -- t[43560] = 7
      "0000111" when "01010101000101001", -- t[43561] = 7
      "0000111" when "01010101000101010", -- t[43562] = 7
      "0000111" when "01010101000101011", -- t[43563] = 7
      "0000111" when "01010101000101100", -- t[43564] = 7
      "0000111" when "01010101000101101", -- t[43565] = 7
      "0000111" when "01010101000101110", -- t[43566] = 7
      "0000111" when "01010101000101111", -- t[43567] = 7
      "0000111" when "01010101000110000", -- t[43568] = 7
      "0000111" when "01010101000110001", -- t[43569] = 7
      "0000111" when "01010101000110010", -- t[43570] = 7
      "0000111" when "01010101000110011", -- t[43571] = 7
      "0000111" when "01010101000110100", -- t[43572] = 7
      "0000111" when "01010101000110101", -- t[43573] = 7
      "0000111" when "01010101000110110", -- t[43574] = 7
      "0000111" when "01010101000110111", -- t[43575] = 7
      "0000111" when "01010101000111000", -- t[43576] = 7
      "0000111" when "01010101000111001", -- t[43577] = 7
      "0000111" when "01010101000111010", -- t[43578] = 7
      "0000111" when "01010101000111011", -- t[43579] = 7
      "0000111" when "01010101000111100", -- t[43580] = 7
      "0000111" when "01010101000111101", -- t[43581] = 7
      "0000111" when "01010101000111110", -- t[43582] = 7
      "0000111" when "01010101000111111", -- t[43583] = 7
      "0000111" when "01010101001000000", -- t[43584] = 7
      "0000111" when "01010101001000001", -- t[43585] = 7
      "0000111" when "01010101001000010", -- t[43586] = 7
      "0000111" when "01010101001000011", -- t[43587] = 7
      "0000111" when "01010101001000100", -- t[43588] = 7
      "0000111" when "01010101001000101", -- t[43589] = 7
      "0000111" when "01010101001000110", -- t[43590] = 7
      "0000111" when "01010101001000111", -- t[43591] = 7
      "0000111" when "01010101001001000", -- t[43592] = 7
      "0000111" when "01010101001001001", -- t[43593] = 7
      "0000111" when "01010101001001010", -- t[43594] = 7
      "0000111" when "01010101001001011", -- t[43595] = 7
      "0000111" when "01010101001001100", -- t[43596] = 7
      "0000111" when "01010101001001101", -- t[43597] = 7
      "0000111" when "01010101001001110", -- t[43598] = 7
      "0000111" when "01010101001001111", -- t[43599] = 7
      "0000111" when "01010101001010000", -- t[43600] = 7
      "0000111" when "01010101001010001", -- t[43601] = 7
      "0000111" when "01010101001010010", -- t[43602] = 7
      "0000111" when "01010101001010011", -- t[43603] = 7
      "0000111" when "01010101001010100", -- t[43604] = 7
      "0000111" when "01010101001010101", -- t[43605] = 7
      "0000111" when "01010101001010110", -- t[43606] = 7
      "0000111" when "01010101001010111", -- t[43607] = 7
      "0000111" when "01010101001011000", -- t[43608] = 7
      "0000111" when "01010101001011001", -- t[43609] = 7
      "0000111" when "01010101001011010", -- t[43610] = 7
      "0000111" when "01010101001011011", -- t[43611] = 7
      "0000111" when "01010101001011100", -- t[43612] = 7
      "0000111" when "01010101001011101", -- t[43613] = 7
      "0000111" when "01010101001011110", -- t[43614] = 7
      "0000111" when "01010101001011111", -- t[43615] = 7
      "0000111" when "01010101001100000", -- t[43616] = 7
      "0000111" when "01010101001100001", -- t[43617] = 7
      "0000111" when "01010101001100010", -- t[43618] = 7
      "0000111" when "01010101001100011", -- t[43619] = 7
      "0000111" when "01010101001100100", -- t[43620] = 7
      "0000111" when "01010101001100101", -- t[43621] = 7
      "0000111" when "01010101001100110", -- t[43622] = 7
      "0000111" when "01010101001100111", -- t[43623] = 7
      "0000111" when "01010101001101000", -- t[43624] = 7
      "0000111" when "01010101001101001", -- t[43625] = 7
      "0000111" when "01010101001101010", -- t[43626] = 7
      "0000111" when "01010101001101011", -- t[43627] = 7
      "0000111" when "01010101001101100", -- t[43628] = 7
      "0000111" when "01010101001101101", -- t[43629] = 7
      "0000111" when "01010101001101110", -- t[43630] = 7
      "0000111" when "01010101001101111", -- t[43631] = 7
      "0000111" when "01010101001110000", -- t[43632] = 7
      "0000111" when "01010101001110001", -- t[43633] = 7
      "0000111" when "01010101001110010", -- t[43634] = 7
      "0000111" when "01010101001110011", -- t[43635] = 7
      "0000111" when "01010101001110100", -- t[43636] = 7
      "0000111" when "01010101001110101", -- t[43637] = 7
      "0000111" when "01010101001110110", -- t[43638] = 7
      "0000111" when "01010101001110111", -- t[43639] = 7
      "0000111" when "01010101001111000", -- t[43640] = 7
      "0000111" when "01010101001111001", -- t[43641] = 7
      "0000111" when "01010101001111010", -- t[43642] = 7
      "0000111" when "01010101001111011", -- t[43643] = 7
      "0000111" when "01010101001111100", -- t[43644] = 7
      "0000111" when "01010101001111101", -- t[43645] = 7
      "0000111" when "01010101001111110", -- t[43646] = 7
      "0000111" when "01010101001111111", -- t[43647] = 7
      "0000111" when "01010101010000000", -- t[43648] = 7
      "0000111" when "01010101010000001", -- t[43649] = 7
      "0000111" when "01010101010000010", -- t[43650] = 7
      "0000111" when "01010101010000011", -- t[43651] = 7
      "0000111" when "01010101010000100", -- t[43652] = 7
      "0000111" when "01010101010000101", -- t[43653] = 7
      "0000111" when "01010101010000110", -- t[43654] = 7
      "0000111" when "01010101010000111", -- t[43655] = 7
      "0000111" when "01010101010001000", -- t[43656] = 7
      "0000111" when "01010101010001001", -- t[43657] = 7
      "0000111" when "01010101010001010", -- t[43658] = 7
      "0000111" when "01010101010001011", -- t[43659] = 7
      "0000111" when "01010101010001100", -- t[43660] = 7
      "0000111" when "01010101010001101", -- t[43661] = 7
      "0000111" when "01010101010001110", -- t[43662] = 7
      "0000111" when "01010101010001111", -- t[43663] = 7
      "0000111" when "01010101010010000", -- t[43664] = 7
      "0000111" when "01010101010010001", -- t[43665] = 7
      "0000111" when "01010101010010010", -- t[43666] = 7
      "0000111" when "01010101010010011", -- t[43667] = 7
      "0000111" when "01010101010010100", -- t[43668] = 7
      "0000111" when "01010101010010101", -- t[43669] = 7
      "0000111" when "01010101010010110", -- t[43670] = 7
      "0000111" when "01010101010010111", -- t[43671] = 7
      "0000111" when "01010101010011000", -- t[43672] = 7
      "0000111" when "01010101010011001", -- t[43673] = 7
      "0000111" when "01010101010011010", -- t[43674] = 7
      "0000111" when "01010101010011011", -- t[43675] = 7
      "0000111" when "01010101010011100", -- t[43676] = 7
      "0000111" when "01010101010011101", -- t[43677] = 7
      "0000111" when "01010101010011110", -- t[43678] = 7
      "0000111" when "01010101010011111", -- t[43679] = 7
      "0000111" when "01010101010100000", -- t[43680] = 7
      "0000111" when "01010101010100001", -- t[43681] = 7
      "0000111" when "01010101010100010", -- t[43682] = 7
      "0000111" when "01010101010100011", -- t[43683] = 7
      "0000111" when "01010101010100100", -- t[43684] = 7
      "0000111" when "01010101010100101", -- t[43685] = 7
      "0000111" when "01010101010100110", -- t[43686] = 7
      "0000111" when "01010101010100111", -- t[43687] = 7
      "0000111" when "01010101010101000", -- t[43688] = 7
      "0000111" when "01010101010101001", -- t[43689] = 7
      "0000111" when "01010101010101010", -- t[43690] = 7
      "0000111" when "01010101010101011", -- t[43691] = 7
      "0000111" when "01010101010101100", -- t[43692] = 7
      "0000111" when "01010101010101101", -- t[43693] = 7
      "0000111" when "01010101010101110", -- t[43694] = 7
      "0000111" when "01010101010101111", -- t[43695] = 7
      "0000111" when "01010101010110000", -- t[43696] = 7
      "0000111" when "01010101010110001", -- t[43697] = 7
      "0000111" when "01010101010110010", -- t[43698] = 7
      "0000111" when "01010101010110011", -- t[43699] = 7
      "0000111" when "01010101010110100", -- t[43700] = 7
      "0000111" when "01010101010110101", -- t[43701] = 7
      "0000111" when "01010101010110110", -- t[43702] = 7
      "0000111" when "01010101010110111", -- t[43703] = 7
      "0000111" when "01010101010111000", -- t[43704] = 7
      "0000111" when "01010101010111001", -- t[43705] = 7
      "0000111" when "01010101010111010", -- t[43706] = 7
      "0000111" when "01010101010111011", -- t[43707] = 7
      "0000111" when "01010101010111100", -- t[43708] = 7
      "0000111" when "01010101010111101", -- t[43709] = 7
      "0000111" when "01010101010111110", -- t[43710] = 7
      "0000111" when "01010101010111111", -- t[43711] = 7
      "0000111" when "01010101011000000", -- t[43712] = 7
      "0000111" when "01010101011000001", -- t[43713] = 7
      "0000111" when "01010101011000010", -- t[43714] = 7
      "0000111" when "01010101011000011", -- t[43715] = 7
      "0000111" when "01010101011000100", -- t[43716] = 7
      "0000111" when "01010101011000101", -- t[43717] = 7
      "0000111" when "01010101011000110", -- t[43718] = 7
      "0000111" when "01010101011000111", -- t[43719] = 7
      "0000111" when "01010101011001000", -- t[43720] = 7
      "0000111" when "01010101011001001", -- t[43721] = 7
      "0000111" when "01010101011001010", -- t[43722] = 7
      "0000111" when "01010101011001011", -- t[43723] = 7
      "0000111" when "01010101011001100", -- t[43724] = 7
      "0000111" when "01010101011001101", -- t[43725] = 7
      "0000111" when "01010101011001110", -- t[43726] = 7
      "0000111" when "01010101011001111", -- t[43727] = 7
      "0000111" when "01010101011010000", -- t[43728] = 7
      "0000111" when "01010101011010001", -- t[43729] = 7
      "0000111" when "01010101011010010", -- t[43730] = 7
      "0000111" when "01010101011010011", -- t[43731] = 7
      "0000111" when "01010101011010100", -- t[43732] = 7
      "0000111" when "01010101011010101", -- t[43733] = 7
      "0000111" when "01010101011010110", -- t[43734] = 7
      "0000111" when "01010101011010111", -- t[43735] = 7
      "0000111" when "01010101011011000", -- t[43736] = 7
      "0000111" when "01010101011011001", -- t[43737] = 7
      "0000111" when "01010101011011010", -- t[43738] = 7
      "0000111" when "01010101011011011", -- t[43739] = 7
      "0000111" when "01010101011011100", -- t[43740] = 7
      "0000111" when "01010101011011101", -- t[43741] = 7
      "0000111" when "01010101011011110", -- t[43742] = 7
      "0000111" when "01010101011011111", -- t[43743] = 7
      "0000111" when "01010101011100000", -- t[43744] = 7
      "0000111" when "01010101011100001", -- t[43745] = 7
      "0000111" when "01010101011100010", -- t[43746] = 7
      "0000111" when "01010101011100011", -- t[43747] = 7
      "0000111" when "01010101011100100", -- t[43748] = 7
      "0000111" when "01010101011100101", -- t[43749] = 7
      "0000111" when "01010101011100110", -- t[43750] = 7
      "0000111" when "01010101011100111", -- t[43751] = 7
      "0000111" when "01010101011101000", -- t[43752] = 7
      "0000111" when "01010101011101001", -- t[43753] = 7
      "0000111" when "01010101011101010", -- t[43754] = 7
      "0000111" when "01010101011101011", -- t[43755] = 7
      "0000111" when "01010101011101100", -- t[43756] = 7
      "0000111" when "01010101011101101", -- t[43757] = 7
      "0000111" when "01010101011101110", -- t[43758] = 7
      "0000111" when "01010101011101111", -- t[43759] = 7
      "0000111" when "01010101011110000", -- t[43760] = 7
      "0000111" when "01010101011110001", -- t[43761] = 7
      "0000111" when "01010101011110010", -- t[43762] = 7
      "0000111" when "01010101011110011", -- t[43763] = 7
      "0000111" when "01010101011110100", -- t[43764] = 7
      "0000111" when "01010101011110101", -- t[43765] = 7
      "0000111" when "01010101011110110", -- t[43766] = 7
      "0000111" when "01010101011110111", -- t[43767] = 7
      "0000111" when "01010101011111000", -- t[43768] = 7
      "0000111" when "01010101011111001", -- t[43769] = 7
      "0000111" when "01010101011111010", -- t[43770] = 7
      "0000111" when "01010101011111011", -- t[43771] = 7
      "0000111" when "01010101011111100", -- t[43772] = 7
      "0000111" when "01010101011111101", -- t[43773] = 7
      "0000111" when "01010101011111110", -- t[43774] = 7
      "0000111" when "01010101011111111", -- t[43775] = 7
      "0000111" when "01010101100000000", -- t[43776] = 7
      "0000111" when "01010101100000001", -- t[43777] = 7
      "0000111" when "01010101100000010", -- t[43778] = 7
      "0000111" when "01010101100000011", -- t[43779] = 7
      "0000111" when "01010101100000100", -- t[43780] = 7
      "0000111" when "01010101100000101", -- t[43781] = 7
      "0000111" when "01010101100000110", -- t[43782] = 7
      "0000111" when "01010101100000111", -- t[43783] = 7
      "0000111" when "01010101100001000", -- t[43784] = 7
      "0000111" when "01010101100001001", -- t[43785] = 7
      "0000111" when "01010101100001010", -- t[43786] = 7
      "0000111" when "01010101100001011", -- t[43787] = 7
      "0000111" when "01010101100001100", -- t[43788] = 7
      "0000111" when "01010101100001101", -- t[43789] = 7
      "0000111" when "01010101100001110", -- t[43790] = 7
      "0000111" when "01010101100001111", -- t[43791] = 7
      "0000111" when "01010101100010000", -- t[43792] = 7
      "0000111" when "01010101100010001", -- t[43793] = 7
      "0000111" when "01010101100010010", -- t[43794] = 7
      "0000111" when "01010101100010011", -- t[43795] = 7
      "0000111" when "01010101100010100", -- t[43796] = 7
      "0000111" when "01010101100010101", -- t[43797] = 7
      "0000111" when "01010101100010110", -- t[43798] = 7
      "0000111" when "01010101100010111", -- t[43799] = 7
      "0000111" when "01010101100011000", -- t[43800] = 7
      "0000111" when "01010101100011001", -- t[43801] = 7
      "0000111" when "01010101100011010", -- t[43802] = 7
      "0000111" when "01010101100011011", -- t[43803] = 7
      "0000111" when "01010101100011100", -- t[43804] = 7
      "0000111" when "01010101100011101", -- t[43805] = 7
      "0000111" when "01010101100011110", -- t[43806] = 7
      "0000111" when "01010101100011111", -- t[43807] = 7
      "0000111" when "01010101100100000", -- t[43808] = 7
      "0000111" when "01010101100100001", -- t[43809] = 7
      "0000111" when "01010101100100010", -- t[43810] = 7
      "0000111" when "01010101100100011", -- t[43811] = 7
      "0000111" when "01010101100100100", -- t[43812] = 7
      "0000111" when "01010101100100101", -- t[43813] = 7
      "0000111" when "01010101100100110", -- t[43814] = 7
      "0000111" when "01010101100100111", -- t[43815] = 7
      "0000111" when "01010101100101000", -- t[43816] = 7
      "0000111" when "01010101100101001", -- t[43817] = 7
      "0000111" when "01010101100101010", -- t[43818] = 7
      "0000111" when "01010101100101011", -- t[43819] = 7
      "0000111" when "01010101100101100", -- t[43820] = 7
      "0000111" when "01010101100101101", -- t[43821] = 7
      "0000111" when "01010101100101110", -- t[43822] = 7
      "0000111" when "01010101100101111", -- t[43823] = 7
      "0000111" when "01010101100110000", -- t[43824] = 7
      "0000111" when "01010101100110001", -- t[43825] = 7
      "0000111" when "01010101100110010", -- t[43826] = 7
      "0000111" when "01010101100110011", -- t[43827] = 7
      "0000111" when "01010101100110100", -- t[43828] = 7
      "0000111" when "01010101100110101", -- t[43829] = 7
      "0000111" when "01010101100110110", -- t[43830] = 7
      "0000111" when "01010101100110111", -- t[43831] = 7
      "0000111" when "01010101100111000", -- t[43832] = 7
      "0000111" when "01010101100111001", -- t[43833] = 7
      "0000111" when "01010101100111010", -- t[43834] = 7
      "0000111" when "01010101100111011", -- t[43835] = 7
      "0000111" when "01010101100111100", -- t[43836] = 7
      "0000111" when "01010101100111101", -- t[43837] = 7
      "0000111" when "01010101100111110", -- t[43838] = 7
      "0000111" when "01010101100111111", -- t[43839] = 7
      "0000111" when "01010101101000000", -- t[43840] = 7
      "0000111" when "01010101101000001", -- t[43841] = 7
      "0000111" when "01010101101000010", -- t[43842] = 7
      "0000111" when "01010101101000011", -- t[43843] = 7
      "0000111" when "01010101101000100", -- t[43844] = 7
      "0000111" when "01010101101000101", -- t[43845] = 7
      "0000111" when "01010101101000110", -- t[43846] = 7
      "0000111" when "01010101101000111", -- t[43847] = 7
      "0000111" when "01010101101001000", -- t[43848] = 7
      "0000111" when "01010101101001001", -- t[43849] = 7
      "0000111" when "01010101101001010", -- t[43850] = 7
      "0000111" when "01010101101001011", -- t[43851] = 7
      "0000111" when "01010101101001100", -- t[43852] = 7
      "0000111" when "01010101101001101", -- t[43853] = 7
      "0000111" when "01010101101001110", -- t[43854] = 7
      "0000111" when "01010101101001111", -- t[43855] = 7
      "0000111" when "01010101101010000", -- t[43856] = 7
      "0000111" when "01010101101010001", -- t[43857] = 7
      "0000111" when "01010101101010010", -- t[43858] = 7
      "0000111" when "01010101101010011", -- t[43859] = 7
      "0000111" when "01010101101010100", -- t[43860] = 7
      "0000111" when "01010101101010101", -- t[43861] = 7
      "0000111" when "01010101101010110", -- t[43862] = 7
      "0000111" when "01010101101010111", -- t[43863] = 7
      "0000111" when "01010101101011000", -- t[43864] = 7
      "0000111" when "01010101101011001", -- t[43865] = 7
      "0000111" when "01010101101011010", -- t[43866] = 7
      "0000111" when "01010101101011011", -- t[43867] = 7
      "0000111" when "01010101101011100", -- t[43868] = 7
      "0000111" when "01010101101011101", -- t[43869] = 7
      "0000111" when "01010101101011110", -- t[43870] = 7
      "0000111" when "01010101101011111", -- t[43871] = 7
      "0000111" when "01010101101100000", -- t[43872] = 7
      "0000111" when "01010101101100001", -- t[43873] = 7
      "0000111" when "01010101101100010", -- t[43874] = 7
      "0000111" when "01010101101100011", -- t[43875] = 7
      "0000111" when "01010101101100100", -- t[43876] = 7
      "0000111" when "01010101101100101", -- t[43877] = 7
      "0000111" when "01010101101100110", -- t[43878] = 7
      "0000111" when "01010101101100111", -- t[43879] = 7
      "0000111" when "01010101101101000", -- t[43880] = 7
      "0000111" when "01010101101101001", -- t[43881] = 7
      "0000111" when "01010101101101010", -- t[43882] = 7
      "0000111" when "01010101101101011", -- t[43883] = 7
      "0000111" when "01010101101101100", -- t[43884] = 7
      "0000111" when "01010101101101101", -- t[43885] = 7
      "0000111" when "01010101101101110", -- t[43886] = 7
      "0000111" when "01010101101101111", -- t[43887] = 7
      "0000111" when "01010101101110000", -- t[43888] = 7
      "0000111" when "01010101101110001", -- t[43889] = 7
      "0000111" when "01010101101110010", -- t[43890] = 7
      "0000111" when "01010101101110011", -- t[43891] = 7
      "0000111" when "01010101101110100", -- t[43892] = 7
      "0000111" when "01010101101110101", -- t[43893] = 7
      "0000111" when "01010101101110110", -- t[43894] = 7
      "0000111" when "01010101101110111", -- t[43895] = 7
      "0000111" when "01010101101111000", -- t[43896] = 7
      "0000111" when "01010101101111001", -- t[43897] = 7
      "0000111" when "01010101101111010", -- t[43898] = 7
      "0000111" when "01010101101111011", -- t[43899] = 7
      "0000111" when "01010101101111100", -- t[43900] = 7
      "0000111" when "01010101101111101", -- t[43901] = 7
      "0000111" when "01010101101111110", -- t[43902] = 7
      "0000111" when "01010101101111111", -- t[43903] = 7
      "0000111" when "01010101110000000", -- t[43904] = 7
      "0000111" when "01010101110000001", -- t[43905] = 7
      "0000111" when "01010101110000010", -- t[43906] = 7
      "0000111" when "01010101110000011", -- t[43907] = 7
      "0000111" when "01010101110000100", -- t[43908] = 7
      "0000111" when "01010101110000101", -- t[43909] = 7
      "0000111" when "01010101110000110", -- t[43910] = 7
      "0000111" when "01010101110000111", -- t[43911] = 7
      "0000111" when "01010101110001000", -- t[43912] = 7
      "0000111" when "01010101110001001", -- t[43913] = 7
      "0000111" when "01010101110001010", -- t[43914] = 7
      "0000111" when "01010101110001011", -- t[43915] = 7
      "0000111" when "01010101110001100", -- t[43916] = 7
      "0000111" when "01010101110001101", -- t[43917] = 7
      "0000111" when "01010101110001110", -- t[43918] = 7
      "0000111" when "01010101110001111", -- t[43919] = 7
      "0000111" when "01010101110010000", -- t[43920] = 7
      "0000111" when "01010101110010001", -- t[43921] = 7
      "0000111" when "01010101110010010", -- t[43922] = 7
      "0000111" when "01010101110010011", -- t[43923] = 7
      "0000111" when "01010101110010100", -- t[43924] = 7
      "0000111" when "01010101110010101", -- t[43925] = 7
      "0000111" when "01010101110010110", -- t[43926] = 7
      "0000111" when "01010101110010111", -- t[43927] = 7
      "0000111" when "01010101110011000", -- t[43928] = 7
      "0000111" when "01010101110011001", -- t[43929] = 7
      "0000111" when "01010101110011010", -- t[43930] = 7
      "0000111" when "01010101110011011", -- t[43931] = 7
      "0000111" when "01010101110011100", -- t[43932] = 7
      "0000111" when "01010101110011101", -- t[43933] = 7
      "0000111" when "01010101110011110", -- t[43934] = 7
      "0000111" when "01010101110011111", -- t[43935] = 7
      "0000111" when "01010101110100000", -- t[43936] = 7
      "0000111" when "01010101110100001", -- t[43937] = 7
      "0000111" when "01010101110100010", -- t[43938] = 7
      "0000111" when "01010101110100011", -- t[43939] = 7
      "0000111" when "01010101110100100", -- t[43940] = 7
      "0000111" when "01010101110100101", -- t[43941] = 7
      "0000111" when "01010101110100110", -- t[43942] = 7
      "0000111" when "01010101110100111", -- t[43943] = 7
      "0000111" when "01010101110101000", -- t[43944] = 7
      "0000111" when "01010101110101001", -- t[43945] = 7
      "0000111" when "01010101110101010", -- t[43946] = 7
      "0000111" when "01010101110101011", -- t[43947] = 7
      "0000111" when "01010101110101100", -- t[43948] = 7
      "0000111" when "01010101110101101", -- t[43949] = 7
      "0000111" when "01010101110101110", -- t[43950] = 7
      "0000111" when "01010101110101111", -- t[43951] = 7
      "0000111" when "01010101110110000", -- t[43952] = 7
      "0000111" when "01010101110110001", -- t[43953] = 7
      "0000111" when "01010101110110010", -- t[43954] = 7
      "0000111" when "01010101110110011", -- t[43955] = 7
      "0000111" when "01010101110110100", -- t[43956] = 7
      "0000111" when "01010101110110101", -- t[43957] = 7
      "0000111" when "01010101110110110", -- t[43958] = 7
      "0000111" when "01010101110110111", -- t[43959] = 7
      "0000111" when "01010101110111000", -- t[43960] = 7
      "0000111" when "01010101110111001", -- t[43961] = 7
      "0000111" when "01010101110111010", -- t[43962] = 7
      "0000111" when "01010101110111011", -- t[43963] = 7
      "0000111" when "01010101110111100", -- t[43964] = 7
      "0000111" when "01010101110111101", -- t[43965] = 7
      "0000111" when "01010101110111110", -- t[43966] = 7
      "0000111" when "01010101110111111", -- t[43967] = 7
      "0000111" when "01010101111000000", -- t[43968] = 7
      "0000111" when "01010101111000001", -- t[43969] = 7
      "0000111" when "01010101111000010", -- t[43970] = 7
      "0000111" when "01010101111000011", -- t[43971] = 7
      "0000111" when "01010101111000100", -- t[43972] = 7
      "0000111" when "01010101111000101", -- t[43973] = 7
      "0000111" when "01010101111000110", -- t[43974] = 7
      "0000111" when "01010101111000111", -- t[43975] = 7
      "0000111" when "01010101111001000", -- t[43976] = 7
      "0000111" when "01010101111001001", -- t[43977] = 7
      "0000111" when "01010101111001010", -- t[43978] = 7
      "0000111" when "01010101111001011", -- t[43979] = 7
      "0000111" when "01010101111001100", -- t[43980] = 7
      "0000111" when "01010101111001101", -- t[43981] = 7
      "0000111" when "01010101111001110", -- t[43982] = 7
      "0000111" when "01010101111001111", -- t[43983] = 7
      "0000111" when "01010101111010000", -- t[43984] = 7
      "0000111" when "01010101111010001", -- t[43985] = 7
      "0000111" when "01010101111010010", -- t[43986] = 7
      "0000111" when "01010101111010011", -- t[43987] = 7
      "0000111" when "01010101111010100", -- t[43988] = 7
      "0000111" when "01010101111010101", -- t[43989] = 7
      "0000111" when "01010101111010110", -- t[43990] = 7
      "0000111" when "01010101111010111", -- t[43991] = 7
      "0000111" when "01010101111011000", -- t[43992] = 7
      "0000111" when "01010101111011001", -- t[43993] = 7
      "0000111" when "01010101111011010", -- t[43994] = 7
      "0000111" when "01010101111011011", -- t[43995] = 7
      "0000111" when "01010101111011100", -- t[43996] = 7
      "0000111" when "01010101111011101", -- t[43997] = 7
      "0000111" when "01010101111011110", -- t[43998] = 7
      "0000111" when "01010101111011111", -- t[43999] = 7
      "0000111" when "01010101111100000", -- t[44000] = 7
      "0000111" when "01010101111100001", -- t[44001] = 7
      "0000111" when "01010101111100010", -- t[44002] = 7
      "0000111" when "01010101111100011", -- t[44003] = 7
      "0000111" when "01010101111100100", -- t[44004] = 7
      "0000111" when "01010101111100101", -- t[44005] = 7
      "0000111" when "01010101111100110", -- t[44006] = 7
      "0000111" when "01010101111100111", -- t[44007] = 7
      "0000111" when "01010101111101000", -- t[44008] = 7
      "0000111" when "01010101111101001", -- t[44009] = 7
      "0000111" when "01010101111101010", -- t[44010] = 7
      "0000111" when "01010101111101011", -- t[44011] = 7
      "0000111" when "01010101111101100", -- t[44012] = 7
      "0000111" when "01010101111101101", -- t[44013] = 7
      "0000111" when "01010101111101110", -- t[44014] = 7
      "0000111" when "01010101111101111", -- t[44015] = 7
      "0000111" when "01010101111110000", -- t[44016] = 7
      "0000111" when "01010101111110001", -- t[44017] = 7
      "0000111" when "01010101111110010", -- t[44018] = 7
      "0000111" when "01010101111110011", -- t[44019] = 7
      "0000111" when "01010101111110100", -- t[44020] = 7
      "0000111" when "01010101111110101", -- t[44021] = 7
      "0000111" when "01010101111110110", -- t[44022] = 7
      "0000111" when "01010101111110111", -- t[44023] = 7
      "0000111" when "01010101111111000", -- t[44024] = 7
      "0000111" when "01010101111111001", -- t[44025] = 7
      "0000111" when "01010101111111010", -- t[44026] = 7
      "0000111" when "01010101111111011", -- t[44027] = 7
      "0000111" when "01010101111111100", -- t[44028] = 7
      "0000111" when "01010101111111101", -- t[44029] = 7
      "0000111" when "01010101111111110", -- t[44030] = 7
      "0000111" when "01010101111111111", -- t[44031] = 7
      "0000111" when "01010110000000000", -- t[44032] = 7
      "0000111" when "01010110000000001", -- t[44033] = 7
      "0000111" when "01010110000000010", -- t[44034] = 7
      "0000111" when "01010110000000011", -- t[44035] = 7
      "0000111" when "01010110000000100", -- t[44036] = 7
      "0000111" when "01010110000000101", -- t[44037] = 7
      "0000111" when "01010110000000110", -- t[44038] = 7
      "0000111" when "01010110000000111", -- t[44039] = 7
      "0000111" when "01010110000001000", -- t[44040] = 7
      "0000111" when "01010110000001001", -- t[44041] = 7
      "0000111" when "01010110000001010", -- t[44042] = 7
      "0000111" when "01010110000001011", -- t[44043] = 7
      "0000111" when "01010110000001100", -- t[44044] = 7
      "0000111" when "01010110000001101", -- t[44045] = 7
      "0000111" when "01010110000001110", -- t[44046] = 7
      "0000111" when "01010110000001111", -- t[44047] = 7
      "0000111" when "01010110000010000", -- t[44048] = 7
      "0000111" when "01010110000010001", -- t[44049] = 7
      "0000111" when "01010110000010010", -- t[44050] = 7
      "0000111" when "01010110000010011", -- t[44051] = 7
      "0000111" when "01010110000010100", -- t[44052] = 7
      "0000111" when "01010110000010101", -- t[44053] = 7
      "0001000" when "01010110000010110", -- t[44054] = 8
      "0001000" when "01010110000010111", -- t[44055] = 8
      "0001000" when "01010110000011000", -- t[44056] = 8
      "0001000" when "01010110000011001", -- t[44057] = 8
      "0001000" when "01010110000011010", -- t[44058] = 8
      "0001000" when "01010110000011011", -- t[44059] = 8
      "0001000" when "01010110000011100", -- t[44060] = 8
      "0001000" when "01010110000011101", -- t[44061] = 8
      "0001000" when "01010110000011110", -- t[44062] = 8
      "0001000" when "01010110000011111", -- t[44063] = 8
      "0001000" when "01010110000100000", -- t[44064] = 8
      "0001000" when "01010110000100001", -- t[44065] = 8
      "0001000" when "01010110000100010", -- t[44066] = 8
      "0001000" when "01010110000100011", -- t[44067] = 8
      "0001000" when "01010110000100100", -- t[44068] = 8
      "0001000" when "01010110000100101", -- t[44069] = 8
      "0001000" when "01010110000100110", -- t[44070] = 8
      "0001000" when "01010110000100111", -- t[44071] = 8
      "0001000" when "01010110000101000", -- t[44072] = 8
      "0001000" when "01010110000101001", -- t[44073] = 8
      "0001000" when "01010110000101010", -- t[44074] = 8
      "0001000" when "01010110000101011", -- t[44075] = 8
      "0001000" when "01010110000101100", -- t[44076] = 8
      "0001000" when "01010110000101101", -- t[44077] = 8
      "0001000" when "01010110000101110", -- t[44078] = 8
      "0001000" when "01010110000101111", -- t[44079] = 8
      "0001000" when "01010110000110000", -- t[44080] = 8
      "0001000" when "01010110000110001", -- t[44081] = 8
      "0001000" when "01010110000110010", -- t[44082] = 8
      "0001000" when "01010110000110011", -- t[44083] = 8
      "0001000" when "01010110000110100", -- t[44084] = 8
      "0001000" when "01010110000110101", -- t[44085] = 8
      "0001000" when "01010110000110110", -- t[44086] = 8
      "0001000" when "01010110000110111", -- t[44087] = 8
      "0001000" when "01010110000111000", -- t[44088] = 8
      "0001000" when "01010110000111001", -- t[44089] = 8
      "0001000" when "01010110000111010", -- t[44090] = 8
      "0001000" when "01010110000111011", -- t[44091] = 8
      "0001000" when "01010110000111100", -- t[44092] = 8
      "0001000" when "01010110000111101", -- t[44093] = 8
      "0001000" when "01010110000111110", -- t[44094] = 8
      "0001000" when "01010110000111111", -- t[44095] = 8
      "0001000" when "01010110001000000", -- t[44096] = 8
      "0001000" when "01010110001000001", -- t[44097] = 8
      "0001000" when "01010110001000010", -- t[44098] = 8
      "0001000" when "01010110001000011", -- t[44099] = 8
      "0001000" when "01010110001000100", -- t[44100] = 8
      "0001000" when "01010110001000101", -- t[44101] = 8
      "0001000" when "01010110001000110", -- t[44102] = 8
      "0001000" when "01010110001000111", -- t[44103] = 8
      "0001000" when "01010110001001000", -- t[44104] = 8
      "0001000" when "01010110001001001", -- t[44105] = 8
      "0001000" when "01010110001001010", -- t[44106] = 8
      "0001000" when "01010110001001011", -- t[44107] = 8
      "0001000" when "01010110001001100", -- t[44108] = 8
      "0001000" when "01010110001001101", -- t[44109] = 8
      "0001000" when "01010110001001110", -- t[44110] = 8
      "0001000" when "01010110001001111", -- t[44111] = 8
      "0001000" when "01010110001010000", -- t[44112] = 8
      "0001000" when "01010110001010001", -- t[44113] = 8
      "0001000" when "01010110001010010", -- t[44114] = 8
      "0001000" when "01010110001010011", -- t[44115] = 8
      "0001000" when "01010110001010100", -- t[44116] = 8
      "0001000" when "01010110001010101", -- t[44117] = 8
      "0001000" when "01010110001010110", -- t[44118] = 8
      "0001000" when "01010110001010111", -- t[44119] = 8
      "0001000" when "01010110001011000", -- t[44120] = 8
      "0001000" when "01010110001011001", -- t[44121] = 8
      "0001000" when "01010110001011010", -- t[44122] = 8
      "0001000" when "01010110001011011", -- t[44123] = 8
      "0001000" when "01010110001011100", -- t[44124] = 8
      "0001000" when "01010110001011101", -- t[44125] = 8
      "0001000" when "01010110001011110", -- t[44126] = 8
      "0001000" when "01010110001011111", -- t[44127] = 8
      "0001000" when "01010110001100000", -- t[44128] = 8
      "0001000" when "01010110001100001", -- t[44129] = 8
      "0001000" when "01010110001100010", -- t[44130] = 8
      "0001000" when "01010110001100011", -- t[44131] = 8
      "0001000" when "01010110001100100", -- t[44132] = 8
      "0001000" when "01010110001100101", -- t[44133] = 8
      "0001000" when "01010110001100110", -- t[44134] = 8
      "0001000" when "01010110001100111", -- t[44135] = 8
      "0001000" when "01010110001101000", -- t[44136] = 8
      "0001000" when "01010110001101001", -- t[44137] = 8
      "0001000" when "01010110001101010", -- t[44138] = 8
      "0001000" when "01010110001101011", -- t[44139] = 8
      "0001000" when "01010110001101100", -- t[44140] = 8
      "0001000" when "01010110001101101", -- t[44141] = 8
      "0001000" when "01010110001101110", -- t[44142] = 8
      "0001000" when "01010110001101111", -- t[44143] = 8
      "0001000" when "01010110001110000", -- t[44144] = 8
      "0001000" when "01010110001110001", -- t[44145] = 8
      "0001000" when "01010110001110010", -- t[44146] = 8
      "0001000" when "01010110001110011", -- t[44147] = 8
      "0001000" when "01010110001110100", -- t[44148] = 8
      "0001000" when "01010110001110101", -- t[44149] = 8
      "0001000" when "01010110001110110", -- t[44150] = 8
      "0001000" when "01010110001110111", -- t[44151] = 8
      "0001000" when "01010110001111000", -- t[44152] = 8
      "0001000" when "01010110001111001", -- t[44153] = 8
      "0001000" when "01010110001111010", -- t[44154] = 8
      "0001000" when "01010110001111011", -- t[44155] = 8
      "0001000" when "01010110001111100", -- t[44156] = 8
      "0001000" when "01010110001111101", -- t[44157] = 8
      "0001000" when "01010110001111110", -- t[44158] = 8
      "0001000" when "01010110001111111", -- t[44159] = 8
      "0001000" when "01010110010000000", -- t[44160] = 8
      "0001000" when "01010110010000001", -- t[44161] = 8
      "0001000" when "01010110010000010", -- t[44162] = 8
      "0001000" when "01010110010000011", -- t[44163] = 8
      "0001000" when "01010110010000100", -- t[44164] = 8
      "0001000" when "01010110010000101", -- t[44165] = 8
      "0001000" when "01010110010000110", -- t[44166] = 8
      "0001000" when "01010110010000111", -- t[44167] = 8
      "0001000" when "01010110010001000", -- t[44168] = 8
      "0001000" when "01010110010001001", -- t[44169] = 8
      "0001000" when "01010110010001010", -- t[44170] = 8
      "0001000" when "01010110010001011", -- t[44171] = 8
      "0001000" when "01010110010001100", -- t[44172] = 8
      "0001000" when "01010110010001101", -- t[44173] = 8
      "0001000" when "01010110010001110", -- t[44174] = 8
      "0001000" when "01010110010001111", -- t[44175] = 8
      "0001000" when "01010110010010000", -- t[44176] = 8
      "0001000" when "01010110010010001", -- t[44177] = 8
      "0001000" when "01010110010010010", -- t[44178] = 8
      "0001000" when "01010110010010011", -- t[44179] = 8
      "0001000" when "01010110010010100", -- t[44180] = 8
      "0001000" when "01010110010010101", -- t[44181] = 8
      "0001000" when "01010110010010110", -- t[44182] = 8
      "0001000" when "01010110010010111", -- t[44183] = 8
      "0001000" when "01010110010011000", -- t[44184] = 8
      "0001000" when "01010110010011001", -- t[44185] = 8
      "0001000" when "01010110010011010", -- t[44186] = 8
      "0001000" when "01010110010011011", -- t[44187] = 8
      "0001000" when "01010110010011100", -- t[44188] = 8
      "0001000" when "01010110010011101", -- t[44189] = 8
      "0001000" when "01010110010011110", -- t[44190] = 8
      "0001000" when "01010110010011111", -- t[44191] = 8
      "0001000" when "01010110010100000", -- t[44192] = 8
      "0001000" when "01010110010100001", -- t[44193] = 8
      "0001000" when "01010110010100010", -- t[44194] = 8
      "0001000" when "01010110010100011", -- t[44195] = 8
      "0001000" when "01010110010100100", -- t[44196] = 8
      "0001000" when "01010110010100101", -- t[44197] = 8
      "0001000" when "01010110010100110", -- t[44198] = 8
      "0001000" when "01010110010100111", -- t[44199] = 8
      "0001000" when "01010110010101000", -- t[44200] = 8
      "0001000" when "01010110010101001", -- t[44201] = 8
      "0001000" when "01010110010101010", -- t[44202] = 8
      "0001000" when "01010110010101011", -- t[44203] = 8
      "0001000" when "01010110010101100", -- t[44204] = 8
      "0001000" when "01010110010101101", -- t[44205] = 8
      "0001000" when "01010110010101110", -- t[44206] = 8
      "0001000" when "01010110010101111", -- t[44207] = 8
      "0001000" when "01010110010110000", -- t[44208] = 8
      "0001000" when "01010110010110001", -- t[44209] = 8
      "0001000" when "01010110010110010", -- t[44210] = 8
      "0001000" when "01010110010110011", -- t[44211] = 8
      "0001000" when "01010110010110100", -- t[44212] = 8
      "0001000" when "01010110010110101", -- t[44213] = 8
      "0001000" when "01010110010110110", -- t[44214] = 8
      "0001000" when "01010110010110111", -- t[44215] = 8
      "0001000" when "01010110010111000", -- t[44216] = 8
      "0001000" when "01010110010111001", -- t[44217] = 8
      "0001000" when "01010110010111010", -- t[44218] = 8
      "0001000" when "01010110010111011", -- t[44219] = 8
      "0001000" when "01010110010111100", -- t[44220] = 8
      "0001000" when "01010110010111101", -- t[44221] = 8
      "0001000" when "01010110010111110", -- t[44222] = 8
      "0001000" when "01010110010111111", -- t[44223] = 8
      "0001000" when "01010110011000000", -- t[44224] = 8
      "0001000" when "01010110011000001", -- t[44225] = 8
      "0001000" when "01010110011000010", -- t[44226] = 8
      "0001000" when "01010110011000011", -- t[44227] = 8
      "0001000" when "01010110011000100", -- t[44228] = 8
      "0001000" when "01010110011000101", -- t[44229] = 8
      "0001000" when "01010110011000110", -- t[44230] = 8
      "0001000" when "01010110011000111", -- t[44231] = 8
      "0001000" when "01010110011001000", -- t[44232] = 8
      "0001000" when "01010110011001001", -- t[44233] = 8
      "0001000" when "01010110011001010", -- t[44234] = 8
      "0001000" when "01010110011001011", -- t[44235] = 8
      "0001000" when "01010110011001100", -- t[44236] = 8
      "0001000" when "01010110011001101", -- t[44237] = 8
      "0001000" when "01010110011001110", -- t[44238] = 8
      "0001000" when "01010110011001111", -- t[44239] = 8
      "0001000" when "01010110011010000", -- t[44240] = 8
      "0001000" when "01010110011010001", -- t[44241] = 8
      "0001000" when "01010110011010010", -- t[44242] = 8
      "0001000" when "01010110011010011", -- t[44243] = 8
      "0001000" when "01010110011010100", -- t[44244] = 8
      "0001000" when "01010110011010101", -- t[44245] = 8
      "0001000" when "01010110011010110", -- t[44246] = 8
      "0001000" when "01010110011010111", -- t[44247] = 8
      "0001000" when "01010110011011000", -- t[44248] = 8
      "0001000" when "01010110011011001", -- t[44249] = 8
      "0001000" when "01010110011011010", -- t[44250] = 8
      "0001000" when "01010110011011011", -- t[44251] = 8
      "0001000" when "01010110011011100", -- t[44252] = 8
      "0001000" when "01010110011011101", -- t[44253] = 8
      "0001000" when "01010110011011110", -- t[44254] = 8
      "0001000" when "01010110011011111", -- t[44255] = 8
      "0001000" when "01010110011100000", -- t[44256] = 8
      "0001000" when "01010110011100001", -- t[44257] = 8
      "0001000" when "01010110011100010", -- t[44258] = 8
      "0001000" when "01010110011100011", -- t[44259] = 8
      "0001000" when "01010110011100100", -- t[44260] = 8
      "0001000" when "01010110011100101", -- t[44261] = 8
      "0001000" when "01010110011100110", -- t[44262] = 8
      "0001000" when "01010110011100111", -- t[44263] = 8
      "0001000" when "01010110011101000", -- t[44264] = 8
      "0001000" when "01010110011101001", -- t[44265] = 8
      "0001000" when "01010110011101010", -- t[44266] = 8
      "0001000" when "01010110011101011", -- t[44267] = 8
      "0001000" when "01010110011101100", -- t[44268] = 8
      "0001000" when "01010110011101101", -- t[44269] = 8
      "0001000" when "01010110011101110", -- t[44270] = 8
      "0001000" when "01010110011101111", -- t[44271] = 8
      "0001000" when "01010110011110000", -- t[44272] = 8
      "0001000" when "01010110011110001", -- t[44273] = 8
      "0001000" when "01010110011110010", -- t[44274] = 8
      "0001000" when "01010110011110011", -- t[44275] = 8
      "0001000" when "01010110011110100", -- t[44276] = 8
      "0001000" when "01010110011110101", -- t[44277] = 8
      "0001000" when "01010110011110110", -- t[44278] = 8
      "0001000" when "01010110011110111", -- t[44279] = 8
      "0001000" when "01010110011111000", -- t[44280] = 8
      "0001000" when "01010110011111001", -- t[44281] = 8
      "0001000" when "01010110011111010", -- t[44282] = 8
      "0001000" when "01010110011111011", -- t[44283] = 8
      "0001000" when "01010110011111100", -- t[44284] = 8
      "0001000" when "01010110011111101", -- t[44285] = 8
      "0001000" when "01010110011111110", -- t[44286] = 8
      "0001000" when "01010110011111111", -- t[44287] = 8
      "0001000" when "01010110100000000", -- t[44288] = 8
      "0001000" when "01010110100000001", -- t[44289] = 8
      "0001000" when "01010110100000010", -- t[44290] = 8
      "0001000" when "01010110100000011", -- t[44291] = 8
      "0001000" when "01010110100000100", -- t[44292] = 8
      "0001000" when "01010110100000101", -- t[44293] = 8
      "0001000" when "01010110100000110", -- t[44294] = 8
      "0001000" when "01010110100000111", -- t[44295] = 8
      "0001000" when "01010110100001000", -- t[44296] = 8
      "0001000" when "01010110100001001", -- t[44297] = 8
      "0001000" when "01010110100001010", -- t[44298] = 8
      "0001000" when "01010110100001011", -- t[44299] = 8
      "0001000" when "01010110100001100", -- t[44300] = 8
      "0001000" when "01010110100001101", -- t[44301] = 8
      "0001000" when "01010110100001110", -- t[44302] = 8
      "0001000" when "01010110100001111", -- t[44303] = 8
      "0001000" when "01010110100010000", -- t[44304] = 8
      "0001000" when "01010110100010001", -- t[44305] = 8
      "0001000" when "01010110100010010", -- t[44306] = 8
      "0001000" when "01010110100010011", -- t[44307] = 8
      "0001000" when "01010110100010100", -- t[44308] = 8
      "0001000" when "01010110100010101", -- t[44309] = 8
      "0001000" when "01010110100010110", -- t[44310] = 8
      "0001000" when "01010110100010111", -- t[44311] = 8
      "0001000" when "01010110100011000", -- t[44312] = 8
      "0001000" when "01010110100011001", -- t[44313] = 8
      "0001000" when "01010110100011010", -- t[44314] = 8
      "0001000" when "01010110100011011", -- t[44315] = 8
      "0001000" when "01010110100011100", -- t[44316] = 8
      "0001000" when "01010110100011101", -- t[44317] = 8
      "0001000" when "01010110100011110", -- t[44318] = 8
      "0001000" when "01010110100011111", -- t[44319] = 8
      "0001000" when "01010110100100000", -- t[44320] = 8
      "0001000" when "01010110100100001", -- t[44321] = 8
      "0001000" when "01010110100100010", -- t[44322] = 8
      "0001000" when "01010110100100011", -- t[44323] = 8
      "0001000" when "01010110100100100", -- t[44324] = 8
      "0001000" when "01010110100100101", -- t[44325] = 8
      "0001000" when "01010110100100110", -- t[44326] = 8
      "0001000" when "01010110100100111", -- t[44327] = 8
      "0001000" when "01010110100101000", -- t[44328] = 8
      "0001000" when "01010110100101001", -- t[44329] = 8
      "0001000" when "01010110100101010", -- t[44330] = 8
      "0001000" when "01010110100101011", -- t[44331] = 8
      "0001000" when "01010110100101100", -- t[44332] = 8
      "0001000" when "01010110100101101", -- t[44333] = 8
      "0001000" when "01010110100101110", -- t[44334] = 8
      "0001000" when "01010110100101111", -- t[44335] = 8
      "0001000" when "01010110100110000", -- t[44336] = 8
      "0001000" when "01010110100110001", -- t[44337] = 8
      "0001000" when "01010110100110010", -- t[44338] = 8
      "0001000" when "01010110100110011", -- t[44339] = 8
      "0001000" when "01010110100110100", -- t[44340] = 8
      "0001000" when "01010110100110101", -- t[44341] = 8
      "0001000" when "01010110100110110", -- t[44342] = 8
      "0001000" when "01010110100110111", -- t[44343] = 8
      "0001000" when "01010110100111000", -- t[44344] = 8
      "0001000" when "01010110100111001", -- t[44345] = 8
      "0001000" when "01010110100111010", -- t[44346] = 8
      "0001000" when "01010110100111011", -- t[44347] = 8
      "0001000" when "01010110100111100", -- t[44348] = 8
      "0001000" when "01010110100111101", -- t[44349] = 8
      "0001000" when "01010110100111110", -- t[44350] = 8
      "0001000" when "01010110100111111", -- t[44351] = 8
      "0001000" when "01010110101000000", -- t[44352] = 8
      "0001000" when "01010110101000001", -- t[44353] = 8
      "0001000" when "01010110101000010", -- t[44354] = 8
      "0001000" when "01010110101000011", -- t[44355] = 8
      "0001000" when "01010110101000100", -- t[44356] = 8
      "0001000" when "01010110101000101", -- t[44357] = 8
      "0001000" when "01010110101000110", -- t[44358] = 8
      "0001000" when "01010110101000111", -- t[44359] = 8
      "0001000" when "01010110101001000", -- t[44360] = 8
      "0001000" when "01010110101001001", -- t[44361] = 8
      "0001000" when "01010110101001010", -- t[44362] = 8
      "0001000" when "01010110101001011", -- t[44363] = 8
      "0001000" when "01010110101001100", -- t[44364] = 8
      "0001000" when "01010110101001101", -- t[44365] = 8
      "0001000" when "01010110101001110", -- t[44366] = 8
      "0001000" when "01010110101001111", -- t[44367] = 8
      "0001000" when "01010110101010000", -- t[44368] = 8
      "0001000" when "01010110101010001", -- t[44369] = 8
      "0001000" when "01010110101010010", -- t[44370] = 8
      "0001000" when "01010110101010011", -- t[44371] = 8
      "0001000" when "01010110101010100", -- t[44372] = 8
      "0001000" when "01010110101010101", -- t[44373] = 8
      "0001000" when "01010110101010110", -- t[44374] = 8
      "0001000" when "01010110101010111", -- t[44375] = 8
      "0001000" when "01010110101011000", -- t[44376] = 8
      "0001000" when "01010110101011001", -- t[44377] = 8
      "0001000" when "01010110101011010", -- t[44378] = 8
      "0001000" when "01010110101011011", -- t[44379] = 8
      "0001000" when "01010110101011100", -- t[44380] = 8
      "0001000" when "01010110101011101", -- t[44381] = 8
      "0001000" when "01010110101011110", -- t[44382] = 8
      "0001000" when "01010110101011111", -- t[44383] = 8
      "0001000" when "01010110101100000", -- t[44384] = 8
      "0001000" when "01010110101100001", -- t[44385] = 8
      "0001000" when "01010110101100010", -- t[44386] = 8
      "0001000" when "01010110101100011", -- t[44387] = 8
      "0001000" when "01010110101100100", -- t[44388] = 8
      "0001000" when "01010110101100101", -- t[44389] = 8
      "0001000" when "01010110101100110", -- t[44390] = 8
      "0001000" when "01010110101100111", -- t[44391] = 8
      "0001000" when "01010110101101000", -- t[44392] = 8
      "0001000" when "01010110101101001", -- t[44393] = 8
      "0001000" when "01010110101101010", -- t[44394] = 8
      "0001000" when "01010110101101011", -- t[44395] = 8
      "0001000" when "01010110101101100", -- t[44396] = 8
      "0001000" when "01010110101101101", -- t[44397] = 8
      "0001000" when "01010110101101110", -- t[44398] = 8
      "0001000" when "01010110101101111", -- t[44399] = 8
      "0001000" when "01010110101110000", -- t[44400] = 8
      "0001000" when "01010110101110001", -- t[44401] = 8
      "0001000" when "01010110101110010", -- t[44402] = 8
      "0001000" when "01010110101110011", -- t[44403] = 8
      "0001000" when "01010110101110100", -- t[44404] = 8
      "0001000" when "01010110101110101", -- t[44405] = 8
      "0001000" when "01010110101110110", -- t[44406] = 8
      "0001000" when "01010110101110111", -- t[44407] = 8
      "0001000" when "01010110101111000", -- t[44408] = 8
      "0001000" when "01010110101111001", -- t[44409] = 8
      "0001000" when "01010110101111010", -- t[44410] = 8
      "0001000" when "01010110101111011", -- t[44411] = 8
      "0001000" when "01010110101111100", -- t[44412] = 8
      "0001000" when "01010110101111101", -- t[44413] = 8
      "0001000" when "01010110101111110", -- t[44414] = 8
      "0001000" when "01010110101111111", -- t[44415] = 8
      "0001000" when "01010110110000000", -- t[44416] = 8
      "0001000" when "01010110110000001", -- t[44417] = 8
      "0001000" when "01010110110000010", -- t[44418] = 8
      "0001000" when "01010110110000011", -- t[44419] = 8
      "0001000" when "01010110110000100", -- t[44420] = 8
      "0001000" when "01010110110000101", -- t[44421] = 8
      "0001000" when "01010110110000110", -- t[44422] = 8
      "0001000" when "01010110110000111", -- t[44423] = 8
      "0001000" when "01010110110001000", -- t[44424] = 8
      "0001000" when "01010110110001001", -- t[44425] = 8
      "0001000" when "01010110110001010", -- t[44426] = 8
      "0001000" when "01010110110001011", -- t[44427] = 8
      "0001000" when "01010110110001100", -- t[44428] = 8
      "0001000" when "01010110110001101", -- t[44429] = 8
      "0001000" when "01010110110001110", -- t[44430] = 8
      "0001000" when "01010110110001111", -- t[44431] = 8
      "0001000" when "01010110110010000", -- t[44432] = 8
      "0001000" when "01010110110010001", -- t[44433] = 8
      "0001000" when "01010110110010010", -- t[44434] = 8
      "0001000" when "01010110110010011", -- t[44435] = 8
      "0001000" when "01010110110010100", -- t[44436] = 8
      "0001000" when "01010110110010101", -- t[44437] = 8
      "0001000" when "01010110110010110", -- t[44438] = 8
      "0001000" when "01010110110010111", -- t[44439] = 8
      "0001000" when "01010110110011000", -- t[44440] = 8
      "0001000" when "01010110110011001", -- t[44441] = 8
      "0001000" when "01010110110011010", -- t[44442] = 8
      "0001000" when "01010110110011011", -- t[44443] = 8
      "0001000" when "01010110110011100", -- t[44444] = 8
      "0001000" when "01010110110011101", -- t[44445] = 8
      "0001000" when "01010110110011110", -- t[44446] = 8
      "0001000" when "01010110110011111", -- t[44447] = 8
      "0001000" when "01010110110100000", -- t[44448] = 8
      "0001000" when "01010110110100001", -- t[44449] = 8
      "0001000" when "01010110110100010", -- t[44450] = 8
      "0001000" when "01010110110100011", -- t[44451] = 8
      "0001000" when "01010110110100100", -- t[44452] = 8
      "0001000" when "01010110110100101", -- t[44453] = 8
      "0001000" when "01010110110100110", -- t[44454] = 8
      "0001000" when "01010110110100111", -- t[44455] = 8
      "0001000" when "01010110110101000", -- t[44456] = 8
      "0001000" when "01010110110101001", -- t[44457] = 8
      "0001000" when "01010110110101010", -- t[44458] = 8
      "0001000" when "01010110110101011", -- t[44459] = 8
      "0001000" when "01010110110101100", -- t[44460] = 8
      "0001000" when "01010110110101101", -- t[44461] = 8
      "0001000" when "01010110110101110", -- t[44462] = 8
      "0001000" when "01010110110101111", -- t[44463] = 8
      "0001000" when "01010110110110000", -- t[44464] = 8
      "0001000" when "01010110110110001", -- t[44465] = 8
      "0001000" when "01010110110110010", -- t[44466] = 8
      "0001000" when "01010110110110011", -- t[44467] = 8
      "0001000" when "01010110110110100", -- t[44468] = 8
      "0001000" when "01010110110110101", -- t[44469] = 8
      "0001000" when "01010110110110110", -- t[44470] = 8
      "0001000" when "01010110110110111", -- t[44471] = 8
      "0001000" when "01010110110111000", -- t[44472] = 8
      "0001000" when "01010110110111001", -- t[44473] = 8
      "0001000" when "01010110110111010", -- t[44474] = 8
      "0001000" when "01010110110111011", -- t[44475] = 8
      "0001000" when "01010110110111100", -- t[44476] = 8
      "0001000" when "01010110110111101", -- t[44477] = 8
      "0001000" when "01010110110111110", -- t[44478] = 8
      "0001000" when "01010110110111111", -- t[44479] = 8
      "0001000" when "01010110111000000", -- t[44480] = 8
      "0001000" when "01010110111000001", -- t[44481] = 8
      "0001000" when "01010110111000010", -- t[44482] = 8
      "0001000" when "01010110111000011", -- t[44483] = 8
      "0001000" when "01010110111000100", -- t[44484] = 8
      "0001000" when "01010110111000101", -- t[44485] = 8
      "0001000" when "01010110111000110", -- t[44486] = 8
      "0001000" when "01010110111000111", -- t[44487] = 8
      "0001000" when "01010110111001000", -- t[44488] = 8
      "0001000" when "01010110111001001", -- t[44489] = 8
      "0001000" when "01010110111001010", -- t[44490] = 8
      "0001000" when "01010110111001011", -- t[44491] = 8
      "0001000" when "01010110111001100", -- t[44492] = 8
      "0001000" when "01010110111001101", -- t[44493] = 8
      "0001000" when "01010110111001110", -- t[44494] = 8
      "0001000" when "01010110111001111", -- t[44495] = 8
      "0001000" when "01010110111010000", -- t[44496] = 8
      "0001000" when "01010110111010001", -- t[44497] = 8
      "0001000" when "01010110111010010", -- t[44498] = 8
      "0001000" when "01010110111010011", -- t[44499] = 8
      "0001000" when "01010110111010100", -- t[44500] = 8
      "0001000" when "01010110111010101", -- t[44501] = 8
      "0001000" when "01010110111010110", -- t[44502] = 8
      "0001000" when "01010110111010111", -- t[44503] = 8
      "0001000" when "01010110111011000", -- t[44504] = 8
      "0001000" when "01010110111011001", -- t[44505] = 8
      "0001000" when "01010110111011010", -- t[44506] = 8
      "0001000" when "01010110111011011", -- t[44507] = 8
      "0001000" when "01010110111011100", -- t[44508] = 8
      "0001000" when "01010110111011101", -- t[44509] = 8
      "0001000" when "01010110111011110", -- t[44510] = 8
      "0001000" when "01010110111011111", -- t[44511] = 8
      "0001000" when "01010110111100000", -- t[44512] = 8
      "0001000" when "01010110111100001", -- t[44513] = 8
      "0001000" when "01010110111100010", -- t[44514] = 8
      "0001000" when "01010110111100011", -- t[44515] = 8
      "0001000" when "01010110111100100", -- t[44516] = 8
      "0001000" when "01010110111100101", -- t[44517] = 8
      "0001000" when "01010110111100110", -- t[44518] = 8
      "0001000" when "01010110111100111", -- t[44519] = 8
      "0001000" when "01010110111101000", -- t[44520] = 8
      "0001000" when "01010110111101001", -- t[44521] = 8
      "0001000" when "01010110111101010", -- t[44522] = 8
      "0001000" when "01010110111101011", -- t[44523] = 8
      "0001000" when "01010110111101100", -- t[44524] = 8
      "0001000" when "01010110111101101", -- t[44525] = 8
      "0001000" when "01010110111101110", -- t[44526] = 8
      "0001000" when "01010110111101111", -- t[44527] = 8
      "0001000" when "01010110111110000", -- t[44528] = 8
      "0001000" when "01010110111110001", -- t[44529] = 8
      "0001000" when "01010110111110010", -- t[44530] = 8
      "0001000" when "01010110111110011", -- t[44531] = 8
      "0001000" when "01010110111110100", -- t[44532] = 8
      "0001000" when "01010110111110101", -- t[44533] = 8
      "0001000" when "01010110111110110", -- t[44534] = 8
      "0001000" when "01010110111110111", -- t[44535] = 8
      "0001000" when "01010110111111000", -- t[44536] = 8
      "0001000" when "01010110111111001", -- t[44537] = 8
      "0001000" when "01010110111111010", -- t[44538] = 8
      "0001000" when "01010110111111011", -- t[44539] = 8
      "0001000" when "01010110111111100", -- t[44540] = 8
      "0001000" when "01010110111111101", -- t[44541] = 8
      "0001000" when "01010110111111110", -- t[44542] = 8
      "0001000" when "01010110111111111", -- t[44543] = 8
      "0001000" when "01010111000000000", -- t[44544] = 8
      "0001000" when "01010111000000001", -- t[44545] = 8
      "0001000" when "01010111000000010", -- t[44546] = 8
      "0001000" when "01010111000000011", -- t[44547] = 8
      "0001000" when "01010111000000100", -- t[44548] = 8
      "0001000" when "01010111000000101", -- t[44549] = 8
      "0001000" when "01010111000000110", -- t[44550] = 8
      "0001000" when "01010111000000111", -- t[44551] = 8
      "0001000" when "01010111000001000", -- t[44552] = 8
      "0001000" when "01010111000001001", -- t[44553] = 8
      "0001000" when "01010111000001010", -- t[44554] = 8
      "0001000" when "01010111000001011", -- t[44555] = 8
      "0001000" when "01010111000001100", -- t[44556] = 8
      "0001000" when "01010111000001101", -- t[44557] = 8
      "0001000" when "01010111000001110", -- t[44558] = 8
      "0001000" when "01010111000001111", -- t[44559] = 8
      "0001000" when "01010111000010000", -- t[44560] = 8
      "0001000" when "01010111000010001", -- t[44561] = 8
      "0001000" when "01010111000010010", -- t[44562] = 8
      "0001000" when "01010111000010011", -- t[44563] = 8
      "0001000" when "01010111000010100", -- t[44564] = 8
      "0001000" when "01010111000010101", -- t[44565] = 8
      "0001000" when "01010111000010110", -- t[44566] = 8
      "0001000" when "01010111000010111", -- t[44567] = 8
      "0001000" when "01010111000011000", -- t[44568] = 8
      "0001000" when "01010111000011001", -- t[44569] = 8
      "0001000" when "01010111000011010", -- t[44570] = 8
      "0001000" when "01010111000011011", -- t[44571] = 8
      "0001000" when "01010111000011100", -- t[44572] = 8
      "0001000" when "01010111000011101", -- t[44573] = 8
      "0001000" when "01010111000011110", -- t[44574] = 8
      "0001000" when "01010111000011111", -- t[44575] = 8
      "0001000" when "01010111000100000", -- t[44576] = 8
      "0001000" when "01010111000100001", -- t[44577] = 8
      "0001000" when "01010111000100010", -- t[44578] = 8
      "0001000" when "01010111000100011", -- t[44579] = 8
      "0001000" when "01010111000100100", -- t[44580] = 8
      "0001000" when "01010111000100101", -- t[44581] = 8
      "0001000" when "01010111000100110", -- t[44582] = 8
      "0001000" when "01010111000100111", -- t[44583] = 8
      "0001000" when "01010111000101000", -- t[44584] = 8
      "0001000" when "01010111000101001", -- t[44585] = 8
      "0001000" when "01010111000101010", -- t[44586] = 8
      "0001000" when "01010111000101011", -- t[44587] = 8
      "0001000" when "01010111000101100", -- t[44588] = 8
      "0001000" when "01010111000101101", -- t[44589] = 8
      "0001000" when "01010111000101110", -- t[44590] = 8
      "0001000" when "01010111000101111", -- t[44591] = 8
      "0001000" when "01010111000110000", -- t[44592] = 8
      "0001000" when "01010111000110001", -- t[44593] = 8
      "0001000" when "01010111000110010", -- t[44594] = 8
      "0001000" when "01010111000110011", -- t[44595] = 8
      "0001000" when "01010111000110100", -- t[44596] = 8
      "0001000" when "01010111000110101", -- t[44597] = 8
      "0001000" when "01010111000110110", -- t[44598] = 8
      "0001000" when "01010111000110111", -- t[44599] = 8
      "0001000" when "01010111000111000", -- t[44600] = 8
      "0001000" when "01010111000111001", -- t[44601] = 8
      "0001000" when "01010111000111010", -- t[44602] = 8
      "0001000" when "01010111000111011", -- t[44603] = 8
      "0001000" when "01010111000111100", -- t[44604] = 8
      "0001000" when "01010111000111101", -- t[44605] = 8
      "0001000" when "01010111000111110", -- t[44606] = 8
      "0001000" when "01010111000111111", -- t[44607] = 8
      "0001000" when "01010111001000000", -- t[44608] = 8
      "0001000" when "01010111001000001", -- t[44609] = 8
      "0001000" when "01010111001000010", -- t[44610] = 8
      "0001000" when "01010111001000011", -- t[44611] = 8
      "0001000" when "01010111001000100", -- t[44612] = 8
      "0001000" when "01010111001000101", -- t[44613] = 8
      "0001000" when "01010111001000110", -- t[44614] = 8
      "0001000" when "01010111001000111", -- t[44615] = 8
      "0001000" when "01010111001001000", -- t[44616] = 8
      "0001000" when "01010111001001001", -- t[44617] = 8
      "0001000" when "01010111001001010", -- t[44618] = 8
      "0001000" when "01010111001001011", -- t[44619] = 8
      "0001000" when "01010111001001100", -- t[44620] = 8
      "0001000" when "01010111001001101", -- t[44621] = 8
      "0001000" when "01010111001001110", -- t[44622] = 8
      "0001000" when "01010111001001111", -- t[44623] = 8
      "0001000" when "01010111001010000", -- t[44624] = 8
      "0001000" when "01010111001010001", -- t[44625] = 8
      "0001000" when "01010111001010010", -- t[44626] = 8
      "0001000" when "01010111001010011", -- t[44627] = 8
      "0001000" when "01010111001010100", -- t[44628] = 8
      "0001000" when "01010111001010101", -- t[44629] = 8
      "0001000" when "01010111001010110", -- t[44630] = 8
      "0001000" when "01010111001010111", -- t[44631] = 8
      "0001000" when "01010111001011000", -- t[44632] = 8
      "0001000" when "01010111001011001", -- t[44633] = 8
      "0001000" when "01010111001011010", -- t[44634] = 8
      "0001000" when "01010111001011011", -- t[44635] = 8
      "0001000" when "01010111001011100", -- t[44636] = 8
      "0001000" when "01010111001011101", -- t[44637] = 8
      "0001000" when "01010111001011110", -- t[44638] = 8
      "0001000" when "01010111001011111", -- t[44639] = 8
      "0001000" when "01010111001100000", -- t[44640] = 8
      "0001000" when "01010111001100001", -- t[44641] = 8
      "0001000" when "01010111001100010", -- t[44642] = 8
      "0001000" when "01010111001100011", -- t[44643] = 8
      "0001000" when "01010111001100100", -- t[44644] = 8
      "0001000" when "01010111001100101", -- t[44645] = 8
      "0001000" when "01010111001100110", -- t[44646] = 8
      "0001000" when "01010111001100111", -- t[44647] = 8
      "0001000" when "01010111001101000", -- t[44648] = 8
      "0001000" when "01010111001101001", -- t[44649] = 8
      "0001000" when "01010111001101010", -- t[44650] = 8
      "0001000" when "01010111001101011", -- t[44651] = 8
      "0001000" when "01010111001101100", -- t[44652] = 8
      "0001000" when "01010111001101101", -- t[44653] = 8
      "0001000" when "01010111001101110", -- t[44654] = 8
      "0001000" when "01010111001101111", -- t[44655] = 8
      "0001000" when "01010111001110000", -- t[44656] = 8
      "0001000" when "01010111001110001", -- t[44657] = 8
      "0001000" when "01010111001110010", -- t[44658] = 8
      "0001000" when "01010111001110011", -- t[44659] = 8
      "0001000" when "01010111001110100", -- t[44660] = 8
      "0001000" when "01010111001110101", -- t[44661] = 8
      "0001000" when "01010111001110110", -- t[44662] = 8
      "0001000" when "01010111001110111", -- t[44663] = 8
      "0001000" when "01010111001111000", -- t[44664] = 8
      "0001000" when "01010111001111001", -- t[44665] = 8
      "0001000" when "01010111001111010", -- t[44666] = 8
      "0001000" when "01010111001111011", -- t[44667] = 8
      "0001000" when "01010111001111100", -- t[44668] = 8
      "0001000" when "01010111001111101", -- t[44669] = 8
      "0001000" when "01010111001111110", -- t[44670] = 8
      "0001000" when "01010111001111111", -- t[44671] = 8
      "0001000" when "01010111010000000", -- t[44672] = 8
      "0001000" when "01010111010000001", -- t[44673] = 8
      "0001000" when "01010111010000010", -- t[44674] = 8
      "0001000" when "01010111010000011", -- t[44675] = 8
      "0001000" when "01010111010000100", -- t[44676] = 8
      "0001000" when "01010111010000101", -- t[44677] = 8
      "0001000" when "01010111010000110", -- t[44678] = 8
      "0001000" when "01010111010000111", -- t[44679] = 8
      "0001000" when "01010111010001000", -- t[44680] = 8
      "0001000" when "01010111010001001", -- t[44681] = 8
      "0001000" when "01010111010001010", -- t[44682] = 8
      "0001000" when "01010111010001011", -- t[44683] = 8
      "0001000" when "01010111010001100", -- t[44684] = 8
      "0001000" when "01010111010001101", -- t[44685] = 8
      "0001000" when "01010111010001110", -- t[44686] = 8
      "0001000" when "01010111010001111", -- t[44687] = 8
      "0001000" when "01010111010010000", -- t[44688] = 8
      "0001000" when "01010111010010001", -- t[44689] = 8
      "0001000" when "01010111010010010", -- t[44690] = 8
      "0001000" when "01010111010010011", -- t[44691] = 8
      "0001000" when "01010111010010100", -- t[44692] = 8
      "0001000" when "01010111010010101", -- t[44693] = 8
      "0001000" when "01010111010010110", -- t[44694] = 8
      "0001000" when "01010111010010111", -- t[44695] = 8
      "0001000" when "01010111010011000", -- t[44696] = 8
      "0001000" when "01010111010011001", -- t[44697] = 8
      "0001000" when "01010111010011010", -- t[44698] = 8
      "0001000" when "01010111010011011", -- t[44699] = 8
      "0001000" when "01010111010011100", -- t[44700] = 8
      "0001000" when "01010111010011101", -- t[44701] = 8
      "0001000" when "01010111010011110", -- t[44702] = 8
      "0001000" when "01010111010011111", -- t[44703] = 8
      "0001000" when "01010111010100000", -- t[44704] = 8
      "0001000" when "01010111010100001", -- t[44705] = 8
      "0001000" when "01010111010100010", -- t[44706] = 8
      "0001000" when "01010111010100011", -- t[44707] = 8
      "0001000" when "01010111010100100", -- t[44708] = 8
      "0001000" when "01010111010100101", -- t[44709] = 8
      "0001000" when "01010111010100110", -- t[44710] = 8
      "0001000" when "01010111010100111", -- t[44711] = 8
      "0001000" when "01010111010101000", -- t[44712] = 8
      "0001000" when "01010111010101001", -- t[44713] = 8
      "0001000" when "01010111010101010", -- t[44714] = 8
      "0001000" when "01010111010101011", -- t[44715] = 8
      "0001000" when "01010111010101100", -- t[44716] = 8
      "0001000" when "01010111010101101", -- t[44717] = 8
      "0001000" when "01010111010101110", -- t[44718] = 8
      "0001000" when "01010111010101111", -- t[44719] = 8
      "0001000" when "01010111010110000", -- t[44720] = 8
      "0001000" when "01010111010110001", -- t[44721] = 8
      "0001000" when "01010111010110010", -- t[44722] = 8
      "0001000" when "01010111010110011", -- t[44723] = 8
      "0001000" when "01010111010110100", -- t[44724] = 8
      "0001000" when "01010111010110101", -- t[44725] = 8
      "0001000" when "01010111010110110", -- t[44726] = 8
      "0001000" when "01010111010110111", -- t[44727] = 8
      "0001000" when "01010111010111000", -- t[44728] = 8
      "0001000" when "01010111010111001", -- t[44729] = 8
      "0001000" when "01010111010111010", -- t[44730] = 8
      "0001000" when "01010111010111011", -- t[44731] = 8
      "0001000" when "01010111010111100", -- t[44732] = 8
      "0001000" when "01010111010111101", -- t[44733] = 8
      "0001000" when "01010111010111110", -- t[44734] = 8
      "0001000" when "01010111010111111", -- t[44735] = 8
      "0001000" when "01010111011000000", -- t[44736] = 8
      "0001000" when "01010111011000001", -- t[44737] = 8
      "0001000" when "01010111011000010", -- t[44738] = 8
      "0001000" when "01010111011000011", -- t[44739] = 8
      "0001000" when "01010111011000100", -- t[44740] = 8
      "0001000" when "01010111011000101", -- t[44741] = 8
      "0001000" when "01010111011000110", -- t[44742] = 8
      "0001000" when "01010111011000111", -- t[44743] = 8
      "0001000" when "01010111011001000", -- t[44744] = 8
      "0001000" when "01010111011001001", -- t[44745] = 8
      "0001000" when "01010111011001010", -- t[44746] = 8
      "0001000" when "01010111011001011", -- t[44747] = 8
      "0001000" when "01010111011001100", -- t[44748] = 8
      "0001000" when "01010111011001101", -- t[44749] = 8
      "0001000" when "01010111011001110", -- t[44750] = 8
      "0001000" when "01010111011001111", -- t[44751] = 8
      "0001000" when "01010111011010000", -- t[44752] = 8
      "0001000" when "01010111011010001", -- t[44753] = 8
      "0001000" when "01010111011010010", -- t[44754] = 8
      "0001000" when "01010111011010011", -- t[44755] = 8
      "0001000" when "01010111011010100", -- t[44756] = 8
      "0001000" when "01010111011010101", -- t[44757] = 8
      "0001000" when "01010111011010110", -- t[44758] = 8
      "0001000" when "01010111011010111", -- t[44759] = 8
      "0001000" when "01010111011011000", -- t[44760] = 8
      "0001000" when "01010111011011001", -- t[44761] = 8
      "0001000" when "01010111011011010", -- t[44762] = 8
      "0001000" when "01010111011011011", -- t[44763] = 8
      "0001000" when "01010111011011100", -- t[44764] = 8
      "0001000" when "01010111011011101", -- t[44765] = 8
      "0001000" when "01010111011011110", -- t[44766] = 8
      "0001000" when "01010111011011111", -- t[44767] = 8
      "0001000" when "01010111011100000", -- t[44768] = 8
      "0001000" when "01010111011100001", -- t[44769] = 8
      "0001000" when "01010111011100010", -- t[44770] = 8
      "0001000" when "01010111011100011", -- t[44771] = 8
      "0001000" when "01010111011100100", -- t[44772] = 8
      "0001000" when "01010111011100101", -- t[44773] = 8
      "0001000" when "01010111011100110", -- t[44774] = 8
      "0001000" when "01010111011100111", -- t[44775] = 8
      "0001000" when "01010111011101000", -- t[44776] = 8
      "0001000" when "01010111011101001", -- t[44777] = 8
      "0001000" when "01010111011101010", -- t[44778] = 8
      "0001000" when "01010111011101011", -- t[44779] = 8
      "0001000" when "01010111011101100", -- t[44780] = 8
      "0001000" when "01010111011101101", -- t[44781] = 8
      "0001000" when "01010111011101110", -- t[44782] = 8
      "0001000" when "01010111011101111", -- t[44783] = 8
      "0001000" when "01010111011110000", -- t[44784] = 8
      "0001000" when "01010111011110001", -- t[44785] = 8
      "0001000" when "01010111011110010", -- t[44786] = 8
      "0001000" when "01010111011110011", -- t[44787] = 8
      "0001000" when "01010111011110100", -- t[44788] = 8
      "0001000" when "01010111011110101", -- t[44789] = 8
      "0001000" when "01010111011110110", -- t[44790] = 8
      "0001000" when "01010111011110111", -- t[44791] = 8
      "0001000" when "01010111011111000", -- t[44792] = 8
      "0001000" when "01010111011111001", -- t[44793] = 8
      "0001000" when "01010111011111010", -- t[44794] = 8
      "0001000" when "01010111011111011", -- t[44795] = 8
      "0001000" when "01010111011111100", -- t[44796] = 8
      "0001000" when "01010111011111101", -- t[44797] = 8
      "0001000" when "01010111011111110", -- t[44798] = 8
      "0001000" when "01010111011111111", -- t[44799] = 8
      "0001000" when "01010111100000000", -- t[44800] = 8
      "0001000" when "01010111100000001", -- t[44801] = 8
      "0001000" when "01010111100000010", -- t[44802] = 8
      "0001000" when "01010111100000011", -- t[44803] = 8
      "0001000" when "01010111100000100", -- t[44804] = 8
      "0001000" when "01010111100000101", -- t[44805] = 8
      "0001000" when "01010111100000110", -- t[44806] = 8
      "0001000" when "01010111100000111", -- t[44807] = 8
      "0001000" when "01010111100001000", -- t[44808] = 8
      "0001000" when "01010111100001001", -- t[44809] = 8
      "0001000" when "01010111100001010", -- t[44810] = 8
      "0001000" when "01010111100001011", -- t[44811] = 8
      "0001000" when "01010111100001100", -- t[44812] = 8
      "0001000" when "01010111100001101", -- t[44813] = 8
      "0001000" when "01010111100001110", -- t[44814] = 8
      "0001000" when "01010111100001111", -- t[44815] = 8
      "0001000" when "01010111100010000", -- t[44816] = 8
      "0001000" when "01010111100010001", -- t[44817] = 8
      "0001000" when "01010111100010010", -- t[44818] = 8
      "0001000" when "01010111100010011", -- t[44819] = 8
      "0001000" when "01010111100010100", -- t[44820] = 8
      "0001000" when "01010111100010101", -- t[44821] = 8
      "0001000" when "01010111100010110", -- t[44822] = 8
      "0001000" when "01010111100010111", -- t[44823] = 8
      "0001000" when "01010111100011000", -- t[44824] = 8
      "0001000" when "01010111100011001", -- t[44825] = 8
      "0001000" when "01010111100011010", -- t[44826] = 8
      "0001000" when "01010111100011011", -- t[44827] = 8
      "0001000" when "01010111100011100", -- t[44828] = 8
      "0001000" when "01010111100011101", -- t[44829] = 8
      "0001000" when "01010111100011110", -- t[44830] = 8
      "0001000" when "01010111100011111", -- t[44831] = 8
      "0001000" when "01010111100100000", -- t[44832] = 8
      "0001000" when "01010111100100001", -- t[44833] = 8
      "0001000" when "01010111100100010", -- t[44834] = 8
      "0001000" when "01010111100100011", -- t[44835] = 8
      "0001000" when "01010111100100100", -- t[44836] = 8
      "0001000" when "01010111100100101", -- t[44837] = 8
      "0001000" when "01010111100100110", -- t[44838] = 8
      "0001000" when "01010111100100111", -- t[44839] = 8
      "0001000" when "01010111100101000", -- t[44840] = 8
      "0001000" when "01010111100101001", -- t[44841] = 8
      "0001000" when "01010111100101010", -- t[44842] = 8
      "0001000" when "01010111100101011", -- t[44843] = 8
      "0001000" when "01010111100101100", -- t[44844] = 8
      "0001000" when "01010111100101101", -- t[44845] = 8
      "0001000" when "01010111100101110", -- t[44846] = 8
      "0001000" when "01010111100101111", -- t[44847] = 8
      "0001000" when "01010111100110000", -- t[44848] = 8
      "0001000" when "01010111100110001", -- t[44849] = 8
      "0001000" when "01010111100110010", -- t[44850] = 8
      "0001000" when "01010111100110011", -- t[44851] = 8
      "0001000" when "01010111100110100", -- t[44852] = 8
      "0001000" when "01010111100110101", -- t[44853] = 8
      "0001000" when "01010111100110110", -- t[44854] = 8
      "0001000" when "01010111100110111", -- t[44855] = 8
      "0001000" when "01010111100111000", -- t[44856] = 8
      "0001000" when "01010111100111001", -- t[44857] = 8
      "0001000" when "01010111100111010", -- t[44858] = 8
      "0001000" when "01010111100111011", -- t[44859] = 8
      "0001000" when "01010111100111100", -- t[44860] = 8
      "0001000" when "01010111100111101", -- t[44861] = 8
      "0001000" when "01010111100111110", -- t[44862] = 8
      "0001000" when "01010111100111111", -- t[44863] = 8
      "0001000" when "01010111101000000", -- t[44864] = 8
      "0001000" when "01010111101000001", -- t[44865] = 8
      "0001000" when "01010111101000010", -- t[44866] = 8
      "0001000" when "01010111101000011", -- t[44867] = 8
      "0001000" when "01010111101000100", -- t[44868] = 8
      "0001000" when "01010111101000101", -- t[44869] = 8
      "0001000" when "01010111101000110", -- t[44870] = 8
      "0001000" when "01010111101000111", -- t[44871] = 8
      "0001000" when "01010111101001000", -- t[44872] = 8
      "0001000" when "01010111101001001", -- t[44873] = 8
      "0001000" when "01010111101001010", -- t[44874] = 8
      "0001000" when "01010111101001011", -- t[44875] = 8
      "0001000" when "01010111101001100", -- t[44876] = 8
      "0001000" when "01010111101001101", -- t[44877] = 8
      "0001000" when "01010111101001110", -- t[44878] = 8
      "0001000" when "01010111101001111", -- t[44879] = 8
      "0001000" when "01010111101010000", -- t[44880] = 8
      "0001000" when "01010111101010001", -- t[44881] = 8
      "0001000" when "01010111101010010", -- t[44882] = 8
      "0001000" when "01010111101010011", -- t[44883] = 8
      "0001000" when "01010111101010100", -- t[44884] = 8
      "0001000" when "01010111101010101", -- t[44885] = 8
      "0001000" when "01010111101010110", -- t[44886] = 8
      "0001000" when "01010111101010111", -- t[44887] = 8
      "0001000" when "01010111101011000", -- t[44888] = 8
      "0001000" when "01010111101011001", -- t[44889] = 8
      "0001000" when "01010111101011010", -- t[44890] = 8
      "0001000" when "01010111101011011", -- t[44891] = 8
      "0001000" when "01010111101011100", -- t[44892] = 8
      "0001000" when "01010111101011101", -- t[44893] = 8
      "0001000" when "01010111101011110", -- t[44894] = 8
      "0001000" when "01010111101011111", -- t[44895] = 8
      "0001000" when "01010111101100000", -- t[44896] = 8
      "0001000" when "01010111101100001", -- t[44897] = 8
      "0001000" when "01010111101100010", -- t[44898] = 8
      "0001000" when "01010111101100011", -- t[44899] = 8
      "0001000" when "01010111101100100", -- t[44900] = 8
      "0001000" when "01010111101100101", -- t[44901] = 8
      "0001000" when "01010111101100110", -- t[44902] = 8
      "0001000" when "01010111101100111", -- t[44903] = 8
      "0001000" when "01010111101101000", -- t[44904] = 8
      "0001000" when "01010111101101001", -- t[44905] = 8
      "0001000" when "01010111101101010", -- t[44906] = 8
      "0001000" when "01010111101101011", -- t[44907] = 8
      "0001000" when "01010111101101100", -- t[44908] = 8
      "0001000" when "01010111101101101", -- t[44909] = 8
      "0001000" when "01010111101101110", -- t[44910] = 8
      "0001000" when "01010111101101111", -- t[44911] = 8
      "0001000" when "01010111101110000", -- t[44912] = 8
      "0001000" when "01010111101110001", -- t[44913] = 8
      "0001000" when "01010111101110010", -- t[44914] = 8
      "0001000" when "01010111101110011", -- t[44915] = 8
      "0001000" when "01010111101110100", -- t[44916] = 8
      "0001000" when "01010111101110101", -- t[44917] = 8
      "0001000" when "01010111101110110", -- t[44918] = 8
      "0001000" when "01010111101110111", -- t[44919] = 8
      "0001000" when "01010111101111000", -- t[44920] = 8
      "0001000" when "01010111101111001", -- t[44921] = 8
      "0001000" when "01010111101111010", -- t[44922] = 8
      "0001000" when "01010111101111011", -- t[44923] = 8
      "0001000" when "01010111101111100", -- t[44924] = 8
      "0001000" when "01010111101111101", -- t[44925] = 8
      "0001000" when "01010111101111110", -- t[44926] = 8
      "0001000" when "01010111101111111", -- t[44927] = 8
      "0001000" when "01010111110000000", -- t[44928] = 8
      "0001000" when "01010111110000001", -- t[44929] = 8
      "0001000" when "01010111110000010", -- t[44930] = 8
      "0001000" when "01010111110000011", -- t[44931] = 8
      "0001000" when "01010111110000100", -- t[44932] = 8
      "0001000" when "01010111110000101", -- t[44933] = 8
      "0001000" when "01010111110000110", -- t[44934] = 8
      "0001000" when "01010111110000111", -- t[44935] = 8
      "0001000" when "01010111110001000", -- t[44936] = 8
      "0001000" when "01010111110001001", -- t[44937] = 8
      "0001000" when "01010111110001010", -- t[44938] = 8
      "0001000" when "01010111110001011", -- t[44939] = 8
      "0001000" when "01010111110001100", -- t[44940] = 8
      "0001000" when "01010111110001101", -- t[44941] = 8
      "0001000" when "01010111110001110", -- t[44942] = 8
      "0001000" when "01010111110001111", -- t[44943] = 8
      "0001000" when "01010111110010000", -- t[44944] = 8
      "0001000" when "01010111110010001", -- t[44945] = 8
      "0001000" when "01010111110010010", -- t[44946] = 8
      "0001000" when "01010111110010011", -- t[44947] = 8
      "0001000" when "01010111110010100", -- t[44948] = 8
      "0001000" when "01010111110010101", -- t[44949] = 8
      "0001000" when "01010111110010110", -- t[44950] = 8
      "0001000" when "01010111110010111", -- t[44951] = 8
      "0001000" when "01010111110011000", -- t[44952] = 8
      "0001000" when "01010111110011001", -- t[44953] = 8
      "0001000" when "01010111110011010", -- t[44954] = 8
      "0001000" when "01010111110011011", -- t[44955] = 8
      "0001000" when "01010111110011100", -- t[44956] = 8
      "0001000" when "01010111110011101", -- t[44957] = 8
      "0001000" when "01010111110011110", -- t[44958] = 8
      "0001000" when "01010111110011111", -- t[44959] = 8
      "0001000" when "01010111110100000", -- t[44960] = 8
      "0001000" when "01010111110100001", -- t[44961] = 8
      "0001000" when "01010111110100010", -- t[44962] = 8
      "0001000" when "01010111110100011", -- t[44963] = 8
      "0001000" when "01010111110100100", -- t[44964] = 8
      "0001000" when "01010111110100101", -- t[44965] = 8
      "0001000" when "01010111110100110", -- t[44966] = 8
      "0001000" when "01010111110100111", -- t[44967] = 8
      "0001000" when "01010111110101000", -- t[44968] = 8
      "0001000" when "01010111110101001", -- t[44969] = 8
      "0001000" when "01010111110101010", -- t[44970] = 8
      "0001000" when "01010111110101011", -- t[44971] = 8
      "0001000" when "01010111110101100", -- t[44972] = 8
      "0001000" when "01010111110101101", -- t[44973] = 8
      "0001000" when "01010111110101110", -- t[44974] = 8
      "0001000" when "01010111110101111", -- t[44975] = 8
      "0001000" when "01010111110110000", -- t[44976] = 8
      "0001000" when "01010111110110001", -- t[44977] = 8
      "0001000" when "01010111110110010", -- t[44978] = 8
      "0001000" when "01010111110110011", -- t[44979] = 8
      "0001000" when "01010111110110100", -- t[44980] = 8
      "0001000" when "01010111110110101", -- t[44981] = 8
      "0001000" when "01010111110110110", -- t[44982] = 8
      "0001000" when "01010111110110111", -- t[44983] = 8
      "0001000" when "01010111110111000", -- t[44984] = 8
      "0001000" when "01010111110111001", -- t[44985] = 8
      "0001000" when "01010111110111010", -- t[44986] = 8
      "0001000" when "01010111110111011", -- t[44987] = 8
      "0001000" when "01010111110111100", -- t[44988] = 8
      "0001000" when "01010111110111101", -- t[44989] = 8
      "0001000" when "01010111110111110", -- t[44990] = 8
      "0001000" when "01010111110111111", -- t[44991] = 8
      "0001000" when "01010111111000000", -- t[44992] = 8
      "0001000" when "01010111111000001", -- t[44993] = 8
      "0001000" when "01010111111000010", -- t[44994] = 8
      "0001000" when "01010111111000011", -- t[44995] = 8
      "0001000" when "01010111111000100", -- t[44996] = 8
      "0001000" when "01010111111000101", -- t[44997] = 8
      "0001000" when "01010111111000110", -- t[44998] = 8
      "0001000" when "01010111111000111", -- t[44999] = 8
      "0001000" when "01010111111001000", -- t[45000] = 8
      "0001000" when "01010111111001001", -- t[45001] = 8
      "0001000" when "01010111111001010", -- t[45002] = 8
      "0001000" when "01010111111001011", -- t[45003] = 8
      "0001000" when "01010111111001100", -- t[45004] = 8
      "0001000" when "01010111111001101", -- t[45005] = 8
      "0001000" when "01010111111001110", -- t[45006] = 8
      "0001000" when "01010111111001111", -- t[45007] = 8
      "0001000" when "01010111111010000", -- t[45008] = 8
      "0001000" when "01010111111010001", -- t[45009] = 8
      "0001000" when "01010111111010010", -- t[45010] = 8
      "0001000" when "01010111111010011", -- t[45011] = 8
      "0001000" when "01010111111010100", -- t[45012] = 8
      "0001000" when "01010111111010101", -- t[45013] = 8
      "0001000" when "01010111111010110", -- t[45014] = 8
      "0001000" when "01010111111010111", -- t[45015] = 8
      "0001000" when "01010111111011000", -- t[45016] = 8
      "0001000" when "01010111111011001", -- t[45017] = 8
      "0001000" when "01010111111011010", -- t[45018] = 8
      "0001000" when "01010111111011011", -- t[45019] = 8
      "0001000" when "01010111111011100", -- t[45020] = 8
      "0001000" when "01010111111011101", -- t[45021] = 8
      "0001000" when "01010111111011110", -- t[45022] = 8
      "0001000" when "01010111111011111", -- t[45023] = 8
      "0001000" when "01010111111100000", -- t[45024] = 8
      "0001000" when "01010111111100001", -- t[45025] = 8
      "0001000" when "01010111111100010", -- t[45026] = 8
      "0001000" when "01010111111100011", -- t[45027] = 8
      "0001000" when "01010111111100100", -- t[45028] = 8
      "0001000" when "01010111111100101", -- t[45029] = 8
      "0001000" when "01010111111100110", -- t[45030] = 8
      "0001000" when "01010111111100111", -- t[45031] = 8
      "0001000" when "01010111111101000", -- t[45032] = 8
      "0001000" when "01010111111101001", -- t[45033] = 8
      "0001000" when "01010111111101010", -- t[45034] = 8
      "0001000" when "01010111111101011", -- t[45035] = 8
      "0001000" when "01010111111101100", -- t[45036] = 8
      "0001000" when "01010111111101101", -- t[45037] = 8
      "0001000" when "01010111111101110", -- t[45038] = 8
      "0001000" when "01010111111101111", -- t[45039] = 8
      "0001000" when "01010111111110000", -- t[45040] = 8
      "0001000" when "01010111111110001", -- t[45041] = 8
      "0001000" when "01010111111110010", -- t[45042] = 8
      "0001000" when "01010111111110011", -- t[45043] = 8
      "0001000" when "01010111111110100", -- t[45044] = 8
      "0001000" when "01010111111110101", -- t[45045] = 8
      "0001000" when "01010111111110110", -- t[45046] = 8
      "0001000" when "01010111111110111", -- t[45047] = 8
      "0001000" when "01010111111111000", -- t[45048] = 8
      "0001000" when "01010111111111001", -- t[45049] = 8
      "0001000" when "01010111111111010", -- t[45050] = 8
      "0001000" when "01010111111111011", -- t[45051] = 8
      "0001000" when "01010111111111100", -- t[45052] = 8
      "0001000" when "01010111111111101", -- t[45053] = 8
      "0001000" when "01010111111111110", -- t[45054] = 8
      "0001000" when "01010111111111111", -- t[45055] = 8
      "0001000" when "01011000000000000", -- t[45056] = 8
      "0001000" when "01011000000000001", -- t[45057] = 8
      "0001000" when "01011000000000010", -- t[45058] = 8
      "0001000" when "01011000000000011", -- t[45059] = 8
      "0001000" when "01011000000000100", -- t[45060] = 8
      "0001000" when "01011000000000101", -- t[45061] = 8
      "0001000" when "01011000000000110", -- t[45062] = 8
      "0001000" when "01011000000000111", -- t[45063] = 8
      "0001000" when "01011000000001000", -- t[45064] = 8
      "0001000" when "01011000000001001", -- t[45065] = 8
      "0001000" when "01011000000001010", -- t[45066] = 8
      "0001000" when "01011000000001011", -- t[45067] = 8
      "0001000" when "01011000000001100", -- t[45068] = 8
      "0001000" when "01011000000001101", -- t[45069] = 8
      "0001000" when "01011000000001110", -- t[45070] = 8
      "0001000" when "01011000000001111", -- t[45071] = 8
      "0001000" when "01011000000010000", -- t[45072] = 8
      "0001000" when "01011000000010001", -- t[45073] = 8
      "0001000" when "01011000000010010", -- t[45074] = 8
      "0001000" when "01011000000010011", -- t[45075] = 8
      "0001000" when "01011000000010100", -- t[45076] = 8
      "0001000" when "01011000000010101", -- t[45077] = 8
      "0001000" when "01011000000010110", -- t[45078] = 8
      "0001000" when "01011000000010111", -- t[45079] = 8
      "0001000" when "01011000000011000", -- t[45080] = 8
      "0001000" when "01011000000011001", -- t[45081] = 8
      "0001000" when "01011000000011010", -- t[45082] = 8
      "0001000" when "01011000000011011", -- t[45083] = 8
      "0001000" when "01011000000011100", -- t[45084] = 8
      "0001000" when "01011000000011101", -- t[45085] = 8
      "0001000" when "01011000000011110", -- t[45086] = 8
      "0001000" when "01011000000011111", -- t[45087] = 8
      "0001000" when "01011000000100000", -- t[45088] = 8
      "0001000" when "01011000000100001", -- t[45089] = 8
      "0001000" when "01011000000100010", -- t[45090] = 8
      "0001000" when "01011000000100011", -- t[45091] = 8
      "0001000" when "01011000000100100", -- t[45092] = 8
      "0001000" when "01011000000100101", -- t[45093] = 8
      "0001000" when "01011000000100110", -- t[45094] = 8
      "0001000" when "01011000000100111", -- t[45095] = 8
      "0001000" when "01011000000101000", -- t[45096] = 8
      "0001000" when "01011000000101001", -- t[45097] = 8
      "0001000" when "01011000000101010", -- t[45098] = 8
      "0001000" when "01011000000101011", -- t[45099] = 8
      "0001000" when "01011000000101100", -- t[45100] = 8
      "0001000" when "01011000000101101", -- t[45101] = 8
      "0001000" when "01011000000101110", -- t[45102] = 8
      "0001000" when "01011000000101111", -- t[45103] = 8
      "0001000" when "01011000000110000", -- t[45104] = 8
      "0001000" when "01011000000110001", -- t[45105] = 8
      "0001000" when "01011000000110010", -- t[45106] = 8
      "0001000" when "01011000000110011", -- t[45107] = 8
      "0001000" when "01011000000110100", -- t[45108] = 8
      "0001000" when "01011000000110101", -- t[45109] = 8
      "0001000" when "01011000000110110", -- t[45110] = 8
      "0001000" when "01011000000110111", -- t[45111] = 8
      "0001000" when "01011000000111000", -- t[45112] = 8
      "0001000" when "01011000000111001", -- t[45113] = 8
      "0001000" when "01011000000111010", -- t[45114] = 8
      "0001000" when "01011000000111011", -- t[45115] = 8
      "0001000" when "01011000000111100", -- t[45116] = 8
      "0001000" when "01011000000111101", -- t[45117] = 8
      "0001000" when "01011000000111110", -- t[45118] = 8
      "0001000" when "01011000000111111", -- t[45119] = 8
      "0001000" when "01011000001000000", -- t[45120] = 8
      "0001000" when "01011000001000001", -- t[45121] = 8
      "0001000" when "01011000001000010", -- t[45122] = 8
      "0001000" when "01011000001000011", -- t[45123] = 8
      "0001000" when "01011000001000100", -- t[45124] = 8
      "0001000" when "01011000001000101", -- t[45125] = 8
      "0001000" when "01011000001000110", -- t[45126] = 8
      "0001000" when "01011000001000111", -- t[45127] = 8
      "0001000" when "01011000001001000", -- t[45128] = 8
      "0001000" when "01011000001001001", -- t[45129] = 8
      "0001000" when "01011000001001010", -- t[45130] = 8
      "0001000" when "01011000001001011", -- t[45131] = 8
      "0001000" when "01011000001001100", -- t[45132] = 8
      "0001000" when "01011000001001101", -- t[45133] = 8
      "0001000" when "01011000001001110", -- t[45134] = 8
      "0001000" when "01011000001001111", -- t[45135] = 8
      "0001000" when "01011000001010000", -- t[45136] = 8
      "0001000" when "01011000001010001", -- t[45137] = 8
      "0001000" when "01011000001010010", -- t[45138] = 8
      "0001000" when "01011000001010011", -- t[45139] = 8
      "0001000" when "01011000001010100", -- t[45140] = 8
      "0001000" when "01011000001010101", -- t[45141] = 8
      "0001000" when "01011000001010110", -- t[45142] = 8
      "0001000" when "01011000001010111", -- t[45143] = 8
      "0001000" when "01011000001011000", -- t[45144] = 8
      "0001000" when "01011000001011001", -- t[45145] = 8
      "0001000" when "01011000001011010", -- t[45146] = 8
      "0001000" when "01011000001011011", -- t[45147] = 8
      "0001000" when "01011000001011100", -- t[45148] = 8
      "0001000" when "01011000001011101", -- t[45149] = 8
      "0001000" when "01011000001011110", -- t[45150] = 8
      "0001000" when "01011000001011111", -- t[45151] = 8
      "0001000" when "01011000001100000", -- t[45152] = 8
      "0001000" when "01011000001100001", -- t[45153] = 8
      "0001000" when "01011000001100010", -- t[45154] = 8
      "0001000" when "01011000001100011", -- t[45155] = 8
      "0001000" when "01011000001100100", -- t[45156] = 8
      "0001000" when "01011000001100101", -- t[45157] = 8
      "0001000" when "01011000001100110", -- t[45158] = 8
      "0001000" when "01011000001100111", -- t[45159] = 8
      "0001000" when "01011000001101000", -- t[45160] = 8
      "0001000" when "01011000001101001", -- t[45161] = 8
      "0001000" when "01011000001101010", -- t[45162] = 8
      "0001000" when "01011000001101011", -- t[45163] = 8
      "0001000" when "01011000001101100", -- t[45164] = 8
      "0001000" when "01011000001101101", -- t[45165] = 8
      "0001000" when "01011000001101110", -- t[45166] = 8
      "0001000" when "01011000001101111", -- t[45167] = 8
      "0001000" when "01011000001110000", -- t[45168] = 8
      "0001000" when "01011000001110001", -- t[45169] = 8
      "0001000" when "01011000001110010", -- t[45170] = 8
      "0001000" when "01011000001110011", -- t[45171] = 8
      "0001000" when "01011000001110100", -- t[45172] = 8
      "0001000" when "01011000001110101", -- t[45173] = 8
      "0001000" when "01011000001110110", -- t[45174] = 8
      "0001000" when "01011000001110111", -- t[45175] = 8
      "0001000" when "01011000001111000", -- t[45176] = 8
      "0001000" when "01011000001111001", -- t[45177] = 8
      "0001000" when "01011000001111010", -- t[45178] = 8
      "0001000" when "01011000001111011", -- t[45179] = 8
      "0001000" when "01011000001111100", -- t[45180] = 8
      "0001000" when "01011000001111101", -- t[45181] = 8
      "0001000" when "01011000001111110", -- t[45182] = 8
      "0001000" when "01011000001111111", -- t[45183] = 8
      "0001000" when "01011000010000000", -- t[45184] = 8
      "0001000" when "01011000010000001", -- t[45185] = 8
      "0001000" when "01011000010000010", -- t[45186] = 8
      "0001000" when "01011000010000011", -- t[45187] = 8
      "0001000" when "01011000010000100", -- t[45188] = 8
      "0001000" when "01011000010000101", -- t[45189] = 8
      "0001000" when "01011000010000110", -- t[45190] = 8
      "0001000" when "01011000010000111", -- t[45191] = 8
      "0001000" when "01011000010001000", -- t[45192] = 8
      "0001000" when "01011000010001001", -- t[45193] = 8
      "0001000" when "01011000010001010", -- t[45194] = 8
      "0001000" when "01011000010001011", -- t[45195] = 8
      "0001000" when "01011000010001100", -- t[45196] = 8
      "0001000" when "01011000010001101", -- t[45197] = 8
      "0001000" when "01011000010001110", -- t[45198] = 8
      "0001000" when "01011000010001111", -- t[45199] = 8
      "0001000" when "01011000010010000", -- t[45200] = 8
      "0001000" when "01011000010010001", -- t[45201] = 8
      "0001000" when "01011000010010010", -- t[45202] = 8
      "0001000" when "01011000010010011", -- t[45203] = 8
      "0001000" when "01011000010010100", -- t[45204] = 8
      "0001000" when "01011000010010101", -- t[45205] = 8
      "0001000" when "01011000010010110", -- t[45206] = 8
      "0001000" when "01011000010010111", -- t[45207] = 8
      "0001000" when "01011000010011000", -- t[45208] = 8
      "0001000" when "01011000010011001", -- t[45209] = 8
      "0001000" when "01011000010011010", -- t[45210] = 8
      "0001000" when "01011000010011011", -- t[45211] = 8
      "0001000" when "01011000010011100", -- t[45212] = 8
      "0001000" when "01011000010011101", -- t[45213] = 8
      "0001000" when "01011000010011110", -- t[45214] = 8
      "0001000" when "01011000010011111", -- t[45215] = 8
      "0001000" when "01011000010100000", -- t[45216] = 8
      "0001000" when "01011000010100001", -- t[45217] = 8
      "0001000" when "01011000010100010", -- t[45218] = 8
      "0001000" when "01011000010100011", -- t[45219] = 8
      "0001000" when "01011000010100100", -- t[45220] = 8
      "0001000" when "01011000010100101", -- t[45221] = 8
      "0001000" when "01011000010100110", -- t[45222] = 8
      "0001000" when "01011000010100111", -- t[45223] = 8
      "0001000" when "01011000010101000", -- t[45224] = 8
      "0001000" when "01011000010101001", -- t[45225] = 8
      "0001000" when "01011000010101010", -- t[45226] = 8
      "0001000" when "01011000010101011", -- t[45227] = 8
      "0001000" when "01011000010101100", -- t[45228] = 8
      "0001000" when "01011000010101101", -- t[45229] = 8
      "0001000" when "01011000010101110", -- t[45230] = 8
      "0001000" when "01011000010101111", -- t[45231] = 8
      "0001000" when "01011000010110000", -- t[45232] = 8
      "0001000" when "01011000010110001", -- t[45233] = 8
      "0001000" when "01011000010110010", -- t[45234] = 8
      "0001000" when "01011000010110011", -- t[45235] = 8
      "0001000" when "01011000010110100", -- t[45236] = 8
      "0001000" when "01011000010110101", -- t[45237] = 8
      "0001000" when "01011000010110110", -- t[45238] = 8
      "0001000" when "01011000010110111", -- t[45239] = 8
      "0001000" when "01011000010111000", -- t[45240] = 8
      "0001000" when "01011000010111001", -- t[45241] = 8
      "0001000" when "01011000010111010", -- t[45242] = 8
      "0001000" when "01011000010111011", -- t[45243] = 8
      "0001000" when "01011000010111100", -- t[45244] = 8
      "0001000" when "01011000010111101", -- t[45245] = 8
      "0001000" when "01011000010111110", -- t[45246] = 8
      "0001000" when "01011000010111111", -- t[45247] = 8
      "0001000" when "01011000011000000", -- t[45248] = 8
      "0001000" when "01011000011000001", -- t[45249] = 8
      "0001000" when "01011000011000010", -- t[45250] = 8
      "0001000" when "01011000011000011", -- t[45251] = 8
      "0001000" when "01011000011000100", -- t[45252] = 8
      "0001000" when "01011000011000101", -- t[45253] = 8
      "0001000" when "01011000011000110", -- t[45254] = 8
      "0001000" when "01011000011000111", -- t[45255] = 8
      "0001000" when "01011000011001000", -- t[45256] = 8
      "0001000" when "01011000011001001", -- t[45257] = 8
      "0001000" when "01011000011001010", -- t[45258] = 8
      "0001000" when "01011000011001011", -- t[45259] = 8
      "0001000" when "01011000011001100", -- t[45260] = 8
      "0001000" when "01011000011001101", -- t[45261] = 8
      "0001000" when "01011000011001110", -- t[45262] = 8
      "0001000" when "01011000011001111", -- t[45263] = 8
      "0001000" when "01011000011010000", -- t[45264] = 8
      "0001000" when "01011000011010001", -- t[45265] = 8
      "0001000" when "01011000011010010", -- t[45266] = 8
      "0001000" when "01011000011010011", -- t[45267] = 8
      "0001000" when "01011000011010100", -- t[45268] = 8
      "0001000" when "01011000011010101", -- t[45269] = 8
      "0001000" when "01011000011010110", -- t[45270] = 8
      "0001000" when "01011000011010111", -- t[45271] = 8
      "0001000" when "01011000011011000", -- t[45272] = 8
      "0001000" when "01011000011011001", -- t[45273] = 8
      "0001000" when "01011000011011010", -- t[45274] = 8
      "0001000" when "01011000011011011", -- t[45275] = 8
      "0001000" when "01011000011011100", -- t[45276] = 8
      "0001000" when "01011000011011101", -- t[45277] = 8
      "0001000" when "01011000011011110", -- t[45278] = 8
      "0001000" when "01011000011011111", -- t[45279] = 8
      "0001000" when "01011000011100000", -- t[45280] = 8
      "0001000" when "01011000011100001", -- t[45281] = 8
      "0001000" when "01011000011100010", -- t[45282] = 8
      "0001000" when "01011000011100011", -- t[45283] = 8
      "0001000" when "01011000011100100", -- t[45284] = 8
      "0001000" when "01011000011100101", -- t[45285] = 8
      "0001000" when "01011000011100110", -- t[45286] = 8
      "0001000" when "01011000011100111", -- t[45287] = 8
      "0001000" when "01011000011101000", -- t[45288] = 8
      "0001000" when "01011000011101001", -- t[45289] = 8
      "0001000" when "01011000011101010", -- t[45290] = 8
      "0001000" when "01011000011101011", -- t[45291] = 8
      "0001000" when "01011000011101100", -- t[45292] = 8
      "0001000" when "01011000011101101", -- t[45293] = 8
      "0001000" when "01011000011101110", -- t[45294] = 8
      "0001000" when "01011000011101111", -- t[45295] = 8
      "0001000" when "01011000011110000", -- t[45296] = 8
      "0001000" when "01011000011110001", -- t[45297] = 8
      "0001000" when "01011000011110010", -- t[45298] = 8
      "0001000" when "01011000011110011", -- t[45299] = 8
      "0001000" when "01011000011110100", -- t[45300] = 8
      "0001000" when "01011000011110101", -- t[45301] = 8
      "0001000" when "01011000011110110", -- t[45302] = 8
      "0001000" when "01011000011110111", -- t[45303] = 8
      "0001000" when "01011000011111000", -- t[45304] = 8
      "0001000" when "01011000011111001", -- t[45305] = 8
      "0001000" when "01011000011111010", -- t[45306] = 8
      "0001000" when "01011000011111011", -- t[45307] = 8
      "0001000" when "01011000011111100", -- t[45308] = 8
      "0001000" when "01011000011111101", -- t[45309] = 8
      "0001000" when "01011000011111110", -- t[45310] = 8
      "0001000" when "01011000011111111", -- t[45311] = 8
      "0001000" when "01011000100000000", -- t[45312] = 8
      "0001000" when "01011000100000001", -- t[45313] = 8
      "0001000" when "01011000100000010", -- t[45314] = 8
      "0001000" when "01011000100000011", -- t[45315] = 8
      "0001000" when "01011000100000100", -- t[45316] = 8
      "0001000" when "01011000100000101", -- t[45317] = 8
      "0001000" when "01011000100000110", -- t[45318] = 8
      "0001000" when "01011000100000111", -- t[45319] = 8
      "0001000" when "01011000100001000", -- t[45320] = 8
      "0001000" when "01011000100001001", -- t[45321] = 8
      "0001000" when "01011000100001010", -- t[45322] = 8
      "0001000" when "01011000100001011", -- t[45323] = 8
      "0001000" when "01011000100001100", -- t[45324] = 8
      "0001000" when "01011000100001101", -- t[45325] = 8
      "0001000" when "01011000100001110", -- t[45326] = 8
      "0001000" when "01011000100001111", -- t[45327] = 8
      "0001000" when "01011000100010000", -- t[45328] = 8
      "0001000" when "01011000100010001", -- t[45329] = 8
      "0001000" when "01011000100010010", -- t[45330] = 8
      "0001000" when "01011000100010011", -- t[45331] = 8
      "0001000" when "01011000100010100", -- t[45332] = 8
      "0001000" when "01011000100010101", -- t[45333] = 8
      "0001000" when "01011000100010110", -- t[45334] = 8
      "0001000" when "01011000100010111", -- t[45335] = 8
      "0001000" when "01011000100011000", -- t[45336] = 8
      "0001000" when "01011000100011001", -- t[45337] = 8
      "0001000" when "01011000100011010", -- t[45338] = 8
      "0001000" when "01011000100011011", -- t[45339] = 8
      "0001000" when "01011000100011100", -- t[45340] = 8
      "0001000" when "01011000100011101", -- t[45341] = 8
      "0001000" when "01011000100011110", -- t[45342] = 8
      "0001000" when "01011000100011111", -- t[45343] = 8
      "0001000" when "01011000100100000", -- t[45344] = 8
      "0001000" when "01011000100100001", -- t[45345] = 8
      "0001000" when "01011000100100010", -- t[45346] = 8
      "0001000" when "01011000100100011", -- t[45347] = 8
      "0001000" when "01011000100100100", -- t[45348] = 8
      "0001000" when "01011000100100101", -- t[45349] = 8
      "0001000" when "01011000100100110", -- t[45350] = 8
      "0001000" when "01011000100100111", -- t[45351] = 8
      "0001000" when "01011000100101000", -- t[45352] = 8
      "0001000" when "01011000100101001", -- t[45353] = 8
      "0001000" when "01011000100101010", -- t[45354] = 8
      "0001000" when "01011000100101011", -- t[45355] = 8
      "0001000" when "01011000100101100", -- t[45356] = 8
      "0001000" when "01011000100101101", -- t[45357] = 8
      "0001000" when "01011000100101110", -- t[45358] = 8
      "0001000" when "01011000100101111", -- t[45359] = 8
      "0001000" when "01011000100110000", -- t[45360] = 8
      "0001000" when "01011000100110001", -- t[45361] = 8
      "0001000" when "01011000100110010", -- t[45362] = 8
      "0001000" when "01011000100110011", -- t[45363] = 8
      "0001000" when "01011000100110100", -- t[45364] = 8
      "0001000" when "01011000100110101", -- t[45365] = 8
      "0001000" when "01011000100110110", -- t[45366] = 8
      "0001000" when "01011000100110111", -- t[45367] = 8
      "0001000" when "01011000100111000", -- t[45368] = 8
      "0001000" when "01011000100111001", -- t[45369] = 8
      "0001000" when "01011000100111010", -- t[45370] = 8
      "0001000" when "01011000100111011", -- t[45371] = 8
      "0001000" when "01011000100111100", -- t[45372] = 8
      "0001000" when "01011000100111101", -- t[45373] = 8
      "0001000" when "01011000100111110", -- t[45374] = 8
      "0001000" when "01011000100111111", -- t[45375] = 8
      "0001000" when "01011000101000000", -- t[45376] = 8
      "0001000" when "01011000101000001", -- t[45377] = 8
      "0001000" when "01011000101000010", -- t[45378] = 8
      "0001000" when "01011000101000011", -- t[45379] = 8
      "0001000" when "01011000101000100", -- t[45380] = 8
      "0001000" when "01011000101000101", -- t[45381] = 8
      "0001000" when "01011000101000110", -- t[45382] = 8
      "0001000" when "01011000101000111", -- t[45383] = 8
      "0001000" when "01011000101001000", -- t[45384] = 8
      "0001000" when "01011000101001001", -- t[45385] = 8
      "0001000" when "01011000101001010", -- t[45386] = 8
      "0001000" when "01011000101001011", -- t[45387] = 8
      "0001000" when "01011000101001100", -- t[45388] = 8
      "0001000" when "01011000101001101", -- t[45389] = 8
      "0001000" when "01011000101001110", -- t[45390] = 8
      "0001000" when "01011000101001111", -- t[45391] = 8
      "0001000" when "01011000101010000", -- t[45392] = 8
      "0001000" when "01011000101010001", -- t[45393] = 8
      "0001000" when "01011000101010010", -- t[45394] = 8
      "0001000" when "01011000101010011", -- t[45395] = 8
      "0001000" when "01011000101010100", -- t[45396] = 8
      "0001000" when "01011000101010101", -- t[45397] = 8
      "0001000" when "01011000101010110", -- t[45398] = 8
      "0001000" when "01011000101010111", -- t[45399] = 8
      "0001000" when "01011000101011000", -- t[45400] = 8
      "0001000" when "01011000101011001", -- t[45401] = 8
      "0001000" when "01011000101011010", -- t[45402] = 8
      "0001000" when "01011000101011011", -- t[45403] = 8
      "0001000" when "01011000101011100", -- t[45404] = 8
      "0001000" when "01011000101011101", -- t[45405] = 8
      "0001000" when "01011000101011110", -- t[45406] = 8
      "0001000" when "01011000101011111", -- t[45407] = 8
      "0001000" when "01011000101100000", -- t[45408] = 8
      "0001000" when "01011000101100001", -- t[45409] = 8
      "0001000" when "01011000101100010", -- t[45410] = 8
      "0001000" when "01011000101100011", -- t[45411] = 8
      "0001000" when "01011000101100100", -- t[45412] = 8
      "0001000" when "01011000101100101", -- t[45413] = 8
      "0001000" when "01011000101100110", -- t[45414] = 8
      "0001000" when "01011000101100111", -- t[45415] = 8
      "0001000" when "01011000101101000", -- t[45416] = 8
      "0001000" when "01011000101101001", -- t[45417] = 8
      "0001000" when "01011000101101010", -- t[45418] = 8
      "0001000" when "01011000101101011", -- t[45419] = 8
      "0001000" when "01011000101101100", -- t[45420] = 8
      "0001000" when "01011000101101101", -- t[45421] = 8
      "0001000" when "01011000101101110", -- t[45422] = 8
      "0001000" when "01011000101101111", -- t[45423] = 8
      "0001000" when "01011000101110000", -- t[45424] = 8
      "0001000" when "01011000101110001", -- t[45425] = 8
      "0001000" when "01011000101110010", -- t[45426] = 8
      "0001000" when "01011000101110011", -- t[45427] = 8
      "0001000" when "01011000101110100", -- t[45428] = 8
      "0001000" when "01011000101110101", -- t[45429] = 8
      "0001000" when "01011000101110110", -- t[45430] = 8
      "0001000" when "01011000101110111", -- t[45431] = 8
      "0001000" when "01011000101111000", -- t[45432] = 8
      "0001000" when "01011000101111001", -- t[45433] = 8
      "0001000" when "01011000101111010", -- t[45434] = 8
      "0001000" when "01011000101111011", -- t[45435] = 8
      "0001000" when "01011000101111100", -- t[45436] = 8
      "0001000" when "01011000101111101", -- t[45437] = 8
      "0001000" when "01011000101111110", -- t[45438] = 8
      "0001000" when "01011000101111111", -- t[45439] = 8
      "0001000" when "01011000110000000", -- t[45440] = 8
      "0001000" when "01011000110000001", -- t[45441] = 8
      "0001000" when "01011000110000010", -- t[45442] = 8
      "0001000" when "01011000110000011", -- t[45443] = 8
      "0001000" when "01011000110000100", -- t[45444] = 8
      "0001000" when "01011000110000101", -- t[45445] = 8
      "0001000" when "01011000110000110", -- t[45446] = 8
      "0001000" when "01011000110000111", -- t[45447] = 8
      "0001000" when "01011000110001000", -- t[45448] = 8
      "0001000" when "01011000110001001", -- t[45449] = 8
      "0001000" when "01011000110001010", -- t[45450] = 8
      "0001000" when "01011000110001011", -- t[45451] = 8
      "0001000" when "01011000110001100", -- t[45452] = 8
      "0001000" when "01011000110001101", -- t[45453] = 8
      "0001000" when "01011000110001110", -- t[45454] = 8
      "0001000" when "01011000110001111", -- t[45455] = 8
      "0001000" when "01011000110010000", -- t[45456] = 8
      "0001000" when "01011000110010001", -- t[45457] = 8
      "0001000" when "01011000110010010", -- t[45458] = 8
      "0001000" when "01011000110010011", -- t[45459] = 8
      "0001000" when "01011000110010100", -- t[45460] = 8
      "0001000" when "01011000110010101", -- t[45461] = 8
      "0001000" when "01011000110010110", -- t[45462] = 8
      "0001000" when "01011000110010111", -- t[45463] = 8
      "0001000" when "01011000110011000", -- t[45464] = 8
      "0001000" when "01011000110011001", -- t[45465] = 8
      "0001000" when "01011000110011010", -- t[45466] = 8
      "0001000" when "01011000110011011", -- t[45467] = 8
      "0001000" when "01011000110011100", -- t[45468] = 8
      "0001000" when "01011000110011101", -- t[45469] = 8
      "0001000" when "01011000110011110", -- t[45470] = 8
      "0001000" when "01011000110011111", -- t[45471] = 8
      "0001000" when "01011000110100000", -- t[45472] = 8
      "0001000" when "01011000110100001", -- t[45473] = 8
      "0001000" when "01011000110100010", -- t[45474] = 8
      "0001000" when "01011000110100011", -- t[45475] = 8
      "0001000" when "01011000110100100", -- t[45476] = 8
      "0001000" when "01011000110100101", -- t[45477] = 8
      "0001000" when "01011000110100110", -- t[45478] = 8
      "0001000" when "01011000110100111", -- t[45479] = 8
      "0001000" when "01011000110101000", -- t[45480] = 8
      "0001000" when "01011000110101001", -- t[45481] = 8
      "0001000" when "01011000110101010", -- t[45482] = 8
      "0001000" when "01011000110101011", -- t[45483] = 8
      "0001000" when "01011000110101100", -- t[45484] = 8
      "0001000" when "01011000110101101", -- t[45485] = 8
      "0001000" when "01011000110101110", -- t[45486] = 8
      "0001000" when "01011000110101111", -- t[45487] = 8
      "0001000" when "01011000110110000", -- t[45488] = 8
      "0001000" when "01011000110110001", -- t[45489] = 8
      "0001000" when "01011000110110010", -- t[45490] = 8
      "0001000" when "01011000110110011", -- t[45491] = 8
      "0001000" when "01011000110110100", -- t[45492] = 8
      "0001000" when "01011000110110101", -- t[45493] = 8
      "0001000" when "01011000110110110", -- t[45494] = 8
      "0001000" when "01011000110110111", -- t[45495] = 8
      "0001000" when "01011000110111000", -- t[45496] = 8
      "0001000" when "01011000110111001", -- t[45497] = 8
      "0001000" when "01011000110111010", -- t[45498] = 8
      "0001000" when "01011000110111011", -- t[45499] = 8
      "0001000" when "01011000110111100", -- t[45500] = 8
      "0001000" when "01011000110111101", -- t[45501] = 8
      "0001000" when "01011000110111110", -- t[45502] = 8
      "0001000" when "01011000110111111", -- t[45503] = 8
      "0001000" when "01011000111000000", -- t[45504] = 8
      "0001000" when "01011000111000001", -- t[45505] = 8
      "0001000" when "01011000111000010", -- t[45506] = 8
      "0001000" when "01011000111000011", -- t[45507] = 8
      "0001000" when "01011000111000100", -- t[45508] = 8
      "0001000" when "01011000111000101", -- t[45509] = 8
      "0001000" when "01011000111000110", -- t[45510] = 8
      "0001000" when "01011000111000111", -- t[45511] = 8
      "0001000" when "01011000111001000", -- t[45512] = 8
      "0001000" when "01011000111001001", -- t[45513] = 8
      "0001000" when "01011000111001010", -- t[45514] = 8
      "0001000" when "01011000111001011", -- t[45515] = 8
      "0001000" when "01011000111001100", -- t[45516] = 8
      "0001000" when "01011000111001101", -- t[45517] = 8
      "0001000" when "01011000111001110", -- t[45518] = 8
      "0001000" when "01011000111001111", -- t[45519] = 8
      "0001000" when "01011000111010000", -- t[45520] = 8
      "0001000" when "01011000111010001", -- t[45521] = 8
      "0001000" when "01011000111010010", -- t[45522] = 8
      "0001000" when "01011000111010011", -- t[45523] = 8
      "0001000" when "01011000111010100", -- t[45524] = 8
      "0001000" when "01011000111010101", -- t[45525] = 8
      "0001000" when "01011000111010110", -- t[45526] = 8
      "0001000" when "01011000111010111", -- t[45527] = 8
      "0001000" when "01011000111011000", -- t[45528] = 8
      "0001000" when "01011000111011001", -- t[45529] = 8
      "0001000" when "01011000111011010", -- t[45530] = 8
      "0001000" when "01011000111011011", -- t[45531] = 8
      "0001000" when "01011000111011100", -- t[45532] = 8
      "0001001" when "01011000111011101", -- t[45533] = 9
      "0001001" when "01011000111011110", -- t[45534] = 9
      "0001001" when "01011000111011111", -- t[45535] = 9
      "0001001" when "01011000111100000", -- t[45536] = 9
      "0001001" when "01011000111100001", -- t[45537] = 9
      "0001001" when "01011000111100010", -- t[45538] = 9
      "0001001" when "01011000111100011", -- t[45539] = 9
      "0001001" when "01011000111100100", -- t[45540] = 9
      "0001001" when "01011000111100101", -- t[45541] = 9
      "0001001" when "01011000111100110", -- t[45542] = 9
      "0001001" when "01011000111100111", -- t[45543] = 9
      "0001001" when "01011000111101000", -- t[45544] = 9
      "0001001" when "01011000111101001", -- t[45545] = 9
      "0001001" when "01011000111101010", -- t[45546] = 9
      "0001001" when "01011000111101011", -- t[45547] = 9
      "0001001" when "01011000111101100", -- t[45548] = 9
      "0001001" when "01011000111101101", -- t[45549] = 9
      "0001001" when "01011000111101110", -- t[45550] = 9
      "0001001" when "01011000111101111", -- t[45551] = 9
      "0001001" when "01011000111110000", -- t[45552] = 9
      "0001001" when "01011000111110001", -- t[45553] = 9
      "0001001" when "01011000111110010", -- t[45554] = 9
      "0001001" when "01011000111110011", -- t[45555] = 9
      "0001001" when "01011000111110100", -- t[45556] = 9
      "0001001" when "01011000111110101", -- t[45557] = 9
      "0001001" when "01011000111110110", -- t[45558] = 9
      "0001001" when "01011000111110111", -- t[45559] = 9
      "0001001" when "01011000111111000", -- t[45560] = 9
      "0001001" when "01011000111111001", -- t[45561] = 9
      "0001001" when "01011000111111010", -- t[45562] = 9
      "0001001" when "01011000111111011", -- t[45563] = 9
      "0001001" when "01011000111111100", -- t[45564] = 9
      "0001001" when "01011000111111101", -- t[45565] = 9
      "0001001" when "01011000111111110", -- t[45566] = 9
      "0001001" when "01011000111111111", -- t[45567] = 9
      "0001001" when "01011001000000000", -- t[45568] = 9
      "0001001" when "01011001000000001", -- t[45569] = 9
      "0001001" when "01011001000000010", -- t[45570] = 9
      "0001001" when "01011001000000011", -- t[45571] = 9
      "0001001" when "01011001000000100", -- t[45572] = 9
      "0001001" when "01011001000000101", -- t[45573] = 9
      "0001001" when "01011001000000110", -- t[45574] = 9
      "0001001" when "01011001000000111", -- t[45575] = 9
      "0001001" when "01011001000001000", -- t[45576] = 9
      "0001001" when "01011001000001001", -- t[45577] = 9
      "0001001" when "01011001000001010", -- t[45578] = 9
      "0001001" when "01011001000001011", -- t[45579] = 9
      "0001001" when "01011001000001100", -- t[45580] = 9
      "0001001" when "01011001000001101", -- t[45581] = 9
      "0001001" when "01011001000001110", -- t[45582] = 9
      "0001001" when "01011001000001111", -- t[45583] = 9
      "0001001" when "01011001000010000", -- t[45584] = 9
      "0001001" when "01011001000010001", -- t[45585] = 9
      "0001001" when "01011001000010010", -- t[45586] = 9
      "0001001" when "01011001000010011", -- t[45587] = 9
      "0001001" when "01011001000010100", -- t[45588] = 9
      "0001001" when "01011001000010101", -- t[45589] = 9
      "0001001" when "01011001000010110", -- t[45590] = 9
      "0001001" when "01011001000010111", -- t[45591] = 9
      "0001001" when "01011001000011000", -- t[45592] = 9
      "0001001" when "01011001000011001", -- t[45593] = 9
      "0001001" when "01011001000011010", -- t[45594] = 9
      "0001001" when "01011001000011011", -- t[45595] = 9
      "0001001" when "01011001000011100", -- t[45596] = 9
      "0001001" when "01011001000011101", -- t[45597] = 9
      "0001001" when "01011001000011110", -- t[45598] = 9
      "0001001" when "01011001000011111", -- t[45599] = 9
      "0001001" when "01011001000100000", -- t[45600] = 9
      "0001001" when "01011001000100001", -- t[45601] = 9
      "0001001" when "01011001000100010", -- t[45602] = 9
      "0001001" when "01011001000100011", -- t[45603] = 9
      "0001001" when "01011001000100100", -- t[45604] = 9
      "0001001" when "01011001000100101", -- t[45605] = 9
      "0001001" when "01011001000100110", -- t[45606] = 9
      "0001001" when "01011001000100111", -- t[45607] = 9
      "0001001" when "01011001000101000", -- t[45608] = 9
      "0001001" when "01011001000101001", -- t[45609] = 9
      "0001001" when "01011001000101010", -- t[45610] = 9
      "0001001" when "01011001000101011", -- t[45611] = 9
      "0001001" when "01011001000101100", -- t[45612] = 9
      "0001001" when "01011001000101101", -- t[45613] = 9
      "0001001" when "01011001000101110", -- t[45614] = 9
      "0001001" when "01011001000101111", -- t[45615] = 9
      "0001001" when "01011001000110000", -- t[45616] = 9
      "0001001" when "01011001000110001", -- t[45617] = 9
      "0001001" when "01011001000110010", -- t[45618] = 9
      "0001001" when "01011001000110011", -- t[45619] = 9
      "0001001" when "01011001000110100", -- t[45620] = 9
      "0001001" when "01011001000110101", -- t[45621] = 9
      "0001001" when "01011001000110110", -- t[45622] = 9
      "0001001" when "01011001000110111", -- t[45623] = 9
      "0001001" when "01011001000111000", -- t[45624] = 9
      "0001001" when "01011001000111001", -- t[45625] = 9
      "0001001" when "01011001000111010", -- t[45626] = 9
      "0001001" when "01011001000111011", -- t[45627] = 9
      "0001001" when "01011001000111100", -- t[45628] = 9
      "0001001" when "01011001000111101", -- t[45629] = 9
      "0001001" when "01011001000111110", -- t[45630] = 9
      "0001001" when "01011001000111111", -- t[45631] = 9
      "0001001" when "01011001001000000", -- t[45632] = 9
      "0001001" when "01011001001000001", -- t[45633] = 9
      "0001001" when "01011001001000010", -- t[45634] = 9
      "0001001" when "01011001001000011", -- t[45635] = 9
      "0001001" when "01011001001000100", -- t[45636] = 9
      "0001001" when "01011001001000101", -- t[45637] = 9
      "0001001" when "01011001001000110", -- t[45638] = 9
      "0001001" when "01011001001000111", -- t[45639] = 9
      "0001001" when "01011001001001000", -- t[45640] = 9
      "0001001" when "01011001001001001", -- t[45641] = 9
      "0001001" when "01011001001001010", -- t[45642] = 9
      "0001001" when "01011001001001011", -- t[45643] = 9
      "0001001" when "01011001001001100", -- t[45644] = 9
      "0001001" when "01011001001001101", -- t[45645] = 9
      "0001001" when "01011001001001110", -- t[45646] = 9
      "0001001" when "01011001001001111", -- t[45647] = 9
      "0001001" when "01011001001010000", -- t[45648] = 9
      "0001001" when "01011001001010001", -- t[45649] = 9
      "0001001" when "01011001001010010", -- t[45650] = 9
      "0001001" when "01011001001010011", -- t[45651] = 9
      "0001001" when "01011001001010100", -- t[45652] = 9
      "0001001" when "01011001001010101", -- t[45653] = 9
      "0001001" when "01011001001010110", -- t[45654] = 9
      "0001001" when "01011001001010111", -- t[45655] = 9
      "0001001" when "01011001001011000", -- t[45656] = 9
      "0001001" when "01011001001011001", -- t[45657] = 9
      "0001001" when "01011001001011010", -- t[45658] = 9
      "0001001" when "01011001001011011", -- t[45659] = 9
      "0001001" when "01011001001011100", -- t[45660] = 9
      "0001001" when "01011001001011101", -- t[45661] = 9
      "0001001" when "01011001001011110", -- t[45662] = 9
      "0001001" when "01011001001011111", -- t[45663] = 9
      "0001001" when "01011001001100000", -- t[45664] = 9
      "0001001" when "01011001001100001", -- t[45665] = 9
      "0001001" when "01011001001100010", -- t[45666] = 9
      "0001001" when "01011001001100011", -- t[45667] = 9
      "0001001" when "01011001001100100", -- t[45668] = 9
      "0001001" when "01011001001100101", -- t[45669] = 9
      "0001001" when "01011001001100110", -- t[45670] = 9
      "0001001" when "01011001001100111", -- t[45671] = 9
      "0001001" when "01011001001101000", -- t[45672] = 9
      "0001001" when "01011001001101001", -- t[45673] = 9
      "0001001" when "01011001001101010", -- t[45674] = 9
      "0001001" when "01011001001101011", -- t[45675] = 9
      "0001001" when "01011001001101100", -- t[45676] = 9
      "0001001" when "01011001001101101", -- t[45677] = 9
      "0001001" when "01011001001101110", -- t[45678] = 9
      "0001001" when "01011001001101111", -- t[45679] = 9
      "0001001" when "01011001001110000", -- t[45680] = 9
      "0001001" when "01011001001110001", -- t[45681] = 9
      "0001001" when "01011001001110010", -- t[45682] = 9
      "0001001" when "01011001001110011", -- t[45683] = 9
      "0001001" when "01011001001110100", -- t[45684] = 9
      "0001001" when "01011001001110101", -- t[45685] = 9
      "0001001" when "01011001001110110", -- t[45686] = 9
      "0001001" when "01011001001110111", -- t[45687] = 9
      "0001001" when "01011001001111000", -- t[45688] = 9
      "0001001" when "01011001001111001", -- t[45689] = 9
      "0001001" when "01011001001111010", -- t[45690] = 9
      "0001001" when "01011001001111011", -- t[45691] = 9
      "0001001" when "01011001001111100", -- t[45692] = 9
      "0001001" when "01011001001111101", -- t[45693] = 9
      "0001001" when "01011001001111110", -- t[45694] = 9
      "0001001" when "01011001001111111", -- t[45695] = 9
      "0001001" when "01011001010000000", -- t[45696] = 9
      "0001001" when "01011001010000001", -- t[45697] = 9
      "0001001" when "01011001010000010", -- t[45698] = 9
      "0001001" when "01011001010000011", -- t[45699] = 9
      "0001001" when "01011001010000100", -- t[45700] = 9
      "0001001" when "01011001010000101", -- t[45701] = 9
      "0001001" when "01011001010000110", -- t[45702] = 9
      "0001001" when "01011001010000111", -- t[45703] = 9
      "0001001" when "01011001010001000", -- t[45704] = 9
      "0001001" when "01011001010001001", -- t[45705] = 9
      "0001001" when "01011001010001010", -- t[45706] = 9
      "0001001" when "01011001010001011", -- t[45707] = 9
      "0001001" when "01011001010001100", -- t[45708] = 9
      "0001001" when "01011001010001101", -- t[45709] = 9
      "0001001" when "01011001010001110", -- t[45710] = 9
      "0001001" when "01011001010001111", -- t[45711] = 9
      "0001001" when "01011001010010000", -- t[45712] = 9
      "0001001" when "01011001010010001", -- t[45713] = 9
      "0001001" when "01011001010010010", -- t[45714] = 9
      "0001001" when "01011001010010011", -- t[45715] = 9
      "0001001" when "01011001010010100", -- t[45716] = 9
      "0001001" when "01011001010010101", -- t[45717] = 9
      "0001001" when "01011001010010110", -- t[45718] = 9
      "0001001" when "01011001010010111", -- t[45719] = 9
      "0001001" when "01011001010011000", -- t[45720] = 9
      "0001001" when "01011001010011001", -- t[45721] = 9
      "0001001" when "01011001010011010", -- t[45722] = 9
      "0001001" when "01011001010011011", -- t[45723] = 9
      "0001001" when "01011001010011100", -- t[45724] = 9
      "0001001" when "01011001010011101", -- t[45725] = 9
      "0001001" when "01011001010011110", -- t[45726] = 9
      "0001001" when "01011001010011111", -- t[45727] = 9
      "0001001" when "01011001010100000", -- t[45728] = 9
      "0001001" when "01011001010100001", -- t[45729] = 9
      "0001001" when "01011001010100010", -- t[45730] = 9
      "0001001" when "01011001010100011", -- t[45731] = 9
      "0001001" when "01011001010100100", -- t[45732] = 9
      "0001001" when "01011001010100101", -- t[45733] = 9
      "0001001" when "01011001010100110", -- t[45734] = 9
      "0001001" when "01011001010100111", -- t[45735] = 9
      "0001001" when "01011001010101000", -- t[45736] = 9
      "0001001" when "01011001010101001", -- t[45737] = 9
      "0001001" when "01011001010101010", -- t[45738] = 9
      "0001001" when "01011001010101011", -- t[45739] = 9
      "0001001" when "01011001010101100", -- t[45740] = 9
      "0001001" when "01011001010101101", -- t[45741] = 9
      "0001001" when "01011001010101110", -- t[45742] = 9
      "0001001" when "01011001010101111", -- t[45743] = 9
      "0001001" when "01011001010110000", -- t[45744] = 9
      "0001001" when "01011001010110001", -- t[45745] = 9
      "0001001" when "01011001010110010", -- t[45746] = 9
      "0001001" when "01011001010110011", -- t[45747] = 9
      "0001001" when "01011001010110100", -- t[45748] = 9
      "0001001" when "01011001010110101", -- t[45749] = 9
      "0001001" when "01011001010110110", -- t[45750] = 9
      "0001001" when "01011001010110111", -- t[45751] = 9
      "0001001" when "01011001010111000", -- t[45752] = 9
      "0001001" when "01011001010111001", -- t[45753] = 9
      "0001001" when "01011001010111010", -- t[45754] = 9
      "0001001" when "01011001010111011", -- t[45755] = 9
      "0001001" when "01011001010111100", -- t[45756] = 9
      "0001001" when "01011001010111101", -- t[45757] = 9
      "0001001" when "01011001010111110", -- t[45758] = 9
      "0001001" when "01011001010111111", -- t[45759] = 9
      "0001001" when "01011001011000000", -- t[45760] = 9
      "0001001" when "01011001011000001", -- t[45761] = 9
      "0001001" when "01011001011000010", -- t[45762] = 9
      "0001001" when "01011001011000011", -- t[45763] = 9
      "0001001" when "01011001011000100", -- t[45764] = 9
      "0001001" when "01011001011000101", -- t[45765] = 9
      "0001001" when "01011001011000110", -- t[45766] = 9
      "0001001" when "01011001011000111", -- t[45767] = 9
      "0001001" when "01011001011001000", -- t[45768] = 9
      "0001001" when "01011001011001001", -- t[45769] = 9
      "0001001" when "01011001011001010", -- t[45770] = 9
      "0001001" when "01011001011001011", -- t[45771] = 9
      "0001001" when "01011001011001100", -- t[45772] = 9
      "0001001" when "01011001011001101", -- t[45773] = 9
      "0001001" when "01011001011001110", -- t[45774] = 9
      "0001001" when "01011001011001111", -- t[45775] = 9
      "0001001" when "01011001011010000", -- t[45776] = 9
      "0001001" when "01011001011010001", -- t[45777] = 9
      "0001001" when "01011001011010010", -- t[45778] = 9
      "0001001" when "01011001011010011", -- t[45779] = 9
      "0001001" when "01011001011010100", -- t[45780] = 9
      "0001001" when "01011001011010101", -- t[45781] = 9
      "0001001" when "01011001011010110", -- t[45782] = 9
      "0001001" when "01011001011010111", -- t[45783] = 9
      "0001001" when "01011001011011000", -- t[45784] = 9
      "0001001" when "01011001011011001", -- t[45785] = 9
      "0001001" when "01011001011011010", -- t[45786] = 9
      "0001001" when "01011001011011011", -- t[45787] = 9
      "0001001" when "01011001011011100", -- t[45788] = 9
      "0001001" when "01011001011011101", -- t[45789] = 9
      "0001001" when "01011001011011110", -- t[45790] = 9
      "0001001" when "01011001011011111", -- t[45791] = 9
      "0001001" when "01011001011100000", -- t[45792] = 9
      "0001001" when "01011001011100001", -- t[45793] = 9
      "0001001" when "01011001011100010", -- t[45794] = 9
      "0001001" when "01011001011100011", -- t[45795] = 9
      "0001001" when "01011001011100100", -- t[45796] = 9
      "0001001" when "01011001011100101", -- t[45797] = 9
      "0001001" when "01011001011100110", -- t[45798] = 9
      "0001001" when "01011001011100111", -- t[45799] = 9
      "0001001" when "01011001011101000", -- t[45800] = 9
      "0001001" when "01011001011101001", -- t[45801] = 9
      "0001001" when "01011001011101010", -- t[45802] = 9
      "0001001" when "01011001011101011", -- t[45803] = 9
      "0001001" when "01011001011101100", -- t[45804] = 9
      "0001001" when "01011001011101101", -- t[45805] = 9
      "0001001" when "01011001011101110", -- t[45806] = 9
      "0001001" when "01011001011101111", -- t[45807] = 9
      "0001001" when "01011001011110000", -- t[45808] = 9
      "0001001" when "01011001011110001", -- t[45809] = 9
      "0001001" when "01011001011110010", -- t[45810] = 9
      "0001001" when "01011001011110011", -- t[45811] = 9
      "0001001" when "01011001011110100", -- t[45812] = 9
      "0001001" when "01011001011110101", -- t[45813] = 9
      "0001001" when "01011001011110110", -- t[45814] = 9
      "0001001" when "01011001011110111", -- t[45815] = 9
      "0001001" when "01011001011111000", -- t[45816] = 9
      "0001001" when "01011001011111001", -- t[45817] = 9
      "0001001" when "01011001011111010", -- t[45818] = 9
      "0001001" when "01011001011111011", -- t[45819] = 9
      "0001001" when "01011001011111100", -- t[45820] = 9
      "0001001" when "01011001011111101", -- t[45821] = 9
      "0001001" when "01011001011111110", -- t[45822] = 9
      "0001001" when "01011001011111111", -- t[45823] = 9
      "0001001" when "01011001100000000", -- t[45824] = 9
      "0001001" when "01011001100000001", -- t[45825] = 9
      "0001001" when "01011001100000010", -- t[45826] = 9
      "0001001" when "01011001100000011", -- t[45827] = 9
      "0001001" when "01011001100000100", -- t[45828] = 9
      "0001001" when "01011001100000101", -- t[45829] = 9
      "0001001" when "01011001100000110", -- t[45830] = 9
      "0001001" when "01011001100000111", -- t[45831] = 9
      "0001001" when "01011001100001000", -- t[45832] = 9
      "0001001" when "01011001100001001", -- t[45833] = 9
      "0001001" when "01011001100001010", -- t[45834] = 9
      "0001001" when "01011001100001011", -- t[45835] = 9
      "0001001" when "01011001100001100", -- t[45836] = 9
      "0001001" when "01011001100001101", -- t[45837] = 9
      "0001001" when "01011001100001110", -- t[45838] = 9
      "0001001" when "01011001100001111", -- t[45839] = 9
      "0001001" when "01011001100010000", -- t[45840] = 9
      "0001001" when "01011001100010001", -- t[45841] = 9
      "0001001" when "01011001100010010", -- t[45842] = 9
      "0001001" when "01011001100010011", -- t[45843] = 9
      "0001001" when "01011001100010100", -- t[45844] = 9
      "0001001" when "01011001100010101", -- t[45845] = 9
      "0001001" when "01011001100010110", -- t[45846] = 9
      "0001001" when "01011001100010111", -- t[45847] = 9
      "0001001" when "01011001100011000", -- t[45848] = 9
      "0001001" when "01011001100011001", -- t[45849] = 9
      "0001001" when "01011001100011010", -- t[45850] = 9
      "0001001" when "01011001100011011", -- t[45851] = 9
      "0001001" when "01011001100011100", -- t[45852] = 9
      "0001001" when "01011001100011101", -- t[45853] = 9
      "0001001" when "01011001100011110", -- t[45854] = 9
      "0001001" when "01011001100011111", -- t[45855] = 9
      "0001001" when "01011001100100000", -- t[45856] = 9
      "0001001" when "01011001100100001", -- t[45857] = 9
      "0001001" when "01011001100100010", -- t[45858] = 9
      "0001001" when "01011001100100011", -- t[45859] = 9
      "0001001" when "01011001100100100", -- t[45860] = 9
      "0001001" when "01011001100100101", -- t[45861] = 9
      "0001001" when "01011001100100110", -- t[45862] = 9
      "0001001" when "01011001100100111", -- t[45863] = 9
      "0001001" when "01011001100101000", -- t[45864] = 9
      "0001001" when "01011001100101001", -- t[45865] = 9
      "0001001" when "01011001100101010", -- t[45866] = 9
      "0001001" when "01011001100101011", -- t[45867] = 9
      "0001001" when "01011001100101100", -- t[45868] = 9
      "0001001" when "01011001100101101", -- t[45869] = 9
      "0001001" when "01011001100101110", -- t[45870] = 9
      "0001001" when "01011001100101111", -- t[45871] = 9
      "0001001" when "01011001100110000", -- t[45872] = 9
      "0001001" when "01011001100110001", -- t[45873] = 9
      "0001001" when "01011001100110010", -- t[45874] = 9
      "0001001" when "01011001100110011", -- t[45875] = 9
      "0001001" when "01011001100110100", -- t[45876] = 9
      "0001001" when "01011001100110101", -- t[45877] = 9
      "0001001" when "01011001100110110", -- t[45878] = 9
      "0001001" when "01011001100110111", -- t[45879] = 9
      "0001001" when "01011001100111000", -- t[45880] = 9
      "0001001" when "01011001100111001", -- t[45881] = 9
      "0001001" when "01011001100111010", -- t[45882] = 9
      "0001001" when "01011001100111011", -- t[45883] = 9
      "0001001" when "01011001100111100", -- t[45884] = 9
      "0001001" when "01011001100111101", -- t[45885] = 9
      "0001001" when "01011001100111110", -- t[45886] = 9
      "0001001" when "01011001100111111", -- t[45887] = 9
      "0001001" when "01011001101000000", -- t[45888] = 9
      "0001001" when "01011001101000001", -- t[45889] = 9
      "0001001" when "01011001101000010", -- t[45890] = 9
      "0001001" when "01011001101000011", -- t[45891] = 9
      "0001001" when "01011001101000100", -- t[45892] = 9
      "0001001" when "01011001101000101", -- t[45893] = 9
      "0001001" when "01011001101000110", -- t[45894] = 9
      "0001001" when "01011001101000111", -- t[45895] = 9
      "0001001" when "01011001101001000", -- t[45896] = 9
      "0001001" when "01011001101001001", -- t[45897] = 9
      "0001001" when "01011001101001010", -- t[45898] = 9
      "0001001" when "01011001101001011", -- t[45899] = 9
      "0001001" when "01011001101001100", -- t[45900] = 9
      "0001001" when "01011001101001101", -- t[45901] = 9
      "0001001" when "01011001101001110", -- t[45902] = 9
      "0001001" when "01011001101001111", -- t[45903] = 9
      "0001001" when "01011001101010000", -- t[45904] = 9
      "0001001" when "01011001101010001", -- t[45905] = 9
      "0001001" when "01011001101010010", -- t[45906] = 9
      "0001001" when "01011001101010011", -- t[45907] = 9
      "0001001" when "01011001101010100", -- t[45908] = 9
      "0001001" when "01011001101010101", -- t[45909] = 9
      "0001001" when "01011001101010110", -- t[45910] = 9
      "0001001" when "01011001101010111", -- t[45911] = 9
      "0001001" when "01011001101011000", -- t[45912] = 9
      "0001001" when "01011001101011001", -- t[45913] = 9
      "0001001" when "01011001101011010", -- t[45914] = 9
      "0001001" when "01011001101011011", -- t[45915] = 9
      "0001001" when "01011001101011100", -- t[45916] = 9
      "0001001" when "01011001101011101", -- t[45917] = 9
      "0001001" when "01011001101011110", -- t[45918] = 9
      "0001001" when "01011001101011111", -- t[45919] = 9
      "0001001" when "01011001101100000", -- t[45920] = 9
      "0001001" when "01011001101100001", -- t[45921] = 9
      "0001001" when "01011001101100010", -- t[45922] = 9
      "0001001" when "01011001101100011", -- t[45923] = 9
      "0001001" when "01011001101100100", -- t[45924] = 9
      "0001001" when "01011001101100101", -- t[45925] = 9
      "0001001" when "01011001101100110", -- t[45926] = 9
      "0001001" when "01011001101100111", -- t[45927] = 9
      "0001001" when "01011001101101000", -- t[45928] = 9
      "0001001" when "01011001101101001", -- t[45929] = 9
      "0001001" when "01011001101101010", -- t[45930] = 9
      "0001001" when "01011001101101011", -- t[45931] = 9
      "0001001" when "01011001101101100", -- t[45932] = 9
      "0001001" when "01011001101101101", -- t[45933] = 9
      "0001001" when "01011001101101110", -- t[45934] = 9
      "0001001" when "01011001101101111", -- t[45935] = 9
      "0001001" when "01011001101110000", -- t[45936] = 9
      "0001001" when "01011001101110001", -- t[45937] = 9
      "0001001" when "01011001101110010", -- t[45938] = 9
      "0001001" when "01011001101110011", -- t[45939] = 9
      "0001001" when "01011001101110100", -- t[45940] = 9
      "0001001" when "01011001101110101", -- t[45941] = 9
      "0001001" when "01011001101110110", -- t[45942] = 9
      "0001001" when "01011001101110111", -- t[45943] = 9
      "0001001" when "01011001101111000", -- t[45944] = 9
      "0001001" when "01011001101111001", -- t[45945] = 9
      "0001001" when "01011001101111010", -- t[45946] = 9
      "0001001" when "01011001101111011", -- t[45947] = 9
      "0001001" when "01011001101111100", -- t[45948] = 9
      "0001001" when "01011001101111101", -- t[45949] = 9
      "0001001" when "01011001101111110", -- t[45950] = 9
      "0001001" when "01011001101111111", -- t[45951] = 9
      "0001001" when "01011001110000000", -- t[45952] = 9
      "0001001" when "01011001110000001", -- t[45953] = 9
      "0001001" when "01011001110000010", -- t[45954] = 9
      "0001001" when "01011001110000011", -- t[45955] = 9
      "0001001" when "01011001110000100", -- t[45956] = 9
      "0001001" when "01011001110000101", -- t[45957] = 9
      "0001001" when "01011001110000110", -- t[45958] = 9
      "0001001" when "01011001110000111", -- t[45959] = 9
      "0001001" when "01011001110001000", -- t[45960] = 9
      "0001001" when "01011001110001001", -- t[45961] = 9
      "0001001" when "01011001110001010", -- t[45962] = 9
      "0001001" when "01011001110001011", -- t[45963] = 9
      "0001001" when "01011001110001100", -- t[45964] = 9
      "0001001" when "01011001110001101", -- t[45965] = 9
      "0001001" when "01011001110001110", -- t[45966] = 9
      "0001001" when "01011001110001111", -- t[45967] = 9
      "0001001" when "01011001110010000", -- t[45968] = 9
      "0001001" when "01011001110010001", -- t[45969] = 9
      "0001001" when "01011001110010010", -- t[45970] = 9
      "0001001" when "01011001110010011", -- t[45971] = 9
      "0001001" when "01011001110010100", -- t[45972] = 9
      "0001001" when "01011001110010101", -- t[45973] = 9
      "0001001" when "01011001110010110", -- t[45974] = 9
      "0001001" when "01011001110010111", -- t[45975] = 9
      "0001001" when "01011001110011000", -- t[45976] = 9
      "0001001" when "01011001110011001", -- t[45977] = 9
      "0001001" when "01011001110011010", -- t[45978] = 9
      "0001001" when "01011001110011011", -- t[45979] = 9
      "0001001" when "01011001110011100", -- t[45980] = 9
      "0001001" when "01011001110011101", -- t[45981] = 9
      "0001001" when "01011001110011110", -- t[45982] = 9
      "0001001" when "01011001110011111", -- t[45983] = 9
      "0001001" when "01011001110100000", -- t[45984] = 9
      "0001001" when "01011001110100001", -- t[45985] = 9
      "0001001" when "01011001110100010", -- t[45986] = 9
      "0001001" when "01011001110100011", -- t[45987] = 9
      "0001001" when "01011001110100100", -- t[45988] = 9
      "0001001" when "01011001110100101", -- t[45989] = 9
      "0001001" when "01011001110100110", -- t[45990] = 9
      "0001001" when "01011001110100111", -- t[45991] = 9
      "0001001" when "01011001110101000", -- t[45992] = 9
      "0001001" when "01011001110101001", -- t[45993] = 9
      "0001001" when "01011001110101010", -- t[45994] = 9
      "0001001" when "01011001110101011", -- t[45995] = 9
      "0001001" when "01011001110101100", -- t[45996] = 9
      "0001001" when "01011001110101101", -- t[45997] = 9
      "0001001" when "01011001110101110", -- t[45998] = 9
      "0001001" when "01011001110101111", -- t[45999] = 9
      "0001001" when "01011001110110000", -- t[46000] = 9
      "0001001" when "01011001110110001", -- t[46001] = 9
      "0001001" when "01011001110110010", -- t[46002] = 9
      "0001001" when "01011001110110011", -- t[46003] = 9
      "0001001" when "01011001110110100", -- t[46004] = 9
      "0001001" when "01011001110110101", -- t[46005] = 9
      "0001001" when "01011001110110110", -- t[46006] = 9
      "0001001" when "01011001110110111", -- t[46007] = 9
      "0001001" when "01011001110111000", -- t[46008] = 9
      "0001001" when "01011001110111001", -- t[46009] = 9
      "0001001" when "01011001110111010", -- t[46010] = 9
      "0001001" when "01011001110111011", -- t[46011] = 9
      "0001001" when "01011001110111100", -- t[46012] = 9
      "0001001" when "01011001110111101", -- t[46013] = 9
      "0001001" when "01011001110111110", -- t[46014] = 9
      "0001001" when "01011001110111111", -- t[46015] = 9
      "0001001" when "01011001111000000", -- t[46016] = 9
      "0001001" when "01011001111000001", -- t[46017] = 9
      "0001001" when "01011001111000010", -- t[46018] = 9
      "0001001" when "01011001111000011", -- t[46019] = 9
      "0001001" when "01011001111000100", -- t[46020] = 9
      "0001001" when "01011001111000101", -- t[46021] = 9
      "0001001" when "01011001111000110", -- t[46022] = 9
      "0001001" when "01011001111000111", -- t[46023] = 9
      "0001001" when "01011001111001000", -- t[46024] = 9
      "0001001" when "01011001111001001", -- t[46025] = 9
      "0001001" when "01011001111001010", -- t[46026] = 9
      "0001001" when "01011001111001011", -- t[46027] = 9
      "0001001" when "01011001111001100", -- t[46028] = 9
      "0001001" when "01011001111001101", -- t[46029] = 9
      "0001001" when "01011001111001110", -- t[46030] = 9
      "0001001" when "01011001111001111", -- t[46031] = 9
      "0001001" when "01011001111010000", -- t[46032] = 9
      "0001001" when "01011001111010001", -- t[46033] = 9
      "0001001" when "01011001111010010", -- t[46034] = 9
      "0001001" when "01011001111010011", -- t[46035] = 9
      "0001001" when "01011001111010100", -- t[46036] = 9
      "0001001" when "01011001111010101", -- t[46037] = 9
      "0001001" when "01011001111010110", -- t[46038] = 9
      "0001001" when "01011001111010111", -- t[46039] = 9
      "0001001" when "01011001111011000", -- t[46040] = 9
      "0001001" when "01011001111011001", -- t[46041] = 9
      "0001001" when "01011001111011010", -- t[46042] = 9
      "0001001" when "01011001111011011", -- t[46043] = 9
      "0001001" when "01011001111011100", -- t[46044] = 9
      "0001001" when "01011001111011101", -- t[46045] = 9
      "0001001" when "01011001111011110", -- t[46046] = 9
      "0001001" when "01011001111011111", -- t[46047] = 9
      "0001001" when "01011001111100000", -- t[46048] = 9
      "0001001" when "01011001111100001", -- t[46049] = 9
      "0001001" when "01011001111100010", -- t[46050] = 9
      "0001001" when "01011001111100011", -- t[46051] = 9
      "0001001" when "01011001111100100", -- t[46052] = 9
      "0001001" when "01011001111100101", -- t[46053] = 9
      "0001001" when "01011001111100110", -- t[46054] = 9
      "0001001" when "01011001111100111", -- t[46055] = 9
      "0001001" when "01011001111101000", -- t[46056] = 9
      "0001001" when "01011001111101001", -- t[46057] = 9
      "0001001" when "01011001111101010", -- t[46058] = 9
      "0001001" when "01011001111101011", -- t[46059] = 9
      "0001001" when "01011001111101100", -- t[46060] = 9
      "0001001" when "01011001111101101", -- t[46061] = 9
      "0001001" when "01011001111101110", -- t[46062] = 9
      "0001001" when "01011001111101111", -- t[46063] = 9
      "0001001" when "01011001111110000", -- t[46064] = 9
      "0001001" when "01011001111110001", -- t[46065] = 9
      "0001001" when "01011001111110010", -- t[46066] = 9
      "0001001" when "01011001111110011", -- t[46067] = 9
      "0001001" when "01011001111110100", -- t[46068] = 9
      "0001001" when "01011001111110101", -- t[46069] = 9
      "0001001" when "01011001111110110", -- t[46070] = 9
      "0001001" when "01011001111110111", -- t[46071] = 9
      "0001001" when "01011001111111000", -- t[46072] = 9
      "0001001" when "01011001111111001", -- t[46073] = 9
      "0001001" when "01011001111111010", -- t[46074] = 9
      "0001001" when "01011001111111011", -- t[46075] = 9
      "0001001" when "01011001111111100", -- t[46076] = 9
      "0001001" when "01011001111111101", -- t[46077] = 9
      "0001001" when "01011001111111110", -- t[46078] = 9
      "0001001" when "01011001111111111", -- t[46079] = 9
      "0001001" when "01011010000000000", -- t[46080] = 9
      "0001001" when "01011010000000001", -- t[46081] = 9
      "0001001" when "01011010000000010", -- t[46082] = 9
      "0001001" when "01011010000000011", -- t[46083] = 9
      "0001001" when "01011010000000100", -- t[46084] = 9
      "0001001" when "01011010000000101", -- t[46085] = 9
      "0001001" when "01011010000000110", -- t[46086] = 9
      "0001001" when "01011010000000111", -- t[46087] = 9
      "0001001" when "01011010000001000", -- t[46088] = 9
      "0001001" when "01011010000001001", -- t[46089] = 9
      "0001001" when "01011010000001010", -- t[46090] = 9
      "0001001" when "01011010000001011", -- t[46091] = 9
      "0001001" when "01011010000001100", -- t[46092] = 9
      "0001001" when "01011010000001101", -- t[46093] = 9
      "0001001" when "01011010000001110", -- t[46094] = 9
      "0001001" when "01011010000001111", -- t[46095] = 9
      "0001001" when "01011010000010000", -- t[46096] = 9
      "0001001" when "01011010000010001", -- t[46097] = 9
      "0001001" when "01011010000010010", -- t[46098] = 9
      "0001001" when "01011010000010011", -- t[46099] = 9
      "0001001" when "01011010000010100", -- t[46100] = 9
      "0001001" when "01011010000010101", -- t[46101] = 9
      "0001001" when "01011010000010110", -- t[46102] = 9
      "0001001" when "01011010000010111", -- t[46103] = 9
      "0001001" when "01011010000011000", -- t[46104] = 9
      "0001001" when "01011010000011001", -- t[46105] = 9
      "0001001" when "01011010000011010", -- t[46106] = 9
      "0001001" when "01011010000011011", -- t[46107] = 9
      "0001001" when "01011010000011100", -- t[46108] = 9
      "0001001" when "01011010000011101", -- t[46109] = 9
      "0001001" when "01011010000011110", -- t[46110] = 9
      "0001001" when "01011010000011111", -- t[46111] = 9
      "0001001" when "01011010000100000", -- t[46112] = 9
      "0001001" when "01011010000100001", -- t[46113] = 9
      "0001001" when "01011010000100010", -- t[46114] = 9
      "0001001" when "01011010000100011", -- t[46115] = 9
      "0001001" when "01011010000100100", -- t[46116] = 9
      "0001001" when "01011010000100101", -- t[46117] = 9
      "0001001" when "01011010000100110", -- t[46118] = 9
      "0001001" when "01011010000100111", -- t[46119] = 9
      "0001001" when "01011010000101000", -- t[46120] = 9
      "0001001" when "01011010000101001", -- t[46121] = 9
      "0001001" when "01011010000101010", -- t[46122] = 9
      "0001001" when "01011010000101011", -- t[46123] = 9
      "0001001" when "01011010000101100", -- t[46124] = 9
      "0001001" when "01011010000101101", -- t[46125] = 9
      "0001001" when "01011010000101110", -- t[46126] = 9
      "0001001" when "01011010000101111", -- t[46127] = 9
      "0001001" when "01011010000110000", -- t[46128] = 9
      "0001001" when "01011010000110001", -- t[46129] = 9
      "0001001" when "01011010000110010", -- t[46130] = 9
      "0001001" when "01011010000110011", -- t[46131] = 9
      "0001001" when "01011010000110100", -- t[46132] = 9
      "0001001" when "01011010000110101", -- t[46133] = 9
      "0001001" when "01011010000110110", -- t[46134] = 9
      "0001001" when "01011010000110111", -- t[46135] = 9
      "0001001" when "01011010000111000", -- t[46136] = 9
      "0001001" when "01011010000111001", -- t[46137] = 9
      "0001001" when "01011010000111010", -- t[46138] = 9
      "0001001" when "01011010000111011", -- t[46139] = 9
      "0001001" when "01011010000111100", -- t[46140] = 9
      "0001001" when "01011010000111101", -- t[46141] = 9
      "0001001" when "01011010000111110", -- t[46142] = 9
      "0001001" when "01011010000111111", -- t[46143] = 9
      "0001001" when "01011010001000000", -- t[46144] = 9
      "0001001" when "01011010001000001", -- t[46145] = 9
      "0001001" when "01011010001000010", -- t[46146] = 9
      "0001001" when "01011010001000011", -- t[46147] = 9
      "0001001" when "01011010001000100", -- t[46148] = 9
      "0001001" when "01011010001000101", -- t[46149] = 9
      "0001001" when "01011010001000110", -- t[46150] = 9
      "0001001" when "01011010001000111", -- t[46151] = 9
      "0001001" when "01011010001001000", -- t[46152] = 9
      "0001001" when "01011010001001001", -- t[46153] = 9
      "0001001" when "01011010001001010", -- t[46154] = 9
      "0001001" when "01011010001001011", -- t[46155] = 9
      "0001001" when "01011010001001100", -- t[46156] = 9
      "0001001" when "01011010001001101", -- t[46157] = 9
      "0001001" when "01011010001001110", -- t[46158] = 9
      "0001001" when "01011010001001111", -- t[46159] = 9
      "0001001" when "01011010001010000", -- t[46160] = 9
      "0001001" when "01011010001010001", -- t[46161] = 9
      "0001001" when "01011010001010010", -- t[46162] = 9
      "0001001" when "01011010001010011", -- t[46163] = 9
      "0001001" when "01011010001010100", -- t[46164] = 9
      "0001001" when "01011010001010101", -- t[46165] = 9
      "0001001" when "01011010001010110", -- t[46166] = 9
      "0001001" when "01011010001010111", -- t[46167] = 9
      "0001001" when "01011010001011000", -- t[46168] = 9
      "0001001" when "01011010001011001", -- t[46169] = 9
      "0001001" when "01011010001011010", -- t[46170] = 9
      "0001001" when "01011010001011011", -- t[46171] = 9
      "0001001" when "01011010001011100", -- t[46172] = 9
      "0001001" when "01011010001011101", -- t[46173] = 9
      "0001001" when "01011010001011110", -- t[46174] = 9
      "0001001" when "01011010001011111", -- t[46175] = 9
      "0001001" when "01011010001100000", -- t[46176] = 9
      "0001001" when "01011010001100001", -- t[46177] = 9
      "0001001" when "01011010001100010", -- t[46178] = 9
      "0001001" when "01011010001100011", -- t[46179] = 9
      "0001001" when "01011010001100100", -- t[46180] = 9
      "0001001" when "01011010001100101", -- t[46181] = 9
      "0001001" when "01011010001100110", -- t[46182] = 9
      "0001001" when "01011010001100111", -- t[46183] = 9
      "0001001" when "01011010001101000", -- t[46184] = 9
      "0001001" when "01011010001101001", -- t[46185] = 9
      "0001001" when "01011010001101010", -- t[46186] = 9
      "0001001" when "01011010001101011", -- t[46187] = 9
      "0001001" when "01011010001101100", -- t[46188] = 9
      "0001001" when "01011010001101101", -- t[46189] = 9
      "0001001" when "01011010001101110", -- t[46190] = 9
      "0001001" when "01011010001101111", -- t[46191] = 9
      "0001001" when "01011010001110000", -- t[46192] = 9
      "0001001" when "01011010001110001", -- t[46193] = 9
      "0001001" when "01011010001110010", -- t[46194] = 9
      "0001001" when "01011010001110011", -- t[46195] = 9
      "0001001" when "01011010001110100", -- t[46196] = 9
      "0001001" when "01011010001110101", -- t[46197] = 9
      "0001001" when "01011010001110110", -- t[46198] = 9
      "0001001" when "01011010001110111", -- t[46199] = 9
      "0001001" when "01011010001111000", -- t[46200] = 9
      "0001001" when "01011010001111001", -- t[46201] = 9
      "0001001" when "01011010001111010", -- t[46202] = 9
      "0001001" when "01011010001111011", -- t[46203] = 9
      "0001001" when "01011010001111100", -- t[46204] = 9
      "0001001" when "01011010001111101", -- t[46205] = 9
      "0001001" when "01011010001111110", -- t[46206] = 9
      "0001001" when "01011010001111111", -- t[46207] = 9
      "0001001" when "01011010010000000", -- t[46208] = 9
      "0001001" when "01011010010000001", -- t[46209] = 9
      "0001001" when "01011010010000010", -- t[46210] = 9
      "0001001" when "01011010010000011", -- t[46211] = 9
      "0001001" when "01011010010000100", -- t[46212] = 9
      "0001001" when "01011010010000101", -- t[46213] = 9
      "0001001" when "01011010010000110", -- t[46214] = 9
      "0001001" when "01011010010000111", -- t[46215] = 9
      "0001001" when "01011010010001000", -- t[46216] = 9
      "0001001" when "01011010010001001", -- t[46217] = 9
      "0001001" when "01011010010001010", -- t[46218] = 9
      "0001001" when "01011010010001011", -- t[46219] = 9
      "0001001" when "01011010010001100", -- t[46220] = 9
      "0001001" when "01011010010001101", -- t[46221] = 9
      "0001001" when "01011010010001110", -- t[46222] = 9
      "0001001" when "01011010010001111", -- t[46223] = 9
      "0001001" when "01011010010010000", -- t[46224] = 9
      "0001001" when "01011010010010001", -- t[46225] = 9
      "0001001" when "01011010010010010", -- t[46226] = 9
      "0001001" when "01011010010010011", -- t[46227] = 9
      "0001001" when "01011010010010100", -- t[46228] = 9
      "0001001" when "01011010010010101", -- t[46229] = 9
      "0001001" when "01011010010010110", -- t[46230] = 9
      "0001001" when "01011010010010111", -- t[46231] = 9
      "0001001" when "01011010010011000", -- t[46232] = 9
      "0001001" when "01011010010011001", -- t[46233] = 9
      "0001001" when "01011010010011010", -- t[46234] = 9
      "0001001" when "01011010010011011", -- t[46235] = 9
      "0001001" when "01011010010011100", -- t[46236] = 9
      "0001001" when "01011010010011101", -- t[46237] = 9
      "0001001" when "01011010010011110", -- t[46238] = 9
      "0001001" when "01011010010011111", -- t[46239] = 9
      "0001001" when "01011010010100000", -- t[46240] = 9
      "0001001" when "01011010010100001", -- t[46241] = 9
      "0001001" when "01011010010100010", -- t[46242] = 9
      "0001001" when "01011010010100011", -- t[46243] = 9
      "0001001" when "01011010010100100", -- t[46244] = 9
      "0001001" when "01011010010100101", -- t[46245] = 9
      "0001001" when "01011010010100110", -- t[46246] = 9
      "0001001" when "01011010010100111", -- t[46247] = 9
      "0001001" when "01011010010101000", -- t[46248] = 9
      "0001001" when "01011010010101001", -- t[46249] = 9
      "0001001" when "01011010010101010", -- t[46250] = 9
      "0001001" when "01011010010101011", -- t[46251] = 9
      "0001001" when "01011010010101100", -- t[46252] = 9
      "0001001" when "01011010010101101", -- t[46253] = 9
      "0001001" when "01011010010101110", -- t[46254] = 9
      "0001001" when "01011010010101111", -- t[46255] = 9
      "0001001" when "01011010010110000", -- t[46256] = 9
      "0001001" when "01011010010110001", -- t[46257] = 9
      "0001001" when "01011010010110010", -- t[46258] = 9
      "0001001" when "01011010010110011", -- t[46259] = 9
      "0001001" when "01011010010110100", -- t[46260] = 9
      "0001001" when "01011010010110101", -- t[46261] = 9
      "0001001" when "01011010010110110", -- t[46262] = 9
      "0001001" when "01011010010110111", -- t[46263] = 9
      "0001001" when "01011010010111000", -- t[46264] = 9
      "0001001" when "01011010010111001", -- t[46265] = 9
      "0001001" when "01011010010111010", -- t[46266] = 9
      "0001001" when "01011010010111011", -- t[46267] = 9
      "0001001" when "01011010010111100", -- t[46268] = 9
      "0001001" when "01011010010111101", -- t[46269] = 9
      "0001001" when "01011010010111110", -- t[46270] = 9
      "0001001" when "01011010010111111", -- t[46271] = 9
      "0001001" when "01011010011000000", -- t[46272] = 9
      "0001001" when "01011010011000001", -- t[46273] = 9
      "0001001" when "01011010011000010", -- t[46274] = 9
      "0001001" when "01011010011000011", -- t[46275] = 9
      "0001001" when "01011010011000100", -- t[46276] = 9
      "0001001" when "01011010011000101", -- t[46277] = 9
      "0001001" when "01011010011000110", -- t[46278] = 9
      "0001001" when "01011010011000111", -- t[46279] = 9
      "0001001" when "01011010011001000", -- t[46280] = 9
      "0001001" when "01011010011001001", -- t[46281] = 9
      "0001001" when "01011010011001010", -- t[46282] = 9
      "0001001" when "01011010011001011", -- t[46283] = 9
      "0001001" when "01011010011001100", -- t[46284] = 9
      "0001001" when "01011010011001101", -- t[46285] = 9
      "0001001" when "01011010011001110", -- t[46286] = 9
      "0001001" when "01011010011001111", -- t[46287] = 9
      "0001001" when "01011010011010000", -- t[46288] = 9
      "0001001" when "01011010011010001", -- t[46289] = 9
      "0001001" when "01011010011010010", -- t[46290] = 9
      "0001001" when "01011010011010011", -- t[46291] = 9
      "0001001" when "01011010011010100", -- t[46292] = 9
      "0001001" when "01011010011010101", -- t[46293] = 9
      "0001001" when "01011010011010110", -- t[46294] = 9
      "0001001" when "01011010011010111", -- t[46295] = 9
      "0001001" when "01011010011011000", -- t[46296] = 9
      "0001001" when "01011010011011001", -- t[46297] = 9
      "0001001" when "01011010011011010", -- t[46298] = 9
      "0001001" when "01011010011011011", -- t[46299] = 9
      "0001001" when "01011010011011100", -- t[46300] = 9
      "0001001" when "01011010011011101", -- t[46301] = 9
      "0001001" when "01011010011011110", -- t[46302] = 9
      "0001001" when "01011010011011111", -- t[46303] = 9
      "0001001" when "01011010011100000", -- t[46304] = 9
      "0001001" when "01011010011100001", -- t[46305] = 9
      "0001001" when "01011010011100010", -- t[46306] = 9
      "0001001" when "01011010011100011", -- t[46307] = 9
      "0001001" when "01011010011100100", -- t[46308] = 9
      "0001001" when "01011010011100101", -- t[46309] = 9
      "0001001" when "01011010011100110", -- t[46310] = 9
      "0001001" when "01011010011100111", -- t[46311] = 9
      "0001001" when "01011010011101000", -- t[46312] = 9
      "0001001" when "01011010011101001", -- t[46313] = 9
      "0001001" when "01011010011101010", -- t[46314] = 9
      "0001001" when "01011010011101011", -- t[46315] = 9
      "0001001" when "01011010011101100", -- t[46316] = 9
      "0001001" when "01011010011101101", -- t[46317] = 9
      "0001001" when "01011010011101110", -- t[46318] = 9
      "0001001" when "01011010011101111", -- t[46319] = 9
      "0001001" when "01011010011110000", -- t[46320] = 9
      "0001001" when "01011010011110001", -- t[46321] = 9
      "0001001" when "01011010011110010", -- t[46322] = 9
      "0001001" when "01011010011110011", -- t[46323] = 9
      "0001001" when "01011010011110100", -- t[46324] = 9
      "0001001" when "01011010011110101", -- t[46325] = 9
      "0001001" when "01011010011110110", -- t[46326] = 9
      "0001001" when "01011010011110111", -- t[46327] = 9
      "0001001" when "01011010011111000", -- t[46328] = 9
      "0001001" when "01011010011111001", -- t[46329] = 9
      "0001001" when "01011010011111010", -- t[46330] = 9
      "0001001" when "01011010011111011", -- t[46331] = 9
      "0001001" when "01011010011111100", -- t[46332] = 9
      "0001001" when "01011010011111101", -- t[46333] = 9
      "0001001" when "01011010011111110", -- t[46334] = 9
      "0001001" when "01011010011111111", -- t[46335] = 9
      "0001001" when "01011010100000000", -- t[46336] = 9
      "0001001" when "01011010100000001", -- t[46337] = 9
      "0001001" when "01011010100000010", -- t[46338] = 9
      "0001001" when "01011010100000011", -- t[46339] = 9
      "0001001" when "01011010100000100", -- t[46340] = 9
      "0001001" when "01011010100000101", -- t[46341] = 9
      "0001001" when "01011010100000110", -- t[46342] = 9
      "0001001" when "01011010100000111", -- t[46343] = 9
      "0001001" when "01011010100001000", -- t[46344] = 9
      "0001001" when "01011010100001001", -- t[46345] = 9
      "0001001" when "01011010100001010", -- t[46346] = 9
      "0001001" when "01011010100001011", -- t[46347] = 9
      "0001001" when "01011010100001100", -- t[46348] = 9
      "0001001" when "01011010100001101", -- t[46349] = 9
      "0001001" when "01011010100001110", -- t[46350] = 9
      "0001001" when "01011010100001111", -- t[46351] = 9
      "0001001" when "01011010100010000", -- t[46352] = 9
      "0001001" when "01011010100010001", -- t[46353] = 9
      "0001001" when "01011010100010010", -- t[46354] = 9
      "0001001" when "01011010100010011", -- t[46355] = 9
      "0001001" when "01011010100010100", -- t[46356] = 9
      "0001001" when "01011010100010101", -- t[46357] = 9
      "0001001" when "01011010100010110", -- t[46358] = 9
      "0001001" when "01011010100010111", -- t[46359] = 9
      "0001001" when "01011010100011000", -- t[46360] = 9
      "0001001" when "01011010100011001", -- t[46361] = 9
      "0001001" when "01011010100011010", -- t[46362] = 9
      "0001001" when "01011010100011011", -- t[46363] = 9
      "0001001" when "01011010100011100", -- t[46364] = 9
      "0001001" when "01011010100011101", -- t[46365] = 9
      "0001001" when "01011010100011110", -- t[46366] = 9
      "0001001" when "01011010100011111", -- t[46367] = 9
      "0001001" when "01011010100100000", -- t[46368] = 9
      "0001001" when "01011010100100001", -- t[46369] = 9
      "0001001" when "01011010100100010", -- t[46370] = 9
      "0001001" when "01011010100100011", -- t[46371] = 9
      "0001001" when "01011010100100100", -- t[46372] = 9
      "0001001" when "01011010100100101", -- t[46373] = 9
      "0001001" when "01011010100100110", -- t[46374] = 9
      "0001001" when "01011010100100111", -- t[46375] = 9
      "0001001" when "01011010100101000", -- t[46376] = 9
      "0001001" when "01011010100101001", -- t[46377] = 9
      "0001001" when "01011010100101010", -- t[46378] = 9
      "0001001" when "01011010100101011", -- t[46379] = 9
      "0001001" when "01011010100101100", -- t[46380] = 9
      "0001001" when "01011010100101101", -- t[46381] = 9
      "0001001" when "01011010100101110", -- t[46382] = 9
      "0001001" when "01011010100101111", -- t[46383] = 9
      "0001001" when "01011010100110000", -- t[46384] = 9
      "0001001" when "01011010100110001", -- t[46385] = 9
      "0001001" when "01011010100110010", -- t[46386] = 9
      "0001001" when "01011010100110011", -- t[46387] = 9
      "0001001" when "01011010100110100", -- t[46388] = 9
      "0001001" when "01011010100110101", -- t[46389] = 9
      "0001001" when "01011010100110110", -- t[46390] = 9
      "0001001" when "01011010100110111", -- t[46391] = 9
      "0001001" when "01011010100111000", -- t[46392] = 9
      "0001001" when "01011010100111001", -- t[46393] = 9
      "0001001" when "01011010100111010", -- t[46394] = 9
      "0001001" when "01011010100111011", -- t[46395] = 9
      "0001001" when "01011010100111100", -- t[46396] = 9
      "0001001" when "01011010100111101", -- t[46397] = 9
      "0001001" when "01011010100111110", -- t[46398] = 9
      "0001001" when "01011010100111111", -- t[46399] = 9
      "0001001" when "01011010101000000", -- t[46400] = 9
      "0001001" when "01011010101000001", -- t[46401] = 9
      "0001001" when "01011010101000010", -- t[46402] = 9
      "0001001" when "01011010101000011", -- t[46403] = 9
      "0001001" when "01011010101000100", -- t[46404] = 9
      "0001001" when "01011010101000101", -- t[46405] = 9
      "0001001" when "01011010101000110", -- t[46406] = 9
      "0001001" when "01011010101000111", -- t[46407] = 9
      "0001001" when "01011010101001000", -- t[46408] = 9
      "0001001" when "01011010101001001", -- t[46409] = 9
      "0001001" when "01011010101001010", -- t[46410] = 9
      "0001001" when "01011010101001011", -- t[46411] = 9
      "0001001" when "01011010101001100", -- t[46412] = 9
      "0001001" when "01011010101001101", -- t[46413] = 9
      "0001001" when "01011010101001110", -- t[46414] = 9
      "0001001" when "01011010101001111", -- t[46415] = 9
      "0001001" when "01011010101010000", -- t[46416] = 9
      "0001001" when "01011010101010001", -- t[46417] = 9
      "0001001" when "01011010101010010", -- t[46418] = 9
      "0001001" when "01011010101010011", -- t[46419] = 9
      "0001001" when "01011010101010100", -- t[46420] = 9
      "0001001" when "01011010101010101", -- t[46421] = 9
      "0001001" when "01011010101010110", -- t[46422] = 9
      "0001001" when "01011010101010111", -- t[46423] = 9
      "0001001" when "01011010101011000", -- t[46424] = 9
      "0001001" when "01011010101011001", -- t[46425] = 9
      "0001001" when "01011010101011010", -- t[46426] = 9
      "0001001" when "01011010101011011", -- t[46427] = 9
      "0001001" when "01011010101011100", -- t[46428] = 9
      "0001001" when "01011010101011101", -- t[46429] = 9
      "0001001" when "01011010101011110", -- t[46430] = 9
      "0001001" when "01011010101011111", -- t[46431] = 9
      "0001001" when "01011010101100000", -- t[46432] = 9
      "0001001" when "01011010101100001", -- t[46433] = 9
      "0001001" when "01011010101100010", -- t[46434] = 9
      "0001001" when "01011010101100011", -- t[46435] = 9
      "0001001" when "01011010101100100", -- t[46436] = 9
      "0001001" when "01011010101100101", -- t[46437] = 9
      "0001001" when "01011010101100110", -- t[46438] = 9
      "0001001" when "01011010101100111", -- t[46439] = 9
      "0001001" when "01011010101101000", -- t[46440] = 9
      "0001001" when "01011010101101001", -- t[46441] = 9
      "0001001" when "01011010101101010", -- t[46442] = 9
      "0001001" when "01011010101101011", -- t[46443] = 9
      "0001001" when "01011010101101100", -- t[46444] = 9
      "0001001" when "01011010101101101", -- t[46445] = 9
      "0001001" when "01011010101101110", -- t[46446] = 9
      "0001001" when "01011010101101111", -- t[46447] = 9
      "0001001" when "01011010101110000", -- t[46448] = 9
      "0001001" when "01011010101110001", -- t[46449] = 9
      "0001001" when "01011010101110010", -- t[46450] = 9
      "0001001" when "01011010101110011", -- t[46451] = 9
      "0001001" when "01011010101110100", -- t[46452] = 9
      "0001001" when "01011010101110101", -- t[46453] = 9
      "0001001" when "01011010101110110", -- t[46454] = 9
      "0001001" when "01011010101110111", -- t[46455] = 9
      "0001001" when "01011010101111000", -- t[46456] = 9
      "0001001" when "01011010101111001", -- t[46457] = 9
      "0001001" when "01011010101111010", -- t[46458] = 9
      "0001001" when "01011010101111011", -- t[46459] = 9
      "0001001" when "01011010101111100", -- t[46460] = 9
      "0001001" when "01011010101111101", -- t[46461] = 9
      "0001001" when "01011010101111110", -- t[46462] = 9
      "0001001" when "01011010101111111", -- t[46463] = 9
      "0001001" when "01011010110000000", -- t[46464] = 9
      "0001001" when "01011010110000001", -- t[46465] = 9
      "0001001" when "01011010110000010", -- t[46466] = 9
      "0001001" when "01011010110000011", -- t[46467] = 9
      "0001001" when "01011010110000100", -- t[46468] = 9
      "0001001" when "01011010110000101", -- t[46469] = 9
      "0001001" when "01011010110000110", -- t[46470] = 9
      "0001001" when "01011010110000111", -- t[46471] = 9
      "0001001" when "01011010110001000", -- t[46472] = 9
      "0001001" when "01011010110001001", -- t[46473] = 9
      "0001001" when "01011010110001010", -- t[46474] = 9
      "0001001" when "01011010110001011", -- t[46475] = 9
      "0001001" when "01011010110001100", -- t[46476] = 9
      "0001001" when "01011010110001101", -- t[46477] = 9
      "0001001" when "01011010110001110", -- t[46478] = 9
      "0001001" when "01011010110001111", -- t[46479] = 9
      "0001001" when "01011010110010000", -- t[46480] = 9
      "0001001" when "01011010110010001", -- t[46481] = 9
      "0001001" when "01011010110010010", -- t[46482] = 9
      "0001001" when "01011010110010011", -- t[46483] = 9
      "0001001" when "01011010110010100", -- t[46484] = 9
      "0001001" when "01011010110010101", -- t[46485] = 9
      "0001001" when "01011010110010110", -- t[46486] = 9
      "0001001" when "01011010110010111", -- t[46487] = 9
      "0001001" when "01011010110011000", -- t[46488] = 9
      "0001001" when "01011010110011001", -- t[46489] = 9
      "0001001" when "01011010110011010", -- t[46490] = 9
      "0001001" when "01011010110011011", -- t[46491] = 9
      "0001001" when "01011010110011100", -- t[46492] = 9
      "0001001" when "01011010110011101", -- t[46493] = 9
      "0001001" when "01011010110011110", -- t[46494] = 9
      "0001001" when "01011010110011111", -- t[46495] = 9
      "0001001" when "01011010110100000", -- t[46496] = 9
      "0001001" when "01011010110100001", -- t[46497] = 9
      "0001001" when "01011010110100010", -- t[46498] = 9
      "0001001" when "01011010110100011", -- t[46499] = 9
      "0001001" when "01011010110100100", -- t[46500] = 9
      "0001001" when "01011010110100101", -- t[46501] = 9
      "0001001" when "01011010110100110", -- t[46502] = 9
      "0001001" when "01011010110100111", -- t[46503] = 9
      "0001001" when "01011010110101000", -- t[46504] = 9
      "0001001" when "01011010110101001", -- t[46505] = 9
      "0001001" when "01011010110101010", -- t[46506] = 9
      "0001001" when "01011010110101011", -- t[46507] = 9
      "0001001" when "01011010110101100", -- t[46508] = 9
      "0001001" when "01011010110101101", -- t[46509] = 9
      "0001001" when "01011010110101110", -- t[46510] = 9
      "0001001" when "01011010110101111", -- t[46511] = 9
      "0001001" when "01011010110110000", -- t[46512] = 9
      "0001001" when "01011010110110001", -- t[46513] = 9
      "0001001" when "01011010110110010", -- t[46514] = 9
      "0001001" when "01011010110110011", -- t[46515] = 9
      "0001001" when "01011010110110100", -- t[46516] = 9
      "0001001" when "01011010110110101", -- t[46517] = 9
      "0001001" when "01011010110110110", -- t[46518] = 9
      "0001001" when "01011010110110111", -- t[46519] = 9
      "0001001" when "01011010110111000", -- t[46520] = 9
      "0001001" when "01011010110111001", -- t[46521] = 9
      "0001001" when "01011010110111010", -- t[46522] = 9
      "0001001" when "01011010110111011", -- t[46523] = 9
      "0001001" when "01011010110111100", -- t[46524] = 9
      "0001001" when "01011010110111101", -- t[46525] = 9
      "0001001" when "01011010110111110", -- t[46526] = 9
      "0001001" when "01011010110111111", -- t[46527] = 9
      "0001001" when "01011010111000000", -- t[46528] = 9
      "0001001" when "01011010111000001", -- t[46529] = 9
      "0001001" when "01011010111000010", -- t[46530] = 9
      "0001001" when "01011010111000011", -- t[46531] = 9
      "0001001" when "01011010111000100", -- t[46532] = 9
      "0001001" when "01011010111000101", -- t[46533] = 9
      "0001001" when "01011010111000110", -- t[46534] = 9
      "0001001" when "01011010111000111", -- t[46535] = 9
      "0001001" when "01011010111001000", -- t[46536] = 9
      "0001001" when "01011010111001001", -- t[46537] = 9
      "0001001" when "01011010111001010", -- t[46538] = 9
      "0001001" when "01011010111001011", -- t[46539] = 9
      "0001001" when "01011010111001100", -- t[46540] = 9
      "0001001" when "01011010111001101", -- t[46541] = 9
      "0001001" when "01011010111001110", -- t[46542] = 9
      "0001001" when "01011010111001111", -- t[46543] = 9
      "0001001" when "01011010111010000", -- t[46544] = 9
      "0001001" when "01011010111010001", -- t[46545] = 9
      "0001001" when "01011010111010010", -- t[46546] = 9
      "0001001" when "01011010111010011", -- t[46547] = 9
      "0001001" when "01011010111010100", -- t[46548] = 9
      "0001001" when "01011010111010101", -- t[46549] = 9
      "0001001" when "01011010111010110", -- t[46550] = 9
      "0001001" when "01011010111010111", -- t[46551] = 9
      "0001001" when "01011010111011000", -- t[46552] = 9
      "0001001" when "01011010111011001", -- t[46553] = 9
      "0001001" when "01011010111011010", -- t[46554] = 9
      "0001001" when "01011010111011011", -- t[46555] = 9
      "0001001" when "01011010111011100", -- t[46556] = 9
      "0001001" when "01011010111011101", -- t[46557] = 9
      "0001001" when "01011010111011110", -- t[46558] = 9
      "0001001" when "01011010111011111", -- t[46559] = 9
      "0001001" when "01011010111100000", -- t[46560] = 9
      "0001001" when "01011010111100001", -- t[46561] = 9
      "0001001" when "01011010111100010", -- t[46562] = 9
      "0001001" when "01011010111100011", -- t[46563] = 9
      "0001001" when "01011010111100100", -- t[46564] = 9
      "0001001" when "01011010111100101", -- t[46565] = 9
      "0001001" when "01011010111100110", -- t[46566] = 9
      "0001001" when "01011010111100111", -- t[46567] = 9
      "0001001" when "01011010111101000", -- t[46568] = 9
      "0001001" when "01011010111101001", -- t[46569] = 9
      "0001001" when "01011010111101010", -- t[46570] = 9
      "0001001" when "01011010111101011", -- t[46571] = 9
      "0001001" when "01011010111101100", -- t[46572] = 9
      "0001001" when "01011010111101101", -- t[46573] = 9
      "0001001" when "01011010111101110", -- t[46574] = 9
      "0001001" when "01011010111101111", -- t[46575] = 9
      "0001001" when "01011010111110000", -- t[46576] = 9
      "0001001" when "01011010111110001", -- t[46577] = 9
      "0001001" when "01011010111110010", -- t[46578] = 9
      "0001001" when "01011010111110011", -- t[46579] = 9
      "0001001" when "01011010111110100", -- t[46580] = 9
      "0001001" when "01011010111110101", -- t[46581] = 9
      "0001001" when "01011010111110110", -- t[46582] = 9
      "0001001" when "01011010111110111", -- t[46583] = 9
      "0001001" when "01011010111111000", -- t[46584] = 9
      "0001001" when "01011010111111001", -- t[46585] = 9
      "0001001" when "01011010111111010", -- t[46586] = 9
      "0001001" when "01011010111111011", -- t[46587] = 9
      "0001001" when "01011010111111100", -- t[46588] = 9
      "0001001" when "01011010111111101", -- t[46589] = 9
      "0001001" when "01011010111111110", -- t[46590] = 9
      "0001001" when "01011010111111111", -- t[46591] = 9
      "0001001" when "01011011000000000", -- t[46592] = 9
      "0001001" when "01011011000000001", -- t[46593] = 9
      "0001001" when "01011011000000010", -- t[46594] = 9
      "0001001" when "01011011000000011", -- t[46595] = 9
      "0001001" when "01011011000000100", -- t[46596] = 9
      "0001001" when "01011011000000101", -- t[46597] = 9
      "0001001" when "01011011000000110", -- t[46598] = 9
      "0001001" when "01011011000000111", -- t[46599] = 9
      "0001001" when "01011011000001000", -- t[46600] = 9
      "0001001" when "01011011000001001", -- t[46601] = 9
      "0001001" when "01011011000001010", -- t[46602] = 9
      "0001001" when "01011011000001011", -- t[46603] = 9
      "0001001" when "01011011000001100", -- t[46604] = 9
      "0001001" when "01011011000001101", -- t[46605] = 9
      "0001001" when "01011011000001110", -- t[46606] = 9
      "0001001" when "01011011000001111", -- t[46607] = 9
      "0001001" when "01011011000010000", -- t[46608] = 9
      "0001001" when "01011011000010001", -- t[46609] = 9
      "0001001" when "01011011000010010", -- t[46610] = 9
      "0001001" when "01011011000010011", -- t[46611] = 9
      "0001001" when "01011011000010100", -- t[46612] = 9
      "0001001" when "01011011000010101", -- t[46613] = 9
      "0001001" when "01011011000010110", -- t[46614] = 9
      "0001001" when "01011011000010111", -- t[46615] = 9
      "0001001" when "01011011000011000", -- t[46616] = 9
      "0001001" when "01011011000011001", -- t[46617] = 9
      "0001001" when "01011011000011010", -- t[46618] = 9
      "0001001" when "01011011000011011", -- t[46619] = 9
      "0001001" when "01011011000011100", -- t[46620] = 9
      "0001001" when "01011011000011101", -- t[46621] = 9
      "0001001" when "01011011000011110", -- t[46622] = 9
      "0001001" when "01011011000011111", -- t[46623] = 9
      "0001001" when "01011011000100000", -- t[46624] = 9
      "0001001" when "01011011000100001", -- t[46625] = 9
      "0001001" when "01011011000100010", -- t[46626] = 9
      "0001001" when "01011011000100011", -- t[46627] = 9
      "0001001" when "01011011000100100", -- t[46628] = 9
      "0001001" when "01011011000100101", -- t[46629] = 9
      "0001001" when "01011011000100110", -- t[46630] = 9
      "0001001" when "01011011000100111", -- t[46631] = 9
      "0001001" when "01011011000101000", -- t[46632] = 9
      "0001001" when "01011011000101001", -- t[46633] = 9
      "0001001" when "01011011000101010", -- t[46634] = 9
      "0001001" when "01011011000101011", -- t[46635] = 9
      "0001001" when "01011011000101100", -- t[46636] = 9
      "0001001" when "01011011000101101", -- t[46637] = 9
      "0001001" when "01011011000101110", -- t[46638] = 9
      "0001001" when "01011011000101111", -- t[46639] = 9
      "0001001" when "01011011000110000", -- t[46640] = 9
      "0001001" when "01011011000110001", -- t[46641] = 9
      "0001001" when "01011011000110010", -- t[46642] = 9
      "0001001" when "01011011000110011", -- t[46643] = 9
      "0001001" when "01011011000110100", -- t[46644] = 9
      "0001001" when "01011011000110101", -- t[46645] = 9
      "0001001" when "01011011000110110", -- t[46646] = 9
      "0001001" when "01011011000110111", -- t[46647] = 9
      "0001001" when "01011011000111000", -- t[46648] = 9
      "0001001" when "01011011000111001", -- t[46649] = 9
      "0001001" when "01011011000111010", -- t[46650] = 9
      "0001001" when "01011011000111011", -- t[46651] = 9
      "0001001" when "01011011000111100", -- t[46652] = 9
      "0001001" when "01011011000111101", -- t[46653] = 9
      "0001001" when "01011011000111110", -- t[46654] = 9
      "0001001" when "01011011000111111", -- t[46655] = 9
      "0001001" when "01011011001000000", -- t[46656] = 9
      "0001001" when "01011011001000001", -- t[46657] = 9
      "0001001" when "01011011001000010", -- t[46658] = 9
      "0001001" when "01011011001000011", -- t[46659] = 9
      "0001001" when "01011011001000100", -- t[46660] = 9
      "0001001" when "01011011001000101", -- t[46661] = 9
      "0001001" when "01011011001000110", -- t[46662] = 9
      "0001001" when "01011011001000111", -- t[46663] = 9
      "0001001" when "01011011001001000", -- t[46664] = 9
      "0001001" when "01011011001001001", -- t[46665] = 9
      "0001001" when "01011011001001010", -- t[46666] = 9
      "0001001" when "01011011001001011", -- t[46667] = 9
      "0001001" when "01011011001001100", -- t[46668] = 9
      "0001001" when "01011011001001101", -- t[46669] = 9
      "0001001" when "01011011001001110", -- t[46670] = 9
      "0001001" when "01011011001001111", -- t[46671] = 9
      "0001001" when "01011011001010000", -- t[46672] = 9
      "0001001" when "01011011001010001", -- t[46673] = 9
      "0001001" when "01011011001010010", -- t[46674] = 9
      "0001001" when "01011011001010011", -- t[46675] = 9
      "0001001" when "01011011001010100", -- t[46676] = 9
      "0001001" when "01011011001010101", -- t[46677] = 9
      "0001001" when "01011011001010110", -- t[46678] = 9
      "0001001" when "01011011001010111", -- t[46679] = 9
      "0001001" when "01011011001011000", -- t[46680] = 9
      "0001001" when "01011011001011001", -- t[46681] = 9
      "0001001" when "01011011001011010", -- t[46682] = 9
      "0001001" when "01011011001011011", -- t[46683] = 9
      "0001001" when "01011011001011100", -- t[46684] = 9
      "0001001" when "01011011001011101", -- t[46685] = 9
      "0001001" when "01011011001011110", -- t[46686] = 9
      "0001001" when "01011011001011111", -- t[46687] = 9
      "0001001" when "01011011001100000", -- t[46688] = 9
      "0001001" when "01011011001100001", -- t[46689] = 9
      "0001001" when "01011011001100010", -- t[46690] = 9
      "0001001" when "01011011001100011", -- t[46691] = 9
      "0001001" when "01011011001100100", -- t[46692] = 9
      "0001001" when "01011011001100101", -- t[46693] = 9
      "0001001" when "01011011001100110", -- t[46694] = 9
      "0001001" when "01011011001100111", -- t[46695] = 9
      "0001001" when "01011011001101000", -- t[46696] = 9
      "0001001" when "01011011001101001", -- t[46697] = 9
      "0001001" when "01011011001101010", -- t[46698] = 9
      "0001001" when "01011011001101011", -- t[46699] = 9
      "0001001" when "01011011001101100", -- t[46700] = 9
      "0001001" when "01011011001101101", -- t[46701] = 9
      "0001001" when "01011011001101110", -- t[46702] = 9
      "0001001" when "01011011001101111", -- t[46703] = 9
      "0001001" when "01011011001110000", -- t[46704] = 9
      "0001001" when "01011011001110001", -- t[46705] = 9
      "0001001" when "01011011001110010", -- t[46706] = 9
      "0001001" when "01011011001110011", -- t[46707] = 9
      "0001001" when "01011011001110100", -- t[46708] = 9
      "0001001" when "01011011001110101", -- t[46709] = 9
      "0001001" when "01011011001110110", -- t[46710] = 9
      "0001001" when "01011011001110111", -- t[46711] = 9
      "0001001" when "01011011001111000", -- t[46712] = 9
      "0001001" when "01011011001111001", -- t[46713] = 9
      "0001001" when "01011011001111010", -- t[46714] = 9
      "0001001" when "01011011001111011", -- t[46715] = 9
      "0001001" when "01011011001111100", -- t[46716] = 9
      "0001001" when "01011011001111101", -- t[46717] = 9
      "0001001" when "01011011001111110", -- t[46718] = 9
      "0001001" when "01011011001111111", -- t[46719] = 9
      "0001001" when "01011011010000000", -- t[46720] = 9
      "0001001" when "01011011010000001", -- t[46721] = 9
      "0001001" when "01011011010000010", -- t[46722] = 9
      "0001001" when "01011011010000011", -- t[46723] = 9
      "0001001" when "01011011010000100", -- t[46724] = 9
      "0001001" when "01011011010000101", -- t[46725] = 9
      "0001001" when "01011011010000110", -- t[46726] = 9
      "0001001" when "01011011010000111", -- t[46727] = 9
      "0001001" when "01011011010001000", -- t[46728] = 9
      "0001001" when "01011011010001001", -- t[46729] = 9
      "0001001" when "01011011010001010", -- t[46730] = 9
      "0001001" when "01011011010001011", -- t[46731] = 9
      "0001001" when "01011011010001100", -- t[46732] = 9
      "0001001" when "01011011010001101", -- t[46733] = 9
      "0001001" when "01011011010001110", -- t[46734] = 9
      "0001001" when "01011011010001111", -- t[46735] = 9
      "0001001" when "01011011010010000", -- t[46736] = 9
      "0001001" when "01011011010010001", -- t[46737] = 9
      "0001001" when "01011011010010010", -- t[46738] = 9
      "0001001" when "01011011010010011", -- t[46739] = 9
      "0001001" when "01011011010010100", -- t[46740] = 9
      "0001001" when "01011011010010101", -- t[46741] = 9
      "0001001" when "01011011010010110", -- t[46742] = 9
      "0001001" when "01011011010010111", -- t[46743] = 9
      "0001001" when "01011011010011000", -- t[46744] = 9
      "0001001" when "01011011010011001", -- t[46745] = 9
      "0001001" when "01011011010011010", -- t[46746] = 9
      "0001001" when "01011011010011011", -- t[46747] = 9
      "0001001" when "01011011010011100", -- t[46748] = 9
      "0001001" when "01011011010011101", -- t[46749] = 9
      "0001001" when "01011011010011110", -- t[46750] = 9
      "0001001" when "01011011010011111", -- t[46751] = 9
      "0001001" when "01011011010100000", -- t[46752] = 9
      "0001001" when "01011011010100001", -- t[46753] = 9
      "0001001" when "01011011010100010", -- t[46754] = 9
      "0001001" when "01011011010100011", -- t[46755] = 9
      "0001001" when "01011011010100100", -- t[46756] = 9
      "0001001" when "01011011010100101", -- t[46757] = 9
      "0001001" when "01011011010100110", -- t[46758] = 9
      "0001001" when "01011011010100111", -- t[46759] = 9
      "0001001" when "01011011010101000", -- t[46760] = 9
      "0001001" when "01011011010101001", -- t[46761] = 9
      "0001001" when "01011011010101010", -- t[46762] = 9
      "0001001" when "01011011010101011", -- t[46763] = 9
      "0001001" when "01011011010101100", -- t[46764] = 9
      "0001001" when "01011011010101101", -- t[46765] = 9
      "0001001" when "01011011010101110", -- t[46766] = 9
      "0001001" when "01011011010101111", -- t[46767] = 9
      "0001001" when "01011011010110000", -- t[46768] = 9
      "0001001" when "01011011010110001", -- t[46769] = 9
      "0001001" when "01011011010110010", -- t[46770] = 9
      "0001001" when "01011011010110011", -- t[46771] = 9
      "0001001" when "01011011010110100", -- t[46772] = 9
      "0001001" when "01011011010110101", -- t[46773] = 9
      "0001001" when "01011011010110110", -- t[46774] = 9
      "0001001" when "01011011010110111", -- t[46775] = 9
      "0001001" when "01011011010111000", -- t[46776] = 9
      "0001001" when "01011011010111001", -- t[46777] = 9
      "0001001" when "01011011010111010", -- t[46778] = 9
      "0001001" when "01011011010111011", -- t[46779] = 9
      "0001001" when "01011011010111100", -- t[46780] = 9
      "0001001" when "01011011010111101", -- t[46781] = 9
      "0001001" when "01011011010111110", -- t[46782] = 9
      "0001001" when "01011011010111111", -- t[46783] = 9
      "0001001" when "01011011011000000", -- t[46784] = 9
      "0001001" when "01011011011000001", -- t[46785] = 9
      "0001001" when "01011011011000010", -- t[46786] = 9
      "0001001" when "01011011011000011", -- t[46787] = 9
      "0001001" when "01011011011000100", -- t[46788] = 9
      "0001001" when "01011011011000101", -- t[46789] = 9
      "0001001" when "01011011011000110", -- t[46790] = 9
      "0001001" when "01011011011000111", -- t[46791] = 9
      "0001001" when "01011011011001000", -- t[46792] = 9
      "0001001" when "01011011011001001", -- t[46793] = 9
      "0001001" when "01011011011001010", -- t[46794] = 9
      "0001001" when "01011011011001011", -- t[46795] = 9
      "0001001" when "01011011011001100", -- t[46796] = 9
      "0001001" when "01011011011001101", -- t[46797] = 9
      "0001001" when "01011011011001110", -- t[46798] = 9
      "0001001" when "01011011011001111", -- t[46799] = 9
      "0001001" when "01011011011010000", -- t[46800] = 9
      "0001001" when "01011011011010001", -- t[46801] = 9
      "0001001" when "01011011011010010", -- t[46802] = 9
      "0001001" when "01011011011010011", -- t[46803] = 9
      "0001001" when "01011011011010100", -- t[46804] = 9
      "0001001" when "01011011011010101", -- t[46805] = 9
      "0001001" when "01011011011010110", -- t[46806] = 9
      "0001001" when "01011011011010111", -- t[46807] = 9
      "0001001" when "01011011011011000", -- t[46808] = 9
      "0001001" when "01011011011011001", -- t[46809] = 9
      "0001001" when "01011011011011010", -- t[46810] = 9
      "0001001" when "01011011011011011", -- t[46811] = 9
      "0001001" when "01011011011011100", -- t[46812] = 9
      "0001001" when "01011011011011101", -- t[46813] = 9
      "0001001" when "01011011011011110", -- t[46814] = 9
      "0001001" when "01011011011011111", -- t[46815] = 9
      "0001001" when "01011011011100000", -- t[46816] = 9
      "0001001" when "01011011011100001", -- t[46817] = 9
      "0001001" when "01011011011100010", -- t[46818] = 9
      "0001001" when "01011011011100011", -- t[46819] = 9
      "0001001" when "01011011011100100", -- t[46820] = 9
      "0001001" when "01011011011100101", -- t[46821] = 9
      "0001001" when "01011011011100110", -- t[46822] = 9
      "0001001" when "01011011011100111", -- t[46823] = 9
      "0001001" when "01011011011101000", -- t[46824] = 9
      "0001001" when "01011011011101001", -- t[46825] = 9
      "0001001" when "01011011011101010", -- t[46826] = 9
      "0001001" when "01011011011101011", -- t[46827] = 9
      "0001001" when "01011011011101100", -- t[46828] = 9
      "0001001" when "01011011011101101", -- t[46829] = 9
      "0001001" when "01011011011101110", -- t[46830] = 9
      "0001001" when "01011011011101111", -- t[46831] = 9
      "0001001" when "01011011011110000", -- t[46832] = 9
      "0001001" when "01011011011110001", -- t[46833] = 9
      "0001001" when "01011011011110010", -- t[46834] = 9
      "0001001" when "01011011011110011", -- t[46835] = 9
      "0001001" when "01011011011110100", -- t[46836] = 9
      "0001001" when "01011011011110101", -- t[46837] = 9
      "0001001" when "01011011011110110", -- t[46838] = 9
      "0001001" when "01011011011110111", -- t[46839] = 9
      "0001001" when "01011011011111000", -- t[46840] = 9
      "0001001" when "01011011011111001", -- t[46841] = 9
      "0001001" when "01011011011111010", -- t[46842] = 9
      "0001001" when "01011011011111011", -- t[46843] = 9
      "0001001" when "01011011011111100", -- t[46844] = 9
      "0001001" when "01011011011111101", -- t[46845] = 9
      "0001001" when "01011011011111110", -- t[46846] = 9
      "0001010" when "01011011011111111", -- t[46847] = 10
      "0001010" when "01011011100000000", -- t[46848] = 10
      "0001010" when "01011011100000001", -- t[46849] = 10
      "0001010" when "01011011100000010", -- t[46850] = 10
      "0001010" when "01011011100000011", -- t[46851] = 10
      "0001010" when "01011011100000100", -- t[46852] = 10
      "0001010" when "01011011100000101", -- t[46853] = 10
      "0001010" when "01011011100000110", -- t[46854] = 10
      "0001010" when "01011011100000111", -- t[46855] = 10
      "0001010" when "01011011100001000", -- t[46856] = 10
      "0001010" when "01011011100001001", -- t[46857] = 10
      "0001010" when "01011011100001010", -- t[46858] = 10
      "0001010" when "01011011100001011", -- t[46859] = 10
      "0001010" when "01011011100001100", -- t[46860] = 10
      "0001010" when "01011011100001101", -- t[46861] = 10
      "0001010" when "01011011100001110", -- t[46862] = 10
      "0001010" when "01011011100001111", -- t[46863] = 10
      "0001010" when "01011011100010000", -- t[46864] = 10
      "0001010" when "01011011100010001", -- t[46865] = 10
      "0001010" when "01011011100010010", -- t[46866] = 10
      "0001010" when "01011011100010011", -- t[46867] = 10
      "0001010" when "01011011100010100", -- t[46868] = 10
      "0001010" when "01011011100010101", -- t[46869] = 10
      "0001010" when "01011011100010110", -- t[46870] = 10
      "0001010" when "01011011100010111", -- t[46871] = 10
      "0001010" when "01011011100011000", -- t[46872] = 10
      "0001010" when "01011011100011001", -- t[46873] = 10
      "0001010" when "01011011100011010", -- t[46874] = 10
      "0001010" when "01011011100011011", -- t[46875] = 10
      "0001010" when "01011011100011100", -- t[46876] = 10
      "0001010" when "01011011100011101", -- t[46877] = 10
      "0001010" when "01011011100011110", -- t[46878] = 10
      "0001010" when "01011011100011111", -- t[46879] = 10
      "0001010" when "01011011100100000", -- t[46880] = 10
      "0001010" when "01011011100100001", -- t[46881] = 10
      "0001010" when "01011011100100010", -- t[46882] = 10
      "0001010" when "01011011100100011", -- t[46883] = 10
      "0001010" when "01011011100100100", -- t[46884] = 10
      "0001010" when "01011011100100101", -- t[46885] = 10
      "0001010" when "01011011100100110", -- t[46886] = 10
      "0001010" when "01011011100100111", -- t[46887] = 10
      "0001010" when "01011011100101000", -- t[46888] = 10
      "0001010" when "01011011100101001", -- t[46889] = 10
      "0001010" when "01011011100101010", -- t[46890] = 10
      "0001010" when "01011011100101011", -- t[46891] = 10
      "0001010" when "01011011100101100", -- t[46892] = 10
      "0001010" when "01011011100101101", -- t[46893] = 10
      "0001010" when "01011011100101110", -- t[46894] = 10
      "0001010" when "01011011100101111", -- t[46895] = 10
      "0001010" when "01011011100110000", -- t[46896] = 10
      "0001010" when "01011011100110001", -- t[46897] = 10
      "0001010" when "01011011100110010", -- t[46898] = 10
      "0001010" when "01011011100110011", -- t[46899] = 10
      "0001010" when "01011011100110100", -- t[46900] = 10
      "0001010" when "01011011100110101", -- t[46901] = 10
      "0001010" when "01011011100110110", -- t[46902] = 10
      "0001010" when "01011011100110111", -- t[46903] = 10
      "0001010" when "01011011100111000", -- t[46904] = 10
      "0001010" when "01011011100111001", -- t[46905] = 10
      "0001010" when "01011011100111010", -- t[46906] = 10
      "0001010" when "01011011100111011", -- t[46907] = 10
      "0001010" when "01011011100111100", -- t[46908] = 10
      "0001010" when "01011011100111101", -- t[46909] = 10
      "0001010" when "01011011100111110", -- t[46910] = 10
      "0001010" when "01011011100111111", -- t[46911] = 10
      "0001010" when "01011011101000000", -- t[46912] = 10
      "0001010" when "01011011101000001", -- t[46913] = 10
      "0001010" when "01011011101000010", -- t[46914] = 10
      "0001010" when "01011011101000011", -- t[46915] = 10
      "0001010" when "01011011101000100", -- t[46916] = 10
      "0001010" when "01011011101000101", -- t[46917] = 10
      "0001010" when "01011011101000110", -- t[46918] = 10
      "0001010" when "01011011101000111", -- t[46919] = 10
      "0001010" when "01011011101001000", -- t[46920] = 10
      "0001010" when "01011011101001001", -- t[46921] = 10
      "0001010" when "01011011101001010", -- t[46922] = 10
      "0001010" when "01011011101001011", -- t[46923] = 10
      "0001010" when "01011011101001100", -- t[46924] = 10
      "0001010" when "01011011101001101", -- t[46925] = 10
      "0001010" when "01011011101001110", -- t[46926] = 10
      "0001010" when "01011011101001111", -- t[46927] = 10
      "0001010" when "01011011101010000", -- t[46928] = 10
      "0001010" when "01011011101010001", -- t[46929] = 10
      "0001010" when "01011011101010010", -- t[46930] = 10
      "0001010" when "01011011101010011", -- t[46931] = 10
      "0001010" when "01011011101010100", -- t[46932] = 10
      "0001010" when "01011011101010101", -- t[46933] = 10
      "0001010" when "01011011101010110", -- t[46934] = 10
      "0001010" when "01011011101010111", -- t[46935] = 10
      "0001010" when "01011011101011000", -- t[46936] = 10
      "0001010" when "01011011101011001", -- t[46937] = 10
      "0001010" when "01011011101011010", -- t[46938] = 10
      "0001010" when "01011011101011011", -- t[46939] = 10
      "0001010" when "01011011101011100", -- t[46940] = 10
      "0001010" when "01011011101011101", -- t[46941] = 10
      "0001010" when "01011011101011110", -- t[46942] = 10
      "0001010" when "01011011101011111", -- t[46943] = 10
      "0001010" when "01011011101100000", -- t[46944] = 10
      "0001010" when "01011011101100001", -- t[46945] = 10
      "0001010" when "01011011101100010", -- t[46946] = 10
      "0001010" when "01011011101100011", -- t[46947] = 10
      "0001010" when "01011011101100100", -- t[46948] = 10
      "0001010" when "01011011101100101", -- t[46949] = 10
      "0001010" when "01011011101100110", -- t[46950] = 10
      "0001010" when "01011011101100111", -- t[46951] = 10
      "0001010" when "01011011101101000", -- t[46952] = 10
      "0001010" when "01011011101101001", -- t[46953] = 10
      "0001010" when "01011011101101010", -- t[46954] = 10
      "0001010" when "01011011101101011", -- t[46955] = 10
      "0001010" when "01011011101101100", -- t[46956] = 10
      "0001010" when "01011011101101101", -- t[46957] = 10
      "0001010" when "01011011101101110", -- t[46958] = 10
      "0001010" when "01011011101101111", -- t[46959] = 10
      "0001010" when "01011011101110000", -- t[46960] = 10
      "0001010" when "01011011101110001", -- t[46961] = 10
      "0001010" when "01011011101110010", -- t[46962] = 10
      "0001010" when "01011011101110011", -- t[46963] = 10
      "0001010" when "01011011101110100", -- t[46964] = 10
      "0001010" when "01011011101110101", -- t[46965] = 10
      "0001010" when "01011011101110110", -- t[46966] = 10
      "0001010" when "01011011101110111", -- t[46967] = 10
      "0001010" when "01011011101111000", -- t[46968] = 10
      "0001010" when "01011011101111001", -- t[46969] = 10
      "0001010" when "01011011101111010", -- t[46970] = 10
      "0001010" when "01011011101111011", -- t[46971] = 10
      "0001010" when "01011011101111100", -- t[46972] = 10
      "0001010" when "01011011101111101", -- t[46973] = 10
      "0001010" when "01011011101111110", -- t[46974] = 10
      "0001010" when "01011011101111111", -- t[46975] = 10
      "0001010" when "01011011110000000", -- t[46976] = 10
      "0001010" when "01011011110000001", -- t[46977] = 10
      "0001010" when "01011011110000010", -- t[46978] = 10
      "0001010" when "01011011110000011", -- t[46979] = 10
      "0001010" when "01011011110000100", -- t[46980] = 10
      "0001010" when "01011011110000101", -- t[46981] = 10
      "0001010" when "01011011110000110", -- t[46982] = 10
      "0001010" when "01011011110000111", -- t[46983] = 10
      "0001010" when "01011011110001000", -- t[46984] = 10
      "0001010" when "01011011110001001", -- t[46985] = 10
      "0001010" when "01011011110001010", -- t[46986] = 10
      "0001010" when "01011011110001011", -- t[46987] = 10
      "0001010" when "01011011110001100", -- t[46988] = 10
      "0001010" when "01011011110001101", -- t[46989] = 10
      "0001010" when "01011011110001110", -- t[46990] = 10
      "0001010" when "01011011110001111", -- t[46991] = 10
      "0001010" when "01011011110010000", -- t[46992] = 10
      "0001010" when "01011011110010001", -- t[46993] = 10
      "0001010" when "01011011110010010", -- t[46994] = 10
      "0001010" when "01011011110010011", -- t[46995] = 10
      "0001010" when "01011011110010100", -- t[46996] = 10
      "0001010" when "01011011110010101", -- t[46997] = 10
      "0001010" when "01011011110010110", -- t[46998] = 10
      "0001010" when "01011011110010111", -- t[46999] = 10
      "0001010" when "01011011110011000", -- t[47000] = 10
      "0001010" when "01011011110011001", -- t[47001] = 10
      "0001010" when "01011011110011010", -- t[47002] = 10
      "0001010" when "01011011110011011", -- t[47003] = 10
      "0001010" when "01011011110011100", -- t[47004] = 10
      "0001010" when "01011011110011101", -- t[47005] = 10
      "0001010" when "01011011110011110", -- t[47006] = 10
      "0001010" when "01011011110011111", -- t[47007] = 10
      "0001010" when "01011011110100000", -- t[47008] = 10
      "0001010" when "01011011110100001", -- t[47009] = 10
      "0001010" when "01011011110100010", -- t[47010] = 10
      "0001010" when "01011011110100011", -- t[47011] = 10
      "0001010" when "01011011110100100", -- t[47012] = 10
      "0001010" when "01011011110100101", -- t[47013] = 10
      "0001010" when "01011011110100110", -- t[47014] = 10
      "0001010" when "01011011110100111", -- t[47015] = 10
      "0001010" when "01011011110101000", -- t[47016] = 10
      "0001010" when "01011011110101001", -- t[47017] = 10
      "0001010" when "01011011110101010", -- t[47018] = 10
      "0001010" when "01011011110101011", -- t[47019] = 10
      "0001010" when "01011011110101100", -- t[47020] = 10
      "0001010" when "01011011110101101", -- t[47021] = 10
      "0001010" when "01011011110101110", -- t[47022] = 10
      "0001010" when "01011011110101111", -- t[47023] = 10
      "0001010" when "01011011110110000", -- t[47024] = 10
      "0001010" when "01011011110110001", -- t[47025] = 10
      "0001010" when "01011011110110010", -- t[47026] = 10
      "0001010" when "01011011110110011", -- t[47027] = 10
      "0001010" when "01011011110110100", -- t[47028] = 10
      "0001010" when "01011011110110101", -- t[47029] = 10
      "0001010" when "01011011110110110", -- t[47030] = 10
      "0001010" when "01011011110110111", -- t[47031] = 10
      "0001010" when "01011011110111000", -- t[47032] = 10
      "0001010" when "01011011110111001", -- t[47033] = 10
      "0001010" when "01011011110111010", -- t[47034] = 10
      "0001010" when "01011011110111011", -- t[47035] = 10
      "0001010" when "01011011110111100", -- t[47036] = 10
      "0001010" when "01011011110111101", -- t[47037] = 10
      "0001010" when "01011011110111110", -- t[47038] = 10
      "0001010" when "01011011110111111", -- t[47039] = 10
      "0001010" when "01011011111000000", -- t[47040] = 10
      "0001010" when "01011011111000001", -- t[47041] = 10
      "0001010" when "01011011111000010", -- t[47042] = 10
      "0001010" when "01011011111000011", -- t[47043] = 10
      "0001010" when "01011011111000100", -- t[47044] = 10
      "0001010" when "01011011111000101", -- t[47045] = 10
      "0001010" when "01011011111000110", -- t[47046] = 10
      "0001010" when "01011011111000111", -- t[47047] = 10
      "0001010" when "01011011111001000", -- t[47048] = 10
      "0001010" when "01011011111001001", -- t[47049] = 10
      "0001010" when "01011011111001010", -- t[47050] = 10
      "0001010" when "01011011111001011", -- t[47051] = 10
      "0001010" when "01011011111001100", -- t[47052] = 10
      "0001010" when "01011011111001101", -- t[47053] = 10
      "0001010" when "01011011111001110", -- t[47054] = 10
      "0001010" when "01011011111001111", -- t[47055] = 10
      "0001010" when "01011011111010000", -- t[47056] = 10
      "0001010" when "01011011111010001", -- t[47057] = 10
      "0001010" when "01011011111010010", -- t[47058] = 10
      "0001010" when "01011011111010011", -- t[47059] = 10
      "0001010" when "01011011111010100", -- t[47060] = 10
      "0001010" when "01011011111010101", -- t[47061] = 10
      "0001010" when "01011011111010110", -- t[47062] = 10
      "0001010" when "01011011111010111", -- t[47063] = 10
      "0001010" when "01011011111011000", -- t[47064] = 10
      "0001010" when "01011011111011001", -- t[47065] = 10
      "0001010" when "01011011111011010", -- t[47066] = 10
      "0001010" when "01011011111011011", -- t[47067] = 10
      "0001010" when "01011011111011100", -- t[47068] = 10
      "0001010" when "01011011111011101", -- t[47069] = 10
      "0001010" when "01011011111011110", -- t[47070] = 10
      "0001010" when "01011011111011111", -- t[47071] = 10
      "0001010" when "01011011111100000", -- t[47072] = 10
      "0001010" when "01011011111100001", -- t[47073] = 10
      "0001010" when "01011011111100010", -- t[47074] = 10
      "0001010" when "01011011111100011", -- t[47075] = 10
      "0001010" when "01011011111100100", -- t[47076] = 10
      "0001010" when "01011011111100101", -- t[47077] = 10
      "0001010" when "01011011111100110", -- t[47078] = 10
      "0001010" when "01011011111100111", -- t[47079] = 10
      "0001010" when "01011011111101000", -- t[47080] = 10
      "0001010" when "01011011111101001", -- t[47081] = 10
      "0001010" when "01011011111101010", -- t[47082] = 10
      "0001010" when "01011011111101011", -- t[47083] = 10
      "0001010" when "01011011111101100", -- t[47084] = 10
      "0001010" when "01011011111101101", -- t[47085] = 10
      "0001010" when "01011011111101110", -- t[47086] = 10
      "0001010" when "01011011111101111", -- t[47087] = 10
      "0001010" when "01011011111110000", -- t[47088] = 10
      "0001010" when "01011011111110001", -- t[47089] = 10
      "0001010" when "01011011111110010", -- t[47090] = 10
      "0001010" when "01011011111110011", -- t[47091] = 10
      "0001010" when "01011011111110100", -- t[47092] = 10
      "0001010" when "01011011111110101", -- t[47093] = 10
      "0001010" when "01011011111110110", -- t[47094] = 10
      "0001010" when "01011011111110111", -- t[47095] = 10
      "0001010" when "01011011111111000", -- t[47096] = 10
      "0001010" when "01011011111111001", -- t[47097] = 10
      "0001010" when "01011011111111010", -- t[47098] = 10
      "0001010" when "01011011111111011", -- t[47099] = 10
      "0001010" when "01011011111111100", -- t[47100] = 10
      "0001010" when "01011011111111101", -- t[47101] = 10
      "0001010" when "01011011111111110", -- t[47102] = 10
      "0001010" when "01011011111111111", -- t[47103] = 10
      "0001010" when "01011100000000000", -- t[47104] = 10
      "0001010" when "01011100000000001", -- t[47105] = 10
      "0001010" when "01011100000000010", -- t[47106] = 10
      "0001010" when "01011100000000011", -- t[47107] = 10
      "0001010" when "01011100000000100", -- t[47108] = 10
      "0001010" when "01011100000000101", -- t[47109] = 10
      "0001010" when "01011100000000110", -- t[47110] = 10
      "0001010" when "01011100000000111", -- t[47111] = 10
      "0001010" when "01011100000001000", -- t[47112] = 10
      "0001010" when "01011100000001001", -- t[47113] = 10
      "0001010" when "01011100000001010", -- t[47114] = 10
      "0001010" when "01011100000001011", -- t[47115] = 10
      "0001010" when "01011100000001100", -- t[47116] = 10
      "0001010" when "01011100000001101", -- t[47117] = 10
      "0001010" when "01011100000001110", -- t[47118] = 10
      "0001010" when "01011100000001111", -- t[47119] = 10
      "0001010" when "01011100000010000", -- t[47120] = 10
      "0001010" when "01011100000010001", -- t[47121] = 10
      "0001010" when "01011100000010010", -- t[47122] = 10
      "0001010" when "01011100000010011", -- t[47123] = 10
      "0001010" when "01011100000010100", -- t[47124] = 10
      "0001010" when "01011100000010101", -- t[47125] = 10
      "0001010" when "01011100000010110", -- t[47126] = 10
      "0001010" when "01011100000010111", -- t[47127] = 10
      "0001010" when "01011100000011000", -- t[47128] = 10
      "0001010" when "01011100000011001", -- t[47129] = 10
      "0001010" when "01011100000011010", -- t[47130] = 10
      "0001010" when "01011100000011011", -- t[47131] = 10
      "0001010" when "01011100000011100", -- t[47132] = 10
      "0001010" when "01011100000011101", -- t[47133] = 10
      "0001010" when "01011100000011110", -- t[47134] = 10
      "0001010" when "01011100000011111", -- t[47135] = 10
      "0001010" when "01011100000100000", -- t[47136] = 10
      "0001010" when "01011100000100001", -- t[47137] = 10
      "0001010" when "01011100000100010", -- t[47138] = 10
      "0001010" when "01011100000100011", -- t[47139] = 10
      "0001010" when "01011100000100100", -- t[47140] = 10
      "0001010" when "01011100000100101", -- t[47141] = 10
      "0001010" when "01011100000100110", -- t[47142] = 10
      "0001010" when "01011100000100111", -- t[47143] = 10
      "0001010" when "01011100000101000", -- t[47144] = 10
      "0001010" when "01011100000101001", -- t[47145] = 10
      "0001010" when "01011100000101010", -- t[47146] = 10
      "0001010" when "01011100000101011", -- t[47147] = 10
      "0001010" when "01011100000101100", -- t[47148] = 10
      "0001010" when "01011100000101101", -- t[47149] = 10
      "0001010" when "01011100000101110", -- t[47150] = 10
      "0001010" when "01011100000101111", -- t[47151] = 10
      "0001010" when "01011100000110000", -- t[47152] = 10
      "0001010" when "01011100000110001", -- t[47153] = 10
      "0001010" when "01011100000110010", -- t[47154] = 10
      "0001010" when "01011100000110011", -- t[47155] = 10
      "0001010" when "01011100000110100", -- t[47156] = 10
      "0001010" when "01011100000110101", -- t[47157] = 10
      "0001010" when "01011100000110110", -- t[47158] = 10
      "0001010" when "01011100000110111", -- t[47159] = 10
      "0001010" when "01011100000111000", -- t[47160] = 10
      "0001010" when "01011100000111001", -- t[47161] = 10
      "0001010" when "01011100000111010", -- t[47162] = 10
      "0001010" when "01011100000111011", -- t[47163] = 10
      "0001010" when "01011100000111100", -- t[47164] = 10
      "0001010" when "01011100000111101", -- t[47165] = 10
      "0001010" when "01011100000111110", -- t[47166] = 10
      "0001010" when "01011100000111111", -- t[47167] = 10
      "0001010" when "01011100001000000", -- t[47168] = 10
      "0001010" when "01011100001000001", -- t[47169] = 10
      "0001010" when "01011100001000010", -- t[47170] = 10
      "0001010" when "01011100001000011", -- t[47171] = 10
      "0001010" when "01011100001000100", -- t[47172] = 10
      "0001010" when "01011100001000101", -- t[47173] = 10
      "0001010" when "01011100001000110", -- t[47174] = 10
      "0001010" when "01011100001000111", -- t[47175] = 10
      "0001010" when "01011100001001000", -- t[47176] = 10
      "0001010" when "01011100001001001", -- t[47177] = 10
      "0001010" when "01011100001001010", -- t[47178] = 10
      "0001010" when "01011100001001011", -- t[47179] = 10
      "0001010" when "01011100001001100", -- t[47180] = 10
      "0001010" when "01011100001001101", -- t[47181] = 10
      "0001010" when "01011100001001110", -- t[47182] = 10
      "0001010" when "01011100001001111", -- t[47183] = 10
      "0001010" when "01011100001010000", -- t[47184] = 10
      "0001010" when "01011100001010001", -- t[47185] = 10
      "0001010" when "01011100001010010", -- t[47186] = 10
      "0001010" when "01011100001010011", -- t[47187] = 10
      "0001010" when "01011100001010100", -- t[47188] = 10
      "0001010" when "01011100001010101", -- t[47189] = 10
      "0001010" when "01011100001010110", -- t[47190] = 10
      "0001010" when "01011100001010111", -- t[47191] = 10
      "0001010" when "01011100001011000", -- t[47192] = 10
      "0001010" when "01011100001011001", -- t[47193] = 10
      "0001010" when "01011100001011010", -- t[47194] = 10
      "0001010" when "01011100001011011", -- t[47195] = 10
      "0001010" when "01011100001011100", -- t[47196] = 10
      "0001010" when "01011100001011101", -- t[47197] = 10
      "0001010" when "01011100001011110", -- t[47198] = 10
      "0001010" when "01011100001011111", -- t[47199] = 10
      "0001010" when "01011100001100000", -- t[47200] = 10
      "0001010" when "01011100001100001", -- t[47201] = 10
      "0001010" when "01011100001100010", -- t[47202] = 10
      "0001010" when "01011100001100011", -- t[47203] = 10
      "0001010" when "01011100001100100", -- t[47204] = 10
      "0001010" when "01011100001100101", -- t[47205] = 10
      "0001010" when "01011100001100110", -- t[47206] = 10
      "0001010" when "01011100001100111", -- t[47207] = 10
      "0001010" when "01011100001101000", -- t[47208] = 10
      "0001010" when "01011100001101001", -- t[47209] = 10
      "0001010" when "01011100001101010", -- t[47210] = 10
      "0001010" when "01011100001101011", -- t[47211] = 10
      "0001010" when "01011100001101100", -- t[47212] = 10
      "0001010" when "01011100001101101", -- t[47213] = 10
      "0001010" when "01011100001101110", -- t[47214] = 10
      "0001010" when "01011100001101111", -- t[47215] = 10
      "0001010" when "01011100001110000", -- t[47216] = 10
      "0001010" when "01011100001110001", -- t[47217] = 10
      "0001010" when "01011100001110010", -- t[47218] = 10
      "0001010" when "01011100001110011", -- t[47219] = 10
      "0001010" when "01011100001110100", -- t[47220] = 10
      "0001010" when "01011100001110101", -- t[47221] = 10
      "0001010" when "01011100001110110", -- t[47222] = 10
      "0001010" when "01011100001110111", -- t[47223] = 10
      "0001010" when "01011100001111000", -- t[47224] = 10
      "0001010" when "01011100001111001", -- t[47225] = 10
      "0001010" when "01011100001111010", -- t[47226] = 10
      "0001010" when "01011100001111011", -- t[47227] = 10
      "0001010" when "01011100001111100", -- t[47228] = 10
      "0001010" when "01011100001111101", -- t[47229] = 10
      "0001010" when "01011100001111110", -- t[47230] = 10
      "0001010" when "01011100001111111", -- t[47231] = 10
      "0001010" when "01011100010000000", -- t[47232] = 10
      "0001010" when "01011100010000001", -- t[47233] = 10
      "0001010" when "01011100010000010", -- t[47234] = 10
      "0001010" when "01011100010000011", -- t[47235] = 10
      "0001010" when "01011100010000100", -- t[47236] = 10
      "0001010" when "01011100010000101", -- t[47237] = 10
      "0001010" when "01011100010000110", -- t[47238] = 10
      "0001010" when "01011100010000111", -- t[47239] = 10
      "0001010" when "01011100010001000", -- t[47240] = 10
      "0001010" when "01011100010001001", -- t[47241] = 10
      "0001010" when "01011100010001010", -- t[47242] = 10
      "0001010" when "01011100010001011", -- t[47243] = 10
      "0001010" when "01011100010001100", -- t[47244] = 10
      "0001010" when "01011100010001101", -- t[47245] = 10
      "0001010" when "01011100010001110", -- t[47246] = 10
      "0001010" when "01011100010001111", -- t[47247] = 10
      "0001010" when "01011100010010000", -- t[47248] = 10
      "0001010" when "01011100010010001", -- t[47249] = 10
      "0001010" when "01011100010010010", -- t[47250] = 10
      "0001010" when "01011100010010011", -- t[47251] = 10
      "0001010" when "01011100010010100", -- t[47252] = 10
      "0001010" when "01011100010010101", -- t[47253] = 10
      "0001010" when "01011100010010110", -- t[47254] = 10
      "0001010" when "01011100010010111", -- t[47255] = 10
      "0001010" when "01011100010011000", -- t[47256] = 10
      "0001010" when "01011100010011001", -- t[47257] = 10
      "0001010" when "01011100010011010", -- t[47258] = 10
      "0001010" when "01011100010011011", -- t[47259] = 10
      "0001010" when "01011100010011100", -- t[47260] = 10
      "0001010" when "01011100010011101", -- t[47261] = 10
      "0001010" when "01011100010011110", -- t[47262] = 10
      "0001010" when "01011100010011111", -- t[47263] = 10
      "0001010" when "01011100010100000", -- t[47264] = 10
      "0001010" when "01011100010100001", -- t[47265] = 10
      "0001010" when "01011100010100010", -- t[47266] = 10
      "0001010" when "01011100010100011", -- t[47267] = 10
      "0001010" when "01011100010100100", -- t[47268] = 10
      "0001010" when "01011100010100101", -- t[47269] = 10
      "0001010" when "01011100010100110", -- t[47270] = 10
      "0001010" when "01011100010100111", -- t[47271] = 10
      "0001010" when "01011100010101000", -- t[47272] = 10
      "0001010" when "01011100010101001", -- t[47273] = 10
      "0001010" when "01011100010101010", -- t[47274] = 10
      "0001010" when "01011100010101011", -- t[47275] = 10
      "0001010" when "01011100010101100", -- t[47276] = 10
      "0001010" when "01011100010101101", -- t[47277] = 10
      "0001010" when "01011100010101110", -- t[47278] = 10
      "0001010" when "01011100010101111", -- t[47279] = 10
      "0001010" when "01011100010110000", -- t[47280] = 10
      "0001010" when "01011100010110001", -- t[47281] = 10
      "0001010" when "01011100010110010", -- t[47282] = 10
      "0001010" when "01011100010110011", -- t[47283] = 10
      "0001010" when "01011100010110100", -- t[47284] = 10
      "0001010" when "01011100010110101", -- t[47285] = 10
      "0001010" when "01011100010110110", -- t[47286] = 10
      "0001010" when "01011100010110111", -- t[47287] = 10
      "0001010" when "01011100010111000", -- t[47288] = 10
      "0001010" when "01011100010111001", -- t[47289] = 10
      "0001010" when "01011100010111010", -- t[47290] = 10
      "0001010" when "01011100010111011", -- t[47291] = 10
      "0001010" when "01011100010111100", -- t[47292] = 10
      "0001010" when "01011100010111101", -- t[47293] = 10
      "0001010" when "01011100010111110", -- t[47294] = 10
      "0001010" when "01011100010111111", -- t[47295] = 10
      "0001010" when "01011100011000000", -- t[47296] = 10
      "0001010" when "01011100011000001", -- t[47297] = 10
      "0001010" when "01011100011000010", -- t[47298] = 10
      "0001010" when "01011100011000011", -- t[47299] = 10
      "0001010" when "01011100011000100", -- t[47300] = 10
      "0001010" when "01011100011000101", -- t[47301] = 10
      "0001010" when "01011100011000110", -- t[47302] = 10
      "0001010" when "01011100011000111", -- t[47303] = 10
      "0001010" when "01011100011001000", -- t[47304] = 10
      "0001010" when "01011100011001001", -- t[47305] = 10
      "0001010" when "01011100011001010", -- t[47306] = 10
      "0001010" when "01011100011001011", -- t[47307] = 10
      "0001010" when "01011100011001100", -- t[47308] = 10
      "0001010" when "01011100011001101", -- t[47309] = 10
      "0001010" when "01011100011001110", -- t[47310] = 10
      "0001010" when "01011100011001111", -- t[47311] = 10
      "0001010" when "01011100011010000", -- t[47312] = 10
      "0001010" when "01011100011010001", -- t[47313] = 10
      "0001010" when "01011100011010010", -- t[47314] = 10
      "0001010" when "01011100011010011", -- t[47315] = 10
      "0001010" when "01011100011010100", -- t[47316] = 10
      "0001010" when "01011100011010101", -- t[47317] = 10
      "0001010" when "01011100011010110", -- t[47318] = 10
      "0001010" when "01011100011010111", -- t[47319] = 10
      "0001010" when "01011100011011000", -- t[47320] = 10
      "0001010" when "01011100011011001", -- t[47321] = 10
      "0001010" when "01011100011011010", -- t[47322] = 10
      "0001010" when "01011100011011011", -- t[47323] = 10
      "0001010" when "01011100011011100", -- t[47324] = 10
      "0001010" when "01011100011011101", -- t[47325] = 10
      "0001010" when "01011100011011110", -- t[47326] = 10
      "0001010" when "01011100011011111", -- t[47327] = 10
      "0001010" when "01011100011100000", -- t[47328] = 10
      "0001010" when "01011100011100001", -- t[47329] = 10
      "0001010" when "01011100011100010", -- t[47330] = 10
      "0001010" when "01011100011100011", -- t[47331] = 10
      "0001010" when "01011100011100100", -- t[47332] = 10
      "0001010" when "01011100011100101", -- t[47333] = 10
      "0001010" when "01011100011100110", -- t[47334] = 10
      "0001010" when "01011100011100111", -- t[47335] = 10
      "0001010" when "01011100011101000", -- t[47336] = 10
      "0001010" when "01011100011101001", -- t[47337] = 10
      "0001010" when "01011100011101010", -- t[47338] = 10
      "0001010" when "01011100011101011", -- t[47339] = 10
      "0001010" when "01011100011101100", -- t[47340] = 10
      "0001010" when "01011100011101101", -- t[47341] = 10
      "0001010" when "01011100011101110", -- t[47342] = 10
      "0001010" when "01011100011101111", -- t[47343] = 10
      "0001010" when "01011100011110000", -- t[47344] = 10
      "0001010" when "01011100011110001", -- t[47345] = 10
      "0001010" when "01011100011110010", -- t[47346] = 10
      "0001010" when "01011100011110011", -- t[47347] = 10
      "0001010" when "01011100011110100", -- t[47348] = 10
      "0001010" when "01011100011110101", -- t[47349] = 10
      "0001010" when "01011100011110110", -- t[47350] = 10
      "0001010" when "01011100011110111", -- t[47351] = 10
      "0001010" when "01011100011111000", -- t[47352] = 10
      "0001010" when "01011100011111001", -- t[47353] = 10
      "0001010" when "01011100011111010", -- t[47354] = 10
      "0001010" when "01011100011111011", -- t[47355] = 10
      "0001010" when "01011100011111100", -- t[47356] = 10
      "0001010" when "01011100011111101", -- t[47357] = 10
      "0001010" when "01011100011111110", -- t[47358] = 10
      "0001010" when "01011100011111111", -- t[47359] = 10
      "0001010" when "01011100100000000", -- t[47360] = 10
      "0001010" when "01011100100000001", -- t[47361] = 10
      "0001010" when "01011100100000010", -- t[47362] = 10
      "0001010" when "01011100100000011", -- t[47363] = 10
      "0001010" when "01011100100000100", -- t[47364] = 10
      "0001010" when "01011100100000101", -- t[47365] = 10
      "0001010" when "01011100100000110", -- t[47366] = 10
      "0001010" when "01011100100000111", -- t[47367] = 10
      "0001010" when "01011100100001000", -- t[47368] = 10
      "0001010" when "01011100100001001", -- t[47369] = 10
      "0001010" when "01011100100001010", -- t[47370] = 10
      "0001010" when "01011100100001011", -- t[47371] = 10
      "0001010" when "01011100100001100", -- t[47372] = 10
      "0001010" when "01011100100001101", -- t[47373] = 10
      "0001010" when "01011100100001110", -- t[47374] = 10
      "0001010" when "01011100100001111", -- t[47375] = 10
      "0001010" when "01011100100010000", -- t[47376] = 10
      "0001010" when "01011100100010001", -- t[47377] = 10
      "0001010" when "01011100100010010", -- t[47378] = 10
      "0001010" when "01011100100010011", -- t[47379] = 10
      "0001010" when "01011100100010100", -- t[47380] = 10
      "0001010" when "01011100100010101", -- t[47381] = 10
      "0001010" when "01011100100010110", -- t[47382] = 10
      "0001010" when "01011100100010111", -- t[47383] = 10
      "0001010" when "01011100100011000", -- t[47384] = 10
      "0001010" when "01011100100011001", -- t[47385] = 10
      "0001010" when "01011100100011010", -- t[47386] = 10
      "0001010" when "01011100100011011", -- t[47387] = 10
      "0001010" when "01011100100011100", -- t[47388] = 10
      "0001010" when "01011100100011101", -- t[47389] = 10
      "0001010" when "01011100100011110", -- t[47390] = 10
      "0001010" when "01011100100011111", -- t[47391] = 10
      "0001010" when "01011100100100000", -- t[47392] = 10
      "0001010" when "01011100100100001", -- t[47393] = 10
      "0001010" when "01011100100100010", -- t[47394] = 10
      "0001010" when "01011100100100011", -- t[47395] = 10
      "0001010" when "01011100100100100", -- t[47396] = 10
      "0001010" when "01011100100100101", -- t[47397] = 10
      "0001010" when "01011100100100110", -- t[47398] = 10
      "0001010" when "01011100100100111", -- t[47399] = 10
      "0001010" when "01011100100101000", -- t[47400] = 10
      "0001010" when "01011100100101001", -- t[47401] = 10
      "0001010" when "01011100100101010", -- t[47402] = 10
      "0001010" when "01011100100101011", -- t[47403] = 10
      "0001010" when "01011100100101100", -- t[47404] = 10
      "0001010" when "01011100100101101", -- t[47405] = 10
      "0001010" when "01011100100101110", -- t[47406] = 10
      "0001010" when "01011100100101111", -- t[47407] = 10
      "0001010" when "01011100100110000", -- t[47408] = 10
      "0001010" when "01011100100110001", -- t[47409] = 10
      "0001010" when "01011100100110010", -- t[47410] = 10
      "0001010" when "01011100100110011", -- t[47411] = 10
      "0001010" when "01011100100110100", -- t[47412] = 10
      "0001010" when "01011100100110101", -- t[47413] = 10
      "0001010" when "01011100100110110", -- t[47414] = 10
      "0001010" when "01011100100110111", -- t[47415] = 10
      "0001010" when "01011100100111000", -- t[47416] = 10
      "0001010" when "01011100100111001", -- t[47417] = 10
      "0001010" when "01011100100111010", -- t[47418] = 10
      "0001010" when "01011100100111011", -- t[47419] = 10
      "0001010" when "01011100100111100", -- t[47420] = 10
      "0001010" when "01011100100111101", -- t[47421] = 10
      "0001010" when "01011100100111110", -- t[47422] = 10
      "0001010" when "01011100100111111", -- t[47423] = 10
      "0001010" when "01011100101000000", -- t[47424] = 10
      "0001010" when "01011100101000001", -- t[47425] = 10
      "0001010" when "01011100101000010", -- t[47426] = 10
      "0001010" when "01011100101000011", -- t[47427] = 10
      "0001010" when "01011100101000100", -- t[47428] = 10
      "0001010" when "01011100101000101", -- t[47429] = 10
      "0001010" when "01011100101000110", -- t[47430] = 10
      "0001010" when "01011100101000111", -- t[47431] = 10
      "0001010" when "01011100101001000", -- t[47432] = 10
      "0001010" when "01011100101001001", -- t[47433] = 10
      "0001010" when "01011100101001010", -- t[47434] = 10
      "0001010" when "01011100101001011", -- t[47435] = 10
      "0001010" when "01011100101001100", -- t[47436] = 10
      "0001010" when "01011100101001101", -- t[47437] = 10
      "0001010" when "01011100101001110", -- t[47438] = 10
      "0001010" when "01011100101001111", -- t[47439] = 10
      "0001010" when "01011100101010000", -- t[47440] = 10
      "0001010" when "01011100101010001", -- t[47441] = 10
      "0001010" when "01011100101010010", -- t[47442] = 10
      "0001010" when "01011100101010011", -- t[47443] = 10
      "0001010" when "01011100101010100", -- t[47444] = 10
      "0001010" when "01011100101010101", -- t[47445] = 10
      "0001010" when "01011100101010110", -- t[47446] = 10
      "0001010" when "01011100101010111", -- t[47447] = 10
      "0001010" when "01011100101011000", -- t[47448] = 10
      "0001010" when "01011100101011001", -- t[47449] = 10
      "0001010" when "01011100101011010", -- t[47450] = 10
      "0001010" when "01011100101011011", -- t[47451] = 10
      "0001010" when "01011100101011100", -- t[47452] = 10
      "0001010" when "01011100101011101", -- t[47453] = 10
      "0001010" when "01011100101011110", -- t[47454] = 10
      "0001010" when "01011100101011111", -- t[47455] = 10
      "0001010" when "01011100101100000", -- t[47456] = 10
      "0001010" when "01011100101100001", -- t[47457] = 10
      "0001010" when "01011100101100010", -- t[47458] = 10
      "0001010" when "01011100101100011", -- t[47459] = 10
      "0001010" when "01011100101100100", -- t[47460] = 10
      "0001010" when "01011100101100101", -- t[47461] = 10
      "0001010" when "01011100101100110", -- t[47462] = 10
      "0001010" when "01011100101100111", -- t[47463] = 10
      "0001010" when "01011100101101000", -- t[47464] = 10
      "0001010" when "01011100101101001", -- t[47465] = 10
      "0001010" when "01011100101101010", -- t[47466] = 10
      "0001010" when "01011100101101011", -- t[47467] = 10
      "0001010" when "01011100101101100", -- t[47468] = 10
      "0001010" when "01011100101101101", -- t[47469] = 10
      "0001010" when "01011100101101110", -- t[47470] = 10
      "0001010" when "01011100101101111", -- t[47471] = 10
      "0001010" when "01011100101110000", -- t[47472] = 10
      "0001010" when "01011100101110001", -- t[47473] = 10
      "0001010" when "01011100101110010", -- t[47474] = 10
      "0001010" when "01011100101110011", -- t[47475] = 10
      "0001010" when "01011100101110100", -- t[47476] = 10
      "0001010" when "01011100101110101", -- t[47477] = 10
      "0001010" when "01011100101110110", -- t[47478] = 10
      "0001010" when "01011100101110111", -- t[47479] = 10
      "0001010" when "01011100101111000", -- t[47480] = 10
      "0001010" when "01011100101111001", -- t[47481] = 10
      "0001010" when "01011100101111010", -- t[47482] = 10
      "0001010" when "01011100101111011", -- t[47483] = 10
      "0001010" when "01011100101111100", -- t[47484] = 10
      "0001010" when "01011100101111101", -- t[47485] = 10
      "0001010" when "01011100101111110", -- t[47486] = 10
      "0001010" when "01011100101111111", -- t[47487] = 10
      "0001010" when "01011100110000000", -- t[47488] = 10
      "0001010" when "01011100110000001", -- t[47489] = 10
      "0001010" when "01011100110000010", -- t[47490] = 10
      "0001010" when "01011100110000011", -- t[47491] = 10
      "0001010" when "01011100110000100", -- t[47492] = 10
      "0001010" when "01011100110000101", -- t[47493] = 10
      "0001010" when "01011100110000110", -- t[47494] = 10
      "0001010" when "01011100110000111", -- t[47495] = 10
      "0001010" when "01011100110001000", -- t[47496] = 10
      "0001010" when "01011100110001001", -- t[47497] = 10
      "0001010" when "01011100110001010", -- t[47498] = 10
      "0001010" when "01011100110001011", -- t[47499] = 10
      "0001010" when "01011100110001100", -- t[47500] = 10
      "0001010" when "01011100110001101", -- t[47501] = 10
      "0001010" when "01011100110001110", -- t[47502] = 10
      "0001010" when "01011100110001111", -- t[47503] = 10
      "0001010" when "01011100110010000", -- t[47504] = 10
      "0001010" when "01011100110010001", -- t[47505] = 10
      "0001010" when "01011100110010010", -- t[47506] = 10
      "0001010" when "01011100110010011", -- t[47507] = 10
      "0001010" when "01011100110010100", -- t[47508] = 10
      "0001010" when "01011100110010101", -- t[47509] = 10
      "0001010" when "01011100110010110", -- t[47510] = 10
      "0001010" when "01011100110010111", -- t[47511] = 10
      "0001010" when "01011100110011000", -- t[47512] = 10
      "0001010" when "01011100110011001", -- t[47513] = 10
      "0001010" when "01011100110011010", -- t[47514] = 10
      "0001010" when "01011100110011011", -- t[47515] = 10
      "0001010" when "01011100110011100", -- t[47516] = 10
      "0001010" when "01011100110011101", -- t[47517] = 10
      "0001010" when "01011100110011110", -- t[47518] = 10
      "0001010" when "01011100110011111", -- t[47519] = 10
      "0001010" when "01011100110100000", -- t[47520] = 10
      "0001010" when "01011100110100001", -- t[47521] = 10
      "0001010" when "01011100110100010", -- t[47522] = 10
      "0001010" when "01011100110100011", -- t[47523] = 10
      "0001010" when "01011100110100100", -- t[47524] = 10
      "0001010" when "01011100110100101", -- t[47525] = 10
      "0001010" when "01011100110100110", -- t[47526] = 10
      "0001010" when "01011100110100111", -- t[47527] = 10
      "0001010" when "01011100110101000", -- t[47528] = 10
      "0001010" when "01011100110101001", -- t[47529] = 10
      "0001010" when "01011100110101010", -- t[47530] = 10
      "0001010" when "01011100110101011", -- t[47531] = 10
      "0001010" when "01011100110101100", -- t[47532] = 10
      "0001010" when "01011100110101101", -- t[47533] = 10
      "0001010" when "01011100110101110", -- t[47534] = 10
      "0001010" when "01011100110101111", -- t[47535] = 10
      "0001010" when "01011100110110000", -- t[47536] = 10
      "0001010" when "01011100110110001", -- t[47537] = 10
      "0001010" when "01011100110110010", -- t[47538] = 10
      "0001010" when "01011100110110011", -- t[47539] = 10
      "0001010" when "01011100110110100", -- t[47540] = 10
      "0001010" when "01011100110110101", -- t[47541] = 10
      "0001010" when "01011100110110110", -- t[47542] = 10
      "0001010" when "01011100110110111", -- t[47543] = 10
      "0001010" when "01011100110111000", -- t[47544] = 10
      "0001010" when "01011100110111001", -- t[47545] = 10
      "0001010" when "01011100110111010", -- t[47546] = 10
      "0001010" when "01011100110111011", -- t[47547] = 10
      "0001010" when "01011100110111100", -- t[47548] = 10
      "0001010" when "01011100110111101", -- t[47549] = 10
      "0001010" when "01011100110111110", -- t[47550] = 10
      "0001010" when "01011100110111111", -- t[47551] = 10
      "0001010" when "01011100111000000", -- t[47552] = 10
      "0001010" when "01011100111000001", -- t[47553] = 10
      "0001010" when "01011100111000010", -- t[47554] = 10
      "0001010" when "01011100111000011", -- t[47555] = 10
      "0001010" when "01011100111000100", -- t[47556] = 10
      "0001010" when "01011100111000101", -- t[47557] = 10
      "0001010" when "01011100111000110", -- t[47558] = 10
      "0001010" when "01011100111000111", -- t[47559] = 10
      "0001010" when "01011100111001000", -- t[47560] = 10
      "0001010" when "01011100111001001", -- t[47561] = 10
      "0001010" when "01011100111001010", -- t[47562] = 10
      "0001010" when "01011100111001011", -- t[47563] = 10
      "0001010" when "01011100111001100", -- t[47564] = 10
      "0001010" when "01011100111001101", -- t[47565] = 10
      "0001010" when "01011100111001110", -- t[47566] = 10
      "0001010" when "01011100111001111", -- t[47567] = 10
      "0001010" when "01011100111010000", -- t[47568] = 10
      "0001010" when "01011100111010001", -- t[47569] = 10
      "0001010" when "01011100111010010", -- t[47570] = 10
      "0001010" when "01011100111010011", -- t[47571] = 10
      "0001010" when "01011100111010100", -- t[47572] = 10
      "0001010" when "01011100111010101", -- t[47573] = 10
      "0001010" when "01011100111010110", -- t[47574] = 10
      "0001010" when "01011100111010111", -- t[47575] = 10
      "0001010" when "01011100111011000", -- t[47576] = 10
      "0001010" when "01011100111011001", -- t[47577] = 10
      "0001010" when "01011100111011010", -- t[47578] = 10
      "0001010" when "01011100111011011", -- t[47579] = 10
      "0001010" when "01011100111011100", -- t[47580] = 10
      "0001010" when "01011100111011101", -- t[47581] = 10
      "0001010" when "01011100111011110", -- t[47582] = 10
      "0001010" when "01011100111011111", -- t[47583] = 10
      "0001010" when "01011100111100000", -- t[47584] = 10
      "0001010" when "01011100111100001", -- t[47585] = 10
      "0001010" when "01011100111100010", -- t[47586] = 10
      "0001010" when "01011100111100011", -- t[47587] = 10
      "0001010" when "01011100111100100", -- t[47588] = 10
      "0001010" when "01011100111100101", -- t[47589] = 10
      "0001010" when "01011100111100110", -- t[47590] = 10
      "0001010" when "01011100111100111", -- t[47591] = 10
      "0001010" when "01011100111101000", -- t[47592] = 10
      "0001010" when "01011100111101001", -- t[47593] = 10
      "0001010" when "01011100111101010", -- t[47594] = 10
      "0001010" when "01011100111101011", -- t[47595] = 10
      "0001010" when "01011100111101100", -- t[47596] = 10
      "0001010" when "01011100111101101", -- t[47597] = 10
      "0001010" when "01011100111101110", -- t[47598] = 10
      "0001010" when "01011100111101111", -- t[47599] = 10
      "0001010" when "01011100111110000", -- t[47600] = 10
      "0001010" when "01011100111110001", -- t[47601] = 10
      "0001010" when "01011100111110010", -- t[47602] = 10
      "0001010" when "01011100111110011", -- t[47603] = 10
      "0001010" when "01011100111110100", -- t[47604] = 10
      "0001010" when "01011100111110101", -- t[47605] = 10
      "0001010" when "01011100111110110", -- t[47606] = 10
      "0001010" when "01011100111110111", -- t[47607] = 10
      "0001010" when "01011100111111000", -- t[47608] = 10
      "0001010" when "01011100111111001", -- t[47609] = 10
      "0001010" when "01011100111111010", -- t[47610] = 10
      "0001010" when "01011100111111011", -- t[47611] = 10
      "0001010" when "01011100111111100", -- t[47612] = 10
      "0001010" when "01011100111111101", -- t[47613] = 10
      "0001010" when "01011100111111110", -- t[47614] = 10
      "0001010" when "01011100111111111", -- t[47615] = 10
      "0001010" when "01011101000000000", -- t[47616] = 10
      "0001010" when "01011101000000001", -- t[47617] = 10
      "0001010" when "01011101000000010", -- t[47618] = 10
      "0001010" when "01011101000000011", -- t[47619] = 10
      "0001010" when "01011101000000100", -- t[47620] = 10
      "0001010" when "01011101000000101", -- t[47621] = 10
      "0001010" when "01011101000000110", -- t[47622] = 10
      "0001010" when "01011101000000111", -- t[47623] = 10
      "0001010" when "01011101000001000", -- t[47624] = 10
      "0001010" when "01011101000001001", -- t[47625] = 10
      "0001010" when "01011101000001010", -- t[47626] = 10
      "0001010" when "01011101000001011", -- t[47627] = 10
      "0001010" when "01011101000001100", -- t[47628] = 10
      "0001010" when "01011101000001101", -- t[47629] = 10
      "0001010" when "01011101000001110", -- t[47630] = 10
      "0001010" when "01011101000001111", -- t[47631] = 10
      "0001010" when "01011101000010000", -- t[47632] = 10
      "0001010" when "01011101000010001", -- t[47633] = 10
      "0001010" when "01011101000010010", -- t[47634] = 10
      "0001010" when "01011101000010011", -- t[47635] = 10
      "0001010" when "01011101000010100", -- t[47636] = 10
      "0001010" when "01011101000010101", -- t[47637] = 10
      "0001010" when "01011101000010110", -- t[47638] = 10
      "0001010" when "01011101000010111", -- t[47639] = 10
      "0001010" when "01011101000011000", -- t[47640] = 10
      "0001010" when "01011101000011001", -- t[47641] = 10
      "0001010" when "01011101000011010", -- t[47642] = 10
      "0001010" when "01011101000011011", -- t[47643] = 10
      "0001010" when "01011101000011100", -- t[47644] = 10
      "0001010" when "01011101000011101", -- t[47645] = 10
      "0001010" when "01011101000011110", -- t[47646] = 10
      "0001010" when "01011101000011111", -- t[47647] = 10
      "0001010" when "01011101000100000", -- t[47648] = 10
      "0001010" when "01011101000100001", -- t[47649] = 10
      "0001010" when "01011101000100010", -- t[47650] = 10
      "0001010" when "01011101000100011", -- t[47651] = 10
      "0001010" when "01011101000100100", -- t[47652] = 10
      "0001010" when "01011101000100101", -- t[47653] = 10
      "0001010" when "01011101000100110", -- t[47654] = 10
      "0001010" when "01011101000100111", -- t[47655] = 10
      "0001010" when "01011101000101000", -- t[47656] = 10
      "0001010" when "01011101000101001", -- t[47657] = 10
      "0001010" when "01011101000101010", -- t[47658] = 10
      "0001010" when "01011101000101011", -- t[47659] = 10
      "0001010" when "01011101000101100", -- t[47660] = 10
      "0001010" when "01011101000101101", -- t[47661] = 10
      "0001010" when "01011101000101110", -- t[47662] = 10
      "0001010" when "01011101000101111", -- t[47663] = 10
      "0001010" when "01011101000110000", -- t[47664] = 10
      "0001010" when "01011101000110001", -- t[47665] = 10
      "0001010" when "01011101000110010", -- t[47666] = 10
      "0001010" when "01011101000110011", -- t[47667] = 10
      "0001010" when "01011101000110100", -- t[47668] = 10
      "0001010" when "01011101000110101", -- t[47669] = 10
      "0001010" when "01011101000110110", -- t[47670] = 10
      "0001010" when "01011101000110111", -- t[47671] = 10
      "0001010" when "01011101000111000", -- t[47672] = 10
      "0001010" when "01011101000111001", -- t[47673] = 10
      "0001010" when "01011101000111010", -- t[47674] = 10
      "0001010" when "01011101000111011", -- t[47675] = 10
      "0001010" when "01011101000111100", -- t[47676] = 10
      "0001010" when "01011101000111101", -- t[47677] = 10
      "0001010" when "01011101000111110", -- t[47678] = 10
      "0001010" when "01011101000111111", -- t[47679] = 10
      "0001010" when "01011101001000000", -- t[47680] = 10
      "0001010" when "01011101001000001", -- t[47681] = 10
      "0001010" when "01011101001000010", -- t[47682] = 10
      "0001010" when "01011101001000011", -- t[47683] = 10
      "0001010" when "01011101001000100", -- t[47684] = 10
      "0001010" when "01011101001000101", -- t[47685] = 10
      "0001010" when "01011101001000110", -- t[47686] = 10
      "0001010" when "01011101001000111", -- t[47687] = 10
      "0001010" when "01011101001001000", -- t[47688] = 10
      "0001010" when "01011101001001001", -- t[47689] = 10
      "0001010" when "01011101001001010", -- t[47690] = 10
      "0001010" when "01011101001001011", -- t[47691] = 10
      "0001010" when "01011101001001100", -- t[47692] = 10
      "0001010" when "01011101001001101", -- t[47693] = 10
      "0001010" when "01011101001001110", -- t[47694] = 10
      "0001010" when "01011101001001111", -- t[47695] = 10
      "0001010" when "01011101001010000", -- t[47696] = 10
      "0001010" when "01011101001010001", -- t[47697] = 10
      "0001010" when "01011101001010010", -- t[47698] = 10
      "0001010" when "01011101001010011", -- t[47699] = 10
      "0001010" when "01011101001010100", -- t[47700] = 10
      "0001010" when "01011101001010101", -- t[47701] = 10
      "0001010" when "01011101001010110", -- t[47702] = 10
      "0001010" when "01011101001010111", -- t[47703] = 10
      "0001010" when "01011101001011000", -- t[47704] = 10
      "0001010" when "01011101001011001", -- t[47705] = 10
      "0001010" when "01011101001011010", -- t[47706] = 10
      "0001010" when "01011101001011011", -- t[47707] = 10
      "0001010" when "01011101001011100", -- t[47708] = 10
      "0001010" when "01011101001011101", -- t[47709] = 10
      "0001010" when "01011101001011110", -- t[47710] = 10
      "0001010" when "01011101001011111", -- t[47711] = 10
      "0001010" when "01011101001100000", -- t[47712] = 10
      "0001010" when "01011101001100001", -- t[47713] = 10
      "0001010" when "01011101001100010", -- t[47714] = 10
      "0001010" when "01011101001100011", -- t[47715] = 10
      "0001010" when "01011101001100100", -- t[47716] = 10
      "0001010" when "01011101001100101", -- t[47717] = 10
      "0001010" when "01011101001100110", -- t[47718] = 10
      "0001010" when "01011101001100111", -- t[47719] = 10
      "0001010" when "01011101001101000", -- t[47720] = 10
      "0001010" when "01011101001101001", -- t[47721] = 10
      "0001010" when "01011101001101010", -- t[47722] = 10
      "0001010" when "01011101001101011", -- t[47723] = 10
      "0001010" when "01011101001101100", -- t[47724] = 10
      "0001010" when "01011101001101101", -- t[47725] = 10
      "0001010" when "01011101001101110", -- t[47726] = 10
      "0001010" when "01011101001101111", -- t[47727] = 10
      "0001010" when "01011101001110000", -- t[47728] = 10
      "0001010" when "01011101001110001", -- t[47729] = 10
      "0001010" when "01011101001110010", -- t[47730] = 10
      "0001010" when "01011101001110011", -- t[47731] = 10
      "0001010" when "01011101001110100", -- t[47732] = 10
      "0001010" when "01011101001110101", -- t[47733] = 10
      "0001010" when "01011101001110110", -- t[47734] = 10
      "0001010" when "01011101001110111", -- t[47735] = 10
      "0001010" when "01011101001111000", -- t[47736] = 10
      "0001010" when "01011101001111001", -- t[47737] = 10
      "0001010" when "01011101001111010", -- t[47738] = 10
      "0001010" when "01011101001111011", -- t[47739] = 10
      "0001010" when "01011101001111100", -- t[47740] = 10
      "0001010" when "01011101001111101", -- t[47741] = 10
      "0001010" when "01011101001111110", -- t[47742] = 10
      "0001010" when "01011101001111111", -- t[47743] = 10
      "0001010" when "01011101010000000", -- t[47744] = 10
      "0001010" when "01011101010000001", -- t[47745] = 10
      "0001010" when "01011101010000010", -- t[47746] = 10
      "0001010" when "01011101010000011", -- t[47747] = 10
      "0001010" when "01011101010000100", -- t[47748] = 10
      "0001010" when "01011101010000101", -- t[47749] = 10
      "0001010" when "01011101010000110", -- t[47750] = 10
      "0001010" when "01011101010000111", -- t[47751] = 10
      "0001010" when "01011101010001000", -- t[47752] = 10
      "0001010" when "01011101010001001", -- t[47753] = 10
      "0001010" when "01011101010001010", -- t[47754] = 10
      "0001010" when "01011101010001011", -- t[47755] = 10
      "0001010" when "01011101010001100", -- t[47756] = 10
      "0001010" when "01011101010001101", -- t[47757] = 10
      "0001010" when "01011101010001110", -- t[47758] = 10
      "0001010" when "01011101010001111", -- t[47759] = 10
      "0001010" when "01011101010010000", -- t[47760] = 10
      "0001010" when "01011101010010001", -- t[47761] = 10
      "0001010" when "01011101010010010", -- t[47762] = 10
      "0001010" when "01011101010010011", -- t[47763] = 10
      "0001010" when "01011101010010100", -- t[47764] = 10
      "0001010" when "01011101010010101", -- t[47765] = 10
      "0001010" when "01011101010010110", -- t[47766] = 10
      "0001010" when "01011101010010111", -- t[47767] = 10
      "0001010" when "01011101010011000", -- t[47768] = 10
      "0001010" when "01011101010011001", -- t[47769] = 10
      "0001010" when "01011101010011010", -- t[47770] = 10
      "0001010" when "01011101010011011", -- t[47771] = 10
      "0001010" when "01011101010011100", -- t[47772] = 10
      "0001010" when "01011101010011101", -- t[47773] = 10
      "0001010" when "01011101010011110", -- t[47774] = 10
      "0001010" when "01011101010011111", -- t[47775] = 10
      "0001010" when "01011101010100000", -- t[47776] = 10
      "0001010" when "01011101010100001", -- t[47777] = 10
      "0001010" when "01011101010100010", -- t[47778] = 10
      "0001010" when "01011101010100011", -- t[47779] = 10
      "0001010" when "01011101010100100", -- t[47780] = 10
      "0001010" when "01011101010100101", -- t[47781] = 10
      "0001010" when "01011101010100110", -- t[47782] = 10
      "0001010" when "01011101010100111", -- t[47783] = 10
      "0001010" when "01011101010101000", -- t[47784] = 10
      "0001010" when "01011101010101001", -- t[47785] = 10
      "0001010" when "01011101010101010", -- t[47786] = 10
      "0001010" when "01011101010101011", -- t[47787] = 10
      "0001010" when "01011101010101100", -- t[47788] = 10
      "0001010" when "01011101010101101", -- t[47789] = 10
      "0001010" when "01011101010101110", -- t[47790] = 10
      "0001010" when "01011101010101111", -- t[47791] = 10
      "0001010" when "01011101010110000", -- t[47792] = 10
      "0001010" when "01011101010110001", -- t[47793] = 10
      "0001010" when "01011101010110010", -- t[47794] = 10
      "0001010" when "01011101010110011", -- t[47795] = 10
      "0001010" when "01011101010110100", -- t[47796] = 10
      "0001010" when "01011101010110101", -- t[47797] = 10
      "0001010" when "01011101010110110", -- t[47798] = 10
      "0001010" when "01011101010110111", -- t[47799] = 10
      "0001010" when "01011101010111000", -- t[47800] = 10
      "0001010" when "01011101010111001", -- t[47801] = 10
      "0001010" when "01011101010111010", -- t[47802] = 10
      "0001010" when "01011101010111011", -- t[47803] = 10
      "0001010" when "01011101010111100", -- t[47804] = 10
      "0001010" when "01011101010111101", -- t[47805] = 10
      "0001010" when "01011101010111110", -- t[47806] = 10
      "0001010" when "01011101010111111", -- t[47807] = 10
      "0001010" when "01011101011000000", -- t[47808] = 10
      "0001010" when "01011101011000001", -- t[47809] = 10
      "0001010" when "01011101011000010", -- t[47810] = 10
      "0001010" when "01011101011000011", -- t[47811] = 10
      "0001010" when "01011101011000100", -- t[47812] = 10
      "0001010" when "01011101011000101", -- t[47813] = 10
      "0001010" when "01011101011000110", -- t[47814] = 10
      "0001010" when "01011101011000111", -- t[47815] = 10
      "0001010" when "01011101011001000", -- t[47816] = 10
      "0001010" when "01011101011001001", -- t[47817] = 10
      "0001010" when "01011101011001010", -- t[47818] = 10
      "0001010" when "01011101011001011", -- t[47819] = 10
      "0001010" when "01011101011001100", -- t[47820] = 10
      "0001010" when "01011101011001101", -- t[47821] = 10
      "0001010" when "01011101011001110", -- t[47822] = 10
      "0001010" when "01011101011001111", -- t[47823] = 10
      "0001010" when "01011101011010000", -- t[47824] = 10
      "0001010" when "01011101011010001", -- t[47825] = 10
      "0001010" when "01011101011010010", -- t[47826] = 10
      "0001010" when "01011101011010011", -- t[47827] = 10
      "0001010" when "01011101011010100", -- t[47828] = 10
      "0001010" when "01011101011010101", -- t[47829] = 10
      "0001010" when "01011101011010110", -- t[47830] = 10
      "0001010" when "01011101011010111", -- t[47831] = 10
      "0001010" when "01011101011011000", -- t[47832] = 10
      "0001010" when "01011101011011001", -- t[47833] = 10
      "0001010" when "01011101011011010", -- t[47834] = 10
      "0001010" when "01011101011011011", -- t[47835] = 10
      "0001010" when "01011101011011100", -- t[47836] = 10
      "0001010" when "01011101011011101", -- t[47837] = 10
      "0001010" when "01011101011011110", -- t[47838] = 10
      "0001010" when "01011101011011111", -- t[47839] = 10
      "0001010" when "01011101011100000", -- t[47840] = 10
      "0001010" when "01011101011100001", -- t[47841] = 10
      "0001010" when "01011101011100010", -- t[47842] = 10
      "0001010" when "01011101011100011", -- t[47843] = 10
      "0001010" when "01011101011100100", -- t[47844] = 10
      "0001010" when "01011101011100101", -- t[47845] = 10
      "0001010" when "01011101011100110", -- t[47846] = 10
      "0001010" when "01011101011100111", -- t[47847] = 10
      "0001010" when "01011101011101000", -- t[47848] = 10
      "0001010" when "01011101011101001", -- t[47849] = 10
      "0001010" when "01011101011101010", -- t[47850] = 10
      "0001010" when "01011101011101011", -- t[47851] = 10
      "0001010" when "01011101011101100", -- t[47852] = 10
      "0001010" when "01011101011101101", -- t[47853] = 10
      "0001010" when "01011101011101110", -- t[47854] = 10
      "0001010" when "01011101011101111", -- t[47855] = 10
      "0001010" when "01011101011110000", -- t[47856] = 10
      "0001010" when "01011101011110001", -- t[47857] = 10
      "0001010" when "01011101011110010", -- t[47858] = 10
      "0001010" when "01011101011110011", -- t[47859] = 10
      "0001010" when "01011101011110100", -- t[47860] = 10
      "0001010" when "01011101011110101", -- t[47861] = 10
      "0001010" when "01011101011110110", -- t[47862] = 10
      "0001010" when "01011101011110111", -- t[47863] = 10
      "0001010" when "01011101011111000", -- t[47864] = 10
      "0001010" when "01011101011111001", -- t[47865] = 10
      "0001010" when "01011101011111010", -- t[47866] = 10
      "0001010" when "01011101011111011", -- t[47867] = 10
      "0001010" when "01011101011111100", -- t[47868] = 10
      "0001010" when "01011101011111101", -- t[47869] = 10
      "0001010" when "01011101011111110", -- t[47870] = 10
      "0001010" when "01011101011111111", -- t[47871] = 10
      "0001010" when "01011101100000000", -- t[47872] = 10
      "0001010" when "01011101100000001", -- t[47873] = 10
      "0001010" when "01011101100000010", -- t[47874] = 10
      "0001010" when "01011101100000011", -- t[47875] = 10
      "0001010" when "01011101100000100", -- t[47876] = 10
      "0001010" when "01011101100000101", -- t[47877] = 10
      "0001010" when "01011101100000110", -- t[47878] = 10
      "0001010" when "01011101100000111", -- t[47879] = 10
      "0001010" when "01011101100001000", -- t[47880] = 10
      "0001010" when "01011101100001001", -- t[47881] = 10
      "0001010" when "01011101100001010", -- t[47882] = 10
      "0001010" when "01011101100001011", -- t[47883] = 10
      "0001010" when "01011101100001100", -- t[47884] = 10
      "0001010" when "01011101100001101", -- t[47885] = 10
      "0001010" when "01011101100001110", -- t[47886] = 10
      "0001010" when "01011101100001111", -- t[47887] = 10
      "0001010" when "01011101100010000", -- t[47888] = 10
      "0001010" when "01011101100010001", -- t[47889] = 10
      "0001010" when "01011101100010010", -- t[47890] = 10
      "0001010" when "01011101100010011", -- t[47891] = 10
      "0001010" when "01011101100010100", -- t[47892] = 10
      "0001010" when "01011101100010101", -- t[47893] = 10
      "0001010" when "01011101100010110", -- t[47894] = 10
      "0001010" when "01011101100010111", -- t[47895] = 10
      "0001010" when "01011101100011000", -- t[47896] = 10
      "0001010" when "01011101100011001", -- t[47897] = 10
      "0001010" when "01011101100011010", -- t[47898] = 10
      "0001010" when "01011101100011011", -- t[47899] = 10
      "0001010" when "01011101100011100", -- t[47900] = 10
      "0001010" when "01011101100011101", -- t[47901] = 10
      "0001010" when "01011101100011110", -- t[47902] = 10
      "0001010" when "01011101100011111", -- t[47903] = 10
      "0001010" when "01011101100100000", -- t[47904] = 10
      "0001010" when "01011101100100001", -- t[47905] = 10
      "0001010" when "01011101100100010", -- t[47906] = 10
      "0001010" when "01011101100100011", -- t[47907] = 10
      "0001010" when "01011101100100100", -- t[47908] = 10
      "0001010" when "01011101100100101", -- t[47909] = 10
      "0001010" when "01011101100100110", -- t[47910] = 10
      "0001010" when "01011101100100111", -- t[47911] = 10
      "0001010" when "01011101100101000", -- t[47912] = 10
      "0001010" when "01011101100101001", -- t[47913] = 10
      "0001010" when "01011101100101010", -- t[47914] = 10
      "0001010" when "01011101100101011", -- t[47915] = 10
      "0001010" when "01011101100101100", -- t[47916] = 10
      "0001010" when "01011101100101101", -- t[47917] = 10
      "0001010" when "01011101100101110", -- t[47918] = 10
      "0001010" when "01011101100101111", -- t[47919] = 10
      "0001010" when "01011101100110000", -- t[47920] = 10
      "0001010" when "01011101100110001", -- t[47921] = 10
      "0001010" when "01011101100110010", -- t[47922] = 10
      "0001010" when "01011101100110011", -- t[47923] = 10
      "0001010" when "01011101100110100", -- t[47924] = 10
      "0001010" when "01011101100110101", -- t[47925] = 10
      "0001010" when "01011101100110110", -- t[47926] = 10
      "0001010" when "01011101100110111", -- t[47927] = 10
      "0001010" when "01011101100111000", -- t[47928] = 10
      "0001010" when "01011101100111001", -- t[47929] = 10
      "0001010" when "01011101100111010", -- t[47930] = 10
      "0001010" when "01011101100111011", -- t[47931] = 10
      "0001010" when "01011101100111100", -- t[47932] = 10
      "0001010" when "01011101100111101", -- t[47933] = 10
      "0001010" when "01011101100111110", -- t[47934] = 10
      "0001010" when "01011101100111111", -- t[47935] = 10
      "0001010" when "01011101101000000", -- t[47936] = 10
      "0001010" when "01011101101000001", -- t[47937] = 10
      "0001010" when "01011101101000010", -- t[47938] = 10
      "0001010" when "01011101101000011", -- t[47939] = 10
      "0001010" when "01011101101000100", -- t[47940] = 10
      "0001010" when "01011101101000101", -- t[47941] = 10
      "0001010" when "01011101101000110", -- t[47942] = 10
      "0001010" when "01011101101000111", -- t[47943] = 10
      "0001010" when "01011101101001000", -- t[47944] = 10
      "0001010" when "01011101101001001", -- t[47945] = 10
      "0001010" when "01011101101001010", -- t[47946] = 10
      "0001010" when "01011101101001011", -- t[47947] = 10
      "0001010" when "01011101101001100", -- t[47948] = 10
      "0001010" when "01011101101001101", -- t[47949] = 10
      "0001010" when "01011101101001110", -- t[47950] = 10
      "0001010" when "01011101101001111", -- t[47951] = 10
      "0001010" when "01011101101010000", -- t[47952] = 10
      "0001010" when "01011101101010001", -- t[47953] = 10
      "0001010" when "01011101101010010", -- t[47954] = 10
      "0001010" when "01011101101010011", -- t[47955] = 10
      "0001010" when "01011101101010100", -- t[47956] = 10
      "0001010" when "01011101101010101", -- t[47957] = 10
      "0001010" when "01011101101010110", -- t[47958] = 10
      "0001010" when "01011101101010111", -- t[47959] = 10
      "0001010" when "01011101101011000", -- t[47960] = 10
      "0001010" when "01011101101011001", -- t[47961] = 10
      "0001010" when "01011101101011010", -- t[47962] = 10
      "0001010" when "01011101101011011", -- t[47963] = 10
      "0001010" when "01011101101011100", -- t[47964] = 10
      "0001010" when "01011101101011101", -- t[47965] = 10
      "0001010" when "01011101101011110", -- t[47966] = 10
      "0001010" when "01011101101011111", -- t[47967] = 10
      "0001010" when "01011101101100000", -- t[47968] = 10
      "0001010" when "01011101101100001", -- t[47969] = 10
      "0001010" when "01011101101100010", -- t[47970] = 10
      "0001010" when "01011101101100011", -- t[47971] = 10
      "0001010" when "01011101101100100", -- t[47972] = 10
      "0001010" when "01011101101100101", -- t[47973] = 10
      "0001010" when "01011101101100110", -- t[47974] = 10
      "0001010" when "01011101101100111", -- t[47975] = 10
      "0001010" when "01011101101101000", -- t[47976] = 10
      "0001010" when "01011101101101001", -- t[47977] = 10
      "0001010" when "01011101101101010", -- t[47978] = 10
      "0001010" when "01011101101101011", -- t[47979] = 10
      "0001010" when "01011101101101100", -- t[47980] = 10
      "0001010" when "01011101101101101", -- t[47981] = 10
      "0001010" when "01011101101101110", -- t[47982] = 10
      "0001010" when "01011101101101111", -- t[47983] = 10
      "0001010" when "01011101101110000", -- t[47984] = 10
      "0001010" when "01011101101110001", -- t[47985] = 10
      "0001010" when "01011101101110010", -- t[47986] = 10
      "0001010" when "01011101101110011", -- t[47987] = 10
      "0001010" when "01011101101110100", -- t[47988] = 10
      "0001010" when "01011101101110101", -- t[47989] = 10
      "0001010" when "01011101101110110", -- t[47990] = 10
      "0001010" when "01011101101110111", -- t[47991] = 10
      "0001010" when "01011101101111000", -- t[47992] = 10
      "0001010" when "01011101101111001", -- t[47993] = 10
      "0001010" when "01011101101111010", -- t[47994] = 10
      "0001010" when "01011101101111011", -- t[47995] = 10
      "0001010" when "01011101101111100", -- t[47996] = 10
      "0001010" when "01011101101111101", -- t[47997] = 10
      "0001010" when "01011101101111110", -- t[47998] = 10
      "0001010" when "01011101101111111", -- t[47999] = 10
      "0001010" when "01011101110000000", -- t[48000] = 10
      "0001010" when "01011101110000001", -- t[48001] = 10
      "0001010" when "01011101110000010", -- t[48002] = 10
      "0001010" when "01011101110000011", -- t[48003] = 10
      "0001010" when "01011101110000100", -- t[48004] = 10
      "0001010" when "01011101110000101", -- t[48005] = 10
      "0001010" when "01011101110000110", -- t[48006] = 10
      "0001010" when "01011101110000111", -- t[48007] = 10
      "0001010" when "01011101110001000", -- t[48008] = 10
      "0001010" when "01011101110001001", -- t[48009] = 10
      "0001010" when "01011101110001010", -- t[48010] = 10
      "0001010" when "01011101110001011", -- t[48011] = 10
      "0001010" when "01011101110001100", -- t[48012] = 10
      "0001010" when "01011101110001101", -- t[48013] = 10
      "0001010" when "01011101110001110", -- t[48014] = 10
      "0001010" when "01011101110001111", -- t[48015] = 10
      "0001010" when "01011101110010000", -- t[48016] = 10
      "0001010" when "01011101110010001", -- t[48017] = 10
      "0001010" when "01011101110010010", -- t[48018] = 10
      "0001010" when "01011101110010011", -- t[48019] = 10
      "0001010" when "01011101110010100", -- t[48020] = 10
      "0001010" when "01011101110010101", -- t[48021] = 10
      "0001010" when "01011101110010110", -- t[48022] = 10
      "0001010" when "01011101110010111", -- t[48023] = 10
      "0001010" when "01011101110011000", -- t[48024] = 10
      "0001010" when "01011101110011001", -- t[48025] = 10
      "0001010" when "01011101110011010", -- t[48026] = 10
      "0001010" when "01011101110011011", -- t[48027] = 10
      "0001010" when "01011101110011100", -- t[48028] = 10
      "0001011" when "01011101110011101", -- t[48029] = 11
      "0001011" when "01011101110011110", -- t[48030] = 11
      "0001011" when "01011101110011111", -- t[48031] = 11
      "0001011" when "01011101110100000", -- t[48032] = 11
      "0001011" when "01011101110100001", -- t[48033] = 11
      "0001011" when "01011101110100010", -- t[48034] = 11
      "0001011" when "01011101110100011", -- t[48035] = 11
      "0001011" when "01011101110100100", -- t[48036] = 11
      "0001011" when "01011101110100101", -- t[48037] = 11
      "0001011" when "01011101110100110", -- t[48038] = 11
      "0001011" when "01011101110100111", -- t[48039] = 11
      "0001011" when "01011101110101000", -- t[48040] = 11
      "0001011" when "01011101110101001", -- t[48041] = 11
      "0001011" when "01011101110101010", -- t[48042] = 11
      "0001011" when "01011101110101011", -- t[48043] = 11
      "0001011" when "01011101110101100", -- t[48044] = 11
      "0001011" when "01011101110101101", -- t[48045] = 11
      "0001011" when "01011101110101110", -- t[48046] = 11
      "0001011" when "01011101110101111", -- t[48047] = 11
      "0001011" when "01011101110110000", -- t[48048] = 11
      "0001011" when "01011101110110001", -- t[48049] = 11
      "0001011" when "01011101110110010", -- t[48050] = 11
      "0001011" when "01011101110110011", -- t[48051] = 11
      "0001011" when "01011101110110100", -- t[48052] = 11
      "0001011" when "01011101110110101", -- t[48053] = 11
      "0001011" when "01011101110110110", -- t[48054] = 11
      "0001011" when "01011101110110111", -- t[48055] = 11
      "0001011" when "01011101110111000", -- t[48056] = 11
      "0001011" when "01011101110111001", -- t[48057] = 11
      "0001011" when "01011101110111010", -- t[48058] = 11
      "0001011" when "01011101110111011", -- t[48059] = 11
      "0001011" when "01011101110111100", -- t[48060] = 11
      "0001011" when "01011101110111101", -- t[48061] = 11
      "0001011" when "01011101110111110", -- t[48062] = 11
      "0001011" when "01011101110111111", -- t[48063] = 11
      "0001011" when "01011101111000000", -- t[48064] = 11
      "0001011" when "01011101111000001", -- t[48065] = 11
      "0001011" when "01011101111000010", -- t[48066] = 11
      "0001011" when "01011101111000011", -- t[48067] = 11
      "0001011" when "01011101111000100", -- t[48068] = 11
      "0001011" when "01011101111000101", -- t[48069] = 11
      "0001011" when "01011101111000110", -- t[48070] = 11
      "0001011" when "01011101111000111", -- t[48071] = 11
      "0001011" when "01011101111001000", -- t[48072] = 11
      "0001011" when "01011101111001001", -- t[48073] = 11
      "0001011" when "01011101111001010", -- t[48074] = 11
      "0001011" when "01011101111001011", -- t[48075] = 11
      "0001011" when "01011101111001100", -- t[48076] = 11
      "0001011" when "01011101111001101", -- t[48077] = 11
      "0001011" when "01011101111001110", -- t[48078] = 11
      "0001011" when "01011101111001111", -- t[48079] = 11
      "0001011" when "01011101111010000", -- t[48080] = 11
      "0001011" when "01011101111010001", -- t[48081] = 11
      "0001011" when "01011101111010010", -- t[48082] = 11
      "0001011" when "01011101111010011", -- t[48083] = 11
      "0001011" when "01011101111010100", -- t[48084] = 11
      "0001011" when "01011101111010101", -- t[48085] = 11
      "0001011" when "01011101111010110", -- t[48086] = 11
      "0001011" when "01011101111010111", -- t[48087] = 11
      "0001011" when "01011101111011000", -- t[48088] = 11
      "0001011" when "01011101111011001", -- t[48089] = 11
      "0001011" when "01011101111011010", -- t[48090] = 11
      "0001011" when "01011101111011011", -- t[48091] = 11
      "0001011" when "01011101111011100", -- t[48092] = 11
      "0001011" when "01011101111011101", -- t[48093] = 11
      "0001011" when "01011101111011110", -- t[48094] = 11
      "0001011" when "01011101111011111", -- t[48095] = 11
      "0001011" when "01011101111100000", -- t[48096] = 11
      "0001011" when "01011101111100001", -- t[48097] = 11
      "0001011" when "01011101111100010", -- t[48098] = 11
      "0001011" when "01011101111100011", -- t[48099] = 11
      "0001011" when "01011101111100100", -- t[48100] = 11
      "0001011" when "01011101111100101", -- t[48101] = 11
      "0001011" when "01011101111100110", -- t[48102] = 11
      "0001011" when "01011101111100111", -- t[48103] = 11
      "0001011" when "01011101111101000", -- t[48104] = 11
      "0001011" when "01011101111101001", -- t[48105] = 11
      "0001011" when "01011101111101010", -- t[48106] = 11
      "0001011" when "01011101111101011", -- t[48107] = 11
      "0001011" when "01011101111101100", -- t[48108] = 11
      "0001011" when "01011101111101101", -- t[48109] = 11
      "0001011" when "01011101111101110", -- t[48110] = 11
      "0001011" when "01011101111101111", -- t[48111] = 11
      "0001011" when "01011101111110000", -- t[48112] = 11
      "0001011" when "01011101111110001", -- t[48113] = 11
      "0001011" when "01011101111110010", -- t[48114] = 11
      "0001011" when "01011101111110011", -- t[48115] = 11
      "0001011" when "01011101111110100", -- t[48116] = 11
      "0001011" when "01011101111110101", -- t[48117] = 11
      "0001011" when "01011101111110110", -- t[48118] = 11
      "0001011" when "01011101111110111", -- t[48119] = 11
      "0001011" when "01011101111111000", -- t[48120] = 11
      "0001011" when "01011101111111001", -- t[48121] = 11
      "0001011" when "01011101111111010", -- t[48122] = 11
      "0001011" when "01011101111111011", -- t[48123] = 11
      "0001011" when "01011101111111100", -- t[48124] = 11
      "0001011" when "01011101111111101", -- t[48125] = 11
      "0001011" when "01011101111111110", -- t[48126] = 11
      "0001011" when "01011101111111111", -- t[48127] = 11
      "0001011" when "01011110000000000", -- t[48128] = 11
      "0001011" when "01011110000000001", -- t[48129] = 11
      "0001011" when "01011110000000010", -- t[48130] = 11
      "0001011" when "01011110000000011", -- t[48131] = 11
      "0001011" when "01011110000000100", -- t[48132] = 11
      "0001011" when "01011110000000101", -- t[48133] = 11
      "0001011" when "01011110000000110", -- t[48134] = 11
      "0001011" when "01011110000000111", -- t[48135] = 11
      "0001011" when "01011110000001000", -- t[48136] = 11
      "0001011" when "01011110000001001", -- t[48137] = 11
      "0001011" when "01011110000001010", -- t[48138] = 11
      "0001011" when "01011110000001011", -- t[48139] = 11
      "0001011" when "01011110000001100", -- t[48140] = 11
      "0001011" when "01011110000001101", -- t[48141] = 11
      "0001011" when "01011110000001110", -- t[48142] = 11
      "0001011" when "01011110000001111", -- t[48143] = 11
      "0001011" when "01011110000010000", -- t[48144] = 11
      "0001011" when "01011110000010001", -- t[48145] = 11
      "0001011" when "01011110000010010", -- t[48146] = 11
      "0001011" when "01011110000010011", -- t[48147] = 11
      "0001011" when "01011110000010100", -- t[48148] = 11
      "0001011" when "01011110000010101", -- t[48149] = 11
      "0001011" when "01011110000010110", -- t[48150] = 11
      "0001011" when "01011110000010111", -- t[48151] = 11
      "0001011" when "01011110000011000", -- t[48152] = 11
      "0001011" when "01011110000011001", -- t[48153] = 11
      "0001011" when "01011110000011010", -- t[48154] = 11
      "0001011" when "01011110000011011", -- t[48155] = 11
      "0001011" when "01011110000011100", -- t[48156] = 11
      "0001011" when "01011110000011101", -- t[48157] = 11
      "0001011" when "01011110000011110", -- t[48158] = 11
      "0001011" when "01011110000011111", -- t[48159] = 11
      "0001011" when "01011110000100000", -- t[48160] = 11
      "0001011" when "01011110000100001", -- t[48161] = 11
      "0001011" when "01011110000100010", -- t[48162] = 11
      "0001011" when "01011110000100011", -- t[48163] = 11
      "0001011" when "01011110000100100", -- t[48164] = 11
      "0001011" when "01011110000100101", -- t[48165] = 11
      "0001011" when "01011110000100110", -- t[48166] = 11
      "0001011" when "01011110000100111", -- t[48167] = 11
      "0001011" when "01011110000101000", -- t[48168] = 11
      "0001011" when "01011110000101001", -- t[48169] = 11
      "0001011" when "01011110000101010", -- t[48170] = 11
      "0001011" when "01011110000101011", -- t[48171] = 11
      "0001011" when "01011110000101100", -- t[48172] = 11
      "0001011" when "01011110000101101", -- t[48173] = 11
      "0001011" when "01011110000101110", -- t[48174] = 11
      "0001011" when "01011110000101111", -- t[48175] = 11
      "0001011" when "01011110000110000", -- t[48176] = 11
      "0001011" when "01011110000110001", -- t[48177] = 11
      "0001011" when "01011110000110010", -- t[48178] = 11
      "0001011" when "01011110000110011", -- t[48179] = 11
      "0001011" when "01011110000110100", -- t[48180] = 11
      "0001011" when "01011110000110101", -- t[48181] = 11
      "0001011" when "01011110000110110", -- t[48182] = 11
      "0001011" when "01011110000110111", -- t[48183] = 11
      "0001011" when "01011110000111000", -- t[48184] = 11
      "0001011" when "01011110000111001", -- t[48185] = 11
      "0001011" when "01011110000111010", -- t[48186] = 11
      "0001011" when "01011110000111011", -- t[48187] = 11
      "0001011" when "01011110000111100", -- t[48188] = 11
      "0001011" when "01011110000111101", -- t[48189] = 11
      "0001011" when "01011110000111110", -- t[48190] = 11
      "0001011" when "01011110000111111", -- t[48191] = 11
      "0001011" when "01011110001000000", -- t[48192] = 11
      "0001011" when "01011110001000001", -- t[48193] = 11
      "0001011" when "01011110001000010", -- t[48194] = 11
      "0001011" when "01011110001000011", -- t[48195] = 11
      "0001011" when "01011110001000100", -- t[48196] = 11
      "0001011" when "01011110001000101", -- t[48197] = 11
      "0001011" when "01011110001000110", -- t[48198] = 11
      "0001011" when "01011110001000111", -- t[48199] = 11
      "0001011" when "01011110001001000", -- t[48200] = 11
      "0001011" when "01011110001001001", -- t[48201] = 11
      "0001011" when "01011110001001010", -- t[48202] = 11
      "0001011" when "01011110001001011", -- t[48203] = 11
      "0001011" when "01011110001001100", -- t[48204] = 11
      "0001011" when "01011110001001101", -- t[48205] = 11
      "0001011" when "01011110001001110", -- t[48206] = 11
      "0001011" when "01011110001001111", -- t[48207] = 11
      "0001011" when "01011110001010000", -- t[48208] = 11
      "0001011" when "01011110001010001", -- t[48209] = 11
      "0001011" when "01011110001010010", -- t[48210] = 11
      "0001011" when "01011110001010011", -- t[48211] = 11
      "0001011" when "01011110001010100", -- t[48212] = 11
      "0001011" when "01011110001010101", -- t[48213] = 11
      "0001011" when "01011110001010110", -- t[48214] = 11
      "0001011" when "01011110001010111", -- t[48215] = 11
      "0001011" when "01011110001011000", -- t[48216] = 11
      "0001011" when "01011110001011001", -- t[48217] = 11
      "0001011" when "01011110001011010", -- t[48218] = 11
      "0001011" when "01011110001011011", -- t[48219] = 11
      "0001011" when "01011110001011100", -- t[48220] = 11
      "0001011" when "01011110001011101", -- t[48221] = 11
      "0001011" when "01011110001011110", -- t[48222] = 11
      "0001011" when "01011110001011111", -- t[48223] = 11
      "0001011" when "01011110001100000", -- t[48224] = 11
      "0001011" when "01011110001100001", -- t[48225] = 11
      "0001011" when "01011110001100010", -- t[48226] = 11
      "0001011" when "01011110001100011", -- t[48227] = 11
      "0001011" when "01011110001100100", -- t[48228] = 11
      "0001011" when "01011110001100101", -- t[48229] = 11
      "0001011" when "01011110001100110", -- t[48230] = 11
      "0001011" when "01011110001100111", -- t[48231] = 11
      "0001011" when "01011110001101000", -- t[48232] = 11
      "0001011" when "01011110001101001", -- t[48233] = 11
      "0001011" when "01011110001101010", -- t[48234] = 11
      "0001011" when "01011110001101011", -- t[48235] = 11
      "0001011" when "01011110001101100", -- t[48236] = 11
      "0001011" when "01011110001101101", -- t[48237] = 11
      "0001011" when "01011110001101110", -- t[48238] = 11
      "0001011" when "01011110001101111", -- t[48239] = 11
      "0001011" when "01011110001110000", -- t[48240] = 11
      "0001011" when "01011110001110001", -- t[48241] = 11
      "0001011" when "01011110001110010", -- t[48242] = 11
      "0001011" when "01011110001110011", -- t[48243] = 11
      "0001011" when "01011110001110100", -- t[48244] = 11
      "0001011" when "01011110001110101", -- t[48245] = 11
      "0001011" when "01011110001110110", -- t[48246] = 11
      "0001011" when "01011110001110111", -- t[48247] = 11
      "0001011" when "01011110001111000", -- t[48248] = 11
      "0001011" when "01011110001111001", -- t[48249] = 11
      "0001011" when "01011110001111010", -- t[48250] = 11
      "0001011" when "01011110001111011", -- t[48251] = 11
      "0001011" when "01011110001111100", -- t[48252] = 11
      "0001011" when "01011110001111101", -- t[48253] = 11
      "0001011" when "01011110001111110", -- t[48254] = 11
      "0001011" when "01011110001111111", -- t[48255] = 11
      "0001011" when "01011110010000000", -- t[48256] = 11
      "0001011" when "01011110010000001", -- t[48257] = 11
      "0001011" when "01011110010000010", -- t[48258] = 11
      "0001011" when "01011110010000011", -- t[48259] = 11
      "0001011" when "01011110010000100", -- t[48260] = 11
      "0001011" when "01011110010000101", -- t[48261] = 11
      "0001011" when "01011110010000110", -- t[48262] = 11
      "0001011" when "01011110010000111", -- t[48263] = 11
      "0001011" when "01011110010001000", -- t[48264] = 11
      "0001011" when "01011110010001001", -- t[48265] = 11
      "0001011" when "01011110010001010", -- t[48266] = 11
      "0001011" when "01011110010001011", -- t[48267] = 11
      "0001011" when "01011110010001100", -- t[48268] = 11
      "0001011" when "01011110010001101", -- t[48269] = 11
      "0001011" when "01011110010001110", -- t[48270] = 11
      "0001011" when "01011110010001111", -- t[48271] = 11
      "0001011" when "01011110010010000", -- t[48272] = 11
      "0001011" when "01011110010010001", -- t[48273] = 11
      "0001011" when "01011110010010010", -- t[48274] = 11
      "0001011" when "01011110010010011", -- t[48275] = 11
      "0001011" when "01011110010010100", -- t[48276] = 11
      "0001011" when "01011110010010101", -- t[48277] = 11
      "0001011" when "01011110010010110", -- t[48278] = 11
      "0001011" when "01011110010010111", -- t[48279] = 11
      "0001011" when "01011110010011000", -- t[48280] = 11
      "0001011" when "01011110010011001", -- t[48281] = 11
      "0001011" when "01011110010011010", -- t[48282] = 11
      "0001011" when "01011110010011011", -- t[48283] = 11
      "0001011" when "01011110010011100", -- t[48284] = 11
      "0001011" when "01011110010011101", -- t[48285] = 11
      "0001011" when "01011110010011110", -- t[48286] = 11
      "0001011" when "01011110010011111", -- t[48287] = 11
      "0001011" when "01011110010100000", -- t[48288] = 11
      "0001011" when "01011110010100001", -- t[48289] = 11
      "0001011" when "01011110010100010", -- t[48290] = 11
      "0001011" when "01011110010100011", -- t[48291] = 11
      "0001011" when "01011110010100100", -- t[48292] = 11
      "0001011" when "01011110010100101", -- t[48293] = 11
      "0001011" when "01011110010100110", -- t[48294] = 11
      "0001011" when "01011110010100111", -- t[48295] = 11
      "0001011" when "01011110010101000", -- t[48296] = 11
      "0001011" when "01011110010101001", -- t[48297] = 11
      "0001011" when "01011110010101010", -- t[48298] = 11
      "0001011" when "01011110010101011", -- t[48299] = 11
      "0001011" when "01011110010101100", -- t[48300] = 11
      "0001011" when "01011110010101101", -- t[48301] = 11
      "0001011" when "01011110010101110", -- t[48302] = 11
      "0001011" when "01011110010101111", -- t[48303] = 11
      "0001011" when "01011110010110000", -- t[48304] = 11
      "0001011" when "01011110010110001", -- t[48305] = 11
      "0001011" when "01011110010110010", -- t[48306] = 11
      "0001011" when "01011110010110011", -- t[48307] = 11
      "0001011" when "01011110010110100", -- t[48308] = 11
      "0001011" when "01011110010110101", -- t[48309] = 11
      "0001011" when "01011110010110110", -- t[48310] = 11
      "0001011" when "01011110010110111", -- t[48311] = 11
      "0001011" when "01011110010111000", -- t[48312] = 11
      "0001011" when "01011110010111001", -- t[48313] = 11
      "0001011" when "01011110010111010", -- t[48314] = 11
      "0001011" when "01011110010111011", -- t[48315] = 11
      "0001011" when "01011110010111100", -- t[48316] = 11
      "0001011" when "01011110010111101", -- t[48317] = 11
      "0001011" when "01011110010111110", -- t[48318] = 11
      "0001011" when "01011110010111111", -- t[48319] = 11
      "0001011" when "01011110011000000", -- t[48320] = 11
      "0001011" when "01011110011000001", -- t[48321] = 11
      "0001011" when "01011110011000010", -- t[48322] = 11
      "0001011" when "01011110011000011", -- t[48323] = 11
      "0001011" when "01011110011000100", -- t[48324] = 11
      "0001011" when "01011110011000101", -- t[48325] = 11
      "0001011" when "01011110011000110", -- t[48326] = 11
      "0001011" when "01011110011000111", -- t[48327] = 11
      "0001011" when "01011110011001000", -- t[48328] = 11
      "0001011" when "01011110011001001", -- t[48329] = 11
      "0001011" when "01011110011001010", -- t[48330] = 11
      "0001011" when "01011110011001011", -- t[48331] = 11
      "0001011" when "01011110011001100", -- t[48332] = 11
      "0001011" when "01011110011001101", -- t[48333] = 11
      "0001011" when "01011110011001110", -- t[48334] = 11
      "0001011" when "01011110011001111", -- t[48335] = 11
      "0001011" when "01011110011010000", -- t[48336] = 11
      "0001011" when "01011110011010001", -- t[48337] = 11
      "0001011" when "01011110011010010", -- t[48338] = 11
      "0001011" when "01011110011010011", -- t[48339] = 11
      "0001011" when "01011110011010100", -- t[48340] = 11
      "0001011" when "01011110011010101", -- t[48341] = 11
      "0001011" when "01011110011010110", -- t[48342] = 11
      "0001011" when "01011110011010111", -- t[48343] = 11
      "0001011" when "01011110011011000", -- t[48344] = 11
      "0001011" when "01011110011011001", -- t[48345] = 11
      "0001011" when "01011110011011010", -- t[48346] = 11
      "0001011" when "01011110011011011", -- t[48347] = 11
      "0001011" when "01011110011011100", -- t[48348] = 11
      "0001011" when "01011110011011101", -- t[48349] = 11
      "0001011" when "01011110011011110", -- t[48350] = 11
      "0001011" when "01011110011011111", -- t[48351] = 11
      "0001011" when "01011110011100000", -- t[48352] = 11
      "0001011" when "01011110011100001", -- t[48353] = 11
      "0001011" when "01011110011100010", -- t[48354] = 11
      "0001011" when "01011110011100011", -- t[48355] = 11
      "0001011" when "01011110011100100", -- t[48356] = 11
      "0001011" when "01011110011100101", -- t[48357] = 11
      "0001011" when "01011110011100110", -- t[48358] = 11
      "0001011" when "01011110011100111", -- t[48359] = 11
      "0001011" when "01011110011101000", -- t[48360] = 11
      "0001011" when "01011110011101001", -- t[48361] = 11
      "0001011" when "01011110011101010", -- t[48362] = 11
      "0001011" when "01011110011101011", -- t[48363] = 11
      "0001011" when "01011110011101100", -- t[48364] = 11
      "0001011" when "01011110011101101", -- t[48365] = 11
      "0001011" when "01011110011101110", -- t[48366] = 11
      "0001011" when "01011110011101111", -- t[48367] = 11
      "0001011" when "01011110011110000", -- t[48368] = 11
      "0001011" when "01011110011110001", -- t[48369] = 11
      "0001011" when "01011110011110010", -- t[48370] = 11
      "0001011" when "01011110011110011", -- t[48371] = 11
      "0001011" when "01011110011110100", -- t[48372] = 11
      "0001011" when "01011110011110101", -- t[48373] = 11
      "0001011" when "01011110011110110", -- t[48374] = 11
      "0001011" when "01011110011110111", -- t[48375] = 11
      "0001011" when "01011110011111000", -- t[48376] = 11
      "0001011" when "01011110011111001", -- t[48377] = 11
      "0001011" when "01011110011111010", -- t[48378] = 11
      "0001011" when "01011110011111011", -- t[48379] = 11
      "0001011" when "01011110011111100", -- t[48380] = 11
      "0001011" when "01011110011111101", -- t[48381] = 11
      "0001011" when "01011110011111110", -- t[48382] = 11
      "0001011" when "01011110011111111", -- t[48383] = 11
      "0001011" when "01011110100000000", -- t[48384] = 11
      "0001011" when "01011110100000001", -- t[48385] = 11
      "0001011" when "01011110100000010", -- t[48386] = 11
      "0001011" when "01011110100000011", -- t[48387] = 11
      "0001011" when "01011110100000100", -- t[48388] = 11
      "0001011" when "01011110100000101", -- t[48389] = 11
      "0001011" when "01011110100000110", -- t[48390] = 11
      "0001011" when "01011110100000111", -- t[48391] = 11
      "0001011" when "01011110100001000", -- t[48392] = 11
      "0001011" when "01011110100001001", -- t[48393] = 11
      "0001011" when "01011110100001010", -- t[48394] = 11
      "0001011" when "01011110100001011", -- t[48395] = 11
      "0001011" when "01011110100001100", -- t[48396] = 11
      "0001011" when "01011110100001101", -- t[48397] = 11
      "0001011" when "01011110100001110", -- t[48398] = 11
      "0001011" when "01011110100001111", -- t[48399] = 11
      "0001011" when "01011110100010000", -- t[48400] = 11
      "0001011" when "01011110100010001", -- t[48401] = 11
      "0001011" when "01011110100010010", -- t[48402] = 11
      "0001011" when "01011110100010011", -- t[48403] = 11
      "0001011" when "01011110100010100", -- t[48404] = 11
      "0001011" when "01011110100010101", -- t[48405] = 11
      "0001011" when "01011110100010110", -- t[48406] = 11
      "0001011" when "01011110100010111", -- t[48407] = 11
      "0001011" when "01011110100011000", -- t[48408] = 11
      "0001011" when "01011110100011001", -- t[48409] = 11
      "0001011" when "01011110100011010", -- t[48410] = 11
      "0001011" when "01011110100011011", -- t[48411] = 11
      "0001011" when "01011110100011100", -- t[48412] = 11
      "0001011" when "01011110100011101", -- t[48413] = 11
      "0001011" when "01011110100011110", -- t[48414] = 11
      "0001011" when "01011110100011111", -- t[48415] = 11
      "0001011" when "01011110100100000", -- t[48416] = 11
      "0001011" when "01011110100100001", -- t[48417] = 11
      "0001011" when "01011110100100010", -- t[48418] = 11
      "0001011" when "01011110100100011", -- t[48419] = 11
      "0001011" when "01011110100100100", -- t[48420] = 11
      "0001011" when "01011110100100101", -- t[48421] = 11
      "0001011" when "01011110100100110", -- t[48422] = 11
      "0001011" when "01011110100100111", -- t[48423] = 11
      "0001011" when "01011110100101000", -- t[48424] = 11
      "0001011" when "01011110100101001", -- t[48425] = 11
      "0001011" when "01011110100101010", -- t[48426] = 11
      "0001011" when "01011110100101011", -- t[48427] = 11
      "0001011" when "01011110100101100", -- t[48428] = 11
      "0001011" when "01011110100101101", -- t[48429] = 11
      "0001011" when "01011110100101110", -- t[48430] = 11
      "0001011" when "01011110100101111", -- t[48431] = 11
      "0001011" when "01011110100110000", -- t[48432] = 11
      "0001011" when "01011110100110001", -- t[48433] = 11
      "0001011" when "01011110100110010", -- t[48434] = 11
      "0001011" when "01011110100110011", -- t[48435] = 11
      "0001011" when "01011110100110100", -- t[48436] = 11
      "0001011" when "01011110100110101", -- t[48437] = 11
      "0001011" when "01011110100110110", -- t[48438] = 11
      "0001011" when "01011110100110111", -- t[48439] = 11
      "0001011" when "01011110100111000", -- t[48440] = 11
      "0001011" when "01011110100111001", -- t[48441] = 11
      "0001011" when "01011110100111010", -- t[48442] = 11
      "0001011" when "01011110100111011", -- t[48443] = 11
      "0001011" when "01011110100111100", -- t[48444] = 11
      "0001011" when "01011110100111101", -- t[48445] = 11
      "0001011" when "01011110100111110", -- t[48446] = 11
      "0001011" when "01011110100111111", -- t[48447] = 11
      "0001011" when "01011110101000000", -- t[48448] = 11
      "0001011" when "01011110101000001", -- t[48449] = 11
      "0001011" when "01011110101000010", -- t[48450] = 11
      "0001011" when "01011110101000011", -- t[48451] = 11
      "0001011" when "01011110101000100", -- t[48452] = 11
      "0001011" when "01011110101000101", -- t[48453] = 11
      "0001011" when "01011110101000110", -- t[48454] = 11
      "0001011" when "01011110101000111", -- t[48455] = 11
      "0001011" when "01011110101001000", -- t[48456] = 11
      "0001011" when "01011110101001001", -- t[48457] = 11
      "0001011" when "01011110101001010", -- t[48458] = 11
      "0001011" when "01011110101001011", -- t[48459] = 11
      "0001011" when "01011110101001100", -- t[48460] = 11
      "0001011" when "01011110101001101", -- t[48461] = 11
      "0001011" when "01011110101001110", -- t[48462] = 11
      "0001011" when "01011110101001111", -- t[48463] = 11
      "0001011" when "01011110101010000", -- t[48464] = 11
      "0001011" when "01011110101010001", -- t[48465] = 11
      "0001011" when "01011110101010010", -- t[48466] = 11
      "0001011" when "01011110101010011", -- t[48467] = 11
      "0001011" when "01011110101010100", -- t[48468] = 11
      "0001011" when "01011110101010101", -- t[48469] = 11
      "0001011" when "01011110101010110", -- t[48470] = 11
      "0001011" when "01011110101010111", -- t[48471] = 11
      "0001011" when "01011110101011000", -- t[48472] = 11
      "0001011" when "01011110101011001", -- t[48473] = 11
      "0001011" when "01011110101011010", -- t[48474] = 11
      "0001011" when "01011110101011011", -- t[48475] = 11
      "0001011" when "01011110101011100", -- t[48476] = 11
      "0001011" when "01011110101011101", -- t[48477] = 11
      "0001011" when "01011110101011110", -- t[48478] = 11
      "0001011" when "01011110101011111", -- t[48479] = 11
      "0001011" when "01011110101100000", -- t[48480] = 11
      "0001011" when "01011110101100001", -- t[48481] = 11
      "0001011" when "01011110101100010", -- t[48482] = 11
      "0001011" when "01011110101100011", -- t[48483] = 11
      "0001011" when "01011110101100100", -- t[48484] = 11
      "0001011" when "01011110101100101", -- t[48485] = 11
      "0001011" when "01011110101100110", -- t[48486] = 11
      "0001011" when "01011110101100111", -- t[48487] = 11
      "0001011" when "01011110101101000", -- t[48488] = 11
      "0001011" when "01011110101101001", -- t[48489] = 11
      "0001011" when "01011110101101010", -- t[48490] = 11
      "0001011" when "01011110101101011", -- t[48491] = 11
      "0001011" when "01011110101101100", -- t[48492] = 11
      "0001011" when "01011110101101101", -- t[48493] = 11
      "0001011" when "01011110101101110", -- t[48494] = 11
      "0001011" when "01011110101101111", -- t[48495] = 11
      "0001011" when "01011110101110000", -- t[48496] = 11
      "0001011" when "01011110101110001", -- t[48497] = 11
      "0001011" when "01011110101110010", -- t[48498] = 11
      "0001011" when "01011110101110011", -- t[48499] = 11
      "0001011" when "01011110101110100", -- t[48500] = 11
      "0001011" when "01011110101110101", -- t[48501] = 11
      "0001011" when "01011110101110110", -- t[48502] = 11
      "0001011" when "01011110101110111", -- t[48503] = 11
      "0001011" when "01011110101111000", -- t[48504] = 11
      "0001011" when "01011110101111001", -- t[48505] = 11
      "0001011" when "01011110101111010", -- t[48506] = 11
      "0001011" when "01011110101111011", -- t[48507] = 11
      "0001011" when "01011110101111100", -- t[48508] = 11
      "0001011" when "01011110101111101", -- t[48509] = 11
      "0001011" when "01011110101111110", -- t[48510] = 11
      "0001011" when "01011110101111111", -- t[48511] = 11
      "0001011" when "01011110110000000", -- t[48512] = 11
      "0001011" when "01011110110000001", -- t[48513] = 11
      "0001011" when "01011110110000010", -- t[48514] = 11
      "0001011" when "01011110110000011", -- t[48515] = 11
      "0001011" when "01011110110000100", -- t[48516] = 11
      "0001011" when "01011110110000101", -- t[48517] = 11
      "0001011" when "01011110110000110", -- t[48518] = 11
      "0001011" when "01011110110000111", -- t[48519] = 11
      "0001011" when "01011110110001000", -- t[48520] = 11
      "0001011" when "01011110110001001", -- t[48521] = 11
      "0001011" when "01011110110001010", -- t[48522] = 11
      "0001011" when "01011110110001011", -- t[48523] = 11
      "0001011" when "01011110110001100", -- t[48524] = 11
      "0001011" when "01011110110001101", -- t[48525] = 11
      "0001011" when "01011110110001110", -- t[48526] = 11
      "0001011" when "01011110110001111", -- t[48527] = 11
      "0001011" when "01011110110010000", -- t[48528] = 11
      "0001011" when "01011110110010001", -- t[48529] = 11
      "0001011" when "01011110110010010", -- t[48530] = 11
      "0001011" when "01011110110010011", -- t[48531] = 11
      "0001011" when "01011110110010100", -- t[48532] = 11
      "0001011" when "01011110110010101", -- t[48533] = 11
      "0001011" when "01011110110010110", -- t[48534] = 11
      "0001011" when "01011110110010111", -- t[48535] = 11
      "0001011" when "01011110110011000", -- t[48536] = 11
      "0001011" when "01011110110011001", -- t[48537] = 11
      "0001011" when "01011110110011010", -- t[48538] = 11
      "0001011" when "01011110110011011", -- t[48539] = 11
      "0001011" when "01011110110011100", -- t[48540] = 11
      "0001011" when "01011110110011101", -- t[48541] = 11
      "0001011" when "01011110110011110", -- t[48542] = 11
      "0001011" when "01011110110011111", -- t[48543] = 11
      "0001011" when "01011110110100000", -- t[48544] = 11
      "0001011" when "01011110110100001", -- t[48545] = 11
      "0001011" when "01011110110100010", -- t[48546] = 11
      "0001011" when "01011110110100011", -- t[48547] = 11
      "0001011" when "01011110110100100", -- t[48548] = 11
      "0001011" when "01011110110100101", -- t[48549] = 11
      "0001011" when "01011110110100110", -- t[48550] = 11
      "0001011" when "01011110110100111", -- t[48551] = 11
      "0001011" when "01011110110101000", -- t[48552] = 11
      "0001011" when "01011110110101001", -- t[48553] = 11
      "0001011" when "01011110110101010", -- t[48554] = 11
      "0001011" when "01011110110101011", -- t[48555] = 11
      "0001011" when "01011110110101100", -- t[48556] = 11
      "0001011" when "01011110110101101", -- t[48557] = 11
      "0001011" when "01011110110101110", -- t[48558] = 11
      "0001011" when "01011110110101111", -- t[48559] = 11
      "0001011" when "01011110110110000", -- t[48560] = 11
      "0001011" when "01011110110110001", -- t[48561] = 11
      "0001011" when "01011110110110010", -- t[48562] = 11
      "0001011" when "01011110110110011", -- t[48563] = 11
      "0001011" when "01011110110110100", -- t[48564] = 11
      "0001011" when "01011110110110101", -- t[48565] = 11
      "0001011" when "01011110110110110", -- t[48566] = 11
      "0001011" when "01011110110110111", -- t[48567] = 11
      "0001011" when "01011110110111000", -- t[48568] = 11
      "0001011" when "01011110110111001", -- t[48569] = 11
      "0001011" when "01011110110111010", -- t[48570] = 11
      "0001011" when "01011110110111011", -- t[48571] = 11
      "0001011" when "01011110110111100", -- t[48572] = 11
      "0001011" when "01011110110111101", -- t[48573] = 11
      "0001011" when "01011110110111110", -- t[48574] = 11
      "0001011" when "01011110110111111", -- t[48575] = 11
      "0001011" when "01011110111000000", -- t[48576] = 11
      "0001011" when "01011110111000001", -- t[48577] = 11
      "0001011" when "01011110111000010", -- t[48578] = 11
      "0001011" when "01011110111000011", -- t[48579] = 11
      "0001011" when "01011110111000100", -- t[48580] = 11
      "0001011" when "01011110111000101", -- t[48581] = 11
      "0001011" when "01011110111000110", -- t[48582] = 11
      "0001011" when "01011110111000111", -- t[48583] = 11
      "0001011" when "01011110111001000", -- t[48584] = 11
      "0001011" when "01011110111001001", -- t[48585] = 11
      "0001011" when "01011110111001010", -- t[48586] = 11
      "0001011" when "01011110111001011", -- t[48587] = 11
      "0001011" when "01011110111001100", -- t[48588] = 11
      "0001011" when "01011110111001101", -- t[48589] = 11
      "0001011" when "01011110111001110", -- t[48590] = 11
      "0001011" when "01011110111001111", -- t[48591] = 11
      "0001011" when "01011110111010000", -- t[48592] = 11
      "0001011" when "01011110111010001", -- t[48593] = 11
      "0001011" when "01011110111010010", -- t[48594] = 11
      "0001011" when "01011110111010011", -- t[48595] = 11
      "0001011" when "01011110111010100", -- t[48596] = 11
      "0001011" when "01011110111010101", -- t[48597] = 11
      "0001011" when "01011110111010110", -- t[48598] = 11
      "0001011" when "01011110111010111", -- t[48599] = 11
      "0001011" when "01011110111011000", -- t[48600] = 11
      "0001011" when "01011110111011001", -- t[48601] = 11
      "0001011" when "01011110111011010", -- t[48602] = 11
      "0001011" when "01011110111011011", -- t[48603] = 11
      "0001011" when "01011110111011100", -- t[48604] = 11
      "0001011" when "01011110111011101", -- t[48605] = 11
      "0001011" when "01011110111011110", -- t[48606] = 11
      "0001011" when "01011110111011111", -- t[48607] = 11
      "0001011" when "01011110111100000", -- t[48608] = 11
      "0001011" when "01011110111100001", -- t[48609] = 11
      "0001011" when "01011110111100010", -- t[48610] = 11
      "0001011" when "01011110111100011", -- t[48611] = 11
      "0001011" when "01011110111100100", -- t[48612] = 11
      "0001011" when "01011110111100101", -- t[48613] = 11
      "0001011" when "01011110111100110", -- t[48614] = 11
      "0001011" when "01011110111100111", -- t[48615] = 11
      "0001011" when "01011110111101000", -- t[48616] = 11
      "0001011" when "01011110111101001", -- t[48617] = 11
      "0001011" when "01011110111101010", -- t[48618] = 11
      "0001011" when "01011110111101011", -- t[48619] = 11
      "0001011" when "01011110111101100", -- t[48620] = 11
      "0001011" when "01011110111101101", -- t[48621] = 11
      "0001011" when "01011110111101110", -- t[48622] = 11
      "0001011" when "01011110111101111", -- t[48623] = 11
      "0001011" when "01011110111110000", -- t[48624] = 11
      "0001011" when "01011110111110001", -- t[48625] = 11
      "0001011" when "01011110111110010", -- t[48626] = 11
      "0001011" when "01011110111110011", -- t[48627] = 11
      "0001011" when "01011110111110100", -- t[48628] = 11
      "0001011" when "01011110111110101", -- t[48629] = 11
      "0001011" when "01011110111110110", -- t[48630] = 11
      "0001011" when "01011110111110111", -- t[48631] = 11
      "0001011" when "01011110111111000", -- t[48632] = 11
      "0001011" when "01011110111111001", -- t[48633] = 11
      "0001011" when "01011110111111010", -- t[48634] = 11
      "0001011" when "01011110111111011", -- t[48635] = 11
      "0001011" when "01011110111111100", -- t[48636] = 11
      "0001011" when "01011110111111101", -- t[48637] = 11
      "0001011" when "01011110111111110", -- t[48638] = 11
      "0001011" when "01011110111111111", -- t[48639] = 11
      "0001011" when "01011111000000000", -- t[48640] = 11
      "0001011" when "01011111000000001", -- t[48641] = 11
      "0001011" when "01011111000000010", -- t[48642] = 11
      "0001011" when "01011111000000011", -- t[48643] = 11
      "0001011" when "01011111000000100", -- t[48644] = 11
      "0001011" when "01011111000000101", -- t[48645] = 11
      "0001011" when "01011111000000110", -- t[48646] = 11
      "0001011" when "01011111000000111", -- t[48647] = 11
      "0001011" when "01011111000001000", -- t[48648] = 11
      "0001011" when "01011111000001001", -- t[48649] = 11
      "0001011" when "01011111000001010", -- t[48650] = 11
      "0001011" when "01011111000001011", -- t[48651] = 11
      "0001011" when "01011111000001100", -- t[48652] = 11
      "0001011" when "01011111000001101", -- t[48653] = 11
      "0001011" when "01011111000001110", -- t[48654] = 11
      "0001011" when "01011111000001111", -- t[48655] = 11
      "0001011" when "01011111000010000", -- t[48656] = 11
      "0001011" when "01011111000010001", -- t[48657] = 11
      "0001011" when "01011111000010010", -- t[48658] = 11
      "0001011" when "01011111000010011", -- t[48659] = 11
      "0001011" when "01011111000010100", -- t[48660] = 11
      "0001011" when "01011111000010101", -- t[48661] = 11
      "0001011" when "01011111000010110", -- t[48662] = 11
      "0001011" when "01011111000010111", -- t[48663] = 11
      "0001011" when "01011111000011000", -- t[48664] = 11
      "0001011" when "01011111000011001", -- t[48665] = 11
      "0001011" when "01011111000011010", -- t[48666] = 11
      "0001011" when "01011111000011011", -- t[48667] = 11
      "0001011" when "01011111000011100", -- t[48668] = 11
      "0001011" when "01011111000011101", -- t[48669] = 11
      "0001011" when "01011111000011110", -- t[48670] = 11
      "0001011" when "01011111000011111", -- t[48671] = 11
      "0001011" when "01011111000100000", -- t[48672] = 11
      "0001011" when "01011111000100001", -- t[48673] = 11
      "0001011" when "01011111000100010", -- t[48674] = 11
      "0001011" when "01011111000100011", -- t[48675] = 11
      "0001011" when "01011111000100100", -- t[48676] = 11
      "0001011" when "01011111000100101", -- t[48677] = 11
      "0001011" when "01011111000100110", -- t[48678] = 11
      "0001011" when "01011111000100111", -- t[48679] = 11
      "0001011" when "01011111000101000", -- t[48680] = 11
      "0001011" when "01011111000101001", -- t[48681] = 11
      "0001011" when "01011111000101010", -- t[48682] = 11
      "0001011" when "01011111000101011", -- t[48683] = 11
      "0001011" when "01011111000101100", -- t[48684] = 11
      "0001011" when "01011111000101101", -- t[48685] = 11
      "0001011" when "01011111000101110", -- t[48686] = 11
      "0001011" when "01011111000101111", -- t[48687] = 11
      "0001011" when "01011111000110000", -- t[48688] = 11
      "0001011" when "01011111000110001", -- t[48689] = 11
      "0001011" when "01011111000110010", -- t[48690] = 11
      "0001011" when "01011111000110011", -- t[48691] = 11
      "0001011" when "01011111000110100", -- t[48692] = 11
      "0001011" when "01011111000110101", -- t[48693] = 11
      "0001011" when "01011111000110110", -- t[48694] = 11
      "0001011" when "01011111000110111", -- t[48695] = 11
      "0001011" when "01011111000111000", -- t[48696] = 11
      "0001011" when "01011111000111001", -- t[48697] = 11
      "0001011" when "01011111000111010", -- t[48698] = 11
      "0001011" when "01011111000111011", -- t[48699] = 11
      "0001011" when "01011111000111100", -- t[48700] = 11
      "0001011" when "01011111000111101", -- t[48701] = 11
      "0001011" when "01011111000111110", -- t[48702] = 11
      "0001011" when "01011111000111111", -- t[48703] = 11
      "0001011" when "01011111001000000", -- t[48704] = 11
      "0001011" when "01011111001000001", -- t[48705] = 11
      "0001011" when "01011111001000010", -- t[48706] = 11
      "0001011" when "01011111001000011", -- t[48707] = 11
      "0001011" when "01011111001000100", -- t[48708] = 11
      "0001011" when "01011111001000101", -- t[48709] = 11
      "0001011" when "01011111001000110", -- t[48710] = 11
      "0001011" when "01011111001000111", -- t[48711] = 11
      "0001011" when "01011111001001000", -- t[48712] = 11
      "0001011" when "01011111001001001", -- t[48713] = 11
      "0001011" when "01011111001001010", -- t[48714] = 11
      "0001011" when "01011111001001011", -- t[48715] = 11
      "0001011" when "01011111001001100", -- t[48716] = 11
      "0001011" when "01011111001001101", -- t[48717] = 11
      "0001011" when "01011111001001110", -- t[48718] = 11
      "0001011" when "01011111001001111", -- t[48719] = 11
      "0001011" when "01011111001010000", -- t[48720] = 11
      "0001011" when "01011111001010001", -- t[48721] = 11
      "0001011" when "01011111001010010", -- t[48722] = 11
      "0001011" when "01011111001010011", -- t[48723] = 11
      "0001011" when "01011111001010100", -- t[48724] = 11
      "0001011" when "01011111001010101", -- t[48725] = 11
      "0001011" when "01011111001010110", -- t[48726] = 11
      "0001011" when "01011111001010111", -- t[48727] = 11
      "0001011" when "01011111001011000", -- t[48728] = 11
      "0001011" when "01011111001011001", -- t[48729] = 11
      "0001011" when "01011111001011010", -- t[48730] = 11
      "0001011" when "01011111001011011", -- t[48731] = 11
      "0001011" when "01011111001011100", -- t[48732] = 11
      "0001011" when "01011111001011101", -- t[48733] = 11
      "0001011" when "01011111001011110", -- t[48734] = 11
      "0001011" when "01011111001011111", -- t[48735] = 11
      "0001011" when "01011111001100000", -- t[48736] = 11
      "0001011" when "01011111001100001", -- t[48737] = 11
      "0001011" when "01011111001100010", -- t[48738] = 11
      "0001011" when "01011111001100011", -- t[48739] = 11
      "0001011" when "01011111001100100", -- t[48740] = 11
      "0001011" when "01011111001100101", -- t[48741] = 11
      "0001011" when "01011111001100110", -- t[48742] = 11
      "0001011" when "01011111001100111", -- t[48743] = 11
      "0001011" when "01011111001101000", -- t[48744] = 11
      "0001011" when "01011111001101001", -- t[48745] = 11
      "0001011" when "01011111001101010", -- t[48746] = 11
      "0001011" when "01011111001101011", -- t[48747] = 11
      "0001011" when "01011111001101100", -- t[48748] = 11
      "0001011" when "01011111001101101", -- t[48749] = 11
      "0001011" when "01011111001101110", -- t[48750] = 11
      "0001011" when "01011111001101111", -- t[48751] = 11
      "0001011" when "01011111001110000", -- t[48752] = 11
      "0001011" when "01011111001110001", -- t[48753] = 11
      "0001011" when "01011111001110010", -- t[48754] = 11
      "0001011" when "01011111001110011", -- t[48755] = 11
      "0001011" when "01011111001110100", -- t[48756] = 11
      "0001011" when "01011111001110101", -- t[48757] = 11
      "0001011" when "01011111001110110", -- t[48758] = 11
      "0001011" when "01011111001110111", -- t[48759] = 11
      "0001011" when "01011111001111000", -- t[48760] = 11
      "0001011" when "01011111001111001", -- t[48761] = 11
      "0001011" when "01011111001111010", -- t[48762] = 11
      "0001011" when "01011111001111011", -- t[48763] = 11
      "0001011" when "01011111001111100", -- t[48764] = 11
      "0001011" when "01011111001111101", -- t[48765] = 11
      "0001011" when "01011111001111110", -- t[48766] = 11
      "0001011" when "01011111001111111", -- t[48767] = 11
      "0001011" when "01011111010000000", -- t[48768] = 11
      "0001011" when "01011111010000001", -- t[48769] = 11
      "0001011" when "01011111010000010", -- t[48770] = 11
      "0001011" when "01011111010000011", -- t[48771] = 11
      "0001011" when "01011111010000100", -- t[48772] = 11
      "0001011" when "01011111010000101", -- t[48773] = 11
      "0001011" when "01011111010000110", -- t[48774] = 11
      "0001011" when "01011111010000111", -- t[48775] = 11
      "0001011" when "01011111010001000", -- t[48776] = 11
      "0001011" when "01011111010001001", -- t[48777] = 11
      "0001011" when "01011111010001010", -- t[48778] = 11
      "0001011" when "01011111010001011", -- t[48779] = 11
      "0001011" when "01011111010001100", -- t[48780] = 11
      "0001011" when "01011111010001101", -- t[48781] = 11
      "0001011" when "01011111010001110", -- t[48782] = 11
      "0001011" when "01011111010001111", -- t[48783] = 11
      "0001011" when "01011111010010000", -- t[48784] = 11
      "0001011" when "01011111010010001", -- t[48785] = 11
      "0001011" when "01011111010010010", -- t[48786] = 11
      "0001011" when "01011111010010011", -- t[48787] = 11
      "0001011" when "01011111010010100", -- t[48788] = 11
      "0001011" when "01011111010010101", -- t[48789] = 11
      "0001011" when "01011111010010110", -- t[48790] = 11
      "0001011" when "01011111010010111", -- t[48791] = 11
      "0001011" when "01011111010011000", -- t[48792] = 11
      "0001011" when "01011111010011001", -- t[48793] = 11
      "0001011" when "01011111010011010", -- t[48794] = 11
      "0001011" when "01011111010011011", -- t[48795] = 11
      "0001011" when "01011111010011100", -- t[48796] = 11
      "0001011" when "01011111010011101", -- t[48797] = 11
      "0001011" when "01011111010011110", -- t[48798] = 11
      "0001011" when "01011111010011111", -- t[48799] = 11
      "0001011" when "01011111010100000", -- t[48800] = 11
      "0001011" when "01011111010100001", -- t[48801] = 11
      "0001011" when "01011111010100010", -- t[48802] = 11
      "0001011" when "01011111010100011", -- t[48803] = 11
      "0001011" when "01011111010100100", -- t[48804] = 11
      "0001011" when "01011111010100101", -- t[48805] = 11
      "0001011" when "01011111010100110", -- t[48806] = 11
      "0001011" when "01011111010100111", -- t[48807] = 11
      "0001011" when "01011111010101000", -- t[48808] = 11
      "0001011" when "01011111010101001", -- t[48809] = 11
      "0001011" when "01011111010101010", -- t[48810] = 11
      "0001011" when "01011111010101011", -- t[48811] = 11
      "0001011" when "01011111010101100", -- t[48812] = 11
      "0001011" when "01011111010101101", -- t[48813] = 11
      "0001011" when "01011111010101110", -- t[48814] = 11
      "0001011" when "01011111010101111", -- t[48815] = 11
      "0001011" when "01011111010110000", -- t[48816] = 11
      "0001011" when "01011111010110001", -- t[48817] = 11
      "0001011" when "01011111010110010", -- t[48818] = 11
      "0001011" when "01011111010110011", -- t[48819] = 11
      "0001011" when "01011111010110100", -- t[48820] = 11
      "0001011" when "01011111010110101", -- t[48821] = 11
      "0001011" when "01011111010110110", -- t[48822] = 11
      "0001011" when "01011111010110111", -- t[48823] = 11
      "0001011" when "01011111010111000", -- t[48824] = 11
      "0001011" when "01011111010111001", -- t[48825] = 11
      "0001011" when "01011111010111010", -- t[48826] = 11
      "0001011" when "01011111010111011", -- t[48827] = 11
      "0001011" when "01011111010111100", -- t[48828] = 11
      "0001011" when "01011111010111101", -- t[48829] = 11
      "0001011" when "01011111010111110", -- t[48830] = 11
      "0001011" when "01011111010111111", -- t[48831] = 11
      "0001011" when "01011111011000000", -- t[48832] = 11
      "0001011" when "01011111011000001", -- t[48833] = 11
      "0001011" when "01011111011000010", -- t[48834] = 11
      "0001011" when "01011111011000011", -- t[48835] = 11
      "0001011" when "01011111011000100", -- t[48836] = 11
      "0001011" when "01011111011000101", -- t[48837] = 11
      "0001011" when "01011111011000110", -- t[48838] = 11
      "0001011" when "01011111011000111", -- t[48839] = 11
      "0001011" when "01011111011001000", -- t[48840] = 11
      "0001011" when "01011111011001001", -- t[48841] = 11
      "0001011" when "01011111011001010", -- t[48842] = 11
      "0001011" when "01011111011001011", -- t[48843] = 11
      "0001011" when "01011111011001100", -- t[48844] = 11
      "0001011" when "01011111011001101", -- t[48845] = 11
      "0001011" when "01011111011001110", -- t[48846] = 11
      "0001011" when "01011111011001111", -- t[48847] = 11
      "0001011" when "01011111011010000", -- t[48848] = 11
      "0001011" when "01011111011010001", -- t[48849] = 11
      "0001011" when "01011111011010010", -- t[48850] = 11
      "0001011" when "01011111011010011", -- t[48851] = 11
      "0001011" when "01011111011010100", -- t[48852] = 11
      "0001011" when "01011111011010101", -- t[48853] = 11
      "0001011" when "01011111011010110", -- t[48854] = 11
      "0001011" when "01011111011010111", -- t[48855] = 11
      "0001011" when "01011111011011000", -- t[48856] = 11
      "0001011" when "01011111011011001", -- t[48857] = 11
      "0001011" when "01011111011011010", -- t[48858] = 11
      "0001011" when "01011111011011011", -- t[48859] = 11
      "0001011" when "01011111011011100", -- t[48860] = 11
      "0001011" when "01011111011011101", -- t[48861] = 11
      "0001011" when "01011111011011110", -- t[48862] = 11
      "0001011" when "01011111011011111", -- t[48863] = 11
      "0001011" when "01011111011100000", -- t[48864] = 11
      "0001011" when "01011111011100001", -- t[48865] = 11
      "0001011" when "01011111011100010", -- t[48866] = 11
      "0001011" when "01011111011100011", -- t[48867] = 11
      "0001011" when "01011111011100100", -- t[48868] = 11
      "0001011" when "01011111011100101", -- t[48869] = 11
      "0001011" when "01011111011100110", -- t[48870] = 11
      "0001011" when "01011111011100111", -- t[48871] = 11
      "0001011" when "01011111011101000", -- t[48872] = 11
      "0001011" when "01011111011101001", -- t[48873] = 11
      "0001011" when "01011111011101010", -- t[48874] = 11
      "0001011" when "01011111011101011", -- t[48875] = 11
      "0001011" when "01011111011101100", -- t[48876] = 11
      "0001011" when "01011111011101101", -- t[48877] = 11
      "0001011" when "01011111011101110", -- t[48878] = 11
      "0001011" when "01011111011101111", -- t[48879] = 11
      "0001011" when "01011111011110000", -- t[48880] = 11
      "0001011" when "01011111011110001", -- t[48881] = 11
      "0001011" when "01011111011110010", -- t[48882] = 11
      "0001011" when "01011111011110011", -- t[48883] = 11
      "0001011" when "01011111011110100", -- t[48884] = 11
      "0001011" when "01011111011110101", -- t[48885] = 11
      "0001011" when "01011111011110110", -- t[48886] = 11
      "0001011" when "01011111011110111", -- t[48887] = 11
      "0001011" when "01011111011111000", -- t[48888] = 11
      "0001011" when "01011111011111001", -- t[48889] = 11
      "0001011" when "01011111011111010", -- t[48890] = 11
      "0001011" when "01011111011111011", -- t[48891] = 11
      "0001011" when "01011111011111100", -- t[48892] = 11
      "0001011" when "01011111011111101", -- t[48893] = 11
      "0001011" when "01011111011111110", -- t[48894] = 11
      "0001011" when "01011111011111111", -- t[48895] = 11
      "0001011" when "01011111100000000", -- t[48896] = 11
      "0001011" when "01011111100000001", -- t[48897] = 11
      "0001011" when "01011111100000010", -- t[48898] = 11
      "0001011" when "01011111100000011", -- t[48899] = 11
      "0001011" when "01011111100000100", -- t[48900] = 11
      "0001011" when "01011111100000101", -- t[48901] = 11
      "0001011" when "01011111100000110", -- t[48902] = 11
      "0001011" when "01011111100000111", -- t[48903] = 11
      "0001011" when "01011111100001000", -- t[48904] = 11
      "0001011" when "01011111100001001", -- t[48905] = 11
      "0001011" when "01011111100001010", -- t[48906] = 11
      "0001011" when "01011111100001011", -- t[48907] = 11
      "0001011" when "01011111100001100", -- t[48908] = 11
      "0001011" when "01011111100001101", -- t[48909] = 11
      "0001011" when "01011111100001110", -- t[48910] = 11
      "0001011" when "01011111100001111", -- t[48911] = 11
      "0001011" when "01011111100010000", -- t[48912] = 11
      "0001011" when "01011111100010001", -- t[48913] = 11
      "0001011" when "01011111100010010", -- t[48914] = 11
      "0001011" when "01011111100010011", -- t[48915] = 11
      "0001011" when "01011111100010100", -- t[48916] = 11
      "0001011" when "01011111100010101", -- t[48917] = 11
      "0001011" when "01011111100010110", -- t[48918] = 11
      "0001011" when "01011111100010111", -- t[48919] = 11
      "0001011" when "01011111100011000", -- t[48920] = 11
      "0001011" when "01011111100011001", -- t[48921] = 11
      "0001011" when "01011111100011010", -- t[48922] = 11
      "0001011" when "01011111100011011", -- t[48923] = 11
      "0001011" when "01011111100011100", -- t[48924] = 11
      "0001011" when "01011111100011101", -- t[48925] = 11
      "0001011" when "01011111100011110", -- t[48926] = 11
      "0001011" when "01011111100011111", -- t[48927] = 11
      "0001011" when "01011111100100000", -- t[48928] = 11
      "0001011" when "01011111100100001", -- t[48929] = 11
      "0001011" when "01011111100100010", -- t[48930] = 11
      "0001011" when "01011111100100011", -- t[48931] = 11
      "0001011" when "01011111100100100", -- t[48932] = 11
      "0001011" when "01011111100100101", -- t[48933] = 11
      "0001011" when "01011111100100110", -- t[48934] = 11
      "0001011" when "01011111100100111", -- t[48935] = 11
      "0001011" when "01011111100101000", -- t[48936] = 11
      "0001011" when "01011111100101001", -- t[48937] = 11
      "0001011" when "01011111100101010", -- t[48938] = 11
      "0001011" when "01011111100101011", -- t[48939] = 11
      "0001011" when "01011111100101100", -- t[48940] = 11
      "0001011" when "01011111100101101", -- t[48941] = 11
      "0001011" when "01011111100101110", -- t[48942] = 11
      "0001011" when "01011111100101111", -- t[48943] = 11
      "0001011" when "01011111100110000", -- t[48944] = 11
      "0001011" when "01011111100110001", -- t[48945] = 11
      "0001011" when "01011111100110010", -- t[48946] = 11
      "0001011" when "01011111100110011", -- t[48947] = 11
      "0001011" when "01011111100110100", -- t[48948] = 11
      "0001011" when "01011111100110101", -- t[48949] = 11
      "0001011" when "01011111100110110", -- t[48950] = 11
      "0001011" when "01011111100110111", -- t[48951] = 11
      "0001011" when "01011111100111000", -- t[48952] = 11
      "0001011" when "01011111100111001", -- t[48953] = 11
      "0001011" when "01011111100111010", -- t[48954] = 11
      "0001011" when "01011111100111011", -- t[48955] = 11
      "0001011" when "01011111100111100", -- t[48956] = 11
      "0001011" when "01011111100111101", -- t[48957] = 11
      "0001011" when "01011111100111110", -- t[48958] = 11
      "0001011" when "01011111100111111", -- t[48959] = 11
      "0001011" when "01011111101000000", -- t[48960] = 11
      "0001011" when "01011111101000001", -- t[48961] = 11
      "0001011" when "01011111101000010", -- t[48962] = 11
      "0001011" when "01011111101000011", -- t[48963] = 11
      "0001011" when "01011111101000100", -- t[48964] = 11
      "0001011" when "01011111101000101", -- t[48965] = 11
      "0001011" when "01011111101000110", -- t[48966] = 11
      "0001011" when "01011111101000111", -- t[48967] = 11
      "0001011" when "01011111101001000", -- t[48968] = 11
      "0001011" when "01011111101001001", -- t[48969] = 11
      "0001011" when "01011111101001010", -- t[48970] = 11
      "0001011" when "01011111101001011", -- t[48971] = 11
      "0001011" when "01011111101001100", -- t[48972] = 11
      "0001011" when "01011111101001101", -- t[48973] = 11
      "0001011" when "01011111101001110", -- t[48974] = 11
      "0001011" when "01011111101001111", -- t[48975] = 11
      "0001011" when "01011111101010000", -- t[48976] = 11
      "0001011" when "01011111101010001", -- t[48977] = 11
      "0001011" when "01011111101010010", -- t[48978] = 11
      "0001011" when "01011111101010011", -- t[48979] = 11
      "0001011" when "01011111101010100", -- t[48980] = 11
      "0001011" when "01011111101010101", -- t[48981] = 11
      "0001011" when "01011111101010110", -- t[48982] = 11
      "0001011" when "01011111101010111", -- t[48983] = 11
      "0001011" when "01011111101011000", -- t[48984] = 11
      "0001011" when "01011111101011001", -- t[48985] = 11
      "0001011" when "01011111101011010", -- t[48986] = 11
      "0001011" when "01011111101011011", -- t[48987] = 11
      "0001011" when "01011111101011100", -- t[48988] = 11
      "0001011" when "01011111101011101", -- t[48989] = 11
      "0001011" when "01011111101011110", -- t[48990] = 11
      "0001011" when "01011111101011111", -- t[48991] = 11
      "0001011" when "01011111101100000", -- t[48992] = 11
      "0001011" when "01011111101100001", -- t[48993] = 11
      "0001011" when "01011111101100010", -- t[48994] = 11
      "0001011" when "01011111101100011", -- t[48995] = 11
      "0001011" when "01011111101100100", -- t[48996] = 11
      "0001011" when "01011111101100101", -- t[48997] = 11
      "0001011" when "01011111101100110", -- t[48998] = 11
      "0001011" when "01011111101100111", -- t[48999] = 11
      "0001011" when "01011111101101000", -- t[49000] = 11
      "0001011" when "01011111101101001", -- t[49001] = 11
      "0001011" when "01011111101101010", -- t[49002] = 11
      "0001011" when "01011111101101011", -- t[49003] = 11
      "0001011" when "01011111101101100", -- t[49004] = 11
      "0001011" when "01011111101101101", -- t[49005] = 11
      "0001011" when "01011111101101110", -- t[49006] = 11
      "0001011" when "01011111101101111", -- t[49007] = 11
      "0001011" when "01011111101110000", -- t[49008] = 11
      "0001011" when "01011111101110001", -- t[49009] = 11
      "0001011" when "01011111101110010", -- t[49010] = 11
      "0001011" when "01011111101110011", -- t[49011] = 11
      "0001011" when "01011111101110100", -- t[49012] = 11
      "0001011" when "01011111101110101", -- t[49013] = 11
      "0001011" when "01011111101110110", -- t[49014] = 11
      "0001011" when "01011111101110111", -- t[49015] = 11
      "0001011" when "01011111101111000", -- t[49016] = 11
      "0001011" when "01011111101111001", -- t[49017] = 11
      "0001011" when "01011111101111010", -- t[49018] = 11
      "0001011" when "01011111101111011", -- t[49019] = 11
      "0001011" when "01011111101111100", -- t[49020] = 11
      "0001011" when "01011111101111101", -- t[49021] = 11
      "0001011" when "01011111101111110", -- t[49022] = 11
      "0001011" when "01011111101111111", -- t[49023] = 11
      "0001011" when "01011111110000000", -- t[49024] = 11
      "0001011" when "01011111110000001", -- t[49025] = 11
      "0001011" when "01011111110000010", -- t[49026] = 11
      "0001011" when "01011111110000011", -- t[49027] = 11
      "0001011" when "01011111110000100", -- t[49028] = 11
      "0001011" when "01011111110000101", -- t[49029] = 11
      "0001011" when "01011111110000110", -- t[49030] = 11
      "0001011" when "01011111110000111", -- t[49031] = 11
      "0001011" when "01011111110001000", -- t[49032] = 11
      "0001011" when "01011111110001001", -- t[49033] = 11
      "0001011" when "01011111110001010", -- t[49034] = 11
      "0001011" when "01011111110001011", -- t[49035] = 11
      "0001011" when "01011111110001100", -- t[49036] = 11
      "0001011" when "01011111110001101", -- t[49037] = 11
      "0001011" when "01011111110001110", -- t[49038] = 11
      "0001011" when "01011111110001111", -- t[49039] = 11
      "0001011" when "01011111110010000", -- t[49040] = 11
      "0001011" when "01011111110010001", -- t[49041] = 11
      "0001011" when "01011111110010010", -- t[49042] = 11
      "0001011" when "01011111110010011", -- t[49043] = 11
      "0001011" when "01011111110010100", -- t[49044] = 11
      "0001011" when "01011111110010101", -- t[49045] = 11
      "0001011" when "01011111110010110", -- t[49046] = 11
      "0001011" when "01011111110010111", -- t[49047] = 11
      "0001011" when "01011111110011000", -- t[49048] = 11
      "0001011" when "01011111110011001", -- t[49049] = 11
      "0001011" when "01011111110011010", -- t[49050] = 11
      "0001011" when "01011111110011011", -- t[49051] = 11
      "0001011" when "01011111110011100", -- t[49052] = 11
      "0001011" when "01011111110011101", -- t[49053] = 11
      "0001011" when "01011111110011110", -- t[49054] = 11
      "0001011" when "01011111110011111", -- t[49055] = 11
      "0001011" when "01011111110100000", -- t[49056] = 11
      "0001011" when "01011111110100001", -- t[49057] = 11
      "0001011" when "01011111110100010", -- t[49058] = 11
      "0001011" when "01011111110100011", -- t[49059] = 11
      "0001011" when "01011111110100100", -- t[49060] = 11
      "0001011" when "01011111110100101", -- t[49061] = 11
      "0001011" when "01011111110100110", -- t[49062] = 11
      "0001011" when "01011111110100111", -- t[49063] = 11
      "0001011" when "01011111110101000", -- t[49064] = 11
      "0001011" when "01011111110101001", -- t[49065] = 11
      "0001011" when "01011111110101010", -- t[49066] = 11
      "0001011" when "01011111110101011", -- t[49067] = 11
      "0001011" when "01011111110101100", -- t[49068] = 11
      "0001011" when "01011111110101101", -- t[49069] = 11
      "0001011" when "01011111110101110", -- t[49070] = 11
      "0001011" when "01011111110101111", -- t[49071] = 11
      "0001011" when "01011111110110000", -- t[49072] = 11
      "0001011" when "01011111110110001", -- t[49073] = 11
      "0001011" when "01011111110110010", -- t[49074] = 11
      "0001011" when "01011111110110011", -- t[49075] = 11
      "0001011" when "01011111110110100", -- t[49076] = 11
      "0001011" when "01011111110110101", -- t[49077] = 11
      "0001011" when "01011111110110110", -- t[49078] = 11
      "0001011" when "01011111110110111", -- t[49079] = 11
      "0001011" when "01011111110111000", -- t[49080] = 11
      "0001011" when "01011111110111001", -- t[49081] = 11
      "0001011" when "01011111110111010", -- t[49082] = 11
      "0001011" when "01011111110111011", -- t[49083] = 11
      "0001011" when "01011111110111100", -- t[49084] = 11
      "0001011" when "01011111110111101", -- t[49085] = 11
      "0001011" when "01011111110111110", -- t[49086] = 11
      "0001011" when "01011111110111111", -- t[49087] = 11
      "0001011" when "01011111111000000", -- t[49088] = 11
      "0001011" when "01011111111000001", -- t[49089] = 11
      "0001011" when "01011111111000010", -- t[49090] = 11
      "0001011" when "01011111111000011", -- t[49091] = 11
      "0001011" when "01011111111000100", -- t[49092] = 11
      "0001011" when "01011111111000101", -- t[49093] = 11
      "0001011" when "01011111111000110", -- t[49094] = 11
      "0001011" when "01011111111000111", -- t[49095] = 11
      "0001011" when "01011111111001000", -- t[49096] = 11
      "0001011" when "01011111111001001", -- t[49097] = 11
      "0001011" when "01011111111001010", -- t[49098] = 11
      "0001011" when "01011111111001011", -- t[49099] = 11
      "0001011" when "01011111111001100", -- t[49100] = 11
      "0001011" when "01011111111001101", -- t[49101] = 11
      "0001011" when "01011111111001110", -- t[49102] = 11
      "0001011" when "01011111111001111", -- t[49103] = 11
      "0001100" when "01011111111010000", -- t[49104] = 12
      "0001100" when "01011111111010001", -- t[49105] = 12
      "0001100" when "01011111111010010", -- t[49106] = 12
      "0001100" when "01011111111010011", -- t[49107] = 12
      "0001100" when "01011111111010100", -- t[49108] = 12
      "0001100" when "01011111111010101", -- t[49109] = 12
      "0001100" when "01011111111010110", -- t[49110] = 12
      "0001100" when "01011111111010111", -- t[49111] = 12
      "0001100" when "01011111111011000", -- t[49112] = 12
      "0001100" when "01011111111011001", -- t[49113] = 12
      "0001100" when "01011111111011010", -- t[49114] = 12
      "0001100" when "01011111111011011", -- t[49115] = 12
      "0001100" when "01011111111011100", -- t[49116] = 12
      "0001100" when "01011111111011101", -- t[49117] = 12
      "0001100" when "01011111111011110", -- t[49118] = 12
      "0001100" when "01011111111011111", -- t[49119] = 12
      "0001100" when "01011111111100000", -- t[49120] = 12
      "0001100" when "01011111111100001", -- t[49121] = 12
      "0001100" when "01011111111100010", -- t[49122] = 12
      "0001100" when "01011111111100011", -- t[49123] = 12
      "0001100" when "01011111111100100", -- t[49124] = 12
      "0001100" when "01011111111100101", -- t[49125] = 12
      "0001100" when "01011111111100110", -- t[49126] = 12
      "0001100" when "01011111111100111", -- t[49127] = 12
      "0001100" when "01011111111101000", -- t[49128] = 12
      "0001100" when "01011111111101001", -- t[49129] = 12
      "0001100" when "01011111111101010", -- t[49130] = 12
      "0001100" when "01011111111101011", -- t[49131] = 12
      "0001100" when "01011111111101100", -- t[49132] = 12
      "0001100" when "01011111111101101", -- t[49133] = 12
      "0001100" when "01011111111101110", -- t[49134] = 12
      "0001100" when "01011111111101111", -- t[49135] = 12
      "0001100" when "01011111111110000", -- t[49136] = 12
      "0001100" when "01011111111110001", -- t[49137] = 12
      "0001100" when "01011111111110010", -- t[49138] = 12
      "0001100" when "01011111111110011", -- t[49139] = 12
      "0001100" when "01011111111110100", -- t[49140] = 12
      "0001100" when "01011111111110101", -- t[49141] = 12
      "0001100" when "01011111111110110", -- t[49142] = 12
      "0001100" when "01011111111110111", -- t[49143] = 12
      "0001100" when "01011111111111000", -- t[49144] = 12
      "0001100" when "01011111111111001", -- t[49145] = 12
      "0001100" when "01011111111111010", -- t[49146] = 12
      "0001100" when "01011111111111011", -- t[49147] = 12
      "0001100" when "01011111111111100", -- t[49148] = 12
      "0001100" when "01011111111111101", -- t[49149] = 12
      "0001100" when "01011111111111110", -- t[49150] = 12
      "0001100" when "01011111111111111", -- t[49151] = 12
      "0001100" when "01100000000000000", -- t[49152] = 12
      "0001100" when "01100000000000001", -- t[49153] = 12
      "0001100" when "01100000000000010", -- t[49154] = 12
      "0001100" when "01100000000000011", -- t[49155] = 12
      "0001100" when "01100000000000100", -- t[49156] = 12
      "0001100" when "01100000000000101", -- t[49157] = 12
      "0001100" when "01100000000000110", -- t[49158] = 12
      "0001100" when "01100000000000111", -- t[49159] = 12
      "0001100" when "01100000000001000", -- t[49160] = 12
      "0001100" when "01100000000001001", -- t[49161] = 12
      "0001100" when "01100000000001010", -- t[49162] = 12
      "0001100" when "01100000000001011", -- t[49163] = 12
      "0001100" when "01100000000001100", -- t[49164] = 12
      "0001100" when "01100000000001101", -- t[49165] = 12
      "0001100" when "01100000000001110", -- t[49166] = 12
      "0001100" when "01100000000001111", -- t[49167] = 12
      "0001100" when "01100000000010000", -- t[49168] = 12
      "0001100" when "01100000000010001", -- t[49169] = 12
      "0001100" when "01100000000010010", -- t[49170] = 12
      "0001100" when "01100000000010011", -- t[49171] = 12
      "0001100" when "01100000000010100", -- t[49172] = 12
      "0001100" when "01100000000010101", -- t[49173] = 12
      "0001100" when "01100000000010110", -- t[49174] = 12
      "0001100" when "01100000000010111", -- t[49175] = 12
      "0001100" when "01100000000011000", -- t[49176] = 12
      "0001100" when "01100000000011001", -- t[49177] = 12
      "0001100" when "01100000000011010", -- t[49178] = 12
      "0001100" when "01100000000011011", -- t[49179] = 12
      "0001100" when "01100000000011100", -- t[49180] = 12
      "0001100" when "01100000000011101", -- t[49181] = 12
      "0001100" when "01100000000011110", -- t[49182] = 12
      "0001100" when "01100000000011111", -- t[49183] = 12
      "0001100" when "01100000000100000", -- t[49184] = 12
      "0001100" when "01100000000100001", -- t[49185] = 12
      "0001100" when "01100000000100010", -- t[49186] = 12
      "0001100" when "01100000000100011", -- t[49187] = 12
      "0001100" when "01100000000100100", -- t[49188] = 12
      "0001100" when "01100000000100101", -- t[49189] = 12
      "0001100" when "01100000000100110", -- t[49190] = 12
      "0001100" when "01100000000100111", -- t[49191] = 12
      "0001100" when "01100000000101000", -- t[49192] = 12
      "0001100" when "01100000000101001", -- t[49193] = 12
      "0001100" when "01100000000101010", -- t[49194] = 12
      "0001100" when "01100000000101011", -- t[49195] = 12
      "0001100" when "01100000000101100", -- t[49196] = 12
      "0001100" when "01100000000101101", -- t[49197] = 12
      "0001100" when "01100000000101110", -- t[49198] = 12
      "0001100" when "01100000000101111", -- t[49199] = 12
      "0001100" when "01100000000110000", -- t[49200] = 12
      "0001100" when "01100000000110001", -- t[49201] = 12
      "0001100" when "01100000000110010", -- t[49202] = 12
      "0001100" when "01100000000110011", -- t[49203] = 12
      "0001100" when "01100000000110100", -- t[49204] = 12
      "0001100" when "01100000000110101", -- t[49205] = 12
      "0001100" when "01100000000110110", -- t[49206] = 12
      "0001100" when "01100000000110111", -- t[49207] = 12
      "0001100" when "01100000000111000", -- t[49208] = 12
      "0001100" when "01100000000111001", -- t[49209] = 12
      "0001100" when "01100000000111010", -- t[49210] = 12
      "0001100" when "01100000000111011", -- t[49211] = 12
      "0001100" when "01100000000111100", -- t[49212] = 12
      "0001100" when "01100000000111101", -- t[49213] = 12
      "0001100" when "01100000000111110", -- t[49214] = 12
      "0001100" when "01100000000111111", -- t[49215] = 12
      "0001100" when "01100000001000000", -- t[49216] = 12
      "0001100" when "01100000001000001", -- t[49217] = 12
      "0001100" when "01100000001000010", -- t[49218] = 12
      "0001100" when "01100000001000011", -- t[49219] = 12
      "0001100" when "01100000001000100", -- t[49220] = 12
      "0001100" when "01100000001000101", -- t[49221] = 12
      "0001100" when "01100000001000110", -- t[49222] = 12
      "0001100" when "01100000001000111", -- t[49223] = 12
      "0001100" when "01100000001001000", -- t[49224] = 12
      "0001100" when "01100000001001001", -- t[49225] = 12
      "0001100" when "01100000001001010", -- t[49226] = 12
      "0001100" when "01100000001001011", -- t[49227] = 12
      "0001100" when "01100000001001100", -- t[49228] = 12
      "0001100" when "01100000001001101", -- t[49229] = 12
      "0001100" when "01100000001001110", -- t[49230] = 12
      "0001100" when "01100000001001111", -- t[49231] = 12
      "0001100" when "01100000001010000", -- t[49232] = 12
      "0001100" when "01100000001010001", -- t[49233] = 12
      "0001100" when "01100000001010010", -- t[49234] = 12
      "0001100" when "01100000001010011", -- t[49235] = 12
      "0001100" when "01100000001010100", -- t[49236] = 12
      "0001100" when "01100000001010101", -- t[49237] = 12
      "0001100" when "01100000001010110", -- t[49238] = 12
      "0001100" when "01100000001010111", -- t[49239] = 12
      "0001100" when "01100000001011000", -- t[49240] = 12
      "0001100" when "01100000001011001", -- t[49241] = 12
      "0001100" when "01100000001011010", -- t[49242] = 12
      "0001100" when "01100000001011011", -- t[49243] = 12
      "0001100" when "01100000001011100", -- t[49244] = 12
      "0001100" when "01100000001011101", -- t[49245] = 12
      "0001100" when "01100000001011110", -- t[49246] = 12
      "0001100" when "01100000001011111", -- t[49247] = 12
      "0001100" when "01100000001100000", -- t[49248] = 12
      "0001100" when "01100000001100001", -- t[49249] = 12
      "0001100" when "01100000001100010", -- t[49250] = 12
      "0001100" when "01100000001100011", -- t[49251] = 12
      "0001100" when "01100000001100100", -- t[49252] = 12
      "0001100" when "01100000001100101", -- t[49253] = 12
      "0001100" when "01100000001100110", -- t[49254] = 12
      "0001100" when "01100000001100111", -- t[49255] = 12
      "0001100" when "01100000001101000", -- t[49256] = 12
      "0001100" when "01100000001101001", -- t[49257] = 12
      "0001100" when "01100000001101010", -- t[49258] = 12
      "0001100" when "01100000001101011", -- t[49259] = 12
      "0001100" when "01100000001101100", -- t[49260] = 12
      "0001100" when "01100000001101101", -- t[49261] = 12
      "0001100" when "01100000001101110", -- t[49262] = 12
      "0001100" when "01100000001101111", -- t[49263] = 12
      "0001100" when "01100000001110000", -- t[49264] = 12
      "0001100" when "01100000001110001", -- t[49265] = 12
      "0001100" when "01100000001110010", -- t[49266] = 12
      "0001100" when "01100000001110011", -- t[49267] = 12
      "0001100" when "01100000001110100", -- t[49268] = 12
      "0001100" when "01100000001110101", -- t[49269] = 12
      "0001100" when "01100000001110110", -- t[49270] = 12
      "0001100" when "01100000001110111", -- t[49271] = 12
      "0001100" when "01100000001111000", -- t[49272] = 12
      "0001100" when "01100000001111001", -- t[49273] = 12
      "0001100" when "01100000001111010", -- t[49274] = 12
      "0001100" when "01100000001111011", -- t[49275] = 12
      "0001100" when "01100000001111100", -- t[49276] = 12
      "0001100" when "01100000001111101", -- t[49277] = 12
      "0001100" when "01100000001111110", -- t[49278] = 12
      "0001100" when "01100000001111111", -- t[49279] = 12
      "0001100" when "01100000010000000", -- t[49280] = 12
      "0001100" when "01100000010000001", -- t[49281] = 12
      "0001100" when "01100000010000010", -- t[49282] = 12
      "0001100" when "01100000010000011", -- t[49283] = 12
      "0001100" when "01100000010000100", -- t[49284] = 12
      "0001100" when "01100000010000101", -- t[49285] = 12
      "0001100" when "01100000010000110", -- t[49286] = 12
      "0001100" when "01100000010000111", -- t[49287] = 12
      "0001100" when "01100000010001000", -- t[49288] = 12
      "0001100" when "01100000010001001", -- t[49289] = 12
      "0001100" when "01100000010001010", -- t[49290] = 12
      "0001100" when "01100000010001011", -- t[49291] = 12
      "0001100" when "01100000010001100", -- t[49292] = 12
      "0001100" when "01100000010001101", -- t[49293] = 12
      "0001100" when "01100000010001110", -- t[49294] = 12
      "0001100" when "01100000010001111", -- t[49295] = 12
      "0001100" when "01100000010010000", -- t[49296] = 12
      "0001100" when "01100000010010001", -- t[49297] = 12
      "0001100" when "01100000010010010", -- t[49298] = 12
      "0001100" when "01100000010010011", -- t[49299] = 12
      "0001100" when "01100000010010100", -- t[49300] = 12
      "0001100" when "01100000010010101", -- t[49301] = 12
      "0001100" when "01100000010010110", -- t[49302] = 12
      "0001100" when "01100000010010111", -- t[49303] = 12
      "0001100" when "01100000010011000", -- t[49304] = 12
      "0001100" when "01100000010011001", -- t[49305] = 12
      "0001100" when "01100000010011010", -- t[49306] = 12
      "0001100" when "01100000010011011", -- t[49307] = 12
      "0001100" when "01100000010011100", -- t[49308] = 12
      "0001100" when "01100000010011101", -- t[49309] = 12
      "0001100" when "01100000010011110", -- t[49310] = 12
      "0001100" when "01100000010011111", -- t[49311] = 12
      "0001100" when "01100000010100000", -- t[49312] = 12
      "0001100" when "01100000010100001", -- t[49313] = 12
      "0001100" when "01100000010100010", -- t[49314] = 12
      "0001100" when "01100000010100011", -- t[49315] = 12
      "0001100" when "01100000010100100", -- t[49316] = 12
      "0001100" when "01100000010100101", -- t[49317] = 12
      "0001100" when "01100000010100110", -- t[49318] = 12
      "0001100" when "01100000010100111", -- t[49319] = 12
      "0001100" when "01100000010101000", -- t[49320] = 12
      "0001100" when "01100000010101001", -- t[49321] = 12
      "0001100" when "01100000010101010", -- t[49322] = 12
      "0001100" when "01100000010101011", -- t[49323] = 12
      "0001100" when "01100000010101100", -- t[49324] = 12
      "0001100" when "01100000010101101", -- t[49325] = 12
      "0001100" when "01100000010101110", -- t[49326] = 12
      "0001100" when "01100000010101111", -- t[49327] = 12
      "0001100" when "01100000010110000", -- t[49328] = 12
      "0001100" when "01100000010110001", -- t[49329] = 12
      "0001100" when "01100000010110010", -- t[49330] = 12
      "0001100" when "01100000010110011", -- t[49331] = 12
      "0001100" when "01100000010110100", -- t[49332] = 12
      "0001100" when "01100000010110101", -- t[49333] = 12
      "0001100" when "01100000010110110", -- t[49334] = 12
      "0001100" when "01100000010110111", -- t[49335] = 12
      "0001100" when "01100000010111000", -- t[49336] = 12
      "0001100" when "01100000010111001", -- t[49337] = 12
      "0001100" when "01100000010111010", -- t[49338] = 12
      "0001100" when "01100000010111011", -- t[49339] = 12
      "0001100" when "01100000010111100", -- t[49340] = 12
      "0001100" when "01100000010111101", -- t[49341] = 12
      "0001100" when "01100000010111110", -- t[49342] = 12
      "0001100" when "01100000010111111", -- t[49343] = 12
      "0001100" when "01100000011000000", -- t[49344] = 12
      "0001100" when "01100000011000001", -- t[49345] = 12
      "0001100" when "01100000011000010", -- t[49346] = 12
      "0001100" when "01100000011000011", -- t[49347] = 12
      "0001100" when "01100000011000100", -- t[49348] = 12
      "0001100" when "01100000011000101", -- t[49349] = 12
      "0001100" when "01100000011000110", -- t[49350] = 12
      "0001100" when "01100000011000111", -- t[49351] = 12
      "0001100" when "01100000011001000", -- t[49352] = 12
      "0001100" when "01100000011001001", -- t[49353] = 12
      "0001100" when "01100000011001010", -- t[49354] = 12
      "0001100" when "01100000011001011", -- t[49355] = 12
      "0001100" when "01100000011001100", -- t[49356] = 12
      "0001100" when "01100000011001101", -- t[49357] = 12
      "0001100" when "01100000011001110", -- t[49358] = 12
      "0001100" when "01100000011001111", -- t[49359] = 12
      "0001100" when "01100000011010000", -- t[49360] = 12
      "0001100" when "01100000011010001", -- t[49361] = 12
      "0001100" when "01100000011010010", -- t[49362] = 12
      "0001100" when "01100000011010011", -- t[49363] = 12
      "0001100" when "01100000011010100", -- t[49364] = 12
      "0001100" when "01100000011010101", -- t[49365] = 12
      "0001100" when "01100000011010110", -- t[49366] = 12
      "0001100" when "01100000011010111", -- t[49367] = 12
      "0001100" when "01100000011011000", -- t[49368] = 12
      "0001100" when "01100000011011001", -- t[49369] = 12
      "0001100" when "01100000011011010", -- t[49370] = 12
      "0001100" when "01100000011011011", -- t[49371] = 12
      "0001100" when "01100000011011100", -- t[49372] = 12
      "0001100" when "01100000011011101", -- t[49373] = 12
      "0001100" when "01100000011011110", -- t[49374] = 12
      "0001100" when "01100000011011111", -- t[49375] = 12
      "0001100" when "01100000011100000", -- t[49376] = 12
      "0001100" when "01100000011100001", -- t[49377] = 12
      "0001100" when "01100000011100010", -- t[49378] = 12
      "0001100" when "01100000011100011", -- t[49379] = 12
      "0001100" when "01100000011100100", -- t[49380] = 12
      "0001100" when "01100000011100101", -- t[49381] = 12
      "0001100" when "01100000011100110", -- t[49382] = 12
      "0001100" when "01100000011100111", -- t[49383] = 12
      "0001100" when "01100000011101000", -- t[49384] = 12
      "0001100" when "01100000011101001", -- t[49385] = 12
      "0001100" when "01100000011101010", -- t[49386] = 12
      "0001100" when "01100000011101011", -- t[49387] = 12
      "0001100" when "01100000011101100", -- t[49388] = 12
      "0001100" when "01100000011101101", -- t[49389] = 12
      "0001100" when "01100000011101110", -- t[49390] = 12
      "0001100" when "01100000011101111", -- t[49391] = 12
      "0001100" when "01100000011110000", -- t[49392] = 12
      "0001100" when "01100000011110001", -- t[49393] = 12
      "0001100" when "01100000011110010", -- t[49394] = 12
      "0001100" when "01100000011110011", -- t[49395] = 12
      "0001100" when "01100000011110100", -- t[49396] = 12
      "0001100" when "01100000011110101", -- t[49397] = 12
      "0001100" when "01100000011110110", -- t[49398] = 12
      "0001100" when "01100000011110111", -- t[49399] = 12
      "0001100" when "01100000011111000", -- t[49400] = 12
      "0001100" when "01100000011111001", -- t[49401] = 12
      "0001100" when "01100000011111010", -- t[49402] = 12
      "0001100" when "01100000011111011", -- t[49403] = 12
      "0001100" when "01100000011111100", -- t[49404] = 12
      "0001100" when "01100000011111101", -- t[49405] = 12
      "0001100" when "01100000011111110", -- t[49406] = 12
      "0001100" when "01100000011111111", -- t[49407] = 12
      "0001100" when "01100000100000000", -- t[49408] = 12
      "0001100" when "01100000100000001", -- t[49409] = 12
      "0001100" when "01100000100000010", -- t[49410] = 12
      "0001100" when "01100000100000011", -- t[49411] = 12
      "0001100" when "01100000100000100", -- t[49412] = 12
      "0001100" when "01100000100000101", -- t[49413] = 12
      "0001100" when "01100000100000110", -- t[49414] = 12
      "0001100" when "01100000100000111", -- t[49415] = 12
      "0001100" when "01100000100001000", -- t[49416] = 12
      "0001100" when "01100000100001001", -- t[49417] = 12
      "0001100" when "01100000100001010", -- t[49418] = 12
      "0001100" when "01100000100001011", -- t[49419] = 12
      "0001100" when "01100000100001100", -- t[49420] = 12
      "0001100" when "01100000100001101", -- t[49421] = 12
      "0001100" when "01100000100001110", -- t[49422] = 12
      "0001100" when "01100000100001111", -- t[49423] = 12
      "0001100" when "01100000100010000", -- t[49424] = 12
      "0001100" when "01100000100010001", -- t[49425] = 12
      "0001100" when "01100000100010010", -- t[49426] = 12
      "0001100" when "01100000100010011", -- t[49427] = 12
      "0001100" when "01100000100010100", -- t[49428] = 12
      "0001100" when "01100000100010101", -- t[49429] = 12
      "0001100" when "01100000100010110", -- t[49430] = 12
      "0001100" when "01100000100010111", -- t[49431] = 12
      "0001100" when "01100000100011000", -- t[49432] = 12
      "0001100" when "01100000100011001", -- t[49433] = 12
      "0001100" when "01100000100011010", -- t[49434] = 12
      "0001100" when "01100000100011011", -- t[49435] = 12
      "0001100" when "01100000100011100", -- t[49436] = 12
      "0001100" when "01100000100011101", -- t[49437] = 12
      "0001100" when "01100000100011110", -- t[49438] = 12
      "0001100" when "01100000100011111", -- t[49439] = 12
      "0001100" when "01100000100100000", -- t[49440] = 12
      "0001100" when "01100000100100001", -- t[49441] = 12
      "0001100" when "01100000100100010", -- t[49442] = 12
      "0001100" when "01100000100100011", -- t[49443] = 12
      "0001100" when "01100000100100100", -- t[49444] = 12
      "0001100" when "01100000100100101", -- t[49445] = 12
      "0001100" when "01100000100100110", -- t[49446] = 12
      "0001100" when "01100000100100111", -- t[49447] = 12
      "0001100" when "01100000100101000", -- t[49448] = 12
      "0001100" when "01100000100101001", -- t[49449] = 12
      "0001100" when "01100000100101010", -- t[49450] = 12
      "0001100" when "01100000100101011", -- t[49451] = 12
      "0001100" when "01100000100101100", -- t[49452] = 12
      "0001100" when "01100000100101101", -- t[49453] = 12
      "0001100" when "01100000100101110", -- t[49454] = 12
      "0001100" when "01100000100101111", -- t[49455] = 12
      "0001100" when "01100000100110000", -- t[49456] = 12
      "0001100" when "01100000100110001", -- t[49457] = 12
      "0001100" when "01100000100110010", -- t[49458] = 12
      "0001100" when "01100000100110011", -- t[49459] = 12
      "0001100" when "01100000100110100", -- t[49460] = 12
      "0001100" when "01100000100110101", -- t[49461] = 12
      "0001100" when "01100000100110110", -- t[49462] = 12
      "0001100" when "01100000100110111", -- t[49463] = 12
      "0001100" when "01100000100111000", -- t[49464] = 12
      "0001100" when "01100000100111001", -- t[49465] = 12
      "0001100" when "01100000100111010", -- t[49466] = 12
      "0001100" when "01100000100111011", -- t[49467] = 12
      "0001100" when "01100000100111100", -- t[49468] = 12
      "0001100" when "01100000100111101", -- t[49469] = 12
      "0001100" when "01100000100111110", -- t[49470] = 12
      "0001100" when "01100000100111111", -- t[49471] = 12
      "0001100" when "01100000101000000", -- t[49472] = 12
      "0001100" when "01100000101000001", -- t[49473] = 12
      "0001100" when "01100000101000010", -- t[49474] = 12
      "0001100" when "01100000101000011", -- t[49475] = 12
      "0001100" when "01100000101000100", -- t[49476] = 12
      "0001100" when "01100000101000101", -- t[49477] = 12
      "0001100" when "01100000101000110", -- t[49478] = 12
      "0001100" when "01100000101000111", -- t[49479] = 12
      "0001100" when "01100000101001000", -- t[49480] = 12
      "0001100" when "01100000101001001", -- t[49481] = 12
      "0001100" when "01100000101001010", -- t[49482] = 12
      "0001100" when "01100000101001011", -- t[49483] = 12
      "0001100" when "01100000101001100", -- t[49484] = 12
      "0001100" when "01100000101001101", -- t[49485] = 12
      "0001100" when "01100000101001110", -- t[49486] = 12
      "0001100" when "01100000101001111", -- t[49487] = 12
      "0001100" when "01100000101010000", -- t[49488] = 12
      "0001100" when "01100000101010001", -- t[49489] = 12
      "0001100" when "01100000101010010", -- t[49490] = 12
      "0001100" when "01100000101010011", -- t[49491] = 12
      "0001100" when "01100000101010100", -- t[49492] = 12
      "0001100" when "01100000101010101", -- t[49493] = 12
      "0001100" when "01100000101010110", -- t[49494] = 12
      "0001100" when "01100000101010111", -- t[49495] = 12
      "0001100" when "01100000101011000", -- t[49496] = 12
      "0001100" when "01100000101011001", -- t[49497] = 12
      "0001100" when "01100000101011010", -- t[49498] = 12
      "0001100" when "01100000101011011", -- t[49499] = 12
      "0001100" when "01100000101011100", -- t[49500] = 12
      "0001100" when "01100000101011101", -- t[49501] = 12
      "0001100" when "01100000101011110", -- t[49502] = 12
      "0001100" when "01100000101011111", -- t[49503] = 12
      "0001100" when "01100000101100000", -- t[49504] = 12
      "0001100" when "01100000101100001", -- t[49505] = 12
      "0001100" when "01100000101100010", -- t[49506] = 12
      "0001100" when "01100000101100011", -- t[49507] = 12
      "0001100" when "01100000101100100", -- t[49508] = 12
      "0001100" when "01100000101100101", -- t[49509] = 12
      "0001100" when "01100000101100110", -- t[49510] = 12
      "0001100" when "01100000101100111", -- t[49511] = 12
      "0001100" when "01100000101101000", -- t[49512] = 12
      "0001100" when "01100000101101001", -- t[49513] = 12
      "0001100" when "01100000101101010", -- t[49514] = 12
      "0001100" when "01100000101101011", -- t[49515] = 12
      "0001100" when "01100000101101100", -- t[49516] = 12
      "0001100" when "01100000101101101", -- t[49517] = 12
      "0001100" when "01100000101101110", -- t[49518] = 12
      "0001100" when "01100000101101111", -- t[49519] = 12
      "0001100" when "01100000101110000", -- t[49520] = 12
      "0001100" when "01100000101110001", -- t[49521] = 12
      "0001100" when "01100000101110010", -- t[49522] = 12
      "0001100" when "01100000101110011", -- t[49523] = 12
      "0001100" when "01100000101110100", -- t[49524] = 12
      "0001100" when "01100000101110101", -- t[49525] = 12
      "0001100" when "01100000101110110", -- t[49526] = 12
      "0001100" when "01100000101110111", -- t[49527] = 12
      "0001100" when "01100000101111000", -- t[49528] = 12
      "0001100" when "01100000101111001", -- t[49529] = 12
      "0001100" when "01100000101111010", -- t[49530] = 12
      "0001100" when "01100000101111011", -- t[49531] = 12
      "0001100" when "01100000101111100", -- t[49532] = 12
      "0001100" when "01100000101111101", -- t[49533] = 12
      "0001100" when "01100000101111110", -- t[49534] = 12
      "0001100" when "01100000101111111", -- t[49535] = 12
      "0001100" when "01100000110000000", -- t[49536] = 12
      "0001100" when "01100000110000001", -- t[49537] = 12
      "0001100" when "01100000110000010", -- t[49538] = 12
      "0001100" when "01100000110000011", -- t[49539] = 12
      "0001100" when "01100000110000100", -- t[49540] = 12
      "0001100" when "01100000110000101", -- t[49541] = 12
      "0001100" when "01100000110000110", -- t[49542] = 12
      "0001100" when "01100000110000111", -- t[49543] = 12
      "0001100" when "01100000110001000", -- t[49544] = 12
      "0001100" when "01100000110001001", -- t[49545] = 12
      "0001100" when "01100000110001010", -- t[49546] = 12
      "0001100" when "01100000110001011", -- t[49547] = 12
      "0001100" when "01100000110001100", -- t[49548] = 12
      "0001100" when "01100000110001101", -- t[49549] = 12
      "0001100" when "01100000110001110", -- t[49550] = 12
      "0001100" when "01100000110001111", -- t[49551] = 12
      "0001100" when "01100000110010000", -- t[49552] = 12
      "0001100" when "01100000110010001", -- t[49553] = 12
      "0001100" when "01100000110010010", -- t[49554] = 12
      "0001100" when "01100000110010011", -- t[49555] = 12
      "0001100" when "01100000110010100", -- t[49556] = 12
      "0001100" when "01100000110010101", -- t[49557] = 12
      "0001100" when "01100000110010110", -- t[49558] = 12
      "0001100" when "01100000110010111", -- t[49559] = 12
      "0001100" when "01100000110011000", -- t[49560] = 12
      "0001100" when "01100000110011001", -- t[49561] = 12
      "0001100" when "01100000110011010", -- t[49562] = 12
      "0001100" when "01100000110011011", -- t[49563] = 12
      "0001100" when "01100000110011100", -- t[49564] = 12
      "0001100" when "01100000110011101", -- t[49565] = 12
      "0001100" when "01100000110011110", -- t[49566] = 12
      "0001100" when "01100000110011111", -- t[49567] = 12
      "0001100" when "01100000110100000", -- t[49568] = 12
      "0001100" when "01100000110100001", -- t[49569] = 12
      "0001100" when "01100000110100010", -- t[49570] = 12
      "0001100" when "01100000110100011", -- t[49571] = 12
      "0001100" when "01100000110100100", -- t[49572] = 12
      "0001100" when "01100000110100101", -- t[49573] = 12
      "0001100" when "01100000110100110", -- t[49574] = 12
      "0001100" when "01100000110100111", -- t[49575] = 12
      "0001100" when "01100000110101000", -- t[49576] = 12
      "0001100" when "01100000110101001", -- t[49577] = 12
      "0001100" when "01100000110101010", -- t[49578] = 12
      "0001100" when "01100000110101011", -- t[49579] = 12
      "0001100" when "01100000110101100", -- t[49580] = 12
      "0001100" when "01100000110101101", -- t[49581] = 12
      "0001100" when "01100000110101110", -- t[49582] = 12
      "0001100" when "01100000110101111", -- t[49583] = 12
      "0001100" when "01100000110110000", -- t[49584] = 12
      "0001100" when "01100000110110001", -- t[49585] = 12
      "0001100" when "01100000110110010", -- t[49586] = 12
      "0001100" when "01100000110110011", -- t[49587] = 12
      "0001100" when "01100000110110100", -- t[49588] = 12
      "0001100" when "01100000110110101", -- t[49589] = 12
      "0001100" when "01100000110110110", -- t[49590] = 12
      "0001100" when "01100000110110111", -- t[49591] = 12
      "0001100" when "01100000110111000", -- t[49592] = 12
      "0001100" when "01100000110111001", -- t[49593] = 12
      "0001100" when "01100000110111010", -- t[49594] = 12
      "0001100" when "01100000110111011", -- t[49595] = 12
      "0001100" when "01100000110111100", -- t[49596] = 12
      "0001100" when "01100000110111101", -- t[49597] = 12
      "0001100" when "01100000110111110", -- t[49598] = 12
      "0001100" when "01100000110111111", -- t[49599] = 12
      "0001100" when "01100000111000000", -- t[49600] = 12
      "0001100" when "01100000111000001", -- t[49601] = 12
      "0001100" when "01100000111000010", -- t[49602] = 12
      "0001100" when "01100000111000011", -- t[49603] = 12
      "0001100" when "01100000111000100", -- t[49604] = 12
      "0001100" when "01100000111000101", -- t[49605] = 12
      "0001100" when "01100000111000110", -- t[49606] = 12
      "0001100" when "01100000111000111", -- t[49607] = 12
      "0001100" when "01100000111001000", -- t[49608] = 12
      "0001100" when "01100000111001001", -- t[49609] = 12
      "0001100" when "01100000111001010", -- t[49610] = 12
      "0001100" when "01100000111001011", -- t[49611] = 12
      "0001100" when "01100000111001100", -- t[49612] = 12
      "0001100" when "01100000111001101", -- t[49613] = 12
      "0001100" when "01100000111001110", -- t[49614] = 12
      "0001100" when "01100000111001111", -- t[49615] = 12
      "0001100" when "01100000111010000", -- t[49616] = 12
      "0001100" when "01100000111010001", -- t[49617] = 12
      "0001100" when "01100000111010010", -- t[49618] = 12
      "0001100" when "01100000111010011", -- t[49619] = 12
      "0001100" when "01100000111010100", -- t[49620] = 12
      "0001100" when "01100000111010101", -- t[49621] = 12
      "0001100" when "01100000111010110", -- t[49622] = 12
      "0001100" when "01100000111010111", -- t[49623] = 12
      "0001100" when "01100000111011000", -- t[49624] = 12
      "0001100" when "01100000111011001", -- t[49625] = 12
      "0001100" when "01100000111011010", -- t[49626] = 12
      "0001100" when "01100000111011011", -- t[49627] = 12
      "0001100" when "01100000111011100", -- t[49628] = 12
      "0001100" when "01100000111011101", -- t[49629] = 12
      "0001100" when "01100000111011110", -- t[49630] = 12
      "0001100" when "01100000111011111", -- t[49631] = 12
      "0001100" when "01100000111100000", -- t[49632] = 12
      "0001100" when "01100000111100001", -- t[49633] = 12
      "0001100" when "01100000111100010", -- t[49634] = 12
      "0001100" when "01100000111100011", -- t[49635] = 12
      "0001100" when "01100000111100100", -- t[49636] = 12
      "0001100" when "01100000111100101", -- t[49637] = 12
      "0001100" when "01100000111100110", -- t[49638] = 12
      "0001100" when "01100000111100111", -- t[49639] = 12
      "0001100" when "01100000111101000", -- t[49640] = 12
      "0001100" when "01100000111101001", -- t[49641] = 12
      "0001100" when "01100000111101010", -- t[49642] = 12
      "0001100" when "01100000111101011", -- t[49643] = 12
      "0001100" when "01100000111101100", -- t[49644] = 12
      "0001100" when "01100000111101101", -- t[49645] = 12
      "0001100" when "01100000111101110", -- t[49646] = 12
      "0001100" when "01100000111101111", -- t[49647] = 12
      "0001100" when "01100000111110000", -- t[49648] = 12
      "0001100" when "01100000111110001", -- t[49649] = 12
      "0001100" when "01100000111110010", -- t[49650] = 12
      "0001100" when "01100000111110011", -- t[49651] = 12
      "0001100" when "01100000111110100", -- t[49652] = 12
      "0001100" when "01100000111110101", -- t[49653] = 12
      "0001100" when "01100000111110110", -- t[49654] = 12
      "0001100" when "01100000111110111", -- t[49655] = 12
      "0001100" when "01100000111111000", -- t[49656] = 12
      "0001100" when "01100000111111001", -- t[49657] = 12
      "0001100" when "01100000111111010", -- t[49658] = 12
      "0001100" when "01100000111111011", -- t[49659] = 12
      "0001100" when "01100000111111100", -- t[49660] = 12
      "0001100" when "01100000111111101", -- t[49661] = 12
      "0001100" when "01100000111111110", -- t[49662] = 12
      "0001100" when "01100000111111111", -- t[49663] = 12
      "0001100" when "01100001000000000", -- t[49664] = 12
      "0001100" when "01100001000000001", -- t[49665] = 12
      "0001100" when "01100001000000010", -- t[49666] = 12
      "0001100" when "01100001000000011", -- t[49667] = 12
      "0001100" when "01100001000000100", -- t[49668] = 12
      "0001100" when "01100001000000101", -- t[49669] = 12
      "0001100" when "01100001000000110", -- t[49670] = 12
      "0001100" when "01100001000000111", -- t[49671] = 12
      "0001100" when "01100001000001000", -- t[49672] = 12
      "0001100" when "01100001000001001", -- t[49673] = 12
      "0001100" when "01100001000001010", -- t[49674] = 12
      "0001100" when "01100001000001011", -- t[49675] = 12
      "0001100" when "01100001000001100", -- t[49676] = 12
      "0001100" when "01100001000001101", -- t[49677] = 12
      "0001100" when "01100001000001110", -- t[49678] = 12
      "0001100" when "01100001000001111", -- t[49679] = 12
      "0001100" when "01100001000010000", -- t[49680] = 12
      "0001100" when "01100001000010001", -- t[49681] = 12
      "0001100" when "01100001000010010", -- t[49682] = 12
      "0001100" when "01100001000010011", -- t[49683] = 12
      "0001100" when "01100001000010100", -- t[49684] = 12
      "0001100" when "01100001000010101", -- t[49685] = 12
      "0001100" when "01100001000010110", -- t[49686] = 12
      "0001100" when "01100001000010111", -- t[49687] = 12
      "0001100" when "01100001000011000", -- t[49688] = 12
      "0001100" when "01100001000011001", -- t[49689] = 12
      "0001100" when "01100001000011010", -- t[49690] = 12
      "0001100" when "01100001000011011", -- t[49691] = 12
      "0001100" when "01100001000011100", -- t[49692] = 12
      "0001100" when "01100001000011101", -- t[49693] = 12
      "0001100" when "01100001000011110", -- t[49694] = 12
      "0001100" when "01100001000011111", -- t[49695] = 12
      "0001100" when "01100001000100000", -- t[49696] = 12
      "0001100" when "01100001000100001", -- t[49697] = 12
      "0001100" when "01100001000100010", -- t[49698] = 12
      "0001100" when "01100001000100011", -- t[49699] = 12
      "0001100" when "01100001000100100", -- t[49700] = 12
      "0001100" when "01100001000100101", -- t[49701] = 12
      "0001100" when "01100001000100110", -- t[49702] = 12
      "0001100" when "01100001000100111", -- t[49703] = 12
      "0001100" when "01100001000101000", -- t[49704] = 12
      "0001100" when "01100001000101001", -- t[49705] = 12
      "0001100" when "01100001000101010", -- t[49706] = 12
      "0001100" when "01100001000101011", -- t[49707] = 12
      "0001100" when "01100001000101100", -- t[49708] = 12
      "0001100" when "01100001000101101", -- t[49709] = 12
      "0001100" when "01100001000101110", -- t[49710] = 12
      "0001100" when "01100001000101111", -- t[49711] = 12
      "0001100" when "01100001000110000", -- t[49712] = 12
      "0001100" when "01100001000110001", -- t[49713] = 12
      "0001100" when "01100001000110010", -- t[49714] = 12
      "0001100" when "01100001000110011", -- t[49715] = 12
      "0001100" when "01100001000110100", -- t[49716] = 12
      "0001100" when "01100001000110101", -- t[49717] = 12
      "0001100" when "01100001000110110", -- t[49718] = 12
      "0001100" when "01100001000110111", -- t[49719] = 12
      "0001100" when "01100001000111000", -- t[49720] = 12
      "0001100" when "01100001000111001", -- t[49721] = 12
      "0001100" when "01100001000111010", -- t[49722] = 12
      "0001100" when "01100001000111011", -- t[49723] = 12
      "0001100" when "01100001000111100", -- t[49724] = 12
      "0001100" when "01100001000111101", -- t[49725] = 12
      "0001100" when "01100001000111110", -- t[49726] = 12
      "0001100" when "01100001000111111", -- t[49727] = 12
      "0001100" when "01100001001000000", -- t[49728] = 12
      "0001100" when "01100001001000001", -- t[49729] = 12
      "0001100" when "01100001001000010", -- t[49730] = 12
      "0001100" when "01100001001000011", -- t[49731] = 12
      "0001100" when "01100001001000100", -- t[49732] = 12
      "0001100" when "01100001001000101", -- t[49733] = 12
      "0001100" when "01100001001000110", -- t[49734] = 12
      "0001100" when "01100001001000111", -- t[49735] = 12
      "0001100" when "01100001001001000", -- t[49736] = 12
      "0001100" when "01100001001001001", -- t[49737] = 12
      "0001100" when "01100001001001010", -- t[49738] = 12
      "0001100" when "01100001001001011", -- t[49739] = 12
      "0001100" when "01100001001001100", -- t[49740] = 12
      "0001100" when "01100001001001101", -- t[49741] = 12
      "0001100" when "01100001001001110", -- t[49742] = 12
      "0001100" when "01100001001001111", -- t[49743] = 12
      "0001100" when "01100001001010000", -- t[49744] = 12
      "0001100" when "01100001001010001", -- t[49745] = 12
      "0001100" when "01100001001010010", -- t[49746] = 12
      "0001100" when "01100001001010011", -- t[49747] = 12
      "0001100" when "01100001001010100", -- t[49748] = 12
      "0001100" when "01100001001010101", -- t[49749] = 12
      "0001100" when "01100001001010110", -- t[49750] = 12
      "0001100" when "01100001001010111", -- t[49751] = 12
      "0001100" when "01100001001011000", -- t[49752] = 12
      "0001100" when "01100001001011001", -- t[49753] = 12
      "0001100" when "01100001001011010", -- t[49754] = 12
      "0001100" when "01100001001011011", -- t[49755] = 12
      "0001100" when "01100001001011100", -- t[49756] = 12
      "0001100" when "01100001001011101", -- t[49757] = 12
      "0001100" when "01100001001011110", -- t[49758] = 12
      "0001100" when "01100001001011111", -- t[49759] = 12
      "0001100" when "01100001001100000", -- t[49760] = 12
      "0001100" when "01100001001100001", -- t[49761] = 12
      "0001100" when "01100001001100010", -- t[49762] = 12
      "0001100" when "01100001001100011", -- t[49763] = 12
      "0001100" when "01100001001100100", -- t[49764] = 12
      "0001100" when "01100001001100101", -- t[49765] = 12
      "0001100" when "01100001001100110", -- t[49766] = 12
      "0001100" when "01100001001100111", -- t[49767] = 12
      "0001100" when "01100001001101000", -- t[49768] = 12
      "0001100" when "01100001001101001", -- t[49769] = 12
      "0001100" when "01100001001101010", -- t[49770] = 12
      "0001100" when "01100001001101011", -- t[49771] = 12
      "0001100" when "01100001001101100", -- t[49772] = 12
      "0001100" when "01100001001101101", -- t[49773] = 12
      "0001100" when "01100001001101110", -- t[49774] = 12
      "0001100" when "01100001001101111", -- t[49775] = 12
      "0001100" when "01100001001110000", -- t[49776] = 12
      "0001100" when "01100001001110001", -- t[49777] = 12
      "0001100" when "01100001001110010", -- t[49778] = 12
      "0001100" when "01100001001110011", -- t[49779] = 12
      "0001100" when "01100001001110100", -- t[49780] = 12
      "0001100" when "01100001001110101", -- t[49781] = 12
      "0001100" when "01100001001110110", -- t[49782] = 12
      "0001100" when "01100001001110111", -- t[49783] = 12
      "0001100" when "01100001001111000", -- t[49784] = 12
      "0001100" when "01100001001111001", -- t[49785] = 12
      "0001100" when "01100001001111010", -- t[49786] = 12
      "0001100" when "01100001001111011", -- t[49787] = 12
      "0001100" when "01100001001111100", -- t[49788] = 12
      "0001100" when "01100001001111101", -- t[49789] = 12
      "0001100" when "01100001001111110", -- t[49790] = 12
      "0001100" when "01100001001111111", -- t[49791] = 12
      "0001100" when "01100001010000000", -- t[49792] = 12
      "0001100" when "01100001010000001", -- t[49793] = 12
      "0001100" when "01100001010000010", -- t[49794] = 12
      "0001100" when "01100001010000011", -- t[49795] = 12
      "0001100" when "01100001010000100", -- t[49796] = 12
      "0001100" when "01100001010000101", -- t[49797] = 12
      "0001100" when "01100001010000110", -- t[49798] = 12
      "0001100" when "01100001010000111", -- t[49799] = 12
      "0001100" when "01100001010001000", -- t[49800] = 12
      "0001100" when "01100001010001001", -- t[49801] = 12
      "0001100" when "01100001010001010", -- t[49802] = 12
      "0001100" when "01100001010001011", -- t[49803] = 12
      "0001100" when "01100001010001100", -- t[49804] = 12
      "0001100" when "01100001010001101", -- t[49805] = 12
      "0001100" when "01100001010001110", -- t[49806] = 12
      "0001100" when "01100001010001111", -- t[49807] = 12
      "0001100" when "01100001010010000", -- t[49808] = 12
      "0001100" when "01100001010010001", -- t[49809] = 12
      "0001100" when "01100001010010010", -- t[49810] = 12
      "0001100" when "01100001010010011", -- t[49811] = 12
      "0001100" when "01100001010010100", -- t[49812] = 12
      "0001100" when "01100001010010101", -- t[49813] = 12
      "0001100" when "01100001010010110", -- t[49814] = 12
      "0001100" when "01100001010010111", -- t[49815] = 12
      "0001100" when "01100001010011000", -- t[49816] = 12
      "0001100" when "01100001010011001", -- t[49817] = 12
      "0001100" when "01100001010011010", -- t[49818] = 12
      "0001100" when "01100001010011011", -- t[49819] = 12
      "0001100" when "01100001010011100", -- t[49820] = 12
      "0001100" when "01100001010011101", -- t[49821] = 12
      "0001100" when "01100001010011110", -- t[49822] = 12
      "0001100" when "01100001010011111", -- t[49823] = 12
      "0001100" when "01100001010100000", -- t[49824] = 12
      "0001100" when "01100001010100001", -- t[49825] = 12
      "0001100" when "01100001010100010", -- t[49826] = 12
      "0001100" when "01100001010100011", -- t[49827] = 12
      "0001100" when "01100001010100100", -- t[49828] = 12
      "0001100" when "01100001010100101", -- t[49829] = 12
      "0001100" when "01100001010100110", -- t[49830] = 12
      "0001100" when "01100001010100111", -- t[49831] = 12
      "0001100" when "01100001010101000", -- t[49832] = 12
      "0001100" when "01100001010101001", -- t[49833] = 12
      "0001100" when "01100001010101010", -- t[49834] = 12
      "0001100" when "01100001010101011", -- t[49835] = 12
      "0001100" when "01100001010101100", -- t[49836] = 12
      "0001100" when "01100001010101101", -- t[49837] = 12
      "0001100" when "01100001010101110", -- t[49838] = 12
      "0001100" when "01100001010101111", -- t[49839] = 12
      "0001100" when "01100001010110000", -- t[49840] = 12
      "0001100" when "01100001010110001", -- t[49841] = 12
      "0001100" when "01100001010110010", -- t[49842] = 12
      "0001100" when "01100001010110011", -- t[49843] = 12
      "0001100" when "01100001010110100", -- t[49844] = 12
      "0001100" when "01100001010110101", -- t[49845] = 12
      "0001100" when "01100001010110110", -- t[49846] = 12
      "0001100" when "01100001010110111", -- t[49847] = 12
      "0001100" when "01100001010111000", -- t[49848] = 12
      "0001100" when "01100001010111001", -- t[49849] = 12
      "0001100" when "01100001010111010", -- t[49850] = 12
      "0001100" when "01100001010111011", -- t[49851] = 12
      "0001100" when "01100001010111100", -- t[49852] = 12
      "0001100" when "01100001010111101", -- t[49853] = 12
      "0001100" when "01100001010111110", -- t[49854] = 12
      "0001100" when "01100001010111111", -- t[49855] = 12
      "0001100" when "01100001011000000", -- t[49856] = 12
      "0001100" when "01100001011000001", -- t[49857] = 12
      "0001100" when "01100001011000010", -- t[49858] = 12
      "0001100" when "01100001011000011", -- t[49859] = 12
      "0001100" when "01100001011000100", -- t[49860] = 12
      "0001100" when "01100001011000101", -- t[49861] = 12
      "0001100" when "01100001011000110", -- t[49862] = 12
      "0001100" when "01100001011000111", -- t[49863] = 12
      "0001100" when "01100001011001000", -- t[49864] = 12
      "0001100" when "01100001011001001", -- t[49865] = 12
      "0001100" when "01100001011001010", -- t[49866] = 12
      "0001100" when "01100001011001011", -- t[49867] = 12
      "0001100" when "01100001011001100", -- t[49868] = 12
      "0001100" when "01100001011001101", -- t[49869] = 12
      "0001100" when "01100001011001110", -- t[49870] = 12
      "0001100" when "01100001011001111", -- t[49871] = 12
      "0001100" when "01100001011010000", -- t[49872] = 12
      "0001100" when "01100001011010001", -- t[49873] = 12
      "0001100" when "01100001011010010", -- t[49874] = 12
      "0001100" when "01100001011010011", -- t[49875] = 12
      "0001100" when "01100001011010100", -- t[49876] = 12
      "0001100" when "01100001011010101", -- t[49877] = 12
      "0001100" when "01100001011010110", -- t[49878] = 12
      "0001100" when "01100001011010111", -- t[49879] = 12
      "0001100" when "01100001011011000", -- t[49880] = 12
      "0001100" when "01100001011011001", -- t[49881] = 12
      "0001100" when "01100001011011010", -- t[49882] = 12
      "0001100" when "01100001011011011", -- t[49883] = 12
      "0001100" when "01100001011011100", -- t[49884] = 12
      "0001100" when "01100001011011101", -- t[49885] = 12
      "0001100" when "01100001011011110", -- t[49886] = 12
      "0001100" when "01100001011011111", -- t[49887] = 12
      "0001100" when "01100001011100000", -- t[49888] = 12
      "0001100" when "01100001011100001", -- t[49889] = 12
      "0001100" when "01100001011100010", -- t[49890] = 12
      "0001100" when "01100001011100011", -- t[49891] = 12
      "0001100" when "01100001011100100", -- t[49892] = 12
      "0001100" when "01100001011100101", -- t[49893] = 12
      "0001100" when "01100001011100110", -- t[49894] = 12
      "0001100" when "01100001011100111", -- t[49895] = 12
      "0001100" when "01100001011101000", -- t[49896] = 12
      "0001100" when "01100001011101001", -- t[49897] = 12
      "0001100" when "01100001011101010", -- t[49898] = 12
      "0001100" when "01100001011101011", -- t[49899] = 12
      "0001100" when "01100001011101100", -- t[49900] = 12
      "0001100" when "01100001011101101", -- t[49901] = 12
      "0001100" when "01100001011101110", -- t[49902] = 12
      "0001100" when "01100001011101111", -- t[49903] = 12
      "0001100" when "01100001011110000", -- t[49904] = 12
      "0001100" when "01100001011110001", -- t[49905] = 12
      "0001100" when "01100001011110010", -- t[49906] = 12
      "0001100" when "01100001011110011", -- t[49907] = 12
      "0001100" when "01100001011110100", -- t[49908] = 12
      "0001100" when "01100001011110101", -- t[49909] = 12
      "0001100" when "01100001011110110", -- t[49910] = 12
      "0001100" when "01100001011110111", -- t[49911] = 12
      "0001100" when "01100001011111000", -- t[49912] = 12
      "0001100" when "01100001011111001", -- t[49913] = 12
      "0001100" when "01100001011111010", -- t[49914] = 12
      "0001100" when "01100001011111011", -- t[49915] = 12
      "0001100" when "01100001011111100", -- t[49916] = 12
      "0001100" when "01100001011111101", -- t[49917] = 12
      "0001100" when "01100001011111110", -- t[49918] = 12
      "0001100" when "01100001011111111", -- t[49919] = 12
      "0001100" when "01100001100000000", -- t[49920] = 12
      "0001100" when "01100001100000001", -- t[49921] = 12
      "0001100" when "01100001100000010", -- t[49922] = 12
      "0001100" when "01100001100000011", -- t[49923] = 12
      "0001100" when "01100001100000100", -- t[49924] = 12
      "0001100" when "01100001100000101", -- t[49925] = 12
      "0001100" when "01100001100000110", -- t[49926] = 12
      "0001100" when "01100001100000111", -- t[49927] = 12
      "0001100" when "01100001100001000", -- t[49928] = 12
      "0001100" when "01100001100001001", -- t[49929] = 12
      "0001100" when "01100001100001010", -- t[49930] = 12
      "0001100" when "01100001100001011", -- t[49931] = 12
      "0001100" when "01100001100001100", -- t[49932] = 12
      "0001100" when "01100001100001101", -- t[49933] = 12
      "0001100" when "01100001100001110", -- t[49934] = 12
      "0001100" when "01100001100001111", -- t[49935] = 12
      "0001100" when "01100001100010000", -- t[49936] = 12
      "0001100" when "01100001100010001", -- t[49937] = 12
      "0001100" when "01100001100010010", -- t[49938] = 12
      "0001100" when "01100001100010011", -- t[49939] = 12
      "0001100" when "01100001100010100", -- t[49940] = 12
      "0001100" when "01100001100010101", -- t[49941] = 12
      "0001100" when "01100001100010110", -- t[49942] = 12
      "0001100" when "01100001100010111", -- t[49943] = 12
      "0001100" when "01100001100011000", -- t[49944] = 12
      "0001100" when "01100001100011001", -- t[49945] = 12
      "0001100" when "01100001100011010", -- t[49946] = 12
      "0001100" when "01100001100011011", -- t[49947] = 12
      "0001100" when "01100001100011100", -- t[49948] = 12
      "0001100" when "01100001100011101", -- t[49949] = 12
      "0001100" when "01100001100011110", -- t[49950] = 12
      "0001100" when "01100001100011111", -- t[49951] = 12
      "0001100" when "01100001100100000", -- t[49952] = 12
      "0001100" when "01100001100100001", -- t[49953] = 12
      "0001100" when "01100001100100010", -- t[49954] = 12
      "0001100" when "01100001100100011", -- t[49955] = 12
      "0001100" when "01100001100100100", -- t[49956] = 12
      "0001100" when "01100001100100101", -- t[49957] = 12
      "0001100" when "01100001100100110", -- t[49958] = 12
      "0001100" when "01100001100100111", -- t[49959] = 12
      "0001100" when "01100001100101000", -- t[49960] = 12
      "0001100" when "01100001100101001", -- t[49961] = 12
      "0001100" when "01100001100101010", -- t[49962] = 12
      "0001100" when "01100001100101011", -- t[49963] = 12
      "0001100" when "01100001100101100", -- t[49964] = 12
      "0001100" when "01100001100101101", -- t[49965] = 12
      "0001100" when "01100001100101110", -- t[49966] = 12
      "0001100" when "01100001100101111", -- t[49967] = 12
      "0001100" when "01100001100110000", -- t[49968] = 12
      "0001100" when "01100001100110001", -- t[49969] = 12
      "0001100" when "01100001100110010", -- t[49970] = 12
      "0001100" when "01100001100110011", -- t[49971] = 12
      "0001100" when "01100001100110100", -- t[49972] = 12
      "0001100" when "01100001100110101", -- t[49973] = 12
      "0001100" when "01100001100110110", -- t[49974] = 12
      "0001100" when "01100001100110111", -- t[49975] = 12
      "0001100" when "01100001100111000", -- t[49976] = 12
      "0001100" when "01100001100111001", -- t[49977] = 12
      "0001100" when "01100001100111010", -- t[49978] = 12
      "0001100" when "01100001100111011", -- t[49979] = 12
      "0001100" when "01100001100111100", -- t[49980] = 12
      "0001100" when "01100001100111101", -- t[49981] = 12
      "0001100" when "01100001100111110", -- t[49982] = 12
      "0001100" when "01100001100111111", -- t[49983] = 12
      "0001100" when "01100001101000000", -- t[49984] = 12
      "0001100" when "01100001101000001", -- t[49985] = 12
      "0001100" when "01100001101000010", -- t[49986] = 12
      "0001100" when "01100001101000011", -- t[49987] = 12
      "0001100" when "01100001101000100", -- t[49988] = 12
      "0001100" when "01100001101000101", -- t[49989] = 12
      "0001100" when "01100001101000110", -- t[49990] = 12
      "0001100" when "01100001101000111", -- t[49991] = 12
      "0001100" when "01100001101001000", -- t[49992] = 12
      "0001100" when "01100001101001001", -- t[49993] = 12
      "0001100" when "01100001101001010", -- t[49994] = 12
      "0001100" when "01100001101001011", -- t[49995] = 12
      "0001100" when "01100001101001100", -- t[49996] = 12
      "0001100" when "01100001101001101", -- t[49997] = 12
      "0001100" when "01100001101001110", -- t[49998] = 12
      "0001100" when "01100001101001111", -- t[49999] = 12
      "0001100" when "01100001101010000", -- t[50000] = 12
      "0001100" when "01100001101010001", -- t[50001] = 12
      "0001100" when "01100001101010010", -- t[50002] = 12
      "0001100" when "01100001101010011", -- t[50003] = 12
      "0001100" when "01100001101010100", -- t[50004] = 12
      "0001100" when "01100001101010101", -- t[50005] = 12
      "0001100" when "01100001101010110", -- t[50006] = 12
      "0001100" when "01100001101010111", -- t[50007] = 12
      "0001100" when "01100001101011000", -- t[50008] = 12
      "0001100" when "01100001101011001", -- t[50009] = 12
      "0001100" when "01100001101011010", -- t[50010] = 12
      "0001100" when "01100001101011011", -- t[50011] = 12
      "0001100" when "01100001101011100", -- t[50012] = 12
      "0001100" when "01100001101011101", -- t[50013] = 12
      "0001100" when "01100001101011110", -- t[50014] = 12
      "0001100" when "01100001101011111", -- t[50015] = 12
      "0001100" when "01100001101100000", -- t[50016] = 12
      "0001100" when "01100001101100001", -- t[50017] = 12
      "0001100" when "01100001101100010", -- t[50018] = 12
      "0001100" when "01100001101100011", -- t[50019] = 12
      "0001100" when "01100001101100100", -- t[50020] = 12
      "0001100" when "01100001101100101", -- t[50021] = 12
      "0001100" when "01100001101100110", -- t[50022] = 12
      "0001100" when "01100001101100111", -- t[50023] = 12
      "0001100" when "01100001101101000", -- t[50024] = 12
      "0001100" when "01100001101101001", -- t[50025] = 12
      "0001100" when "01100001101101010", -- t[50026] = 12
      "0001100" when "01100001101101011", -- t[50027] = 12
      "0001100" when "01100001101101100", -- t[50028] = 12
      "0001100" when "01100001101101101", -- t[50029] = 12
      "0001100" when "01100001101101110", -- t[50030] = 12
      "0001100" when "01100001101101111", -- t[50031] = 12
      "0001100" when "01100001101110000", -- t[50032] = 12
      "0001100" when "01100001101110001", -- t[50033] = 12
      "0001100" when "01100001101110010", -- t[50034] = 12
      "0001100" when "01100001101110011", -- t[50035] = 12
      "0001100" when "01100001101110100", -- t[50036] = 12
      "0001100" when "01100001101110101", -- t[50037] = 12
      "0001100" when "01100001101110110", -- t[50038] = 12
      "0001100" when "01100001101110111", -- t[50039] = 12
      "0001100" when "01100001101111000", -- t[50040] = 12
      "0001100" when "01100001101111001", -- t[50041] = 12
      "0001100" when "01100001101111010", -- t[50042] = 12
      "0001100" when "01100001101111011", -- t[50043] = 12
      "0001100" when "01100001101111100", -- t[50044] = 12
      "0001100" when "01100001101111101", -- t[50045] = 12
      "0001100" when "01100001101111110", -- t[50046] = 12
      "0001100" when "01100001101111111", -- t[50047] = 12
      "0001100" when "01100001110000000", -- t[50048] = 12
      "0001100" when "01100001110000001", -- t[50049] = 12
      "0001100" when "01100001110000010", -- t[50050] = 12
      "0001100" when "01100001110000011", -- t[50051] = 12
      "0001100" when "01100001110000100", -- t[50052] = 12
      "0001100" when "01100001110000101", -- t[50053] = 12
      "0001100" when "01100001110000110", -- t[50054] = 12
      "0001100" when "01100001110000111", -- t[50055] = 12
      "0001100" when "01100001110001000", -- t[50056] = 12
      "0001100" when "01100001110001001", -- t[50057] = 12
      "0001100" when "01100001110001010", -- t[50058] = 12
      "0001100" when "01100001110001011", -- t[50059] = 12
      "0001100" when "01100001110001100", -- t[50060] = 12
      "0001100" when "01100001110001101", -- t[50061] = 12
      "0001100" when "01100001110001110", -- t[50062] = 12
      "0001100" when "01100001110001111", -- t[50063] = 12
      "0001100" when "01100001110010000", -- t[50064] = 12
      "0001100" when "01100001110010001", -- t[50065] = 12
      "0001100" when "01100001110010010", -- t[50066] = 12
      "0001100" when "01100001110010011", -- t[50067] = 12
      "0001100" when "01100001110010100", -- t[50068] = 12
      "0001100" when "01100001110010101", -- t[50069] = 12
      "0001100" when "01100001110010110", -- t[50070] = 12
      "0001100" when "01100001110010111", -- t[50071] = 12
      "0001100" when "01100001110011000", -- t[50072] = 12
      "0001100" when "01100001110011001", -- t[50073] = 12
      "0001100" when "01100001110011010", -- t[50074] = 12
      "0001100" when "01100001110011011", -- t[50075] = 12
      "0001100" when "01100001110011100", -- t[50076] = 12
      "0001100" when "01100001110011101", -- t[50077] = 12
      "0001100" when "01100001110011110", -- t[50078] = 12
      "0001100" when "01100001110011111", -- t[50079] = 12
      "0001100" when "01100001110100000", -- t[50080] = 12
      "0001100" when "01100001110100001", -- t[50081] = 12
      "0001100" when "01100001110100010", -- t[50082] = 12
      "0001100" when "01100001110100011", -- t[50083] = 12
      "0001100" when "01100001110100100", -- t[50084] = 12
      "0001100" when "01100001110100101", -- t[50085] = 12
      "0001100" when "01100001110100110", -- t[50086] = 12
      "0001100" when "01100001110100111", -- t[50087] = 12
      "0001100" when "01100001110101000", -- t[50088] = 12
      "0001101" when "01100001110101001", -- t[50089] = 13
      "0001101" when "01100001110101010", -- t[50090] = 13
      "0001101" when "01100001110101011", -- t[50091] = 13
      "0001101" when "01100001110101100", -- t[50092] = 13
      "0001101" when "01100001110101101", -- t[50093] = 13
      "0001101" when "01100001110101110", -- t[50094] = 13
      "0001101" when "01100001110101111", -- t[50095] = 13
      "0001101" when "01100001110110000", -- t[50096] = 13
      "0001101" when "01100001110110001", -- t[50097] = 13
      "0001101" when "01100001110110010", -- t[50098] = 13
      "0001101" when "01100001110110011", -- t[50099] = 13
      "0001101" when "01100001110110100", -- t[50100] = 13
      "0001101" when "01100001110110101", -- t[50101] = 13
      "0001101" when "01100001110110110", -- t[50102] = 13
      "0001101" when "01100001110110111", -- t[50103] = 13
      "0001101" when "01100001110111000", -- t[50104] = 13
      "0001101" when "01100001110111001", -- t[50105] = 13
      "0001101" when "01100001110111010", -- t[50106] = 13
      "0001101" when "01100001110111011", -- t[50107] = 13
      "0001101" when "01100001110111100", -- t[50108] = 13
      "0001101" when "01100001110111101", -- t[50109] = 13
      "0001101" when "01100001110111110", -- t[50110] = 13
      "0001101" when "01100001110111111", -- t[50111] = 13
      "0001101" when "01100001111000000", -- t[50112] = 13
      "0001101" when "01100001111000001", -- t[50113] = 13
      "0001101" when "01100001111000010", -- t[50114] = 13
      "0001101" when "01100001111000011", -- t[50115] = 13
      "0001101" when "01100001111000100", -- t[50116] = 13
      "0001101" when "01100001111000101", -- t[50117] = 13
      "0001101" when "01100001111000110", -- t[50118] = 13
      "0001101" when "01100001111000111", -- t[50119] = 13
      "0001101" when "01100001111001000", -- t[50120] = 13
      "0001101" when "01100001111001001", -- t[50121] = 13
      "0001101" when "01100001111001010", -- t[50122] = 13
      "0001101" when "01100001111001011", -- t[50123] = 13
      "0001101" when "01100001111001100", -- t[50124] = 13
      "0001101" when "01100001111001101", -- t[50125] = 13
      "0001101" when "01100001111001110", -- t[50126] = 13
      "0001101" when "01100001111001111", -- t[50127] = 13
      "0001101" when "01100001111010000", -- t[50128] = 13
      "0001101" when "01100001111010001", -- t[50129] = 13
      "0001101" when "01100001111010010", -- t[50130] = 13
      "0001101" when "01100001111010011", -- t[50131] = 13
      "0001101" when "01100001111010100", -- t[50132] = 13
      "0001101" when "01100001111010101", -- t[50133] = 13
      "0001101" when "01100001111010110", -- t[50134] = 13
      "0001101" when "01100001111010111", -- t[50135] = 13
      "0001101" when "01100001111011000", -- t[50136] = 13
      "0001101" when "01100001111011001", -- t[50137] = 13
      "0001101" when "01100001111011010", -- t[50138] = 13
      "0001101" when "01100001111011011", -- t[50139] = 13
      "0001101" when "01100001111011100", -- t[50140] = 13
      "0001101" when "01100001111011101", -- t[50141] = 13
      "0001101" when "01100001111011110", -- t[50142] = 13
      "0001101" when "01100001111011111", -- t[50143] = 13
      "0001101" when "01100001111100000", -- t[50144] = 13
      "0001101" when "01100001111100001", -- t[50145] = 13
      "0001101" when "01100001111100010", -- t[50146] = 13
      "0001101" when "01100001111100011", -- t[50147] = 13
      "0001101" when "01100001111100100", -- t[50148] = 13
      "0001101" when "01100001111100101", -- t[50149] = 13
      "0001101" when "01100001111100110", -- t[50150] = 13
      "0001101" when "01100001111100111", -- t[50151] = 13
      "0001101" when "01100001111101000", -- t[50152] = 13
      "0001101" when "01100001111101001", -- t[50153] = 13
      "0001101" when "01100001111101010", -- t[50154] = 13
      "0001101" when "01100001111101011", -- t[50155] = 13
      "0001101" when "01100001111101100", -- t[50156] = 13
      "0001101" when "01100001111101101", -- t[50157] = 13
      "0001101" when "01100001111101110", -- t[50158] = 13
      "0001101" when "01100001111101111", -- t[50159] = 13
      "0001101" when "01100001111110000", -- t[50160] = 13
      "0001101" when "01100001111110001", -- t[50161] = 13
      "0001101" when "01100001111110010", -- t[50162] = 13
      "0001101" when "01100001111110011", -- t[50163] = 13
      "0001101" when "01100001111110100", -- t[50164] = 13
      "0001101" when "01100001111110101", -- t[50165] = 13
      "0001101" when "01100001111110110", -- t[50166] = 13
      "0001101" when "01100001111110111", -- t[50167] = 13
      "0001101" when "01100001111111000", -- t[50168] = 13
      "0001101" when "01100001111111001", -- t[50169] = 13
      "0001101" when "01100001111111010", -- t[50170] = 13
      "0001101" when "01100001111111011", -- t[50171] = 13
      "0001101" when "01100001111111100", -- t[50172] = 13
      "0001101" when "01100001111111101", -- t[50173] = 13
      "0001101" when "01100001111111110", -- t[50174] = 13
      "0001101" when "01100001111111111", -- t[50175] = 13
      "0001101" when "01100010000000000", -- t[50176] = 13
      "0001101" when "01100010000000001", -- t[50177] = 13
      "0001101" when "01100010000000010", -- t[50178] = 13
      "0001101" when "01100010000000011", -- t[50179] = 13
      "0001101" when "01100010000000100", -- t[50180] = 13
      "0001101" when "01100010000000101", -- t[50181] = 13
      "0001101" when "01100010000000110", -- t[50182] = 13
      "0001101" when "01100010000000111", -- t[50183] = 13
      "0001101" when "01100010000001000", -- t[50184] = 13
      "0001101" when "01100010000001001", -- t[50185] = 13
      "0001101" when "01100010000001010", -- t[50186] = 13
      "0001101" when "01100010000001011", -- t[50187] = 13
      "0001101" when "01100010000001100", -- t[50188] = 13
      "0001101" when "01100010000001101", -- t[50189] = 13
      "0001101" when "01100010000001110", -- t[50190] = 13
      "0001101" when "01100010000001111", -- t[50191] = 13
      "0001101" when "01100010000010000", -- t[50192] = 13
      "0001101" when "01100010000010001", -- t[50193] = 13
      "0001101" when "01100010000010010", -- t[50194] = 13
      "0001101" when "01100010000010011", -- t[50195] = 13
      "0001101" when "01100010000010100", -- t[50196] = 13
      "0001101" when "01100010000010101", -- t[50197] = 13
      "0001101" when "01100010000010110", -- t[50198] = 13
      "0001101" when "01100010000010111", -- t[50199] = 13
      "0001101" when "01100010000011000", -- t[50200] = 13
      "0001101" when "01100010000011001", -- t[50201] = 13
      "0001101" when "01100010000011010", -- t[50202] = 13
      "0001101" when "01100010000011011", -- t[50203] = 13
      "0001101" when "01100010000011100", -- t[50204] = 13
      "0001101" when "01100010000011101", -- t[50205] = 13
      "0001101" when "01100010000011110", -- t[50206] = 13
      "0001101" when "01100010000011111", -- t[50207] = 13
      "0001101" when "01100010000100000", -- t[50208] = 13
      "0001101" when "01100010000100001", -- t[50209] = 13
      "0001101" when "01100010000100010", -- t[50210] = 13
      "0001101" when "01100010000100011", -- t[50211] = 13
      "0001101" when "01100010000100100", -- t[50212] = 13
      "0001101" when "01100010000100101", -- t[50213] = 13
      "0001101" when "01100010000100110", -- t[50214] = 13
      "0001101" when "01100010000100111", -- t[50215] = 13
      "0001101" when "01100010000101000", -- t[50216] = 13
      "0001101" when "01100010000101001", -- t[50217] = 13
      "0001101" when "01100010000101010", -- t[50218] = 13
      "0001101" when "01100010000101011", -- t[50219] = 13
      "0001101" when "01100010000101100", -- t[50220] = 13
      "0001101" when "01100010000101101", -- t[50221] = 13
      "0001101" when "01100010000101110", -- t[50222] = 13
      "0001101" when "01100010000101111", -- t[50223] = 13
      "0001101" when "01100010000110000", -- t[50224] = 13
      "0001101" when "01100010000110001", -- t[50225] = 13
      "0001101" when "01100010000110010", -- t[50226] = 13
      "0001101" when "01100010000110011", -- t[50227] = 13
      "0001101" when "01100010000110100", -- t[50228] = 13
      "0001101" when "01100010000110101", -- t[50229] = 13
      "0001101" when "01100010000110110", -- t[50230] = 13
      "0001101" when "01100010000110111", -- t[50231] = 13
      "0001101" when "01100010000111000", -- t[50232] = 13
      "0001101" when "01100010000111001", -- t[50233] = 13
      "0001101" when "01100010000111010", -- t[50234] = 13
      "0001101" when "01100010000111011", -- t[50235] = 13
      "0001101" when "01100010000111100", -- t[50236] = 13
      "0001101" when "01100010000111101", -- t[50237] = 13
      "0001101" when "01100010000111110", -- t[50238] = 13
      "0001101" when "01100010000111111", -- t[50239] = 13
      "0001101" when "01100010001000000", -- t[50240] = 13
      "0001101" when "01100010001000001", -- t[50241] = 13
      "0001101" when "01100010001000010", -- t[50242] = 13
      "0001101" when "01100010001000011", -- t[50243] = 13
      "0001101" when "01100010001000100", -- t[50244] = 13
      "0001101" when "01100010001000101", -- t[50245] = 13
      "0001101" when "01100010001000110", -- t[50246] = 13
      "0001101" when "01100010001000111", -- t[50247] = 13
      "0001101" when "01100010001001000", -- t[50248] = 13
      "0001101" when "01100010001001001", -- t[50249] = 13
      "0001101" when "01100010001001010", -- t[50250] = 13
      "0001101" when "01100010001001011", -- t[50251] = 13
      "0001101" when "01100010001001100", -- t[50252] = 13
      "0001101" when "01100010001001101", -- t[50253] = 13
      "0001101" when "01100010001001110", -- t[50254] = 13
      "0001101" when "01100010001001111", -- t[50255] = 13
      "0001101" when "01100010001010000", -- t[50256] = 13
      "0001101" when "01100010001010001", -- t[50257] = 13
      "0001101" when "01100010001010010", -- t[50258] = 13
      "0001101" when "01100010001010011", -- t[50259] = 13
      "0001101" when "01100010001010100", -- t[50260] = 13
      "0001101" when "01100010001010101", -- t[50261] = 13
      "0001101" when "01100010001010110", -- t[50262] = 13
      "0001101" when "01100010001010111", -- t[50263] = 13
      "0001101" when "01100010001011000", -- t[50264] = 13
      "0001101" when "01100010001011001", -- t[50265] = 13
      "0001101" when "01100010001011010", -- t[50266] = 13
      "0001101" when "01100010001011011", -- t[50267] = 13
      "0001101" when "01100010001011100", -- t[50268] = 13
      "0001101" when "01100010001011101", -- t[50269] = 13
      "0001101" when "01100010001011110", -- t[50270] = 13
      "0001101" when "01100010001011111", -- t[50271] = 13
      "0001101" when "01100010001100000", -- t[50272] = 13
      "0001101" when "01100010001100001", -- t[50273] = 13
      "0001101" when "01100010001100010", -- t[50274] = 13
      "0001101" when "01100010001100011", -- t[50275] = 13
      "0001101" when "01100010001100100", -- t[50276] = 13
      "0001101" when "01100010001100101", -- t[50277] = 13
      "0001101" when "01100010001100110", -- t[50278] = 13
      "0001101" when "01100010001100111", -- t[50279] = 13
      "0001101" when "01100010001101000", -- t[50280] = 13
      "0001101" when "01100010001101001", -- t[50281] = 13
      "0001101" when "01100010001101010", -- t[50282] = 13
      "0001101" when "01100010001101011", -- t[50283] = 13
      "0001101" when "01100010001101100", -- t[50284] = 13
      "0001101" when "01100010001101101", -- t[50285] = 13
      "0001101" when "01100010001101110", -- t[50286] = 13
      "0001101" when "01100010001101111", -- t[50287] = 13
      "0001101" when "01100010001110000", -- t[50288] = 13
      "0001101" when "01100010001110001", -- t[50289] = 13
      "0001101" when "01100010001110010", -- t[50290] = 13
      "0001101" when "01100010001110011", -- t[50291] = 13
      "0001101" when "01100010001110100", -- t[50292] = 13
      "0001101" when "01100010001110101", -- t[50293] = 13
      "0001101" when "01100010001110110", -- t[50294] = 13
      "0001101" when "01100010001110111", -- t[50295] = 13
      "0001101" when "01100010001111000", -- t[50296] = 13
      "0001101" when "01100010001111001", -- t[50297] = 13
      "0001101" when "01100010001111010", -- t[50298] = 13
      "0001101" when "01100010001111011", -- t[50299] = 13
      "0001101" when "01100010001111100", -- t[50300] = 13
      "0001101" when "01100010001111101", -- t[50301] = 13
      "0001101" when "01100010001111110", -- t[50302] = 13
      "0001101" when "01100010001111111", -- t[50303] = 13
      "0001101" when "01100010010000000", -- t[50304] = 13
      "0001101" when "01100010010000001", -- t[50305] = 13
      "0001101" when "01100010010000010", -- t[50306] = 13
      "0001101" when "01100010010000011", -- t[50307] = 13
      "0001101" when "01100010010000100", -- t[50308] = 13
      "0001101" when "01100010010000101", -- t[50309] = 13
      "0001101" when "01100010010000110", -- t[50310] = 13
      "0001101" when "01100010010000111", -- t[50311] = 13
      "0001101" when "01100010010001000", -- t[50312] = 13
      "0001101" when "01100010010001001", -- t[50313] = 13
      "0001101" when "01100010010001010", -- t[50314] = 13
      "0001101" when "01100010010001011", -- t[50315] = 13
      "0001101" when "01100010010001100", -- t[50316] = 13
      "0001101" when "01100010010001101", -- t[50317] = 13
      "0001101" when "01100010010001110", -- t[50318] = 13
      "0001101" when "01100010010001111", -- t[50319] = 13
      "0001101" when "01100010010010000", -- t[50320] = 13
      "0001101" when "01100010010010001", -- t[50321] = 13
      "0001101" when "01100010010010010", -- t[50322] = 13
      "0001101" when "01100010010010011", -- t[50323] = 13
      "0001101" when "01100010010010100", -- t[50324] = 13
      "0001101" when "01100010010010101", -- t[50325] = 13
      "0001101" when "01100010010010110", -- t[50326] = 13
      "0001101" when "01100010010010111", -- t[50327] = 13
      "0001101" when "01100010010011000", -- t[50328] = 13
      "0001101" when "01100010010011001", -- t[50329] = 13
      "0001101" when "01100010010011010", -- t[50330] = 13
      "0001101" when "01100010010011011", -- t[50331] = 13
      "0001101" when "01100010010011100", -- t[50332] = 13
      "0001101" when "01100010010011101", -- t[50333] = 13
      "0001101" when "01100010010011110", -- t[50334] = 13
      "0001101" when "01100010010011111", -- t[50335] = 13
      "0001101" when "01100010010100000", -- t[50336] = 13
      "0001101" when "01100010010100001", -- t[50337] = 13
      "0001101" when "01100010010100010", -- t[50338] = 13
      "0001101" when "01100010010100011", -- t[50339] = 13
      "0001101" when "01100010010100100", -- t[50340] = 13
      "0001101" when "01100010010100101", -- t[50341] = 13
      "0001101" when "01100010010100110", -- t[50342] = 13
      "0001101" when "01100010010100111", -- t[50343] = 13
      "0001101" when "01100010010101000", -- t[50344] = 13
      "0001101" when "01100010010101001", -- t[50345] = 13
      "0001101" when "01100010010101010", -- t[50346] = 13
      "0001101" when "01100010010101011", -- t[50347] = 13
      "0001101" when "01100010010101100", -- t[50348] = 13
      "0001101" when "01100010010101101", -- t[50349] = 13
      "0001101" when "01100010010101110", -- t[50350] = 13
      "0001101" when "01100010010101111", -- t[50351] = 13
      "0001101" when "01100010010110000", -- t[50352] = 13
      "0001101" when "01100010010110001", -- t[50353] = 13
      "0001101" when "01100010010110010", -- t[50354] = 13
      "0001101" when "01100010010110011", -- t[50355] = 13
      "0001101" when "01100010010110100", -- t[50356] = 13
      "0001101" when "01100010010110101", -- t[50357] = 13
      "0001101" when "01100010010110110", -- t[50358] = 13
      "0001101" when "01100010010110111", -- t[50359] = 13
      "0001101" when "01100010010111000", -- t[50360] = 13
      "0001101" when "01100010010111001", -- t[50361] = 13
      "0001101" when "01100010010111010", -- t[50362] = 13
      "0001101" when "01100010010111011", -- t[50363] = 13
      "0001101" when "01100010010111100", -- t[50364] = 13
      "0001101" when "01100010010111101", -- t[50365] = 13
      "0001101" when "01100010010111110", -- t[50366] = 13
      "0001101" when "01100010010111111", -- t[50367] = 13
      "0001101" when "01100010011000000", -- t[50368] = 13
      "0001101" when "01100010011000001", -- t[50369] = 13
      "0001101" when "01100010011000010", -- t[50370] = 13
      "0001101" when "01100010011000011", -- t[50371] = 13
      "0001101" when "01100010011000100", -- t[50372] = 13
      "0001101" when "01100010011000101", -- t[50373] = 13
      "0001101" when "01100010011000110", -- t[50374] = 13
      "0001101" when "01100010011000111", -- t[50375] = 13
      "0001101" when "01100010011001000", -- t[50376] = 13
      "0001101" when "01100010011001001", -- t[50377] = 13
      "0001101" when "01100010011001010", -- t[50378] = 13
      "0001101" when "01100010011001011", -- t[50379] = 13
      "0001101" when "01100010011001100", -- t[50380] = 13
      "0001101" when "01100010011001101", -- t[50381] = 13
      "0001101" when "01100010011001110", -- t[50382] = 13
      "0001101" when "01100010011001111", -- t[50383] = 13
      "0001101" when "01100010011010000", -- t[50384] = 13
      "0001101" when "01100010011010001", -- t[50385] = 13
      "0001101" when "01100010011010010", -- t[50386] = 13
      "0001101" when "01100010011010011", -- t[50387] = 13
      "0001101" when "01100010011010100", -- t[50388] = 13
      "0001101" when "01100010011010101", -- t[50389] = 13
      "0001101" when "01100010011010110", -- t[50390] = 13
      "0001101" when "01100010011010111", -- t[50391] = 13
      "0001101" when "01100010011011000", -- t[50392] = 13
      "0001101" when "01100010011011001", -- t[50393] = 13
      "0001101" when "01100010011011010", -- t[50394] = 13
      "0001101" when "01100010011011011", -- t[50395] = 13
      "0001101" when "01100010011011100", -- t[50396] = 13
      "0001101" when "01100010011011101", -- t[50397] = 13
      "0001101" when "01100010011011110", -- t[50398] = 13
      "0001101" when "01100010011011111", -- t[50399] = 13
      "0001101" when "01100010011100000", -- t[50400] = 13
      "0001101" when "01100010011100001", -- t[50401] = 13
      "0001101" when "01100010011100010", -- t[50402] = 13
      "0001101" when "01100010011100011", -- t[50403] = 13
      "0001101" when "01100010011100100", -- t[50404] = 13
      "0001101" when "01100010011100101", -- t[50405] = 13
      "0001101" when "01100010011100110", -- t[50406] = 13
      "0001101" when "01100010011100111", -- t[50407] = 13
      "0001101" when "01100010011101000", -- t[50408] = 13
      "0001101" when "01100010011101001", -- t[50409] = 13
      "0001101" when "01100010011101010", -- t[50410] = 13
      "0001101" when "01100010011101011", -- t[50411] = 13
      "0001101" when "01100010011101100", -- t[50412] = 13
      "0001101" when "01100010011101101", -- t[50413] = 13
      "0001101" when "01100010011101110", -- t[50414] = 13
      "0001101" when "01100010011101111", -- t[50415] = 13
      "0001101" when "01100010011110000", -- t[50416] = 13
      "0001101" when "01100010011110001", -- t[50417] = 13
      "0001101" when "01100010011110010", -- t[50418] = 13
      "0001101" when "01100010011110011", -- t[50419] = 13
      "0001101" when "01100010011110100", -- t[50420] = 13
      "0001101" when "01100010011110101", -- t[50421] = 13
      "0001101" when "01100010011110110", -- t[50422] = 13
      "0001101" when "01100010011110111", -- t[50423] = 13
      "0001101" when "01100010011111000", -- t[50424] = 13
      "0001101" when "01100010011111001", -- t[50425] = 13
      "0001101" when "01100010011111010", -- t[50426] = 13
      "0001101" when "01100010011111011", -- t[50427] = 13
      "0001101" when "01100010011111100", -- t[50428] = 13
      "0001101" when "01100010011111101", -- t[50429] = 13
      "0001101" when "01100010011111110", -- t[50430] = 13
      "0001101" when "01100010011111111", -- t[50431] = 13
      "0001101" when "01100010100000000", -- t[50432] = 13
      "0001101" when "01100010100000001", -- t[50433] = 13
      "0001101" when "01100010100000010", -- t[50434] = 13
      "0001101" when "01100010100000011", -- t[50435] = 13
      "0001101" when "01100010100000100", -- t[50436] = 13
      "0001101" when "01100010100000101", -- t[50437] = 13
      "0001101" when "01100010100000110", -- t[50438] = 13
      "0001101" when "01100010100000111", -- t[50439] = 13
      "0001101" when "01100010100001000", -- t[50440] = 13
      "0001101" when "01100010100001001", -- t[50441] = 13
      "0001101" when "01100010100001010", -- t[50442] = 13
      "0001101" when "01100010100001011", -- t[50443] = 13
      "0001101" when "01100010100001100", -- t[50444] = 13
      "0001101" when "01100010100001101", -- t[50445] = 13
      "0001101" when "01100010100001110", -- t[50446] = 13
      "0001101" when "01100010100001111", -- t[50447] = 13
      "0001101" when "01100010100010000", -- t[50448] = 13
      "0001101" when "01100010100010001", -- t[50449] = 13
      "0001101" when "01100010100010010", -- t[50450] = 13
      "0001101" when "01100010100010011", -- t[50451] = 13
      "0001101" when "01100010100010100", -- t[50452] = 13
      "0001101" when "01100010100010101", -- t[50453] = 13
      "0001101" when "01100010100010110", -- t[50454] = 13
      "0001101" when "01100010100010111", -- t[50455] = 13
      "0001101" when "01100010100011000", -- t[50456] = 13
      "0001101" when "01100010100011001", -- t[50457] = 13
      "0001101" when "01100010100011010", -- t[50458] = 13
      "0001101" when "01100010100011011", -- t[50459] = 13
      "0001101" when "01100010100011100", -- t[50460] = 13
      "0001101" when "01100010100011101", -- t[50461] = 13
      "0001101" when "01100010100011110", -- t[50462] = 13
      "0001101" when "01100010100011111", -- t[50463] = 13
      "0001101" when "01100010100100000", -- t[50464] = 13
      "0001101" when "01100010100100001", -- t[50465] = 13
      "0001101" when "01100010100100010", -- t[50466] = 13
      "0001101" when "01100010100100011", -- t[50467] = 13
      "0001101" when "01100010100100100", -- t[50468] = 13
      "0001101" when "01100010100100101", -- t[50469] = 13
      "0001101" when "01100010100100110", -- t[50470] = 13
      "0001101" when "01100010100100111", -- t[50471] = 13
      "0001101" when "01100010100101000", -- t[50472] = 13
      "0001101" when "01100010100101001", -- t[50473] = 13
      "0001101" when "01100010100101010", -- t[50474] = 13
      "0001101" when "01100010100101011", -- t[50475] = 13
      "0001101" when "01100010100101100", -- t[50476] = 13
      "0001101" when "01100010100101101", -- t[50477] = 13
      "0001101" when "01100010100101110", -- t[50478] = 13
      "0001101" when "01100010100101111", -- t[50479] = 13
      "0001101" when "01100010100110000", -- t[50480] = 13
      "0001101" when "01100010100110001", -- t[50481] = 13
      "0001101" when "01100010100110010", -- t[50482] = 13
      "0001101" when "01100010100110011", -- t[50483] = 13
      "0001101" when "01100010100110100", -- t[50484] = 13
      "0001101" when "01100010100110101", -- t[50485] = 13
      "0001101" when "01100010100110110", -- t[50486] = 13
      "0001101" when "01100010100110111", -- t[50487] = 13
      "0001101" when "01100010100111000", -- t[50488] = 13
      "0001101" when "01100010100111001", -- t[50489] = 13
      "0001101" when "01100010100111010", -- t[50490] = 13
      "0001101" when "01100010100111011", -- t[50491] = 13
      "0001101" when "01100010100111100", -- t[50492] = 13
      "0001101" when "01100010100111101", -- t[50493] = 13
      "0001101" when "01100010100111110", -- t[50494] = 13
      "0001101" when "01100010100111111", -- t[50495] = 13
      "0001101" when "01100010101000000", -- t[50496] = 13
      "0001101" when "01100010101000001", -- t[50497] = 13
      "0001101" when "01100010101000010", -- t[50498] = 13
      "0001101" when "01100010101000011", -- t[50499] = 13
      "0001101" when "01100010101000100", -- t[50500] = 13
      "0001101" when "01100010101000101", -- t[50501] = 13
      "0001101" when "01100010101000110", -- t[50502] = 13
      "0001101" when "01100010101000111", -- t[50503] = 13
      "0001101" when "01100010101001000", -- t[50504] = 13
      "0001101" when "01100010101001001", -- t[50505] = 13
      "0001101" when "01100010101001010", -- t[50506] = 13
      "0001101" when "01100010101001011", -- t[50507] = 13
      "0001101" when "01100010101001100", -- t[50508] = 13
      "0001101" when "01100010101001101", -- t[50509] = 13
      "0001101" when "01100010101001110", -- t[50510] = 13
      "0001101" when "01100010101001111", -- t[50511] = 13
      "0001101" when "01100010101010000", -- t[50512] = 13
      "0001101" when "01100010101010001", -- t[50513] = 13
      "0001101" when "01100010101010010", -- t[50514] = 13
      "0001101" when "01100010101010011", -- t[50515] = 13
      "0001101" when "01100010101010100", -- t[50516] = 13
      "0001101" when "01100010101010101", -- t[50517] = 13
      "0001101" when "01100010101010110", -- t[50518] = 13
      "0001101" when "01100010101010111", -- t[50519] = 13
      "0001101" when "01100010101011000", -- t[50520] = 13
      "0001101" when "01100010101011001", -- t[50521] = 13
      "0001101" when "01100010101011010", -- t[50522] = 13
      "0001101" when "01100010101011011", -- t[50523] = 13
      "0001101" when "01100010101011100", -- t[50524] = 13
      "0001101" when "01100010101011101", -- t[50525] = 13
      "0001101" when "01100010101011110", -- t[50526] = 13
      "0001101" when "01100010101011111", -- t[50527] = 13
      "0001101" when "01100010101100000", -- t[50528] = 13
      "0001101" when "01100010101100001", -- t[50529] = 13
      "0001101" when "01100010101100010", -- t[50530] = 13
      "0001101" when "01100010101100011", -- t[50531] = 13
      "0001101" when "01100010101100100", -- t[50532] = 13
      "0001101" when "01100010101100101", -- t[50533] = 13
      "0001101" when "01100010101100110", -- t[50534] = 13
      "0001101" when "01100010101100111", -- t[50535] = 13
      "0001101" when "01100010101101000", -- t[50536] = 13
      "0001101" when "01100010101101001", -- t[50537] = 13
      "0001101" when "01100010101101010", -- t[50538] = 13
      "0001101" when "01100010101101011", -- t[50539] = 13
      "0001101" when "01100010101101100", -- t[50540] = 13
      "0001101" when "01100010101101101", -- t[50541] = 13
      "0001101" when "01100010101101110", -- t[50542] = 13
      "0001101" when "01100010101101111", -- t[50543] = 13
      "0001101" when "01100010101110000", -- t[50544] = 13
      "0001101" when "01100010101110001", -- t[50545] = 13
      "0001101" when "01100010101110010", -- t[50546] = 13
      "0001101" when "01100010101110011", -- t[50547] = 13
      "0001101" when "01100010101110100", -- t[50548] = 13
      "0001101" when "01100010101110101", -- t[50549] = 13
      "0001101" when "01100010101110110", -- t[50550] = 13
      "0001101" when "01100010101110111", -- t[50551] = 13
      "0001101" when "01100010101111000", -- t[50552] = 13
      "0001101" when "01100010101111001", -- t[50553] = 13
      "0001101" when "01100010101111010", -- t[50554] = 13
      "0001101" when "01100010101111011", -- t[50555] = 13
      "0001101" when "01100010101111100", -- t[50556] = 13
      "0001101" when "01100010101111101", -- t[50557] = 13
      "0001101" when "01100010101111110", -- t[50558] = 13
      "0001101" when "01100010101111111", -- t[50559] = 13
      "0001101" when "01100010110000000", -- t[50560] = 13
      "0001101" when "01100010110000001", -- t[50561] = 13
      "0001101" when "01100010110000010", -- t[50562] = 13
      "0001101" when "01100010110000011", -- t[50563] = 13
      "0001101" when "01100010110000100", -- t[50564] = 13
      "0001101" when "01100010110000101", -- t[50565] = 13
      "0001101" when "01100010110000110", -- t[50566] = 13
      "0001101" when "01100010110000111", -- t[50567] = 13
      "0001101" when "01100010110001000", -- t[50568] = 13
      "0001101" when "01100010110001001", -- t[50569] = 13
      "0001101" when "01100010110001010", -- t[50570] = 13
      "0001101" when "01100010110001011", -- t[50571] = 13
      "0001101" when "01100010110001100", -- t[50572] = 13
      "0001101" when "01100010110001101", -- t[50573] = 13
      "0001101" when "01100010110001110", -- t[50574] = 13
      "0001101" when "01100010110001111", -- t[50575] = 13
      "0001101" when "01100010110010000", -- t[50576] = 13
      "0001101" when "01100010110010001", -- t[50577] = 13
      "0001101" when "01100010110010010", -- t[50578] = 13
      "0001101" when "01100010110010011", -- t[50579] = 13
      "0001101" when "01100010110010100", -- t[50580] = 13
      "0001101" when "01100010110010101", -- t[50581] = 13
      "0001101" when "01100010110010110", -- t[50582] = 13
      "0001101" when "01100010110010111", -- t[50583] = 13
      "0001101" when "01100010110011000", -- t[50584] = 13
      "0001101" when "01100010110011001", -- t[50585] = 13
      "0001101" when "01100010110011010", -- t[50586] = 13
      "0001101" when "01100010110011011", -- t[50587] = 13
      "0001101" when "01100010110011100", -- t[50588] = 13
      "0001101" when "01100010110011101", -- t[50589] = 13
      "0001101" when "01100010110011110", -- t[50590] = 13
      "0001101" when "01100010110011111", -- t[50591] = 13
      "0001101" when "01100010110100000", -- t[50592] = 13
      "0001101" when "01100010110100001", -- t[50593] = 13
      "0001101" when "01100010110100010", -- t[50594] = 13
      "0001101" when "01100010110100011", -- t[50595] = 13
      "0001101" when "01100010110100100", -- t[50596] = 13
      "0001101" when "01100010110100101", -- t[50597] = 13
      "0001101" when "01100010110100110", -- t[50598] = 13
      "0001101" when "01100010110100111", -- t[50599] = 13
      "0001101" when "01100010110101000", -- t[50600] = 13
      "0001101" when "01100010110101001", -- t[50601] = 13
      "0001101" when "01100010110101010", -- t[50602] = 13
      "0001101" when "01100010110101011", -- t[50603] = 13
      "0001101" when "01100010110101100", -- t[50604] = 13
      "0001101" when "01100010110101101", -- t[50605] = 13
      "0001101" when "01100010110101110", -- t[50606] = 13
      "0001101" when "01100010110101111", -- t[50607] = 13
      "0001101" when "01100010110110000", -- t[50608] = 13
      "0001101" when "01100010110110001", -- t[50609] = 13
      "0001101" when "01100010110110010", -- t[50610] = 13
      "0001101" when "01100010110110011", -- t[50611] = 13
      "0001101" when "01100010110110100", -- t[50612] = 13
      "0001101" when "01100010110110101", -- t[50613] = 13
      "0001101" when "01100010110110110", -- t[50614] = 13
      "0001101" when "01100010110110111", -- t[50615] = 13
      "0001101" when "01100010110111000", -- t[50616] = 13
      "0001101" when "01100010110111001", -- t[50617] = 13
      "0001101" when "01100010110111010", -- t[50618] = 13
      "0001101" when "01100010110111011", -- t[50619] = 13
      "0001101" when "01100010110111100", -- t[50620] = 13
      "0001101" when "01100010110111101", -- t[50621] = 13
      "0001101" when "01100010110111110", -- t[50622] = 13
      "0001101" when "01100010110111111", -- t[50623] = 13
      "0001101" when "01100010111000000", -- t[50624] = 13
      "0001101" when "01100010111000001", -- t[50625] = 13
      "0001101" when "01100010111000010", -- t[50626] = 13
      "0001101" when "01100010111000011", -- t[50627] = 13
      "0001101" when "01100010111000100", -- t[50628] = 13
      "0001101" when "01100010111000101", -- t[50629] = 13
      "0001101" when "01100010111000110", -- t[50630] = 13
      "0001101" when "01100010111000111", -- t[50631] = 13
      "0001101" when "01100010111001000", -- t[50632] = 13
      "0001101" when "01100010111001001", -- t[50633] = 13
      "0001101" when "01100010111001010", -- t[50634] = 13
      "0001101" when "01100010111001011", -- t[50635] = 13
      "0001101" when "01100010111001100", -- t[50636] = 13
      "0001101" when "01100010111001101", -- t[50637] = 13
      "0001101" when "01100010111001110", -- t[50638] = 13
      "0001101" when "01100010111001111", -- t[50639] = 13
      "0001101" when "01100010111010000", -- t[50640] = 13
      "0001101" when "01100010111010001", -- t[50641] = 13
      "0001101" when "01100010111010010", -- t[50642] = 13
      "0001101" when "01100010111010011", -- t[50643] = 13
      "0001101" when "01100010111010100", -- t[50644] = 13
      "0001101" when "01100010111010101", -- t[50645] = 13
      "0001101" when "01100010111010110", -- t[50646] = 13
      "0001101" when "01100010111010111", -- t[50647] = 13
      "0001101" when "01100010111011000", -- t[50648] = 13
      "0001101" when "01100010111011001", -- t[50649] = 13
      "0001101" when "01100010111011010", -- t[50650] = 13
      "0001101" when "01100010111011011", -- t[50651] = 13
      "0001101" when "01100010111011100", -- t[50652] = 13
      "0001101" when "01100010111011101", -- t[50653] = 13
      "0001101" when "01100010111011110", -- t[50654] = 13
      "0001101" when "01100010111011111", -- t[50655] = 13
      "0001101" when "01100010111100000", -- t[50656] = 13
      "0001101" when "01100010111100001", -- t[50657] = 13
      "0001101" when "01100010111100010", -- t[50658] = 13
      "0001101" when "01100010111100011", -- t[50659] = 13
      "0001101" when "01100010111100100", -- t[50660] = 13
      "0001101" when "01100010111100101", -- t[50661] = 13
      "0001101" when "01100010111100110", -- t[50662] = 13
      "0001101" when "01100010111100111", -- t[50663] = 13
      "0001101" when "01100010111101000", -- t[50664] = 13
      "0001101" when "01100010111101001", -- t[50665] = 13
      "0001101" when "01100010111101010", -- t[50666] = 13
      "0001101" when "01100010111101011", -- t[50667] = 13
      "0001101" when "01100010111101100", -- t[50668] = 13
      "0001101" when "01100010111101101", -- t[50669] = 13
      "0001101" when "01100010111101110", -- t[50670] = 13
      "0001101" when "01100010111101111", -- t[50671] = 13
      "0001101" when "01100010111110000", -- t[50672] = 13
      "0001101" when "01100010111110001", -- t[50673] = 13
      "0001101" when "01100010111110010", -- t[50674] = 13
      "0001101" when "01100010111110011", -- t[50675] = 13
      "0001101" when "01100010111110100", -- t[50676] = 13
      "0001101" when "01100010111110101", -- t[50677] = 13
      "0001101" when "01100010111110110", -- t[50678] = 13
      "0001101" when "01100010111110111", -- t[50679] = 13
      "0001101" when "01100010111111000", -- t[50680] = 13
      "0001101" when "01100010111111001", -- t[50681] = 13
      "0001101" when "01100010111111010", -- t[50682] = 13
      "0001101" when "01100010111111011", -- t[50683] = 13
      "0001101" when "01100010111111100", -- t[50684] = 13
      "0001101" when "01100010111111101", -- t[50685] = 13
      "0001101" when "01100010111111110", -- t[50686] = 13
      "0001101" when "01100010111111111", -- t[50687] = 13
      "0001101" when "01100011000000000", -- t[50688] = 13
      "0001101" when "01100011000000001", -- t[50689] = 13
      "0001101" when "01100011000000010", -- t[50690] = 13
      "0001101" when "01100011000000011", -- t[50691] = 13
      "0001101" when "01100011000000100", -- t[50692] = 13
      "0001101" when "01100011000000101", -- t[50693] = 13
      "0001101" when "01100011000000110", -- t[50694] = 13
      "0001101" when "01100011000000111", -- t[50695] = 13
      "0001101" when "01100011000001000", -- t[50696] = 13
      "0001101" when "01100011000001001", -- t[50697] = 13
      "0001101" when "01100011000001010", -- t[50698] = 13
      "0001101" when "01100011000001011", -- t[50699] = 13
      "0001101" when "01100011000001100", -- t[50700] = 13
      "0001101" when "01100011000001101", -- t[50701] = 13
      "0001101" when "01100011000001110", -- t[50702] = 13
      "0001101" when "01100011000001111", -- t[50703] = 13
      "0001101" when "01100011000010000", -- t[50704] = 13
      "0001101" when "01100011000010001", -- t[50705] = 13
      "0001101" when "01100011000010010", -- t[50706] = 13
      "0001101" when "01100011000010011", -- t[50707] = 13
      "0001101" when "01100011000010100", -- t[50708] = 13
      "0001101" when "01100011000010101", -- t[50709] = 13
      "0001101" when "01100011000010110", -- t[50710] = 13
      "0001101" when "01100011000010111", -- t[50711] = 13
      "0001101" when "01100011000011000", -- t[50712] = 13
      "0001101" when "01100011000011001", -- t[50713] = 13
      "0001101" when "01100011000011010", -- t[50714] = 13
      "0001101" when "01100011000011011", -- t[50715] = 13
      "0001101" when "01100011000011100", -- t[50716] = 13
      "0001101" when "01100011000011101", -- t[50717] = 13
      "0001101" when "01100011000011110", -- t[50718] = 13
      "0001101" when "01100011000011111", -- t[50719] = 13
      "0001101" when "01100011000100000", -- t[50720] = 13
      "0001101" when "01100011000100001", -- t[50721] = 13
      "0001101" when "01100011000100010", -- t[50722] = 13
      "0001101" when "01100011000100011", -- t[50723] = 13
      "0001101" when "01100011000100100", -- t[50724] = 13
      "0001101" when "01100011000100101", -- t[50725] = 13
      "0001101" when "01100011000100110", -- t[50726] = 13
      "0001101" when "01100011000100111", -- t[50727] = 13
      "0001101" when "01100011000101000", -- t[50728] = 13
      "0001101" when "01100011000101001", -- t[50729] = 13
      "0001101" when "01100011000101010", -- t[50730] = 13
      "0001101" when "01100011000101011", -- t[50731] = 13
      "0001101" when "01100011000101100", -- t[50732] = 13
      "0001101" when "01100011000101101", -- t[50733] = 13
      "0001101" when "01100011000101110", -- t[50734] = 13
      "0001101" when "01100011000101111", -- t[50735] = 13
      "0001101" when "01100011000110000", -- t[50736] = 13
      "0001101" when "01100011000110001", -- t[50737] = 13
      "0001101" when "01100011000110010", -- t[50738] = 13
      "0001101" when "01100011000110011", -- t[50739] = 13
      "0001101" when "01100011000110100", -- t[50740] = 13
      "0001101" when "01100011000110101", -- t[50741] = 13
      "0001101" when "01100011000110110", -- t[50742] = 13
      "0001101" when "01100011000110111", -- t[50743] = 13
      "0001101" when "01100011000111000", -- t[50744] = 13
      "0001101" when "01100011000111001", -- t[50745] = 13
      "0001101" when "01100011000111010", -- t[50746] = 13
      "0001101" when "01100011000111011", -- t[50747] = 13
      "0001101" when "01100011000111100", -- t[50748] = 13
      "0001101" when "01100011000111101", -- t[50749] = 13
      "0001101" when "01100011000111110", -- t[50750] = 13
      "0001101" when "01100011000111111", -- t[50751] = 13
      "0001101" when "01100011001000000", -- t[50752] = 13
      "0001101" when "01100011001000001", -- t[50753] = 13
      "0001101" when "01100011001000010", -- t[50754] = 13
      "0001101" when "01100011001000011", -- t[50755] = 13
      "0001101" when "01100011001000100", -- t[50756] = 13
      "0001101" when "01100011001000101", -- t[50757] = 13
      "0001101" when "01100011001000110", -- t[50758] = 13
      "0001101" when "01100011001000111", -- t[50759] = 13
      "0001101" when "01100011001001000", -- t[50760] = 13
      "0001101" when "01100011001001001", -- t[50761] = 13
      "0001101" when "01100011001001010", -- t[50762] = 13
      "0001101" when "01100011001001011", -- t[50763] = 13
      "0001101" when "01100011001001100", -- t[50764] = 13
      "0001101" when "01100011001001101", -- t[50765] = 13
      "0001101" when "01100011001001110", -- t[50766] = 13
      "0001101" when "01100011001001111", -- t[50767] = 13
      "0001101" when "01100011001010000", -- t[50768] = 13
      "0001101" when "01100011001010001", -- t[50769] = 13
      "0001101" when "01100011001010010", -- t[50770] = 13
      "0001101" when "01100011001010011", -- t[50771] = 13
      "0001101" when "01100011001010100", -- t[50772] = 13
      "0001101" when "01100011001010101", -- t[50773] = 13
      "0001101" when "01100011001010110", -- t[50774] = 13
      "0001101" when "01100011001010111", -- t[50775] = 13
      "0001101" when "01100011001011000", -- t[50776] = 13
      "0001101" when "01100011001011001", -- t[50777] = 13
      "0001101" when "01100011001011010", -- t[50778] = 13
      "0001101" when "01100011001011011", -- t[50779] = 13
      "0001101" when "01100011001011100", -- t[50780] = 13
      "0001101" when "01100011001011101", -- t[50781] = 13
      "0001101" when "01100011001011110", -- t[50782] = 13
      "0001101" when "01100011001011111", -- t[50783] = 13
      "0001101" when "01100011001100000", -- t[50784] = 13
      "0001101" when "01100011001100001", -- t[50785] = 13
      "0001101" when "01100011001100010", -- t[50786] = 13
      "0001101" when "01100011001100011", -- t[50787] = 13
      "0001101" when "01100011001100100", -- t[50788] = 13
      "0001101" when "01100011001100101", -- t[50789] = 13
      "0001101" when "01100011001100110", -- t[50790] = 13
      "0001101" when "01100011001100111", -- t[50791] = 13
      "0001101" when "01100011001101000", -- t[50792] = 13
      "0001101" when "01100011001101001", -- t[50793] = 13
      "0001101" when "01100011001101010", -- t[50794] = 13
      "0001101" when "01100011001101011", -- t[50795] = 13
      "0001101" when "01100011001101100", -- t[50796] = 13
      "0001101" when "01100011001101101", -- t[50797] = 13
      "0001101" when "01100011001101110", -- t[50798] = 13
      "0001101" when "01100011001101111", -- t[50799] = 13
      "0001101" when "01100011001110000", -- t[50800] = 13
      "0001101" when "01100011001110001", -- t[50801] = 13
      "0001101" when "01100011001110010", -- t[50802] = 13
      "0001101" when "01100011001110011", -- t[50803] = 13
      "0001101" when "01100011001110100", -- t[50804] = 13
      "0001101" when "01100011001110101", -- t[50805] = 13
      "0001101" when "01100011001110110", -- t[50806] = 13
      "0001101" when "01100011001110111", -- t[50807] = 13
      "0001101" when "01100011001111000", -- t[50808] = 13
      "0001101" when "01100011001111001", -- t[50809] = 13
      "0001101" when "01100011001111010", -- t[50810] = 13
      "0001101" when "01100011001111011", -- t[50811] = 13
      "0001101" when "01100011001111100", -- t[50812] = 13
      "0001101" when "01100011001111101", -- t[50813] = 13
      "0001101" when "01100011001111110", -- t[50814] = 13
      "0001101" when "01100011001111111", -- t[50815] = 13
      "0001101" when "01100011010000000", -- t[50816] = 13
      "0001101" when "01100011010000001", -- t[50817] = 13
      "0001101" when "01100011010000010", -- t[50818] = 13
      "0001101" when "01100011010000011", -- t[50819] = 13
      "0001101" when "01100011010000100", -- t[50820] = 13
      "0001101" when "01100011010000101", -- t[50821] = 13
      "0001101" when "01100011010000110", -- t[50822] = 13
      "0001101" when "01100011010000111", -- t[50823] = 13
      "0001101" when "01100011010001000", -- t[50824] = 13
      "0001101" when "01100011010001001", -- t[50825] = 13
      "0001101" when "01100011010001010", -- t[50826] = 13
      "0001101" when "01100011010001011", -- t[50827] = 13
      "0001101" when "01100011010001100", -- t[50828] = 13
      "0001101" when "01100011010001101", -- t[50829] = 13
      "0001101" when "01100011010001110", -- t[50830] = 13
      "0001101" when "01100011010001111", -- t[50831] = 13
      "0001101" when "01100011010010000", -- t[50832] = 13
      "0001101" when "01100011010010001", -- t[50833] = 13
      "0001101" when "01100011010010010", -- t[50834] = 13
      "0001101" when "01100011010010011", -- t[50835] = 13
      "0001101" when "01100011010010100", -- t[50836] = 13
      "0001101" when "01100011010010101", -- t[50837] = 13
      "0001101" when "01100011010010110", -- t[50838] = 13
      "0001101" when "01100011010010111", -- t[50839] = 13
      "0001101" when "01100011010011000", -- t[50840] = 13
      "0001101" when "01100011010011001", -- t[50841] = 13
      "0001101" when "01100011010011010", -- t[50842] = 13
      "0001101" when "01100011010011011", -- t[50843] = 13
      "0001101" when "01100011010011100", -- t[50844] = 13
      "0001101" when "01100011010011101", -- t[50845] = 13
      "0001101" when "01100011010011110", -- t[50846] = 13
      "0001101" when "01100011010011111", -- t[50847] = 13
      "0001101" when "01100011010100000", -- t[50848] = 13
      "0001101" when "01100011010100001", -- t[50849] = 13
      "0001101" when "01100011010100010", -- t[50850] = 13
      "0001101" when "01100011010100011", -- t[50851] = 13
      "0001101" when "01100011010100100", -- t[50852] = 13
      "0001101" when "01100011010100101", -- t[50853] = 13
      "0001101" when "01100011010100110", -- t[50854] = 13
      "0001101" when "01100011010100111", -- t[50855] = 13
      "0001101" when "01100011010101000", -- t[50856] = 13
      "0001101" when "01100011010101001", -- t[50857] = 13
      "0001101" when "01100011010101010", -- t[50858] = 13
      "0001101" when "01100011010101011", -- t[50859] = 13
      "0001101" when "01100011010101100", -- t[50860] = 13
      "0001101" when "01100011010101101", -- t[50861] = 13
      "0001101" when "01100011010101110", -- t[50862] = 13
      "0001101" when "01100011010101111", -- t[50863] = 13
      "0001101" when "01100011010110000", -- t[50864] = 13
      "0001101" when "01100011010110001", -- t[50865] = 13
      "0001101" when "01100011010110010", -- t[50866] = 13
      "0001101" when "01100011010110011", -- t[50867] = 13
      "0001101" when "01100011010110100", -- t[50868] = 13
      "0001101" when "01100011010110101", -- t[50869] = 13
      "0001101" when "01100011010110110", -- t[50870] = 13
      "0001101" when "01100011010110111", -- t[50871] = 13
      "0001101" when "01100011010111000", -- t[50872] = 13
      "0001101" when "01100011010111001", -- t[50873] = 13
      "0001101" when "01100011010111010", -- t[50874] = 13
      "0001101" when "01100011010111011", -- t[50875] = 13
      "0001101" when "01100011010111100", -- t[50876] = 13
      "0001101" when "01100011010111101", -- t[50877] = 13
      "0001101" when "01100011010111110", -- t[50878] = 13
      "0001101" when "01100011010111111", -- t[50879] = 13
      "0001101" when "01100011011000000", -- t[50880] = 13
      "0001101" when "01100011011000001", -- t[50881] = 13
      "0001101" when "01100011011000010", -- t[50882] = 13
      "0001101" when "01100011011000011", -- t[50883] = 13
      "0001101" when "01100011011000100", -- t[50884] = 13
      "0001101" when "01100011011000101", -- t[50885] = 13
      "0001101" when "01100011011000110", -- t[50886] = 13
      "0001101" when "01100011011000111", -- t[50887] = 13
      "0001101" when "01100011011001000", -- t[50888] = 13
      "0001101" when "01100011011001001", -- t[50889] = 13
      "0001101" when "01100011011001010", -- t[50890] = 13
      "0001101" when "01100011011001011", -- t[50891] = 13
      "0001101" when "01100011011001100", -- t[50892] = 13
      "0001101" when "01100011011001101", -- t[50893] = 13
      "0001101" when "01100011011001110", -- t[50894] = 13
      "0001101" when "01100011011001111", -- t[50895] = 13
      "0001101" when "01100011011010000", -- t[50896] = 13
      "0001101" when "01100011011010001", -- t[50897] = 13
      "0001101" when "01100011011010010", -- t[50898] = 13
      "0001101" when "01100011011010011", -- t[50899] = 13
      "0001101" when "01100011011010100", -- t[50900] = 13
      "0001101" when "01100011011010101", -- t[50901] = 13
      "0001101" when "01100011011010110", -- t[50902] = 13
      "0001101" when "01100011011010111", -- t[50903] = 13
      "0001101" when "01100011011011000", -- t[50904] = 13
      "0001101" when "01100011011011001", -- t[50905] = 13
      "0001101" when "01100011011011010", -- t[50906] = 13
      "0001101" when "01100011011011011", -- t[50907] = 13
      "0001101" when "01100011011011100", -- t[50908] = 13
      "0001101" when "01100011011011101", -- t[50909] = 13
      "0001101" when "01100011011011110", -- t[50910] = 13
      "0001101" when "01100011011011111", -- t[50911] = 13
      "0001101" when "01100011011100000", -- t[50912] = 13
      "0001101" when "01100011011100001", -- t[50913] = 13
      "0001101" when "01100011011100010", -- t[50914] = 13
      "0001101" when "01100011011100011", -- t[50915] = 13
      "0001101" when "01100011011100100", -- t[50916] = 13
      "0001101" when "01100011011100101", -- t[50917] = 13
      "0001101" when "01100011011100110", -- t[50918] = 13
      "0001101" when "01100011011100111", -- t[50919] = 13
      "0001101" when "01100011011101000", -- t[50920] = 13
      "0001101" when "01100011011101001", -- t[50921] = 13
      "0001101" when "01100011011101010", -- t[50922] = 13
      "0001101" when "01100011011101011", -- t[50923] = 13
      "0001101" when "01100011011101100", -- t[50924] = 13
      "0001101" when "01100011011101101", -- t[50925] = 13
      "0001101" when "01100011011101110", -- t[50926] = 13
      "0001101" when "01100011011101111", -- t[50927] = 13
      "0001101" when "01100011011110000", -- t[50928] = 13
      "0001101" when "01100011011110001", -- t[50929] = 13
      "0001101" when "01100011011110010", -- t[50930] = 13
      "0001101" when "01100011011110011", -- t[50931] = 13
      "0001101" when "01100011011110100", -- t[50932] = 13
      "0001101" when "01100011011110101", -- t[50933] = 13
      "0001101" when "01100011011110110", -- t[50934] = 13
      "0001101" when "01100011011110111", -- t[50935] = 13
      "0001101" when "01100011011111000", -- t[50936] = 13
      "0001101" when "01100011011111001", -- t[50937] = 13
      "0001101" when "01100011011111010", -- t[50938] = 13
      "0001101" when "01100011011111011", -- t[50939] = 13
      "0001101" when "01100011011111100", -- t[50940] = 13
      "0001101" when "01100011011111101", -- t[50941] = 13
      "0001101" when "01100011011111110", -- t[50942] = 13
      "0001101" when "01100011011111111", -- t[50943] = 13
      "0001101" when "01100011100000000", -- t[50944] = 13
      "0001101" when "01100011100000001", -- t[50945] = 13
      "0001101" when "01100011100000010", -- t[50946] = 13
      "0001101" when "01100011100000011", -- t[50947] = 13
      "0001101" when "01100011100000100", -- t[50948] = 13
      "0001101" when "01100011100000101", -- t[50949] = 13
      "0001101" when "01100011100000110", -- t[50950] = 13
      "0001101" when "01100011100000111", -- t[50951] = 13
      "0001101" when "01100011100001000", -- t[50952] = 13
      "0001101" when "01100011100001001", -- t[50953] = 13
      "0001101" when "01100011100001010", -- t[50954] = 13
      "0001101" when "01100011100001011", -- t[50955] = 13
      "0001101" when "01100011100001100", -- t[50956] = 13
      "0001101" when "01100011100001101", -- t[50957] = 13
      "0001101" when "01100011100001110", -- t[50958] = 13
      "0001101" when "01100011100001111", -- t[50959] = 13
      "0001101" when "01100011100010000", -- t[50960] = 13
      "0001101" when "01100011100010001", -- t[50961] = 13
      "0001101" when "01100011100010010", -- t[50962] = 13
      "0001101" when "01100011100010011", -- t[50963] = 13
      "0001101" when "01100011100010100", -- t[50964] = 13
      "0001101" when "01100011100010101", -- t[50965] = 13
      "0001101" when "01100011100010110", -- t[50966] = 13
      "0001101" when "01100011100010111", -- t[50967] = 13
      "0001101" when "01100011100011000", -- t[50968] = 13
      "0001101" when "01100011100011001", -- t[50969] = 13
      "0001101" when "01100011100011010", -- t[50970] = 13
      "0001101" when "01100011100011011", -- t[50971] = 13
      "0001101" when "01100011100011100", -- t[50972] = 13
      "0001101" when "01100011100011101", -- t[50973] = 13
      "0001101" when "01100011100011110", -- t[50974] = 13
      "0001101" when "01100011100011111", -- t[50975] = 13
      "0001101" when "01100011100100000", -- t[50976] = 13
      "0001101" when "01100011100100001", -- t[50977] = 13
      "0001101" when "01100011100100010", -- t[50978] = 13
      "0001101" when "01100011100100011", -- t[50979] = 13
      "0001101" when "01100011100100100", -- t[50980] = 13
      "0001101" when "01100011100100101", -- t[50981] = 13
      "0001101" when "01100011100100110", -- t[50982] = 13
      "0001101" when "01100011100100111", -- t[50983] = 13
      "0001101" when "01100011100101000", -- t[50984] = 13
      "0001101" when "01100011100101001", -- t[50985] = 13
      "0001101" when "01100011100101010", -- t[50986] = 13
      "0001101" when "01100011100101011", -- t[50987] = 13
      "0001101" when "01100011100101100", -- t[50988] = 13
      "0001101" when "01100011100101101", -- t[50989] = 13
      "0001101" when "01100011100101110", -- t[50990] = 13
      "0001101" when "01100011100101111", -- t[50991] = 13
      "0001101" when "01100011100110000", -- t[50992] = 13
      "0001101" when "01100011100110001", -- t[50993] = 13
      "0001101" when "01100011100110010", -- t[50994] = 13
      "0001101" when "01100011100110011", -- t[50995] = 13
      "0001101" when "01100011100110100", -- t[50996] = 13
      "0001101" when "01100011100110101", -- t[50997] = 13
      "0001110" when "01100011100110110", -- t[50998] = 14
      "0001110" when "01100011100110111", -- t[50999] = 14
      "0001110" when "01100011100111000", -- t[51000] = 14
      "0001110" when "01100011100111001", -- t[51001] = 14
      "0001110" when "01100011100111010", -- t[51002] = 14
      "0001110" when "01100011100111011", -- t[51003] = 14
      "0001110" when "01100011100111100", -- t[51004] = 14
      "0001110" when "01100011100111101", -- t[51005] = 14
      "0001110" when "01100011100111110", -- t[51006] = 14
      "0001110" when "01100011100111111", -- t[51007] = 14
      "0001110" when "01100011101000000", -- t[51008] = 14
      "0001110" when "01100011101000001", -- t[51009] = 14
      "0001110" when "01100011101000010", -- t[51010] = 14
      "0001110" when "01100011101000011", -- t[51011] = 14
      "0001110" when "01100011101000100", -- t[51012] = 14
      "0001110" when "01100011101000101", -- t[51013] = 14
      "0001110" when "01100011101000110", -- t[51014] = 14
      "0001110" when "01100011101000111", -- t[51015] = 14
      "0001110" when "01100011101001000", -- t[51016] = 14
      "0001110" when "01100011101001001", -- t[51017] = 14
      "0001110" when "01100011101001010", -- t[51018] = 14
      "0001110" when "01100011101001011", -- t[51019] = 14
      "0001110" when "01100011101001100", -- t[51020] = 14
      "0001110" when "01100011101001101", -- t[51021] = 14
      "0001110" when "01100011101001110", -- t[51022] = 14
      "0001110" when "01100011101001111", -- t[51023] = 14
      "0001110" when "01100011101010000", -- t[51024] = 14
      "0001110" when "01100011101010001", -- t[51025] = 14
      "0001110" when "01100011101010010", -- t[51026] = 14
      "0001110" when "01100011101010011", -- t[51027] = 14
      "0001110" when "01100011101010100", -- t[51028] = 14
      "0001110" when "01100011101010101", -- t[51029] = 14
      "0001110" when "01100011101010110", -- t[51030] = 14
      "0001110" when "01100011101010111", -- t[51031] = 14
      "0001110" when "01100011101011000", -- t[51032] = 14
      "0001110" when "01100011101011001", -- t[51033] = 14
      "0001110" when "01100011101011010", -- t[51034] = 14
      "0001110" when "01100011101011011", -- t[51035] = 14
      "0001110" when "01100011101011100", -- t[51036] = 14
      "0001110" when "01100011101011101", -- t[51037] = 14
      "0001110" when "01100011101011110", -- t[51038] = 14
      "0001110" when "01100011101011111", -- t[51039] = 14
      "0001110" when "01100011101100000", -- t[51040] = 14
      "0001110" when "01100011101100001", -- t[51041] = 14
      "0001110" when "01100011101100010", -- t[51042] = 14
      "0001110" when "01100011101100011", -- t[51043] = 14
      "0001110" when "01100011101100100", -- t[51044] = 14
      "0001110" when "01100011101100101", -- t[51045] = 14
      "0001110" when "01100011101100110", -- t[51046] = 14
      "0001110" when "01100011101100111", -- t[51047] = 14
      "0001110" when "01100011101101000", -- t[51048] = 14
      "0001110" when "01100011101101001", -- t[51049] = 14
      "0001110" when "01100011101101010", -- t[51050] = 14
      "0001110" when "01100011101101011", -- t[51051] = 14
      "0001110" when "01100011101101100", -- t[51052] = 14
      "0001110" when "01100011101101101", -- t[51053] = 14
      "0001110" when "01100011101101110", -- t[51054] = 14
      "0001110" when "01100011101101111", -- t[51055] = 14
      "0001110" when "01100011101110000", -- t[51056] = 14
      "0001110" when "01100011101110001", -- t[51057] = 14
      "0001110" when "01100011101110010", -- t[51058] = 14
      "0001110" when "01100011101110011", -- t[51059] = 14
      "0001110" when "01100011101110100", -- t[51060] = 14
      "0001110" when "01100011101110101", -- t[51061] = 14
      "0001110" when "01100011101110110", -- t[51062] = 14
      "0001110" when "01100011101110111", -- t[51063] = 14
      "0001110" when "01100011101111000", -- t[51064] = 14
      "0001110" when "01100011101111001", -- t[51065] = 14
      "0001110" when "01100011101111010", -- t[51066] = 14
      "0001110" when "01100011101111011", -- t[51067] = 14
      "0001110" when "01100011101111100", -- t[51068] = 14
      "0001110" when "01100011101111101", -- t[51069] = 14
      "0001110" when "01100011101111110", -- t[51070] = 14
      "0001110" when "01100011101111111", -- t[51071] = 14
      "0001110" when "01100011110000000", -- t[51072] = 14
      "0001110" when "01100011110000001", -- t[51073] = 14
      "0001110" when "01100011110000010", -- t[51074] = 14
      "0001110" when "01100011110000011", -- t[51075] = 14
      "0001110" when "01100011110000100", -- t[51076] = 14
      "0001110" when "01100011110000101", -- t[51077] = 14
      "0001110" when "01100011110000110", -- t[51078] = 14
      "0001110" when "01100011110000111", -- t[51079] = 14
      "0001110" when "01100011110001000", -- t[51080] = 14
      "0001110" when "01100011110001001", -- t[51081] = 14
      "0001110" when "01100011110001010", -- t[51082] = 14
      "0001110" when "01100011110001011", -- t[51083] = 14
      "0001110" when "01100011110001100", -- t[51084] = 14
      "0001110" when "01100011110001101", -- t[51085] = 14
      "0001110" when "01100011110001110", -- t[51086] = 14
      "0001110" when "01100011110001111", -- t[51087] = 14
      "0001110" when "01100011110010000", -- t[51088] = 14
      "0001110" when "01100011110010001", -- t[51089] = 14
      "0001110" when "01100011110010010", -- t[51090] = 14
      "0001110" when "01100011110010011", -- t[51091] = 14
      "0001110" when "01100011110010100", -- t[51092] = 14
      "0001110" when "01100011110010101", -- t[51093] = 14
      "0001110" when "01100011110010110", -- t[51094] = 14
      "0001110" when "01100011110010111", -- t[51095] = 14
      "0001110" when "01100011110011000", -- t[51096] = 14
      "0001110" when "01100011110011001", -- t[51097] = 14
      "0001110" when "01100011110011010", -- t[51098] = 14
      "0001110" when "01100011110011011", -- t[51099] = 14
      "0001110" when "01100011110011100", -- t[51100] = 14
      "0001110" when "01100011110011101", -- t[51101] = 14
      "0001110" when "01100011110011110", -- t[51102] = 14
      "0001110" when "01100011110011111", -- t[51103] = 14
      "0001110" when "01100011110100000", -- t[51104] = 14
      "0001110" when "01100011110100001", -- t[51105] = 14
      "0001110" when "01100011110100010", -- t[51106] = 14
      "0001110" when "01100011110100011", -- t[51107] = 14
      "0001110" when "01100011110100100", -- t[51108] = 14
      "0001110" when "01100011110100101", -- t[51109] = 14
      "0001110" when "01100011110100110", -- t[51110] = 14
      "0001110" when "01100011110100111", -- t[51111] = 14
      "0001110" when "01100011110101000", -- t[51112] = 14
      "0001110" when "01100011110101001", -- t[51113] = 14
      "0001110" when "01100011110101010", -- t[51114] = 14
      "0001110" when "01100011110101011", -- t[51115] = 14
      "0001110" when "01100011110101100", -- t[51116] = 14
      "0001110" when "01100011110101101", -- t[51117] = 14
      "0001110" when "01100011110101110", -- t[51118] = 14
      "0001110" when "01100011110101111", -- t[51119] = 14
      "0001110" when "01100011110110000", -- t[51120] = 14
      "0001110" when "01100011110110001", -- t[51121] = 14
      "0001110" when "01100011110110010", -- t[51122] = 14
      "0001110" when "01100011110110011", -- t[51123] = 14
      "0001110" when "01100011110110100", -- t[51124] = 14
      "0001110" when "01100011110110101", -- t[51125] = 14
      "0001110" when "01100011110110110", -- t[51126] = 14
      "0001110" when "01100011110110111", -- t[51127] = 14
      "0001110" when "01100011110111000", -- t[51128] = 14
      "0001110" when "01100011110111001", -- t[51129] = 14
      "0001110" when "01100011110111010", -- t[51130] = 14
      "0001110" when "01100011110111011", -- t[51131] = 14
      "0001110" when "01100011110111100", -- t[51132] = 14
      "0001110" when "01100011110111101", -- t[51133] = 14
      "0001110" when "01100011110111110", -- t[51134] = 14
      "0001110" when "01100011110111111", -- t[51135] = 14
      "0001110" when "01100011111000000", -- t[51136] = 14
      "0001110" when "01100011111000001", -- t[51137] = 14
      "0001110" when "01100011111000010", -- t[51138] = 14
      "0001110" when "01100011111000011", -- t[51139] = 14
      "0001110" when "01100011111000100", -- t[51140] = 14
      "0001110" when "01100011111000101", -- t[51141] = 14
      "0001110" when "01100011111000110", -- t[51142] = 14
      "0001110" when "01100011111000111", -- t[51143] = 14
      "0001110" when "01100011111001000", -- t[51144] = 14
      "0001110" when "01100011111001001", -- t[51145] = 14
      "0001110" when "01100011111001010", -- t[51146] = 14
      "0001110" when "01100011111001011", -- t[51147] = 14
      "0001110" when "01100011111001100", -- t[51148] = 14
      "0001110" when "01100011111001101", -- t[51149] = 14
      "0001110" when "01100011111001110", -- t[51150] = 14
      "0001110" when "01100011111001111", -- t[51151] = 14
      "0001110" when "01100011111010000", -- t[51152] = 14
      "0001110" when "01100011111010001", -- t[51153] = 14
      "0001110" when "01100011111010010", -- t[51154] = 14
      "0001110" when "01100011111010011", -- t[51155] = 14
      "0001110" when "01100011111010100", -- t[51156] = 14
      "0001110" when "01100011111010101", -- t[51157] = 14
      "0001110" when "01100011111010110", -- t[51158] = 14
      "0001110" when "01100011111010111", -- t[51159] = 14
      "0001110" when "01100011111011000", -- t[51160] = 14
      "0001110" when "01100011111011001", -- t[51161] = 14
      "0001110" when "01100011111011010", -- t[51162] = 14
      "0001110" when "01100011111011011", -- t[51163] = 14
      "0001110" when "01100011111011100", -- t[51164] = 14
      "0001110" when "01100011111011101", -- t[51165] = 14
      "0001110" when "01100011111011110", -- t[51166] = 14
      "0001110" when "01100011111011111", -- t[51167] = 14
      "0001110" when "01100011111100000", -- t[51168] = 14
      "0001110" when "01100011111100001", -- t[51169] = 14
      "0001110" when "01100011111100010", -- t[51170] = 14
      "0001110" when "01100011111100011", -- t[51171] = 14
      "0001110" when "01100011111100100", -- t[51172] = 14
      "0001110" when "01100011111100101", -- t[51173] = 14
      "0001110" when "01100011111100110", -- t[51174] = 14
      "0001110" when "01100011111100111", -- t[51175] = 14
      "0001110" when "01100011111101000", -- t[51176] = 14
      "0001110" when "01100011111101001", -- t[51177] = 14
      "0001110" when "01100011111101010", -- t[51178] = 14
      "0001110" when "01100011111101011", -- t[51179] = 14
      "0001110" when "01100011111101100", -- t[51180] = 14
      "0001110" when "01100011111101101", -- t[51181] = 14
      "0001110" when "01100011111101110", -- t[51182] = 14
      "0001110" when "01100011111101111", -- t[51183] = 14
      "0001110" when "01100011111110000", -- t[51184] = 14
      "0001110" when "01100011111110001", -- t[51185] = 14
      "0001110" when "01100011111110010", -- t[51186] = 14
      "0001110" when "01100011111110011", -- t[51187] = 14
      "0001110" when "01100011111110100", -- t[51188] = 14
      "0001110" when "01100011111110101", -- t[51189] = 14
      "0001110" when "01100011111110110", -- t[51190] = 14
      "0001110" when "01100011111110111", -- t[51191] = 14
      "0001110" when "01100011111111000", -- t[51192] = 14
      "0001110" when "01100011111111001", -- t[51193] = 14
      "0001110" when "01100011111111010", -- t[51194] = 14
      "0001110" when "01100011111111011", -- t[51195] = 14
      "0001110" when "01100011111111100", -- t[51196] = 14
      "0001110" when "01100011111111101", -- t[51197] = 14
      "0001110" when "01100011111111110", -- t[51198] = 14
      "0001110" when "01100011111111111", -- t[51199] = 14
      "0001110" when "01100100000000000", -- t[51200] = 14
      "0001110" when "01100100000000001", -- t[51201] = 14
      "0001110" when "01100100000000010", -- t[51202] = 14
      "0001110" when "01100100000000011", -- t[51203] = 14
      "0001110" when "01100100000000100", -- t[51204] = 14
      "0001110" when "01100100000000101", -- t[51205] = 14
      "0001110" when "01100100000000110", -- t[51206] = 14
      "0001110" when "01100100000000111", -- t[51207] = 14
      "0001110" when "01100100000001000", -- t[51208] = 14
      "0001110" when "01100100000001001", -- t[51209] = 14
      "0001110" when "01100100000001010", -- t[51210] = 14
      "0001110" when "01100100000001011", -- t[51211] = 14
      "0001110" when "01100100000001100", -- t[51212] = 14
      "0001110" when "01100100000001101", -- t[51213] = 14
      "0001110" when "01100100000001110", -- t[51214] = 14
      "0001110" when "01100100000001111", -- t[51215] = 14
      "0001110" when "01100100000010000", -- t[51216] = 14
      "0001110" when "01100100000010001", -- t[51217] = 14
      "0001110" when "01100100000010010", -- t[51218] = 14
      "0001110" when "01100100000010011", -- t[51219] = 14
      "0001110" when "01100100000010100", -- t[51220] = 14
      "0001110" when "01100100000010101", -- t[51221] = 14
      "0001110" when "01100100000010110", -- t[51222] = 14
      "0001110" when "01100100000010111", -- t[51223] = 14
      "0001110" when "01100100000011000", -- t[51224] = 14
      "0001110" when "01100100000011001", -- t[51225] = 14
      "0001110" when "01100100000011010", -- t[51226] = 14
      "0001110" when "01100100000011011", -- t[51227] = 14
      "0001110" when "01100100000011100", -- t[51228] = 14
      "0001110" when "01100100000011101", -- t[51229] = 14
      "0001110" when "01100100000011110", -- t[51230] = 14
      "0001110" when "01100100000011111", -- t[51231] = 14
      "0001110" when "01100100000100000", -- t[51232] = 14
      "0001110" when "01100100000100001", -- t[51233] = 14
      "0001110" when "01100100000100010", -- t[51234] = 14
      "0001110" when "01100100000100011", -- t[51235] = 14
      "0001110" when "01100100000100100", -- t[51236] = 14
      "0001110" when "01100100000100101", -- t[51237] = 14
      "0001110" when "01100100000100110", -- t[51238] = 14
      "0001110" when "01100100000100111", -- t[51239] = 14
      "0001110" when "01100100000101000", -- t[51240] = 14
      "0001110" when "01100100000101001", -- t[51241] = 14
      "0001110" when "01100100000101010", -- t[51242] = 14
      "0001110" when "01100100000101011", -- t[51243] = 14
      "0001110" when "01100100000101100", -- t[51244] = 14
      "0001110" when "01100100000101101", -- t[51245] = 14
      "0001110" when "01100100000101110", -- t[51246] = 14
      "0001110" when "01100100000101111", -- t[51247] = 14
      "0001110" when "01100100000110000", -- t[51248] = 14
      "0001110" when "01100100000110001", -- t[51249] = 14
      "0001110" when "01100100000110010", -- t[51250] = 14
      "0001110" when "01100100000110011", -- t[51251] = 14
      "0001110" when "01100100000110100", -- t[51252] = 14
      "0001110" when "01100100000110101", -- t[51253] = 14
      "0001110" when "01100100000110110", -- t[51254] = 14
      "0001110" when "01100100000110111", -- t[51255] = 14
      "0001110" when "01100100000111000", -- t[51256] = 14
      "0001110" when "01100100000111001", -- t[51257] = 14
      "0001110" when "01100100000111010", -- t[51258] = 14
      "0001110" when "01100100000111011", -- t[51259] = 14
      "0001110" when "01100100000111100", -- t[51260] = 14
      "0001110" when "01100100000111101", -- t[51261] = 14
      "0001110" when "01100100000111110", -- t[51262] = 14
      "0001110" when "01100100000111111", -- t[51263] = 14
      "0001110" when "01100100001000000", -- t[51264] = 14
      "0001110" when "01100100001000001", -- t[51265] = 14
      "0001110" when "01100100001000010", -- t[51266] = 14
      "0001110" when "01100100001000011", -- t[51267] = 14
      "0001110" when "01100100001000100", -- t[51268] = 14
      "0001110" when "01100100001000101", -- t[51269] = 14
      "0001110" when "01100100001000110", -- t[51270] = 14
      "0001110" when "01100100001000111", -- t[51271] = 14
      "0001110" when "01100100001001000", -- t[51272] = 14
      "0001110" when "01100100001001001", -- t[51273] = 14
      "0001110" when "01100100001001010", -- t[51274] = 14
      "0001110" when "01100100001001011", -- t[51275] = 14
      "0001110" when "01100100001001100", -- t[51276] = 14
      "0001110" when "01100100001001101", -- t[51277] = 14
      "0001110" when "01100100001001110", -- t[51278] = 14
      "0001110" when "01100100001001111", -- t[51279] = 14
      "0001110" when "01100100001010000", -- t[51280] = 14
      "0001110" when "01100100001010001", -- t[51281] = 14
      "0001110" when "01100100001010010", -- t[51282] = 14
      "0001110" when "01100100001010011", -- t[51283] = 14
      "0001110" when "01100100001010100", -- t[51284] = 14
      "0001110" when "01100100001010101", -- t[51285] = 14
      "0001110" when "01100100001010110", -- t[51286] = 14
      "0001110" when "01100100001010111", -- t[51287] = 14
      "0001110" when "01100100001011000", -- t[51288] = 14
      "0001110" when "01100100001011001", -- t[51289] = 14
      "0001110" when "01100100001011010", -- t[51290] = 14
      "0001110" when "01100100001011011", -- t[51291] = 14
      "0001110" when "01100100001011100", -- t[51292] = 14
      "0001110" when "01100100001011101", -- t[51293] = 14
      "0001110" when "01100100001011110", -- t[51294] = 14
      "0001110" when "01100100001011111", -- t[51295] = 14
      "0001110" when "01100100001100000", -- t[51296] = 14
      "0001110" when "01100100001100001", -- t[51297] = 14
      "0001110" when "01100100001100010", -- t[51298] = 14
      "0001110" when "01100100001100011", -- t[51299] = 14
      "0001110" when "01100100001100100", -- t[51300] = 14
      "0001110" when "01100100001100101", -- t[51301] = 14
      "0001110" when "01100100001100110", -- t[51302] = 14
      "0001110" when "01100100001100111", -- t[51303] = 14
      "0001110" when "01100100001101000", -- t[51304] = 14
      "0001110" when "01100100001101001", -- t[51305] = 14
      "0001110" when "01100100001101010", -- t[51306] = 14
      "0001110" when "01100100001101011", -- t[51307] = 14
      "0001110" when "01100100001101100", -- t[51308] = 14
      "0001110" when "01100100001101101", -- t[51309] = 14
      "0001110" when "01100100001101110", -- t[51310] = 14
      "0001110" when "01100100001101111", -- t[51311] = 14
      "0001110" when "01100100001110000", -- t[51312] = 14
      "0001110" when "01100100001110001", -- t[51313] = 14
      "0001110" when "01100100001110010", -- t[51314] = 14
      "0001110" when "01100100001110011", -- t[51315] = 14
      "0001110" when "01100100001110100", -- t[51316] = 14
      "0001110" when "01100100001110101", -- t[51317] = 14
      "0001110" when "01100100001110110", -- t[51318] = 14
      "0001110" when "01100100001110111", -- t[51319] = 14
      "0001110" when "01100100001111000", -- t[51320] = 14
      "0001110" when "01100100001111001", -- t[51321] = 14
      "0001110" when "01100100001111010", -- t[51322] = 14
      "0001110" when "01100100001111011", -- t[51323] = 14
      "0001110" when "01100100001111100", -- t[51324] = 14
      "0001110" when "01100100001111101", -- t[51325] = 14
      "0001110" when "01100100001111110", -- t[51326] = 14
      "0001110" when "01100100001111111", -- t[51327] = 14
      "0001110" when "01100100010000000", -- t[51328] = 14
      "0001110" when "01100100010000001", -- t[51329] = 14
      "0001110" when "01100100010000010", -- t[51330] = 14
      "0001110" when "01100100010000011", -- t[51331] = 14
      "0001110" when "01100100010000100", -- t[51332] = 14
      "0001110" when "01100100010000101", -- t[51333] = 14
      "0001110" when "01100100010000110", -- t[51334] = 14
      "0001110" when "01100100010000111", -- t[51335] = 14
      "0001110" when "01100100010001000", -- t[51336] = 14
      "0001110" when "01100100010001001", -- t[51337] = 14
      "0001110" when "01100100010001010", -- t[51338] = 14
      "0001110" when "01100100010001011", -- t[51339] = 14
      "0001110" when "01100100010001100", -- t[51340] = 14
      "0001110" when "01100100010001101", -- t[51341] = 14
      "0001110" when "01100100010001110", -- t[51342] = 14
      "0001110" when "01100100010001111", -- t[51343] = 14
      "0001110" when "01100100010010000", -- t[51344] = 14
      "0001110" when "01100100010010001", -- t[51345] = 14
      "0001110" when "01100100010010010", -- t[51346] = 14
      "0001110" when "01100100010010011", -- t[51347] = 14
      "0001110" when "01100100010010100", -- t[51348] = 14
      "0001110" when "01100100010010101", -- t[51349] = 14
      "0001110" when "01100100010010110", -- t[51350] = 14
      "0001110" when "01100100010010111", -- t[51351] = 14
      "0001110" when "01100100010011000", -- t[51352] = 14
      "0001110" when "01100100010011001", -- t[51353] = 14
      "0001110" when "01100100010011010", -- t[51354] = 14
      "0001110" when "01100100010011011", -- t[51355] = 14
      "0001110" when "01100100010011100", -- t[51356] = 14
      "0001110" when "01100100010011101", -- t[51357] = 14
      "0001110" when "01100100010011110", -- t[51358] = 14
      "0001110" when "01100100010011111", -- t[51359] = 14
      "0001110" when "01100100010100000", -- t[51360] = 14
      "0001110" when "01100100010100001", -- t[51361] = 14
      "0001110" when "01100100010100010", -- t[51362] = 14
      "0001110" when "01100100010100011", -- t[51363] = 14
      "0001110" when "01100100010100100", -- t[51364] = 14
      "0001110" when "01100100010100101", -- t[51365] = 14
      "0001110" when "01100100010100110", -- t[51366] = 14
      "0001110" when "01100100010100111", -- t[51367] = 14
      "0001110" when "01100100010101000", -- t[51368] = 14
      "0001110" when "01100100010101001", -- t[51369] = 14
      "0001110" when "01100100010101010", -- t[51370] = 14
      "0001110" when "01100100010101011", -- t[51371] = 14
      "0001110" when "01100100010101100", -- t[51372] = 14
      "0001110" when "01100100010101101", -- t[51373] = 14
      "0001110" when "01100100010101110", -- t[51374] = 14
      "0001110" when "01100100010101111", -- t[51375] = 14
      "0001110" when "01100100010110000", -- t[51376] = 14
      "0001110" when "01100100010110001", -- t[51377] = 14
      "0001110" when "01100100010110010", -- t[51378] = 14
      "0001110" when "01100100010110011", -- t[51379] = 14
      "0001110" when "01100100010110100", -- t[51380] = 14
      "0001110" when "01100100010110101", -- t[51381] = 14
      "0001110" when "01100100010110110", -- t[51382] = 14
      "0001110" when "01100100010110111", -- t[51383] = 14
      "0001110" when "01100100010111000", -- t[51384] = 14
      "0001110" when "01100100010111001", -- t[51385] = 14
      "0001110" when "01100100010111010", -- t[51386] = 14
      "0001110" when "01100100010111011", -- t[51387] = 14
      "0001110" when "01100100010111100", -- t[51388] = 14
      "0001110" when "01100100010111101", -- t[51389] = 14
      "0001110" when "01100100010111110", -- t[51390] = 14
      "0001110" when "01100100010111111", -- t[51391] = 14
      "0001110" when "01100100011000000", -- t[51392] = 14
      "0001110" when "01100100011000001", -- t[51393] = 14
      "0001110" when "01100100011000010", -- t[51394] = 14
      "0001110" when "01100100011000011", -- t[51395] = 14
      "0001110" when "01100100011000100", -- t[51396] = 14
      "0001110" when "01100100011000101", -- t[51397] = 14
      "0001110" when "01100100011000110", -- t[51398] = 14
      "0001110" when "01100100011000111", -- t[51399] = 14
      "0001110" when "01100100011001000", -- t[51400] = 14
      "0001110" when "01100100011001001", -- t[51401] = 14
      "0001110" when "01100100011001010", -- t[51402] = 14
      "0001110" when "01100100011001011", -- t[51403] = 14
      "0001110" when "01100100011001100", -- t[51404] = 14
      "0001110" when "01100100011001101", -- t[51405] = 14
      "0001110" when "01100100011001110", -- t[51406] = 14
      "0001110" when "01100100011001111", -- t[51407] = 14
      "0001110" when "01100100011010000", -- t[51408] = 14
      "0001110" when "01100100011010001", -- t[51409] = 14
      "0001110" when "01100100011010010", -- t[51410] = 14
      "0001110" when "01100100011010011", -- t[51411] = 14
      "0001110" when "01100100011010100", -- t[51412] = 14
      "0001110" when "01100100011010101", -- t[51413] = 14
      "0001110" when "01100100011010110", -- t[51414] = 14
      "0001110" when "01100100011010111", -- t[51415] = 14
      "0001110" when "01100100011011000", -- t[51416] = 14
      "0001110" when "01100100011011001", -- t[51417] = 14
      "0001110" when "01100100011011010", -- t[51418] = 14
      "0001110" when "01100100011011011", -- t[51419] = 14
      "0001110" when "01100100011011100", -- t[51420] = 14
      "0001110" when "01100100011011101", -- t[51421] = 14
      "0001110" when "01100100011011110", -- t[51422] = 14
      "0001110" when "01100100011011111", -- t[51423] = 14
      "0001110" when "01100100011100000", -- t[51424] = 14
      "0001110" when "01100100011100001", -- t[51425] = 14
      "0001110" when "01100100011100010", -- t[51426] = 14
      "0001110" when "01100100011100011", -- t[51427] = 14
      "0001110" when "01100100011100100", -- t[51428] = 14
      "0001110" when "01100100011100101", -- t[51429] = 14
      "0001110" when "01100100011100110", -- t[51430] = 14
      "0001110" when "01100100011100111", -- t[51431] = 14
      "0001110" when "01100100011101000", -- t[51432] = 14
      "0001110" when "01100100011101001", -- t[51433] = 14
      "0001110" when "01100100011101010", -- t[51434] = 14
      "0001110" when "01100100011101011", -- t[51435] = 14
      "0001110" when "01100100011101100", -- t[51436] = 14
      "0001110" when "01100100011101101", -- t[51437] = 14
      "0001110" when "01100100011101110", -- t[51438] = 14
      "0001110" when "01100100011101111", -- t[51439] = 14
      "0001110" when "01100100011110000", -- t[51440] = 14
      "0001110" when "01100100011110001", -- t[51441] = 14
      "0001110" when "01100100011110010", -- t[51442] = 14
      "0001110" when "01100100011110011", -- t[51443] = 14
      "0001110" when "01100100011110100", -- t[51444] = 14
      "0001110" when "01100100011110101", -- t[51445] = 14
      "0001110" when "01100100011110110", -- t[51446] = 14
      "0001110" when "01100100011110111", -- t[51447] = 14
      "0001110" when "01100100011111000", -- t[51448] = 14
      "0001110" when "01100100011111001", -- t[51449] = 14
      "0001110" when "01100100011111010", -- t[51450] = 14
      "0001110" when "01100100011111011", -- t[51451] = 14
      "0001110" when "01100100011111100", -- t[51452] = 14
      "0001110" when "01100100011111101", -- t[51453] = 14
      "0001110" when "01100100011111110", -- t[51454] = 14
      "0001110" when "01100100011111111", -- t[51455] = 14
      "0001110" when "01100100100000000", -- t[51456] = 14
      "0001110" when "01100100100000001", -- t[51457] = 14
      "0001110" when "01100100100000010", -- t[51458] = 14
      "0001110" when "01100100100000011", -- t[51459] = 14
      "0001110" when "01100100100000100", -- t[51460] = 14
      "0001110" when "01100100100000101", -- t[51461] = 14
      "0001110" when "01100100100000110", -- t[51462] = 14
      "0001110" when "01100100100000111", -- t[51463] = 14
      "0001110" when "01100100100001000", -- t[51464] = 14
      "0001110" when "01100100100001001", -- t[51465] = 14
      "0001110" when "01100100100001010", -- t[51466] = 14
      "0001110" when "01100100100001011", -- t[51467] = 14
      "0001110" when "01100100100001100", -- t[51468] = 14
      "0001110" when "01100100100001101", -- t[51469] = 14
      "0001110" when "01100100100001110", -- t[51470] = 14
      "0001110" when "01100100100001111", -- t[51471] = 14
      "0001110" when "01100100100010000", -- t[51472] = 14
      "0001110" when "01100100100010001", -- t[51473] = 14
      "0001110" when "01100100100010010", -- t[51474] = 14
      "0001110" when "01100100100010011", -- t[51475] = 14
      "0001110" when "01100100100010100", -- t[51476] = 14
      "0001110" when "01100100100010101", -- t[51477] = 14
      "0001110" when "01100100100010110", -- t[51478] = 14
      "0001110" when "01100100100010111", -- t[51479] = 14
      "0001110" when "01100100100011000", -- t[51480] = 14
      "0001110" when "01100100100011001", -- t[51481] = 14
      "0001110" when "01100100100011010", -- t[51482] = 14
      "0001110" when "01100100100011011", -- t[51483] = 14
      "0001110" when "01100100100011100", -- t[51484] = 14
      "0001110" when "01100100100011101", -- t[51485] = 14
      "0001110" when "01100100100011110", -- t[51486] = 14
      "0001110" when "01100100100011111", -- t[51487] = 14
      "0001110" when "01100100100100000", -- t[51488] = 14
      "0001110" when "01100100100100001", -- t[51489] = 14
      "0001110" when "01100100100100010", -- t[51490] = 14
      "0001110" when "01100100100100011", -- t[51491] = 14
      "0001110" when "01100100100100100", -- t[51492] = 14
      "0001110" when "01100100100100101", -- t[51493] = 14
      "0001110" when "01100100100100110", -- t[51494] = 14
      "0001110" when "01100100100100111", -- t[51495] = 14
      "0001110" when "01100100100101000", -- t[51496] = 14
      "0001110" when "01100100100101001", -- t[51497] = 14
      "0001110" when "01100100100101010", -- t[51498] = 14
      "0001110" when "01100100100101011", -- t[51499] = 14
      "0001110" when "01100100100101100", -- t[51500] = 14
      "0001110" when "01100100100101101", -- t[51501] = 14
      "0001110" when "01100100100101110", -- t[51502] = 14
      "0001110" when "01100100100101111", -- t[51503] = 14
      "0001110" when "01100100100110000", -- t[51504] = 14
      "0001110" when "01100100100110001", -- t[51505] = 14
      "0001110" when "01100100100110010", -- t[51506] = 14
      "0001110" when "01100100100110011", -- t[51507] = 14
      "0001110" when "01100100100110100", -- t[51508] = 14
      "0001110" when "01100100100110101", -- t[51509] = 14
      "0001110" when "01100100100110110", -- t[51510] = 14
      "0001110" when "01100100100110111", -- t[51511] = 14
      "0001110" when "01100100100111000", -- t[51512] = 14
      "0001110" when "01100100100111001", -- t[51513] = 14
      "0001110" when "01100100100111010", -- t[51514] = 14
      "0001110" when "01100100100111011", -- t[51515] = 14
      "0001110" when "01100100100111100", -- t[51516] = 14
      "0001110" when "01100100100111101", -- t[51517] = 14
      "0001110" when "01100100100111110", -- t[51518] = 14
      "0001110" when "01100100100111111", -- t[51519] = 14
      "0001110" when "01100100101000000", -- t[51520] = 14
      "0001110" when "01100100101000001", -- t[51521] = 14
      "0001110" when "01100100101000010", -- t[51522] = 14
      "0001110" when "01100100101000011", -- t[51523] = 14
      "0001110" when "01100100101000100", -- t[51524] = 14
      "0001110" when "01100100101000101", -- t[51525] = 14
      "0001110" when "01100100101000110", -- t[51526] = 14
      "0001110" when "01100100101000111", -- t[51527] = 14
      "0001110" when "01100100101001000", -- t[51528] = 14
      "0001110" when "01100100101001001", -- t[51529] = 14
      "0001110" when "01100100101001010", -- t[51530] = 14
      "0001110" when "01100100101001011", -- t[51531] = 14
      "0001110" when "01100100101001100", -- t[51532] = 14
      "0001110" when "01100100101001101", -- t[51533] = 14
      "0001110" when "01100100101001110", -- t[51534] = 14
      "0001110" when "01100100101001111", -- t[51535] = 14
      "0001110" when "01100100101010000", -- t[51536] = 14
      "0001110" when "01100100101010001", -- t[51537] = 14
      "0001110" when "01100100101010010", -- t[51538] = 14
      "0001110" when "01100100101010011", -- t[51539] = 14
      "0001110" when "01100100101010100", -- t[51540] = 14
      "0001110" when "01100100101010101", -- t[51541] = 14
      "0001110" when "01100100101010110", -- t[51542] = 14
      "0001110" when "01100100101010111", -- t[51543] = 14
      "0001110" when "01100100101011000", -- t[51544] = 14
      "0001110" when "01100100101011001", -- t[51545] = 14
      "0001110" when "01100100101011010", -- t[51546] = 14
      "0001110" when "01100100101011011", -- t[51547] = 14
      "0001110" when "01100100101011100", -- t[51548] = 14
      "0001110" when "01100100101011101", -- t[51549] = 14
      "0001110" when "01100100101011110", -- t[51550] = 14
      "0001110" when "01100100101011111", -- t[51551] = 14
      "0001110" when "01100100101100000", -- t[51552] = 14
      "0001110" when "01100100101100001", -- t[51553] = 14
      "0001110" when "01100100101100010", -- t[51554] = 14
      "0001110" when "01100100101100011", -- t[51555] = 14
      "0001110" when "01100100101100100", -- t[51556] = 14
      "0001110" when "01100100101100101", -- t[51557] = 14
      "0001110" when "01100100101100110", -- t[51558] = 14
      "0001110" when "01100100101100111", -- t[51559] = 14
      "0001110" when "01100100101101000", -- t[51560] = 14
      "0001110" when "01100100101101001", -- t[51561] = 14
      "0001110" when "01100100101101010", -- t[51562] = 14
      "0001110" when "01100100101101011", -- t[51563] = 14
      "0001110" when "01100100101101100", -- t[51564] = 14
      "0001110" when "01100100101101101", -- t[51565] = 14
      "0001110" when "01100100101101110", -- t[51566] = 14
      "0001110" when "01100100101101111", -- t[51567] = 14
      "0001110" when "01100100101110000", -- t[51568] = 14
      "0001110" when "01100100101110001", -- t[51569] = 14
      "0001110" when "01100100101110010", -- t[51570] = 14
      "0001110" when "01100100101110011", -- t[51571] = 14
      "0001110" when "01100100101110100", -- t[51572] = 14
      "0001110" when "01100100101110101", -- t[51573] = 14
      "0001110" when "01100100101110110", -- t[51574] = 14
      "0001110" when "01100100101110111", -- t[51575] = 14
      "0001110" when "01100100101111000", -- t[51576] = 14
      "0001110" when "01100100101111001", -- t[51577] = 14
      "0001110" when "01100100101111010", -- t[51578] = 14
      "0001110" when "01100100101111011", -- t[51579] = 14
      "0001110" when "01100100101111100", -- t[51580] = 14
      "0001110" when "01100100101111101", -- t[51581] = 14
      "0001110" when "01100100101111110", -- t[51582] = 14
      "0001110" when "01100100101111111", -- t[51583] = 14
      "0001110" when "01100100110000000", -- t[51584] = 14
      "0001110" when "01100100110000001", -- t[51585] = 14
      "0001110" when "01100100110000010", -- t[51586] = 14
      "0001110" when "01100100110000011", -- t[51587] = 14
      "0001110" when "01100100110000100", -- t[51588] = 14
      "0001110" when "01100100110000101", -- t[51589] = 14
      "0001110" when "01100100110000110", -- t[51590] = 14
      "0001110" when "01100100110000111", -- t[51591] = 14
      "0001110" when "01100100110001000", -- t[51592] = 14
      "0001110" when "01100100110001001", -- t[51593] = 14
      "0001110" when "01100100110001010", -- t[51594] = 14
      "0001110" when "01100100110001011", -- t[51595] = 14
      "0001110" when "01100100110001100", -- t[51596] = 14
      "0001110" when "01100100110001101", -- t[51597] = 14
      "0001110" when "01100100110001110", -- t[51598] = 14
      "0001110" when "01100100110001111", -- t[51599] = 14
      "0001110" when "01100100110010000", -- t[51600] = 14
      "0001110" when "01100100110010001", -- t[51601] = 14
      "0001110" when "01100100110010010", -- t[51602] = 14
      "0001110" when "01100100110010011", -- t[51603] = 14
      "0001110" when "01100100110010100", -- t[51604] = 14
      "0001110" when "01100100110010101", -- t[51605] = 14
      "0001110" when "01100100110010110", -- t[51606] = 14
      "0001110" when "01100100110010111", -- t[51607] = 14
      "0001110" when "01100100110011000", -- t[51608] = 14
      "0001110" when "01100100110011001", -- t[51609] = 14
      "0001110" when "01100100110011010", -- t[51610] = 14
      "0001110" when "01100100110011011", -- t[51611] = 14
      "0001110" when "01100100110011100", -- t[51612] = 14
      "0001110" when "01100100110011101", -- t[51613] = 14
      "0001110" when "01100100110011110", -- t[51614] = 14
      "0001110" when "01100100110011111", -- t[51615] = 14
      "0001110" when "01100100110100000", -- t[51616] = 14
      "0001110" when "01100100110100001", -- t[51617] = 14
      "0001110" when "01100100110100010", -- t[51618] = 14
      "0001110" when "01100100110100011", -- t[51619] = 14
      "0001110" when "01100100110100100", -- t[51620] = 14
      "0001110" when "01100100110100101", -- t[51621] = 14
      "0001110" when "01100100110100110", -- t[51622] = 14
      "0001110" when "01100100110100111", -- t[51623] = 14
      "0001110" when "01100100110101000", -- t[51624] = 14
      "0001110" when "01100100110101001", -- t[51625] = 14
      "0001110" when "01100100110101010", -- t[51626] = 14
      "0001110" when "01100100110101011", -- t[51627] = 14
      "0001110" when "01100100110101100", -- t[51628] = 14
      "0001110" when "01100100110101101", -- t[51629] = 14
      "0001110" when "01100100110101110", -- t[51630] = 14
      "0001110" when "01100100110101111", -- t[51631] = 14
      "0001110" when "01100100110110000", -- t[51632] = 14
      "0001110" when "01100100110110001", -- t[51633] = 14
      "0001110" when "01100100110110010", -- t[51634] = 14
      "0001110" when "01100100110110011", -- t[51635] = 14
      "0001110" when "01100100110110100", -- t[51636] = 14
      "0001110" when "01100100110110101", -- t[51637] = 14
      "0001110" when "01100100110110110", -- t[51638] = 14
      "0001110" when "01100100110110111", -- t[51639] = 14
      "0001110" when "01100100110111000", -- t[51640] = 14
      "0001110" when "01100100110111001", -- t[51641] = 14
      "0001110" when "01100100110111010", -- t[51642] = 14
      "0001110" when "01100100110111011", -- t[51643] = 14
      "0001110" when "01100100110111100", -- t[51644] = 14
      "0001110" when "01100100110111101", -- t[51645] = 14
      "0001110" when "01100100110111110", -- t[51646] = 14
      "0001110" when "01100100110111111", -- t[51647] = 14
      "0001110" when "01100100111000000", -- t[51648] = 14
      "0001110" when "01100100111000001", -- t[51649] = 14
      "0001110" when "01100100111000010", -- t[51650] = 14
      "0001110" when "01100100111000011", -- t[51651] = 14
      "0001110" when "01100100111000100", -- t[51652] = 14
      "0001110" when "01100100111000101", -- t[51653] = 14
      "0001110" when "01100100111000110", -- t[51654] = 14
      "0001110" when "01100100111000111", -- t[51655] = 14
      "0001110" when "01100100111001000", -- t[51656] = 14
      "0001110" when "01100100111001001", -- t[51657] = 14
      "0001110" when "01100100111001010", -- t[51658] = 14
      "0001110" when "01100100111001011", -- t[51659] = 14
      "0001110" when "01100100111001100", -- t[51660] = 14
      "0001110" when "01100100111001101", -- t[51661] = 14
      "0001110" when "01100100111001110", -- t[51662] = 14
      "0001110" when "01100100111001111", -- t[51663] = 14
      "0001110" when "01100100111010000", -- t[51664] = 14
      "0001110" when "01100100111010001", -- t[51665] = 14
      "0001110" when "01100100111010010", -- t[51666] = 14
      "0001110" when "01100100111010011", -- t[51667] = 14
      "0001110" when "01100100111010100", -- t[51668] = 14
      "0001110" when "01100100111010101", -- t[51669] = 14
      "0001110" when "01100100111010110", -- t[51670] = 14
      "0001110" when "01100100111010111", -- t[51671] = 14
      "0001110" when "01100100111011000", -- t[51672] = 14
      "0001110" when "01100100111011001", -- t[51673] = 14
      "0001110" when "01100100111011010", -- t[51674] = 14
      "0001110" when "01100100111011011", -- t[51675] = 14
      "0001110" when "01100100111011100", -- t[51676] = 14
      "0001110" when "01100100111011101", -- t[51677] = 14
      "0001110" when "01100100111011110", -- t[51678] = 14
      "0001110" when "01100100111011111", -- t[51679] = 14
      "0001110" when "01100100111100000", -- t[51680] = 14
      "0001110" when "01100100111100001", -- t[51681] = 14
      "0001110" when "01100100111100010", -- t[51682] = 14
      "0001110" when "01100100111100011", -- t[51683] = 14
      "0001110" when "01100100111100100", -- t[51684] = 14
      "0001110" when "01100100111100101", -- t[51685] = 14
      "0001110" when "01100100111100110", -- t[51686] = 14
      "0001110" when "01100100111100111", -- t[51687] = 14
      "0001110" when "01100100111101000", -- t[51688] = 14
      "0001110" when "01100100111101001", -- t[51689] = 14
      "0001110" when "01100100111101010", -- t[51690] = 14
      "0001110" when "01100100111101011", -- t[51691] = 14
      "0001110" when "01100100111101100", -- t[51692] = 14
      "0001110" when "01100100111101101", -- t[51693] = 14
      "0001110" when "01100100111101110", -- t[51694] = 14
      "0001110" when "01100100111101111", -- t[51695] = 14
      "0001110" when "01100100111110000", -- t[51696] = 14
      "0001110" when "01100100111110001", -- t[51697] = 14
      "0001110" when "01100100111110010", -- t[51698] = 14
      "0001110" when "01100100111110011", -- t[51699] = 14
      "0001110" when "01100100111110100", -- t[51700] = 14
      "0001110" when "01100100111110101", -- t[51701] = 14
      "0001110" when "01100100111110110", -- t[51702] = 14
      "0001110" when "01100100111110111", -- t[51703] = 14
      "0001110" when "01100100111111000", -- t[51704] = 14
      "0001110" when "01100100111111001", -- t[51705] = 14
      "0001110" when "01100100111111010", -- t[51706] = 14
      "0001110" when "01100100111111011", -- t[51707] = 14
      "0001110" when "01100100111111100", -- t[51708] = 14
      "0001110" when "01100100111111101", -- t[51709] = 14
      "0001110" when "01100100111111110", -- t[51710] = 14
      "0001110" when "01100100111111111", -- t[51711] = 14
      "0001110" when "01100101000000000", -- t[51712] = 14
      "0001110" when "01100101000000001", -- t[51713] = 14
      "0001110" when "01100101000000010", -- t[51714] = 14
      "0001110" when "01100101000000011", -- t[51715] = 14
      "0001110" when "01100101000000100", -- t[51716] = 14
      "0001110" when "01100101000000101", -- t[51717] = 14
      "0001110" when "01100101000000110", -- t[51718] = 14
      "0001110" when "01100101000000111", -- t[51719] = 14
      "0001110" when "01100101000001000", -- t[51720] = 14
      "0001110" when "01100101000001001", -- t[51721] = 14
      "0001110" when "01100101000001010", -- t[51722] = 14
      "0001110" when "01100101000001011", -- t[51723] = 14
      "0001110" when "01100101000001100", -- t[51724] = 14
      "0001110" when "01100101000001101", -- t[51725] = 14
      "0001110" when "01100101000001110", -- t[51726] = 14
      "0001110" when "01100101000001111", -- t[51727] = 14
      "0001110" when "01100101000010000", -- t[51728] = 14
      "0001110" when "01100101000010001", -- t[51729] = 14
      "0001110" when "01100101000010010", -- t[51730] = 14
      "0001110" when "01100101000010011", -- t[51731] = 14
      "0001110" when "01100101000010100", -- t[51732] = 14
      "0001110" when "01100101000010101", -- t[51733] = 14
      "0001110" when "01100101000010110", -- t[51734] = 14
      "0001110" when "01100101000010111", -- t[51735] = 14
      "0001110" when "01100101000011000", -- t[51736] = 14
      "0001110" when "01100101000011001", -- t[51737] = 14
      "0001110" when "01100101000011010", -- t[51738] = 14
      "0001110" when "01100101000011011", -- t[51739] = 14
      "0001110" when "01100101000011100", -- t[51740] = 14
      "0001110" when "01100101000011101", -- t[51741] = 14
      "0001110" when "01100101000011110", -- t[51742] = 14
      "0001110" when "01100101000011111", -- t[51743] = 14
      "0001110" when "01100101000100000", -- t[51744] = 14
      "0001110" when "01100101000100001", -- t[51745] = 14
      "0001110" when "01100101000100010", -- t[51746] = 14
      "0001110" when "01100101000100011", -- t[51747] = 14
      "0001110" when "01100101000100100", -- t[51748] = 14
      "0001110" when "01100101000100101", -- t[51749] = 14
      "0001110" when "01100101000100110", -- t[51750] = 14
      "0001110" when "01100101000100111", -- t[51751] = 14
      "0001110" when "01100101000101000", -- t[51752] = 14
      "0001110" when "01100101000101001", -- t[51753] = 14
      "0001110" when "01100101000101010", -- t[51754] = 14
      "0001110" when "01100101000101011", -- t[51755] = 14
      "0001110" when "01100101000101100", -- t[51756] = 14
      "0001110" when "01100101000101101", -- t[51757] = 14
      "0001110" when "01100101000101110", -- t[51758] = 14
      "0001110" when "01100101000101111", -- t[51759] = 14
      "0001110" when "01100101000110000", -- t[51760] = 14
      "0001110" when "01100101000110001", -- t[51761] = 14
      "0001110" when "01100101000110010", -- t[51762] = 14
      "0001110" when "01100101000110011", -- t[51763] = 14
      "0001110" when "01100101000110100", -- t[51764] = 14
      "0001110" when "01100101000110101", -- t[51765] = 14
      "0001110" when "01100101000110110", -- t[51766] = 14
      "0001110" when "01100101000110111", -- t[51767] = 14
      "0001110" when "01100101000111000", -- t[51768] = 14
      "0001110" when "01100101000111001", -- t[51769] = 14
      "0001110" when "01100101000111010", -- t[51770] = 14
      "0001110" when "01100101000111011", -- t[51771] = 14
      "0001110" when "01100101000111100", -- t[51772] = 14
      "0001110" when "01100101000111101", -- t[51773] = 14
      "0001110" when "01100101000111110", -- t[51774] = 14
      "0001110" when "01100101000111111", -- t[51775] = 14
      "0001110" when "01100101001000000", -- t[51776] = 14
      "0001110" when "01100101001000001", -- t[51777] = 14
      "0001110" when "01100101001000010", -- t[51778] = 14
      "0001110" when "01100101001000011", -- t[51779] = 14
      "0001110" when "01100101001000100", -- t[51780] = 14
      "0001110" when "01100101001000101", -- t[51781] = 14
      "0001110" when "01100101001000110", -- t[51782] = 14
      "0001110" when "01100101001000111", -- t[51783] = 14
      "0001110" when "01100101001001000", -- t[51784] = 14
      "0001110" when "01100101001001001", -- t[51785] = 14
      "0001110" when "01100101001001010", -- t[51786] = 14
      "0001110" when "01100101001001011", -- t[51787] = 14
      "0001110" when "01100101001001100", -- t[51788] = 14
      "0001110" when "01100101001001101", -- t[51789] = 14
      "0001110" when "01100101001001110", -- t[51790] = 14
      "0001110" when "01100101001001111", -- t[51791] = 14
      "0001110" when "01100101001010000", -- t[51792] = 14
      "0001110" when "01100101001010001", -- t[51793] = 14
      "0001110" when "01100101001010010", -- t[51794] = 14
      "0001110" when "01100101001010011", -- t[51795] = 14
      "0001110" when "01100101001010100", -- t[51796] = 14
      "0001110" when "01100101001010101", -- t[51797] = 14
      "0001110" when "01100101001010110", -- t[51798] = 14
      "0001110" when "01100101001010111", -- t[51799] = 14
      "0001110" when "01100101001011000", -- t[51800] = 14
      "0001110" when "01100101001011001", -- t[51801] = 14
      "0001110" when "01100101001011010", -- t[51802] = 14
      "0001110" when "01100101001011011", -- t[51803] = 14
      "0001110" when "01100101001011100", -- t[51804] = 14
      "0001110" when "01100101001011101", -- t[51805] = 14
      "0001110" when "01100101001011110", -- t[51806] = 14
      "0001110" when "01100101001011111", -- t[51807] = 14
      "0001110" when "01100101001100000", -- t[51808] = 14
      "0001110" when "01100101001100001", -- t[51809] = 14
      "0001110" when "01100101001100010", -- t[51810] = 14
      "0001110" when "01100101001100011", -- t[51811] = 14
      "0001110" when "01100101001100100", -- t[51812] = 14
      "0001110" when "01100101001100101", -- t[51813] = 14
      "0001110" when "01100101001100110", -- t[51814] = 14
      "0001110" when "01100101001100111", -- t[51815] = 14
      "0001110" when "01100101001101000", -- t[51816] = 14
      "0001110" when "01100101001101001", -- t[51817] = 14
      "0001110" when "01100101001101010", -- t[51818] = 14
      "0001110" when "01100101001101011", -- t[51819] = 14
      "0001110" when "01100101001101100", -- t[51820] = 14
      "0001110" when "01100101001101101", -- t[51821] = 14
      "0001110" when "01100101001101110", -- t[51822] = 14
      "0001110" when "01100101001101111", -- t[51823] = 14
      "0001110" when "01100101001110000", -- t[51824] = 14
      "0001110" when "01100101001110001", -- t[51825] = 14
      "0001110" when "01100101001110010", -- t[51826] = 14
      "0001110" when "01100101001110011", -- t[51827] = 14
      "0001110" when "01100101001110100", -- t[51828] = 14
      "0001110" when "01100101001110101", -- t[51829] = 14
      "0001110" when "01100101001110110", -- t[51830] = 14
      "0001110" when "01100101001110111", -- t[51831] = 14
      "0001110" when "01100101001111000", -- t[51832] = 14
      "0001110" when "01100101001111001", -- t[51833] = 14
      "0001110" when "01100101001111010", -- t[51834] = 14
      "0001110" when "01100101001111011", -- t[51835] = 14
      "0001110" when "01100101001111100", -- t[51836] = 14
      "0001110" when "01100101001111101", -- t[51837] = 14
      "0001110" when "01100101001111110", -- t[51838] = 14
      "0001110" when "01100101001111111", -- t[51839] = 14
      "0001110" when "01100101010000000", -- t[51840] = 14
      "0001110" when "01100101010000001", -- t[51841] = 14
      "0001111" when "01100101010000010", -- t[51842] = 15
      "0001111" when "01100101010000011", -- t[51843] = 15
      "0001111" when "01100101010000100", -- t[51844] = 15
      "0001111" when "01100101010000101", -- t[51845] = 15
      "0001111" when "01100101010000110", -- t[51846] = 15
      "0001111" when "01100101010000111", -- t[51847] = 15
      "0001111" when "01100101010001000", -- t[51848] = 15
      "0001111" when "01100101010001001", -- t[51849] = 15
      "0001111" when "01100101010001010", -- t[51850] = 15
      "0001111" when "01100101010001011", -- t[51851] = 15
      "0001111" when "01100101010001100", -- t[51852] = 15
      "0001111" when "01100101010001101", -- t[51853] = 15
      "0001111" when "01100101010001110", -- t[51854] = 15
      "0001111" when "01100101010001111", -- t[51855] = 15
      "0001111" when "01100101010010000", -- t[51856] = 15
      "0001111" when "01100101010010001", -- t[51857] = 15
      "0001111" when "01100101010010010", -- t[51858] = 15
      "0001111" when "01100101010010011", -- t[51859] = 15
      "0001111" when "01100101010010100", -- t[51860] = 15
      "0001111" when "01100101010010101", -- t[51861] = 15
      "0001111" when "01100101010010110", -- t[51862] = 15
      "0001111" when "01100101010010111", -- t[51863] = 15
      "0001111" when "01100101010011000", -- t[51864] = 15
      "0001111" when "01100101010011001", -- t[51865] = 15
      "0001111" when "01100101010011010", -- t[51866] = 15
      "0001111" when "01100101010011011", -- t[51867] = 15
      "0001111" when "01100101010011100", -- t[51868] = 15
      "0001111" when "01100101010011101", -- t[51869] = 15
      "0001111" when "01100101010011110", -- t[51870] = 15
      "0001111" when "01100101010011111", -- t[51871] = 15
      "0001111" when "01100101010100000", -- t[51872] = 15
      "0001111" when "01100101010100001", -- t[51873] = 15
      "0001111" when "01100101010100010", -- t[51874] = 15
      "0001111" when "01100101010100011", -- t[51875] = 15
      "0001111" when "01100101010100100", -- t[51876] = 15
      "0001111" when "01100101010100101", -- t[51877] = 15
      "0001111" when "01100101010100110", -- t[51878] = 15
      "0001111" when "01100101010100111", -- t[51879] = 15
      "0001111" when "01100101010101000", -- t[51880] = 15
      "0001111" when "01100101010101001", -- t[51881] = 15
      "0001111" when "01100101010101010", -- t[51882] = 15
      "0001111" when "01100101010101011", -- t[51883] = 15
      "0001111" when "01100101010101100", -- t[51884] = 15
      "0001111" when "01100101010101101", -- t[51885] = 15
      "0001111" when "01100101010101110", -- t[51886] = 15
      "0001111" when "01100101010101111", -- t[51887] = 15
      "0001111" when "01100101010110000", -- t[51888] = 15
      "0001111" when "01100101010110001", -- t[51889] = 15
      "0001111" when "01100101010110010", -- t[51890] = 15
      "0001111" when "01100101010110011", -- t[51891] = 15
      "0001111" when "01100101010110100", -- t[51892] = 15
      "0001111" when "01100101010110101", -- t[51893] = 15
      "0001111" when "01100101010110110", -- t[51894] = 15
      "0001111" when "01100101010110111", -- t[51895] = 15
      "0001111" when "01100101010111000", -- t[51896] = 15
      "0001111" when "01100101010111001", -- t[51897] = 15
      "0001111" when "01100101010111010", -- t[51898] = 15
      "0001111" when "01100101010111011", -- t[51899] = 15
      "0001111" when "01100101010111100", -- t[51900] = 15
      "0001111" when "01100101010111101", -- t[51901] = 15
      "0001111" when "01100101010111110", -- t[51902] = 15
      "0001111" when "01100101010111111", -- t[51903] = 15
      "0001111" when "01100101011000000", -- t[51904] = 15
      "0001111" when "01100101011000001", -- t[51905] = 15
      "0001111" when "01100101011000010", -- t[51906] = 15
      "0001111" when "01100101011000011", -- t[51907] = 15
      "0001111" when "01100101011000100", -- t[51908] = 15
      "0001111" when "01100101011000101", -- t[51909] = 15
      "0001111" when "01100101011000110", -- t[51910] = 15
      "0001111" when "01100101011000111", -- t[51911] = 15
      "0001111" when "01100101011001000", -- t[51912] = 15
      "0001111" when "01100101011001001", -- t[51913] = 15
      "0001111" when "01100101011001010", -- t[51914] = 15
      "0001111" when "01100101011001011", -- t[51915] = 15
      "0001111" when "01100101011001100", -- t[51916] = 15
      "0001111" when "01100101011001101", -- t[51917] = 15
      "0001111" when "01100101011001110", -- t[51918] = 15
      "0001111" when "01100101011001111", -- t[51919] = 15
      "0001111" when "01100101011010000", -- t[51920] = 15
      "0001111" when "01100101011010001", -- t[51921] = 15
      "0001111" when "01100101011010010", -- t[51922] = 15
      "0001111" when "01100101011010011", -- t[51923] = 15
      "0001111" when "01100101011010100", -- t[51924] = 15
      "0001111" when "01100101011010101", -- t[51925] = 15
      "0001111" when "01100101011010110", -- t[51926] = 15
      "0001111" when "01100101011010111", -- t[51927] = 15
      "0001111" when "01100101011011000", -- t[51928] = 15
      "0001111" when "01100101011011001", -- t[51929] = 15
      "0001111" when "01100101011011010", -- t[51930] = 15
      "0001111" when "01100101011011011", -- t[51931] = 15
      "0001111" when "01100101011011100", -- t[51932] = 15
      "0001111" when "01100101011011101", -- t[51933] = 15
      "0001111" when "01100101011011110", -- t[51934] = 15
      "0001111" when "01100101011011111", -- t[51935] = 15
      "0001111" when "01100101011100000", -- t[51936] = 15
      "0001111" when "01100101011100001", -- t[51937] = 15
      "0001111" when "01100101011100010", -- t[51938] = 15
      "0001111" when "01100101011100011", -- t[51939] = 15
      "0001111" when "01100101011100100", -- t[51940] = 15
      "0001111" when "01100101011100101", -- t[51941] = 15
      "0001111" when "01100101011100110", -- t[51942] = 15
      "0001111" when "01100101011100111", -- t[51943] = 15
      "0001111" when "01100101011101000", -- t[51944] = 15
      "0001111" when "01100101011101001", -- t[51945] = 15
      "0001111" when "01100101011101010", -- t[51946] = 15
      "0001111" when "01100101011101011", -- t[51947] = 15
      "0001111" when "01100101011101100", -- t[51948] = 15
      "0001111" when "01100101011101101", -- t[51949] = 15
      "0001111" when "01100101011101110", -- t[51950] = 15
      "0001111" when "01100101011101111", -- t[51951] = 15
      "0001111" when "01100101011110000", -- t[51952] = 15
      "0001111" when "01100101011110001", -- t[51953] = 15
      "0001111" when "01100101011110010", -- t[51954] = 15
      "0001111" when "01100101011110011", -- t[51955] = 15
      "0001111" when "01100101011110100", -- t[51956] = 15
      "0001111" when "01100101011110101", -- t[51957] = 15
      "0001111" when "01100101011110110", -- t[51958] = 15
      "0001111" when "01100101011110111", -- t[51959] = 15
      "0001111" when "01100101011111000", -- t[51960] = 15
      "0001111" when "01100101011111001", -- t[51961] = 15
      "0001111" when "01100101011111010", -- t[51962] = 15
      "0001111" when "01100101011111011", -- t[51963] = 15
      "0001111" when "01100101011111100", -- t[51964] = 15
      "0001111" when "01100101011111101", -- t[51965] = 15
      "0001111" when "01100101011111110", -- t[51966] = 15
      "0001111" when "01100101011111111", -- t[51967] = 15
      "0001111" when "01100101100000000", -- t[51968] = 15
      "0001111" when "01100101100000001", -- t[51969] = 15
      "0001111" when "01100101100000010", -- t[51970] = 15
      "0001111" when "01100101100000011", -- t[51971] = 15
      "0001111" when "01100101100000100", -- t[51972] = 15
      "0001111" when "01100101100000101", -- t[51973] = 15
      "0001111" when "01100101100000110", -- t[51974] = 15
      "0001111" when "01100101100000111", -- t[51975] = 15
      "0001111" when "01100101100001000", -- t[51976] = 15
      "0001111" when "01100101100001001", -- t[51977] = 15
      "0001111" when "01100101100001010", -- t[51978] = 15
      "0001111" when "01100101100001011", -- t[51979] = 15
      "0001111" when "01100101100001100", -- t[51980] = 15
      "0001111" when "01100101100001101", -- t[51981] = 15
      "0001111" when "01100101100001110", -- t[51982] = 15
      "0001111" when "01100101100001111", -- t[51983] = 15
      "0001111" when "01100101100010000", -- t[51984] = 15
      "0001111" when "01100101100010001", -- t[51985] = 15
      "0001111" when "01100101100010010", -- t[51986] = 15
      "0001111" when "01100101100010011", -- t[51987] = 15
      "0001111" when "01100101100010100", -- t[51988] = 15
      "0001111" when "01100101100010101", -- t[51989] = 15
      "0001111" when "01100101100010110", -- t[51990] = 15
      "0001111" when "01100101100010111", -- t[51991] = 15
      "0001111" when "01100101100011000", -- t[51992] = 15
      "0001111" when "01100101100011001", -- t[51993] = 15
      "0001111" when "01100101100011010", -- t[51994] = 15
      "0001111" when "01100101100011011", -- t[51995] = 15
      "0001111" when "01100101100011100", -- t[51996] = 15
      "0001111" when "01100101100011101", -- t[51997] = 15
      "0001111" when "01100101100011110", -- t[51998] = 15
      "0001111" when "01100101100011111", -- t[51999] = 15
      "0001111" when "01100101100100000", -- t[52000] = 15
      "0001111" when "01100101100100001", -- t[52001] = 15
      "0001111" when "01100101100100010", -- t[52002] = 15
      "0001111" when "01100101100100011", -- t[52003] = 15
      "0001111" when "01100101100100100", -- t[52004] = 15
      "0001111" when "01100101100100101", -- t[52005] = 15
      "0001111" when "01100101100100110", -- t[52006] = 15
      "0001111" when "01100101100100111", -- t[52007] = 15
      "0001111" when "01100101100101000", -- t[52008] = 15
      "0001111" when "01100101100101001", -- t[52009] = 15
      "0001111" when "01100101100101010", -- t[52010] = 15
      "0001111" when "01100101100101011", -- t[52011] = 15
      "0001111" when "01100101100101100", -- t[52012] = 15
      "0001111" when "01100101100101101", -- t[52013] = 15
      "0001111" when "01100101100101110", -- t[52014] = 15
      "0001111" when "01100101100101111", -- t[52015] = 15
      "0001111" when "01100101100110000", -- t[52016] = 15
      "0001111" when "01100101100110001", -- t[52017] = 15
      "0001111" when "01100101100110010", -- t[52018] = 15
      "0001111" when "01100101100110011", -- t[52019] = 15
      "0001111" when "01100101100110100", -- t[52020] = 15
      "0001111" when "01100101100110101", -- t[52021] = 15
      "0001111" when "01100101100110110", -- t[52022] = 15
      "0001111" when "01100101100110111", -- t[52023] = 15
      "0001111" when "01100101100111000", -- t[52024] = 15
      "0001111" when "01100101100111001", -- t[52025] = 15
      "0001111" when "01100101100111010", -- t[52026] = 15
      "0001111" when "01100101100111011", -- t[52027] = 15
      "0001111" when "01100101100111100", -- t[52028] = 15
      "0001111" when "01100101100111101", -- t[52029] = 15
      "0001111" when "01100101100111110", -- t[52030] = 15
      "0001111" when "01100101100111111", -- t[52031] = 15
      "0001111" when "01100101101000000", -- t[52032] = 15
      "0001111" when "01100101101000001", -- t[52033] = 15
      "0001111" when "01100101101000010", -- t[52034] = 15
      "0001111" when "01100101101000011", -- t[52035] = 15
      "0001111" when "01100101101000100", -- t[52036] = 15
      "0001111" when "01100101101000101", -- t[52037] = 15
      "0001111" when "01100101101000110", -- t[52038] = 15
      "0001111" when "01100101101000111", -- t[52039] = 15
      "0001111" when "01100101101001000", -- t[52040] = 15
      "0001111" when "01100101101001001", -- t[52041] = 15
      "0001111" when "01100101101001010", -- t[52042] = 15
      "0001111" when "01100101101001011", -- t[52043] = 15
      "0001111" when "01100101101001100", -- t[52044] = 15
      "0001111" when "01100101101001101", -- t[52045] = 15
      "0001111" when "01100101101001110", -- t[52046] = 15
      "0001111" when "01100101101001111", -- t[52047] = 15
      "0001111" when "01100101101010000", -- t[52048] = 15
      "0001111" when "01100101101010001", -- t[52049] = 15
      "0001111" when "01100101101010010", -- t[52050] = 15
      "0001111" when "01100101101010011", -- t[52051] = 15
      "0001111" when "01100101101010100", -- t[52052] = 15
      "0001111" when "01100101101010101", -- t[52053] = 15
      "0001111" when "01100101101010110", -- t[52054] = 15
      "0001111" when "01100101101010111", -- t[52055] = 15
      "0001111" when "01100101101011000", -- t[52056] = 15
      "0001111" when "01100101101011001", -- t[52057] = 15
      "0001111" when "01100101101011010", -- t[52058] = 15
      "0001111" when "01100101101011011", -- t[52059] = 15
      "0001111" when "01100101101011100", -- t[52060] = 15
      "0001111" when "01100101101011101", -- t[52061] = 15
      "0001111" when "01100101101011110", -- t[52062] = 15
      "0001111" when "01100101101011111", -- t[52063] = 15
      "0001111" when "01100101101100000", -- t[52064] = 15
      "0001111" when "01100101101100001", -- t[52065] = 15
      "0001111" when "01100101101100010", -- t[52066] = 15
      "0001111" when "01100101101100011", -- t[52067] = 15
      "0001111" when "01100101101100100", -- t[52068] = 15
      "0001111" when "01100101101100101", -- t[52069] = 15
      "0001111" when "01100101101100110", -- t[52070] = 15
      "0001111" when "01100101101100111", -- t[52071] = 15
      "0001111" when "01100101101101000", -- t[52072] = 15
      "0001111" when "01100101101101001", -- t[52073] = 15
      "0001111" when "01100101101101010", -- t[52074] = 15
      "0001111" when "01100101101101011", -- t[52075] = 15
      "0001111" when "01100101101101100", -- t[52076] = 15
      "0001111" when "01100101101101101", -- t[52077] = 15
      "0001111" when "01100101101101110", -- t[52078] = 15
      "0001111" when "01100101101101111", -- t[52079] = 15
      "0001111" when "01100101101110000", -- t[52080] = 15
      "0001111" when "01100101101110001", -- t[52081] = 15
      "0001111" when "01100101101110010", -- t[52082] = 15
      "0001111" when "01100101101110011", -- t[52083] = 15
      "0001111" when "01100101101110100", -- t[52084] = 15
      "0001111" when "01100101101110101", -- t[52085] = 15
      "0001111" when "01100101101110110", -- t[52086] = 15
      "0001111" when "01100101101110111", -- t[52087] = 15
      "0001111" when "01100101101111000", -- t[52088] = 15
      "0001111" when "01100101101111001", -- t[52089] = 15
      "0001111" when "01100101101111010", -- t[52090] = 15
      "0001111" when "01100101101111011", -- t[52091] = 15
      "0001111" when "01100101101111100", -- t[52092] = 15
      "0001111" when "01100101101111101", -- t[52093] = 15
      "0001111" when "01100101101111110", -- t[52094] = 15
      "0001111" when "01100101101111111", -- t[52095] = 15
      "0001111" when "01100101110000000", -- t[52096] = 15
      "0001111" when "01100101110000001", -- t[52097] = 15
      "0001111" when "01100101110000010", -- t[52098] = 15
      "0001111" when "01100101110000011", -- t[52099] = 15
      "0001111" when "01100101110000100", -- t[52100] = 15
      "0001111" when "01100101110000101", -- t[52101] = 15
      "0001111" when "01100101110000110", -- t[52102] = 15
      "0001111" when "01100101110000111", -- t[52103] = 15
      "0001111" when "01100101110001000", -- t[52104] = 15
      "0001111" when "01100101110001001", -- t[52105] = 15
      "0001111" when "01100101110001010", -- t[52106] = 15
      "0001111" when "01100101110001011", -- t[52107] = 15
      "0001111" when "01100101110001100", -- t[52108] = 15
      "0001111" when "01100101110001101", -- t[52109] = 15
      "0001111" when "01100101110001110", -- t[52110] = 15
      "0001111" when "01100101110001111", -- t[52111] = 15
      "0001111" when "01100101110010000", -- t[52112] = 15
      "0001111" when "01100101110010001", -- t[52113] = 15
      "0001111" when "01100101110010010", -- t[52114] = 15
      "0001111" when "01100101110010011", -- t[52115] = 15
      "0001111" when "01100101110010100", -- t[52116] = 15
      "0001111" when "01100101110010101", -- t[52117] = 15
      "0001111" when "01100101110010110", -- t[52118] = 15
      "0001111" when "01100101110010111", -- t[52119] = 15
      "0001111" when "01100101110011000", -- t[52120] = 15
      "0001111" when "01100101110011001", -- t[52121] = 15
      "0001111" when "01100101110011010", -- t[52122] = 15
      "0001111" when "01100101110011011", -- t[52123] = 15
      "0001111" when "01100101110011100", -- t[52124] = 15
      "0001111" when "01100101110011101", -- t[52125] = 15
      "0001111" when "01100101110011110", -- t[52126] = 15
      "0001111" when "01100101110011111", -- t[52127] = 15
      "0001111" when "01100101110100000", -- t[52128] = 15
      "0001111" when "01100101110100001", -- t[52129] = 15
      "0001111" when "01100101110100010", -- t[52130] = 15
      "0001111" when "01100101110100011", -- t[52131] = 15
      "0001111" when "01100101110100100", -- t[52132] = 15
      "0001111" when "01100101110100101", -- t[52133] = 15
      "0001111" when "01100101110100110", -- t[52134] = 15
      "0001111" when "01100101110100111", -- t[52135] = 15
      "0001111" when "01100101110101000", -- t[52136] = 15
      "0001111" when "01100101110101001", -- t[52137] = 15
      "0001111" when "01100101110101010", -- t[52138] = 15
      "0001111" when "01100101110101011", -- t[52139] = 15
      "0001111" when "01100101110101100", -- t[52140] = 15
      "0001111" when "01100101110101101", -- t[52141] = 15
      "0001111" when "01100101110101110", -- t[52142] = 15
      "0001111" when "01100101110101111", -- t[52143] = 15
      "0001111" when "01100101110110000", -- t[52144] = 15
      "0001111" when "01100101110110001", -- t[52145] = 15
      "0001111" when "01100101110110010", -- t[52146] = 15
      "0001111" when "01100101110110011", -- t[52147] = 15
      "0001111" when "01100101110110100", -- t[52148] = 15
      "0001111" when "01100101110110101", -- t[52149] = 15
      "0001111" when "01100101110110110", -- t[52150] = 15
      "0001111" when "01100101110110111", -- t[52151] = 15
      "0001111" when "01100101110111000", -- t[52152] = 15
      "0001111" when "01100101110111001", -- t[52153] = 15
      "0001111" when "01100101110111010", -- t[52154] = 15
      "0001111" when "01100101110111011", -- t[52155] = 15
      "0001111" when "01100101110111100", -- t[52156] = 15
      "0001111" when "01100101110111101", -- t[52157] = 15
      "0001111" when "01100101110111110", -- t[52158] = 15
      "0001111" when "01100101110111111", -- t[52159] = 15
      "0001111" when "01100101111000000", -- t[52160] = 15
      "0001111" when "01100101111000001", -- t[52161] = 15
      "0001111" when "01100101111000010", -- t[52162] = 15
      "0001111" when "01100101111000011", -- t[52163] = 15
      "0001111" when "01100101111000100", -- t[52164] = 15
      "0001111" when "01100101111000101", -- t[52165] = 15
      "0001111" when "01100101111000110", -- t[52166] = 15
      "0001111" when "01100101111000111", -- t[52167] = 15
      "0001111" when "01100101111001000", -- t[52168] = 15
      "0001111" when "01100101111001001", -- t[52169] = 15
      "0001111" when "01100101111001010", -- t[52170] = 15
      "0001111" when "01100101111001011", -- t[52171] = 15
      "0001111" when "01100101111001100", -- t[52172] = 15
      "0001111" when "01100101111001101", -- t[52173] = 15
      "0001111" when "01100101111001110", -- t[52174] = 15
      "0001111" when "01100101111001111", -- t[52175] = 15
      "0001111" when "01100101111010000", -- t[52176] = 15
      "0001111" when "01100101111010001", -- t[52177] = 15
      "0001111" when "01100101111010010", -- t[52178] = 15
      "0001111" when "01100101111010011", -- t[52179] = 15
      "0001111" when "01100101111010100", -- t[52180] = 15
      "0001111" when "01100101111010101", -- t[52181] = 15
      "0001111" when "01100101111010110", -- t[52182] = 15
      "0001111" when "01100101111010111", -- t[52183] = 15
      "0001111" when "01100101111011000", -- t[52184] = 15
      "0001111" when "01100101111011001", -- t[52185] = 15
      "0001111" when "01100101111011010", -- t[52186] = 15
      "0001111" when "01100101111011011", -- t[52187] = 15
      "0001111" when "01100101111011100", -- t[52188] = 15
      "0001111" when "01100101111011101", -- t[52189] = 15
      "0001111" when "01100101111011110", -- t[52190] = 15
      "0001111" when "01100101111011111", -- t[52191] = 15
      "0001111" when "01100101111100000", -- t[52192] = 15
      "0001111" when "01100101111100001", -- t[52193] = 15
      "0001111" when "01100101111100010", -- t[52194] = 15
      "0001111" when "01100101111100011", -- t[52195] = 15
      "0001111" when "01100101111100100", -- t[52196] = 15
      "0001111" when "01100101111100101", -- t[52197] = 15
      "0001111" when "01100101111100110", -- t[52198] = 15
      "0001111" when "01100101111100111", -- t[52199] = 15
      "0001111" when "01100101111101000", -- t[52200] = 15
      "0001111" when "01100101111101001", -- t[52201] = 15
      "0001111" when "01100101111101010", -- t[52202] = 15
      "0001111" when "01100101111101011", -- t[52203] = 15
      "0001111" when "01100101111101100", -- t[52204] = 15
      "0001111" when "01100101111101101", -- t[52205] = 15
      "0001111" when "01100101111101110", -- t[52206] = 15
      "0001111" when "01100101111101111", -- t[52207] = 15
      "0001111" when "01100101111110000", -- t[52208] = 15
      "0001111" when "01100101111110001", -- t[52209] = 15
      "0001111" when "01100101111110010", -- t[52210] = 15
      "0001111" when "01100101111110011", -- t[52211] = 15
      "0001111" when "01100101111110100", -- t[52212] = 15
      "0001111" when "01100101111110101", -- t[52213] = 15
      "0001111" when "01100101111110110", -- t[52214] = 15
      "0001111" when "01100101111110111", -- t[52215] = 15
      "0001111" when "01100101111111000", -- t[52216] = 15
      "0001111" when "01100101111111001", -- t[52217] = 15
      "0001111" when "01100101111111010", -- t[52218] = 15
      "0001111" when "01100101111111011", -- t[52219] = 15
      "0001111" when "01100101111111100", -- t[52220] = 15
      "0001111" when "01100101111111101", -- t[52221] = 15
      "0001111" when "01100101111111110", -- t[52222] = 15
      "0001111" when "01100101111111111", -- t[52223] = 15
      "0001111" when "01100110000000000", -- t[52224] = 15
      "0001111" when "01100110000000001", -- t[52225] = 15
      "0001111" when "01100110000000010", -- t[52226] = 15
      "0001111" when "01100110000000011", -- t[52227] = 15
      "0001111" when "01100110000000100", -- t[52228] = 15
      "0001111" when "01100110000000101", -- t[52229] = 15
      "0001111" when "01100110000000110", -- t[52230] = 15
      "0001111" when "01100110000000111", -- t[52231] = 15
      "0001111" when "01100110000001000", -- t[52232] = 15
      "0001111" when "01100110000001001", -- t[52233] = 15
      "0001111" when "01100110000001010", -- t[52234] = 15
      "0001111" when "01100110000001011", -- t[52235] = 15
      "0001111" when "01100110000001100", -- t[52236] = 15
      "0001111" when "01100110000001101", -- t[52237] = 15
      "0001111" when "01100110000001110", -- t[52238] = 15
      "0001111" when "01100110000001111", -- t[52239] = 15
      "0001111" when "01100110000010000", -- t[52240] = 15
      "0001111" when "01100110000010001", -- t[52241] = 15
      "0001111" when "01100110000010010", -- t[52242] = 15
      "0001111" when "01100110000010011", -- t[52243] = 15
      "0001111" when "01100110000010100", -- t[52244] = 15
      "0001111" when "01100110000010101", -- t[52245] = 15
      "0001111" when "01100110000010110", -- t[52246] = 15
      "0001111" when "01100110000010111", -- t[52247] = 15
      "0001111" when "01100110000011000", -- t[52248] = 15
      "0001111" when "01100110000011001", -- t[52249] = 15
      "0001111" when "01100110000011010", -- t[52250] = 15
      "0001111" when "01100110000011011", -- t[52251] = 15
      "0001111" when "01100110000011100", -- t[52252] = 15
      "0001111" when "01100110000011101", -- t[52253] = 15
      "0001111" when "01100110000011110", -- t[52254] = 15
      "0001111" when "01100110000011111", -- t[52255] = 15
      "0001111" when "01100110000100000", -- t[52256] = 15
      "0001111" when "01100110000100001", -- t[52257] = 15
      "0001111" when "01100110000100010", -- t[52258] = 15
      "0001111" when "01100110000100011", -- t[52259] = 15
      "0001111" when "01100110000100100", -- t[52260] = 15
      "0001111" when "01100110000100101", -- t[52261] = 15
      "0001111" when "01100110000100110", -- t[52262] = 15
      "0001111" when "01100110000100111", -- t[52263] = 15
      "0001111" when "01100110000101000", -- t[52264] = 15
      "0001111" when "01100110000101001", -- t[52265] = 15
      "0001111" when "01100110000101010", -- t[52266] = 15
      "0001111" when "01100110000101011", -- t[52267] = 15
      "0001111" when "01100110000101100", -- t[52268] = 15
      "0001111" when "01100110000101101", -- t[52269] = 15
      "0001111" when "01100110000101110", -- t[52270] = 15
      "0001111" when "01100110000101111", -- t[52271] = 15
      "0001111" when "01100110000110000", -- t[52272] = 15
      "0001111" when "01100110000110001", -- t[52273] = 15
      "0001111" when "01100110000110010", -- t[52274] = 15
      "0001111" when "01100110000110011", -- t[52275] = 15
      "0001111" when "01100110000110100", -- t[52276] = 15
      "0001111" when "01100110000110101", -- t[52277] = 15
      "0001111" when "01100110000110110", -- t[52278] = 15
      "0001111" when "01100110000110111", -- t[52279] = 15
      "0001111" when "01100110000111000", -- t[52280] = 15
      "0001111" when "01100110000111001", -- t[52281] = 15
      "0001111" when "01100110000111010", -- t[52282] = 15
      "0001111" when "01100110000111011", -- t[52283] = 15
      "0001111" when "01100110000111100", -- t[52284] = 15
      "0001111" when "01100110000111101", -- t[52285] = 15
      "0001111" when "01100110000111110", -- t[52286] = 15
      "0001111" when "01100110000111111", -- t[52287] = 15
      "0001111" when "01100110001000000", -- t[52288] = 15
      "0001111" when "01100110001000001", -- t[52289] = 15
      "0001111" when "01100110001000010", -- t[52290] = 15
      "0001111" when "01100110001000011", -- t[52291] = 15
      "0001111" when "01100110001000100", -- t[52292] = 15
      "0001111" when "01100110001000101", -- t[52293] = 15
      "0001111" when "01100110001000110", -- t[52294] = 15
      "0001111" when "01100110001000111", -- t[52295] = 15
      "0001111" when "01100110001001000", -- t[52296] = 15
      "0001111" when "01100110001001001", -- t[52297] = 15
      "0001111" when "01100110001001010", -- t[52298] = 15
      "0001111" when "01100110001001011", -- t[52299] = 15
      "0001111" when "01100110001001100", -- t[52300] = 15
      "0001111" when "01100110001001101", -- t[52301] = 15
      "0001111" when "01100110001001110", -- t[52302] = 15
      "0001111" when "01100110001001111", -- t[52303] = 15
      "0001111" when "01100110001010000", -- t[52304] = 15
      "0001111" when "01100110001010001", -- t[52305] = 15
      "0001111" when "01100110001010010", -- t[52306] = 15
      "0001111" when "01100110001010011", -- t[52307] = 15
      "0001111" when "01100110001010100", -- t[52308] = 15
      "0001111" when "01100110001010101", -- t[52309] = 15
      "0001111" when "01100110001010110", -- t[52310] = 15
      "0001111" when "01100110001010111", -- t[52311] = 15
      "0001111" when "01100110001011000", -- t[52312] = 15
      "0001111" when "01100110001011001", -- t[52313] = 15
      "0001111" when "01100110001011010", -- t[52314] = 15
      "0001111" when "01100110001011011", -- t[52315] = 15
      "0001111" when "01100110001011100", -- t[52316] = 15
      "0001111" when "01100110001011101", -- t[52317] = 15
      "0001111" when "01100110001011110", -- t[52318] = 15
      "0001111" when "01100110001011111", -- t[52319] = 15
      "0001111" when "01100110001100000", -- t[52320] = 15
      "0001111" when "01100110001100001", -- t[52321] = 15
      "0001111" when "01100110001100010", -- t[52322] = 15
      "0001111" when "01100110001100011", -- t[52323] = 15
      "0001111" when "01100110001100100", -- t[52324] = 15
      "0001111" when "01100110001100101", -- t[52325] = 15
      "0001111" when "01100110001100110", -- t[52326] = 15
      "0001111" when "01100110001100111", -- t[52327] = 15
      "0001111" when "01100110001101000", -- t[52328] = 15
      "0001111" when "01100110001101001", -- t[52329] = 15
      "0001111" when "01100110001101010", -- t[52330] = 15
      "0001111" when "01100110001101011", -- t[52331] = 15
      "0001111" when "01100110001101100", -- t[52332] = 15
      "0001111" when "01100110001101101", -- t[52333] = 15
      "0001111" when "01100110001101110", -- t[52334] = 15
      "0001111" when "01100110001101111", -- t[52335] = 15
      "0001111" when "01100110001110000", -- t[52336] = 15
      "0001111" when "01100110001110001", -- t[52337] = 15
      "0001111" when "01100110001110010", -- t[52338] = 15
      "0001111" when "01100110001110011", -- t[52339] = 15
      "0001111" when "01100110001110100", -- t[52340] = 15
      "0001111" when "01100110001110101", -- t[52341] = 15
      "0001111" when "01100110001110110", -- t[52342] = 15
      "0001111" when "01100110001110111", -- t[52343] = 15
      "0001111" when "01100110001111000", -- t[52344] = 15
      "0001111" when "01100110001111001", -- t[52345] = 15
      "0001111" when "01100110001111010", -- t[52346] = 15
      "0001111" when "01100110001111011", -- t[52347] = 15
      "0001111" when "01100110001111100", -- t[52348] = 15
      "0001111" when "01100110001111101", -- t[52349] = 15
      "0001111" when "01100110001111110", -- t[52350] = 15
      "0001111" when "01100110001111111", -- t[52351] = 15
      "0001111" when "01100110010000000", -- t[52352] = 15
      "0001111" when "01100110010000001", -- t[52353] = 15
      "0001111" when "01100110010000010", -- t[52354] = 15
      "0001111" when "01100110010000011", -- t[52355] = 15
      "0001111" when "01100110010000100", -- t[52356] = 15
      "0001111" when "01100110010000101", -- t[52357] = 15
      "0001111" when "01100110010000110", -- t[52358] = 15
      "0001111" when "01100110010000111", -- t[52359] = 15
      "0001111" when "01100110010001000", -- t[52360] = 15
      "0001111" when "01100110010001001", -- t[52361] = 15
      "0001111" when "01100110010001010", -- t[52362] = 15
      "0001111" when "01100110010001011", -- t[52363] = 15
      "0001111" when "01100110010001100", -- t[52364] = 15
      "0001111" when "01100110010001101", -- t[52365] = 15
      "0001111" when "01100110010001110", -- t[52366] = 15
      "0001111" when "01100110010001111", -- t[52367] = 15
      "0001111" when "01100110010010000", -- t[52368] = 15
      "0001111" when "01100110010010001", -- t[52369] = 15
      "0001111" when "01100110010010010", -- t[52370] = 15
      "0001111" when "01100110010010011", -- t[52371] = 15
      "0001111" when "01100110010010100", -- t[52372] = 15
      "0001111" when "01100110010010101", -- t[52373] = 15
      "0001111" when "01100110010010110", -- t[52374] = 15
      "0001111" when "01100110010010111", -- t[52375] = 15
      "0001111" when "01100110010011000", -- t[52376] = 15
      "0001111" when "01100110010011001", -- t[52377] = 15
      "0001111" when "01100110010011010", -- t[52378] = 15
      "0001111" when "01100110010011011", -- t[52379] = 15
      "0001111" when "01100110010011100", -- t[52380] = 15
      "0001111" when "01100110010011101", -- t[52381] = 15
      "0001111" when "01100110010011110", -- t[52382] = 15
      "0001111" when "01100110010011111", -- t[52383] = 15
      "0001111" when "01100110010100000", -- t[52384] = 15
      "0001111" when "01100110010100001", -- t[52385] = 15
      "0001111" when "01100110010100010", -- t[52386] = 15
      "0001111" when "01100110010100011", -- t[52387] = 15
      "0001111" when "01100110010100100", -- t[52388] = 15
      "0001111" when "01100110010100101", -- t[52389] = 15
      "0001111" when "01100110010100110", -- t[52390] = 15
      "0001111" when "01100110010100111", -- t[52391] = 15
      "0001111" when "01100110010101000", -- t[52392] = 15
      "0001111" when "01100110010101001", -- t[52393] = 15
      "0001111" when "01100110010101010", -- t[52394] = 15
      "0001111" when "01100110010101011", -- t[52395] = 15
      "0001111" when "01100110010101100", -- t[52396] = 15
      "0001111" when "01100110010101101", -- t[52397] = 15
      "0001111" when "01100110010101110", -- t[52398] = 15
      "0001111" when "01100110010101111", -- t[52399] = 15
      "0001111" when "01100110010110000", -- t[52400] = 15
      "0001111" when "01100110010110001", -- t[52401] = 15
      "0001111" when "01100110010110010", -- t[52402] = 15
      "0001111" when "01100110010110011", -- t[52403] = 15
      "0001111" when "01100110010110100", -- t[52404] = 15
      "0001111" when "01100110010110101", -- t[52405] = 15
      "0001111" when "01100110010110110", -- t[52406] = 15
      "0001111" when "01100110010110111", -- t[52407] = 15
      "0001111" when "01100110010111000", -- t[52408] = 15
      "0001111" when "01100110010111001", -- t[52409] = 15
      "0001111" when "01100110010111010", -- t[52410] = 15
      "0001111" when "01100110010111011", -- t[52411] = 15
      "0001111" when "01100110010111100", -- t[52412] = 15
      "0001111" when "01100110010111101", -- t[52413] = 15
      "0001111" when "01100110010111110", -- t[52414] = 15
      "0001111" when "01100110010111111", -- t[52415] = 15
      "0001111" when "01100110011000000", -- t[52416] = 15
      "0001111" when "01100110011000001", -- t[52417] = 15
      "0001111" when "01100110011000010", -- t[52418] = 15
      "0001111" when "01100110011000011", -- t[52419] = 15
      "0001111" when "01100110011000100", -- t[52420] = 15
      "0001111" when "01100110011000101", -- t[52421] = 15
      "0001111" when "01100110011000110", -- t[52422] = 15
      "0001111" when "01100110011000111", -- t[52423] = 15
      "0001111" when "01100110011001000", -- t[52424] = 15
      "0001111" when "01100110011001001", -- t[52425] = 15
      "0001111" when "01100110011001010", -- t[52426] = 15
      "0001111" when "01100110011001011", -- t[52427] = 15
      "0001111" when "01100110011001100", -- t[52428] = 15
      "0001111" when "01100110011001101", -- t[52429] = 15
      "0001111" when "01100110011001110", -- t[52430] = 15
      "0001111" when "01100110011001111", -- t[52431] = 15
      "0001111" when "01100110011010000", -- t[52432] = 15
      "0001111" when "01100110011010001", -- t[52433] = 15
      "0001111" when "01100110011010010", -- t[52434] = 15
      "0001111" when "01100110011010011", -- t[52435] = 15
      "0001111" when "01100110011010100", -- t[52436] = 15
      "0001111" when "01100110011010101", -- t[52437] = 15
      "0001111" when "01100110011010110", -- t[52438] = 15
      "0001111" when "01100110011010111", -- t[52439] = 15
      "0001111" when "01100110011011000", -- t[52440] = 15
      "0001111" when "01100110011011001", -- t[52441] = 15
      "0001111" when "01100110011011010", -- t[52442] = 15
      "0001111" when "01100110011011011", -- t[52443] = 15
      "0001111" when "01100110011011100", -- t[52444] = 15
      "0001111" when "01100110011011101", -- t[52445] = 15
      "0001111" when "01100110011011110", -- t[52446] = 15
      "0001111" when "01100110011011111", -- t[52447] = 15
      "0001111" when "01100110011100000", -- t[52448] = 15
      "0001111" when "01100110011100001", -- t[52449] = 15
      "0001111" when "01100110011100010", -- t[52450] = 15
      "0001111" when "01100110011100011", -- t[52451] = 15
      "0001111" when "01100110011100100", -- t[52452] = 15
      "0001111" when "01100110011100101", -- t[52453] = 15
      "0001111" when "01100110011100110", -- t[52454] = 15
      "0001111" when "01100110011100111", -- t[52455] = 15
      "0001111" when "01100110011101000", -- t[52456] = 15
      "0001111" when "01100110011101001", -- t[52457] = 15
      "0001111" when "01100110011101010", -- t[52458] = 15
      "0001111" when "01100110011101011", -- t[52459] = 15
      "0001111" when "01100110011101100", -- t[52460] = 15
      "0001111" when "01100110011101101", -- t[52461] = 15
      "0001111" when "01100110011101110", -- t[52462] = 15
      "0001111" when "01100110011101111", -- t[52463] = 15
      "0001111" when "01100110011110000", -- t[52464] = 15
      "0001111" when "01100110011110001", -- t[52465] = 15
      "0001111" when "01100110011110010", -- t[52466] = 15
      "0001111" when "01100110011110011", -- t[52467] = 15
      "0001111" when "01100110011110100", -- t[52468] = 15
      "0001111" when "01100110011110101", -- t[52469] = 15
      "0001111" when "01100110011110110", -- t[52470] = 15
      "0001111" when "01100110011110111", -- t[52471] = 15
      "0001111" when "01100110011111000", -- t[52472] = 15
      "0001111" when "01100110011111001", -- t[52473] = 15
      "0001111" when "01100110011111010", -- t[52474] = 15
      "0001111" when "01100110011111011", -- t[52475] = 15
      "0001111" when "01100110011111100", -- t[52476] = 15
      "0001111" when "01100110011111101", -- t[52477] = 15
      "0001111" when "01100110011111110", -- t[52478] = 15
      "0001111" when "01100110011111111", -- t[52479] = 15
      "0001111" when "01100110100000000", -- t[52480] = 15
      "0001111" when "01100110100000001", -- t[52481] = 15
      "0001111" when "01100110100000010", -- t[52482] = 15
      "0001111" when "01100110100000011", -- t[52483] = 15
      "0001111" when "01100110100000100", -- t[52484] = 15
      "0001111" when "01100110100000101", -- t[52485] = 15
      "0001111" when "01100110100000110", -- t[52486] = 15
      "0001111" when "01100110100000111", -- t[52487] = 15
      "0001111" when "01100110100001000", -- t[52488] = 15
      "0001111" when "01100110100001001", -- t[52489] = 15
      "0001111" when "01100110100001010", -- t[52490] = 15
      "0001111" when "01100110100001011", -- t[52491] = 15
      "0001111" when "01100110100001100", -- t[52492] = 15
      "0001111" when "01100110100001101", -- t[52493] = 15
      "0001111" when "01100110100001110", -- t[52494] = 15
      "0001111" when "01100110100001111", -- t[52495] = 15
      "0001111" when "01100110100010000", -- t[52496] = 15
      "0001111" when "01100110100010001", -- t[52497] = 15
      "0001111" when "01100110100010010", -- t[52498] = 15
      "0001111" when "01100110100010011", -- t[52499] = 15
      "0001111" when "01100110100010100", -- t[52500] = 15
      "0001111" when "01100110100010101", -- t[52501] = 15
      "0001111" when "01100110100010110", -- t[52502] = 15
      "0001111" when "01100110100010111", -- t[52503] = 15
      "0001111" when "01100110100011000", -- t[52504] = 15
      "0001111" when "01100110100011001", -- t[52505] = 15
      "0001111" when "01100110100011010", -- t[52506] = 15
      "0001111" when "01100110100011011", -- t[52507] = 15
      "0001111" when "01100110100011100", -- t[52508] = 15
      "0001111" when "01100110100011101", -- t[52509] = 15
      "0001111" when "01100110100011110", -- t[52510] = 15
      "0001111" when "01100110100011111", -- t[52511] = 15
      "0001111" when "01100110100100000", -- t[52512] = 15
      "0001111" when "01100110100100001", -- t[52513] = 15
      "0001111" when "01100110100100010", -- t[52514] = 15
      "0001111" when "01100110100100011", -- t[52515] = 15
      "0001111" when "01100110100100100", -- t[52516] = 15
      "0001111" when "01100110100100101", -- t[52517] = 15
      "0001111" when "01100110100100110", -- t[52518] = 15
      "0001111" when "01100110100100111", -- t[52519] = 15
      "0001111" when "01100110100101000", -- t[52520] = 15
      "0001111" when "01100110100101001", -- t[52521] = 15
      "0001111" when "01100110100101010", -- t[52522] = 15
      "0001111" when "01100110100101011", -- t[52523] = 15
      "0001111" when "01100110100101100", -- t[52524] = 15
      "0001111" when "01100110100101101", -- t[52525] = 15
      "0001111" when "01100110100101110", -- t[52526] = 15
      "0001111" when "01100110100101111", -- t[52527] = 15
      "0001111" when "01100110100110000", -- t[52528] = 15
      "0001111" when "01100110100110001", -- t[52529] = 15
      "0001111" when "01100110100110010", -- t[52530] = 15
      "0001111" when "01100110100110011", -- t[52531] = 15
      "0001111" when "01100110100110100", -- t[52532] = 15
      "0001111" when "01100110100110101", -- t[52533] = 15
      "0001111" when "01100110100110110", -- t[52534] = 15
      "0001111" when "01100110100110111", -- t[52535] = 15
      "0001111" when "01100110100111000", -- t[52536] = 15
      "0001111" when "01100110100111001", -- t[52537] = 15
      "0001111" when "01100110100111010", -- t[52538] = 15
      "0001111" when "01100110100111011", -- t[52539] = 15
      "0001111" when "01100110100111100", -- t[52540] = 15
      "0001111" when "01100110100111101", -- t[52541] = 15
      "0001111" when "01100110100111110", -- t[52542] = 15
      "0001111" when "01100110100111111", -- t[52543] = 15
      "0001111" when "01100110101000000", -- t[52544] = 15
      "0001111" when "01100110101000001", -- t[52545] = 15
      "0001111" when "01100110101000010", -- t[52546] = 15
      "0001111" when "01100110101000011", -- t[52547] = 15
      "0001111" when "01100110101000100", -- t[52548] = 15
      "0001111" when "01100110101000101", -- t[52549] = 15
      "0001111" when "01100110101000110", -- t[52550] = 15
      "0001111" when "01100110101000111", -- t[52551] = 15
      "0001111" when "01100110101001000", -- t[52552] = 15
      "0001111" when "01100110101001001", -- t[52553] = 15
      "0001111" when "01100110101001010", -- t[52554] = 15
      "0001111" when "01100110101001011", -- t[52555] = 15
      "0001111" when "01100110101001100", -- t[52556] = 15
      "0001111" when "01100110101001101", -- t[52557] = 15
      "0001111" when "01100110101001110", -- t[52558] = 15
      "0001111" when "01100110101001111", -- t[52559] = 15
      "0001111" when "01100110101010000", -- t[52560] = 15
      "0001111" when "01100110101010001", -- t[52561] = 15
      "0001111" when "01100110101010010", -- t[52562] = 15
      "0001111" when "01100110101010011", -- t[52563] = 15
      "0001111" when "01100110101010100", -- t[52564] = 15
      "0001111" when "01100110101010101", -- t[52565] = 15
      "0001111" when "01100110101010110", -- t[52566] = 15
      "0001111" when "01100110101010111", -- t[52567] = 15
      "0001111" when "01100110101011000", -- t[52568] = 15
      "0001111" when "01100110101011001", -- t[52569] = 15
      "0001111" when "01100110101011010", -- t[52570] = 15
      "0001111" when "01100110101011011", -- t[52571] = 15
      "0001111" when "01100110101011100", -- t[52572] = 15
      "0001111" when "01100110101011101", -- t[52573] = 15
      "0001111" when "01100110101011110", -- t[52574] = 15
      "0001111" when "01100110101011111", -- t[52575] = 15
      "0001111" when "01100110101100000", -- t[52576] = 15
      "0001111" when "01100110101100001", -- t[52577] = 15
      "0001111" when "01100110101100010", -- t[52578] = 15
      "0001111" when "01100110101100011", -- t[52579] = 15
      "0001111" when "01100110101100100", -- t[52580] = 15
      "0001111" when "01100110101100101", -- t[52581] = 15
      "0001111" when "01100110101100110", -- t[52582] = 15
      "0001111" when "01100110101100111", -- t[52583] = 15
      "0001111" when "01100110101101000", -- t[52584] = 15
      "0001111" when "01100110101101001", -- t[52585] = 15
      "0001111" when "01100110101101010", -- t[52586] = 15
      "0001111" when "01100110101101011", -- t[52587] = 15
      "0001111" when "01100110101101100", -- t[52588] = 15
      "0001111" when "01100110101101101", -- t[52589] = 15
      "0001111" when "01100110101101110", -- t[52590] = 15
      "0001111" when "01100110101101111", -- t[52591] = 15
      "0001111" when "01100110101110000", -- t[52592] = 15
      "0001111" when "01100110101110001", -- t[52593] = 15
      "0001111" when "01100110101110010", -- t[52594] = 15
      "0001111" when "01100110101110011", -- t[52595] = 15
      "0001111" when "01100110101110100", -- t[52596] = 15
      "0001111" when "01100110101110101", -- t[52597] = 15
      "0001111" when "01100110101110110", -- t[52598] = 15
      "0001111" when "01100110101110111", -- t[52599] = 15
      "0001111" when "01100110101111000", -- t[52600] = 15
      "0001111" when "01100110101111001", -- t[52601] = 15
      "0001111" when "01100110101111010", -- t[52602] = 15
      "0001111" when "01100110101111011", -- t[52603] = 15
      "0001111" when "01100110101111100", -- t[52604] = 15
      "0001111" when "01100110101111101", -- t[52605] = 15
      "0001111" when "01100110101111110", -- t[52606] = 15
      "0001111" when "01100110101111111", -- t[52607] = 15
      "0001111" when "01100110110000000", -- t[52608] = 15
      "0001111" when "01100110110000001", -- t[52609] = 15
      "0001111" when "01100110110000010", -- t[52610] = 15
      "0001111" when "01100110110000011", -- t[52611] = 15
      "0001111" when "01100110110000100", -- t[52612] = 15
      "0001111" when "01100110110000101", -- t[52613] = 15
      "0001111" when "01100110110000110", -- t[52614] = 15
      "0001111" when "01100110110000111", -- t[52615] = 15
      "0001111" when "01100110110001000", -- t[52616] = 15
      "0001111" when "01100110110001001", -- t[52617] = 15
      "0001111" when "01100110110001010", -- t[52618] = 15
      "0001111" when "01100110110001011", -- t[52619] = 15
      "0001111" when "01100110110001100", -- t[52620] = 15
      "0001111" when "01100110110001101", -- t[52621] = 15
      "0001111" when "01100110110001110", -- t[52622] = 15
      "0001111" when "01100110110001111", -- t[52623] = 15
      "0001111" when "01100110110010000", -- t[52624] = 15
      "0001111" when "01100110110010001", -- t[52625] = 15
      "0001111" when "01100110110010010", -- t[52626] = 15
      "0001111" when "01100110110010011", -- t[52627] = 15
      "0001111" when "01100110110010100", -- t[52628] = 15
      "0001111" when "01100110110010101", -- t[52629] = 15
      "0010000" when "01100110110010110", -- t[52630] = 16
      "0010000" when "01100110110010111", -- t[52631] = 16
      "0010000" when "01100110110011000", -- t[52632] = 16
      "0010000" when "01100110110011001", -- t[52633] = 16
      "0010000" when "01100110110011010", -- t[52634] = 16
      "0010000" when "01100110110011011", -- t[52635] = 16
      "0010000" when "01100110110011100", -- t[52636] = 16
      "0010000" when "01100110110011101", -- t[52637] = 16
      "0010000" when "01100110110011110", -- t[52638] = 16
      "0010000" when "01100110110011111", -- t[52639] = 16
      "0010000" when "01100110110100000", -- t[52640] = 16
      "0010000" when "01100110110100001", -- t[52641] = 16
      "0010000" when "01100110110100010", -- t[52642] = 16
      "0010000" when "01100110110100011", -- t[52643] = 16
      "0010000" when "01100110110100100", -- t[52644] = 16
      "0010000" when "01100110110100101", -- t[52645] = 16
      "0010000" when "01100110110100110", -- t[52646] = 16
      "0010000" when "01100110110100111", -- t[52647] = 16
      "0010000" when "01100110110101000", -- t[52648] = 16
      "0010000" when "01100110110101001", -- t[52649] = 16
      "0010000" when "01100110110101010", -- t[52650] = 16
      "0010000" when "01100110110101011", -- t[52651] = 16
      "0010000" when "01100110110101100", -- t[52652] = 16
      "0010000" when "01100110110101101", -- t[52653] = 16
      "0010000" when "01100110110101110", -- t[52654] = 16
      "0010000" when "01100110110101111", -- t[52655] = 16
      "0010000" when "01100110110110000", -- t[52656] = 16
      "0010000" when "01100110110110001", -- t[52657] = 16
      "0010000" when "01100110110110010", -- t[52658] = 16
      "0010000" when "01100110110110011", -- t[52659] = 16
      "0010000" when "01100110110110100", -- t[52660] = 16
      "0010000" when "01100110110110101", -- t[52661] = 16
      "0010000" when "01100110110110110", -- t[52662] = 16
      "0010000" when "01100110110110111", -- t[52663] = 16
      "0010000" when "01100110110111000", -- t[52664] = 16
      "0010000" when "01100110110111001", -- t[52665] = 16
      "0010000" when "01100110110111010", -- t[52666] = 16
      "0010000" when "01100110110111011", -- t[52667] = 16
      "0010000" when "01100110110111100", -- t[52668] = 16
      "0010000" when "01100110110111101", -- t[52669] = 16
      "0010000" when "01100110110111110", -- t[52670] = 16
      "0010000" when "01100110110111111", -- t[52671] = 16
      "0010000" when "01100110111000000", -- t[52672] = 16
      "0010000" when "01100110111000001", -- t[52673] = 16
      "0010000" when "01100110111000010", -- t[52674] = 16
      "0010000" when "01100110111000011", -- t[52675] = 16
      "0010000" when "01100110111000100", -- t[52676] = 16
      "0010000" when "01100110111000101", -- t[52677] = 16
      "0010000" when "01100110111000110", -- t[52678] = 16
      "0010000" when "01100110111000111", -- t[52679] = 16
      "0010000" when "01100110111001000", -- t[52680] = 16
      "0010000" when "01100110111001001", -- t[52681] = 16
      "0010000" when "01100110111001010", -- t[52682] = 16
      "0010000" when "01100110111001011", -- t[52683] = 16
      "0010000" when "01100110111001100", -- t[52684] = 16
      "0010000" when "01100110111001101", -- t[52685] = 16
      "0010000" when "01100110111001110", -- t[52686] = 16
      "0010000" when "01100110111001111", -- t[52687] = 16
      "0010000" when "01100110111010000", -- t[52688] = 16
      "0010000" when "01100110111010001", -- t[52689] = 16
      "0010000" when "01100110111010010", -- t[52690] = 16
      "0010000" when "01100110111010011", -- t[52691] = 16
      "0010000" when "01100110111010100", -- t[52692] = 16
      "0010000" when "01100110111010101", -- t[52693] = 16
      "0010000" when "01100110111010110", -- t[52694] = 16
      "0010000" when "01100110111010111", -- t[52695] = 16
      "0010000" when "01100110111011000", -- t[52696] = 16
      "0010000" when "01100110111011001", -- t[52697] = 16
      "0010000" when "01100110111011010", -- t[52698] = 16
      "0010000" when "01100110111011011", -- t[52699] = 16
      "0010000" when "01100110111011100", -- t[52700] = 16
      "0010000" when "01100110111011101", -- t[52701] = 16
      "0010000" when "01100110111011110", -- t[52702] = 16
      "0010000" when "01100110111011111", -- t[52703] = 16
      "0010000" when "01100110111100000", -- t[52704] = 16
      "0010000" when "01100110111100001", -- t[52705] = 16
      "0010000" when "01100110111100010", -- t[52706] = 16
      "0010000" when "01100110111100011", -- t[52707] = 16
      "0010000" when "01100110111100100", -- t[52708] = 16
      "0010000" when "01100110111100101", -- t[52709] = 16
      "0010000" when "01100110111100110", -- t[52710] = 16
      "0010000" when "01100110111100111", -- t[52711] = 16
      "0010000" when "01100110111101000", -- t[52712] = 16
      "0010000" when "01100110111101001", -- t[52713] = 16
      "0010000" when "01100110111101010", -- t[52714] = 16
      "0010000" when "01100110111101011", -- t[52715] = 16
      "0010000" when "01100110111101100", -- t[52716] = 16
      "0010000" when "01100110111101101", -- t[52717] = 16
      "0010000" when "01100110111101110", -- t[52718] = 16
      "0010000" when "01100110111101111", -- t[52719] = 16
      "0010000" when "01100110111110000", -- t[52720] = 16
      "0010000" when "01100110111110001", -- t[52721] = 16
      "0010000" when "01100110111110010", -- t[52722] = 16
      "0010000" when "01100110111110011", -- t[52723] = 16
      "0010000" when "01100110111110100", -- t[52724] = 16
      "0010000" when "01100110111110101", -- t[52725] = 16
      "0010000" when "01100110111110110", -- t[52726] = 16
      "0010000" when "01100110111110111", -- t[52727] = 16
      "0010000" when "01100110111111000", -- t[52728] = 16
      "0010000" when "01100110111111001", -- t[52729] = 16
      "0010000" when "01100110111111010", -- t[52730] = 16
      "0010000" when "01100110111111011", -- t[52731] = 16
      "0010000" when "01100110111111100", -- t[52732] = 16
      "0010000" when "01100110111111101", -- t[52733] = 16
      "0010000" when "01100110111111110", -- t[52734] = 16
      "0010000" when "01100110111111111", -- t[52735] = 16
      "0010000" when "01100111000000000", -- t[52736] = 16
      "0010000" when "01100111000000001", -- t[52737] = 16
      "0010000" when "01100111000000010", -- t[52738] = 16
      "0010000" when "01100111000000011", -- t[52739] = 16
      "0010000" when "01100111000000100", -- t[52740] = 16
      "0010000" when "01100111000000101", -- t[52741] = 16
      "0010000" when "01100111000000110", -- t[52742] = 16
      "0010000" when "01100111000000111", -- t[52743] = 16
      "0010000" when "01100111000001000", -- t[52744] = 16
      "0010000" when "01100111000001001", -- t[52745] = 16
      "0010000" when "01100111000001010", -- t[52746] = 16
      "0010000" when "01100111000001011", -- t[52747] = 16
      "0010000" when "01100111000001100", -- t[52748] = 16
      "0010000" when "01100111000001101", -- t[52749] = 16
      "0010000" when "01100111000001110", -- t[52750] = 16
      "0010000" when "01100111000001111", -- t[52751] = 16
      "0010000" when "01100111000010000", -- t[52752] = 16
      "0010000" when "01100111000010001", -- t[52753] = 16
      "0010000" when "01100111000010010", -- t[52754] = 16
      "0010000" when "01100111000010011", -- t[52755] = 16
      "0010000" when "01100111000010100", -- t[52756] = 16
      "0010000" when "01100111000010101", -- t[52757] = 16
      "0010000" when "01100111000010110", -- t[52758] = 16
      "0010000" when "01100111000010111", -- t[52759] = 16
      "0010000" when "01100111000011000", -- t[52760] = 16
      "0010000" when "01100111000011001", -- t[52761] = 16
      "0010000" when "01100111000011010", -- t[52762] = 16
      "0010000" when "01100111000011011", -- t[52763] = 16
      "0010000" when "01100111000011100", -- t[52764] = 16
      "0010000" when "01100111000011101", -- t[52765] = 16
      "0010000" when "01100111000011110", -- t[52766] = 16
      "0010000" when "01100111000011111", -- t[52767] = 16
      "0010000" when "01100111000100000", -- t[52768] = 16
      "0010000" when "01100111000100001", -- t[52769] = 16
      "0010000" when "01100111000100010", -- t[52770] = 16
      "0010000" when "01100111000100011", -- t[52771] = 16
      "0010000" when "01100111000100100", -- t[52772] = 16
      "0010000" when "01100111000100101", -- t[52773] = 16
      "0010000" when "01100111000100110", -- t[52774] = 16
      "0010000" when "01100111000100111", -- t[52775] = 16
      "0010000" when "01100111000101000", -- t[52776] = 16
      "0010000" when "01100111000101001", -- t[52777] = 16
      "0010000" when "01100111000101010", -- t[52778] = 16
      "0010000" when "01100111000101011", -- t[52779] = 16
      "0010000" when "01100111000101100", -- t[52780] = 16
      "0010000" when "01100111000101101", -- t[52781] = 16
      "0010000" when "01100111000101110", -- t[52782] = 16
      "0010000" when "01100111000101111", -- t[52783] = 16
      "0010000" when "01100111000110000", -- t[52784] = 16
      "0010000" when "01100111000110001", -- t[52785] = 16
      "0010000" when "01100111000110010", -- t[52786] = 16
      "0010000" when "01100111000110011", -- t[52787] = 16
      "0010000" when "01100111000110100", -- t[52788] = 16
      "0010000" when "01100111000110101", -- t[52789] = 16
      "0010000" when "01100111000110110", -- t[52790] = 16
      "0010000" when "01100111000110111", -- t[52791] = 16
      "0010000" when "01100111000111000", -- t[52792] = 16
      "0010000" when "01100111000111001", -- t[52793] = 16
      "0010000" when "01100111000111010", -- t[52794] = 16
      "0010000" when "01100111000111011", -- t[52795] = 16
      "0010000" when "01100111000111100", -- t[52796] = 16
      "0010000" when "01100111000111101", -- t[52797] = 16
      "0010000" when "01100111000111110", -- t[52798] = 16
      "0010000" when "01100111000111111", -- t[52799] = 16
      "0010000" when "01100111001000000", -- t[52800] = 16
      "0010000" when "01100111001000001", -- t[52801] = 16
      "0010000" when "01100111001000010", -- t[52802] = 16
      "0010000" when "01100111001000011", -- t[52803] = 16
      "0010000" when "01100111001000100", -- t[52804] = 16
      "0010000" when "01100111001000101", -- t[52805] = 16
      "0010000" when "01100111001000110", -- t[52806] = 16
      "0010000" when "01100111001000111", -- t[52807] = 16
      "0010000" when "01100111001001000", -- t[52808] = 16
      "0010000" when "01100111001001001", -- t[52809] = 16
      "0010000" when "01100111001001010", -- t[52810] = 16
      "0010000" when "01100111001001011", -- t[52811] = 16
      "0010000" when "01100111001001100", -- t[52812] = 16
      "0010000" when "01100111001001101", -- t[52813] = 16
      "0010000" when "01100111001001110", -- t[52814] = 16
      "0010000" when "01100111001001111", -- t[52815] = 16
      "0010000" when "01100111001010000", -- t[52816] = 16
      "0010000" when "01100111001010001", -- t[52817] = 16
      "0010000" when "01100111001010010", -- t[52818] = 16
      "0010000" when "01100111001010011", -- t[52819] = 16
      "0010000" when "01100111001010100", -- t[52820] = 16
      "0010000" when "01100111001010101", -- t[52821] = 16
      "0010000" when "01100111001010110", -- t[52822] = 16
      "0010000" when "01100111001010111", -- t[52823] = 16
      "0010000" when "01100111001011000", -- t[52824] = 16
      "0010000" when "01100111001011001", -- t[52825] = 16
      "0010000" when "01100111001011010", -- t[52826] = 16
      "0010000" when "01100111001011011", -- t[52827] = 16
      "0010000" when "01100111001011100", -- t[52828] = 16
      "0010000" when "01100111001011101", -- t[52829] = 16
      "0010000" when "01100111001011110", -- t[52830] = 16
      "0010000" when "01100111001011111", -- t[52831] = 16
      "0010000" when "01100111001100000", -- t[52832] = 16
      "0010000" when "01100111001100001", -- t[52833] = 16
      "0010000" when "01100111001100010", -- t[52834] = 16
      "0010000" when "01100111001100011", -- t[52835] = 16
      "0010000" when "01100111001100100", -- t[52836] = 16
      "0010000" when "01100111001100101", -- t[52837] = 16
      "0010000" when "01100111001100110", -- t[52838] = 16
      "0010000" when "01100111001100111", -- t[52839] = 16
      "0010000" when "01100111001101000", -- t[52840] = 16
      "0010000" when "01100111001101001", -- t[52841] = 16
      "0010000" when "01100111001101010", -- t[52842] = 16
      "0010000" when "01100111001101011", -- t[52843] = 16
      "0010000" when "01100111001101100", -- t[52844] = 16
      "0010000" when "01100111001101101", -- t[52845] = 16
      "0010000" when "01100111001101110", -- t[52846] = 16
      "0010000" when "01100111001101111", -- t[52847] = 16
      "0010000" when "01100111001110000", -- t[52848] = 16
      "0010000" when "01100111001110001", -- t[52849] = 16
      "0010000" when "01100111001110010", -- t[52850] = 16
      "0010000" when "01100111001110011", -- t[52851] = 16
      "0010000" when "01100111001110100", -- t[52852] = 16
      "0010000" when "01100111001110101", -- t[52853] = 16
      "0010000" when "01100111001110110", -- t[52854] = 16
      "0010000" when "01100111001110111", -- t[52855] = 16
      "0010000" when "01100111001111000", -- t[52856] = 16
      "0010000" when "01100111001111001", -- t[52857] = 16
      "0010000" when "01100111001111010", -- t[52858] = 16
      "0010000" when "01100111001111011", -- t[52859] = 16
      "0010000" when "01100111001111100", -- t[52860] = 16
      "0010000" when "01100111001111101", -- t[52861] = 16
      "0010000" when "01100111001111110", -- t[52862] = 16
      "0010000" when "01100111001111111", -- t[52863] = 16
      "0010000" when "01100111010000000", -- t[52864] = 16
      "0010000" when "01100111010000001", -- t[52865] = 16
      "0010000" when "01100111010000010", -- t[52866] = 16
      "0010000" when "01100111010000011", -- t[52867] = 16
      "0010000" when "01100111010000100", -- t[52868] = 16
      "0010000" when "01100111010000101", -- t[52869] = 16
      "0010000" when "01100111010000110", -- t[52870] = 16
      "0010000" when "01100111010000111", -- t[52871] = 16
      "0010000" when "01100111010001000", -- t[52872] = 16
      "0010000" when "01100111010001001", -- t[52873] = 16
      "0010000" when "01100111010001010", -- t[52874] = 16
      "0010000" when "01100111010001011", -- t[52875] = 16
      "0010000" when "01100111010001100", -- t[52876] = 16
      "0010000" when "01100111010001101", -- t[52877] = 16
      "0010000" when "01100111010001110", -- t[52878] = 16
      "0010000" when "01100111010001111", -- t[52879] = 16
      "0010000" when "01100111010010000", -- t[52880] = 16
      "0010000" when "01100111010010001", -- t[52881] = 16
      "0010000" when "01100111010010010", -- t[52882] = 16
      "0010000" when "01100111010010011", -- t[52883] = 16
      "0010000" when "01100111010010100", -- t[52884] = 16
      "0010000" when "01100111010010101", -- t[52885] = 16
      "0010000" when "01100111010010110", -- t[52886] = 16
      "0010000" when "01100111010010111", -- t[52887] = 16
      "0010000" when "01100111010011000", -- t[52888] = 16
      "0010000" when "01100111010011001", -- t[52889] = 16
      "0010000" when "01100111010011010", -- t[52890] = 16
      "0010000" when "01100111010011011", -- t[52891] = 16
      "0010000" when "01100111010011100", -- t[52892] = 16
      "0010000" when "01100111010011101", -- t[52893] = 16
      "0010000" when "01100111010011110", -- t[52894] = 16
      "0010000" when "01100111010011111", -- t[52895] = 16
      "0010000" when "01100111010100000", -- t[52896] = 16
      "0010000" when "01100111010100001", -- t[52897] = 16
      "0010000" when "01100111010100010", -- t[52898] = 16
      "0010000" when "01100111010100011", -- t[52899] = 16
      "0010000" when "01100111010100100", -- t[52900] = 16
      "0010000" when "01100111010100101", -- t[52901] = 16
      "0010000" when "01100111010100110", -- t[52902] = 16
      "0010000" when "01100111010100111", -- t[52903] = 16
      "0010000" when "01100111010101000", -- t[52904] = 16
      "0010000" when "01100111010101001", -- t[52905] = 16
      "0010000" when "01100111010101010", -- t[52906] = 16
      "0010000" when "01100111010101011", -- t[52907] = 16
      "0010000" when "01100111010101100", -- t[52908] = 16
      "0010000" when "01100111010101101", -- t[52909] = 16
      "0010000" when "01100111010101110", -- t[52910] = 16
      "0010000" when "01100111010101111", -- t[52911] = 16
      "0010000" when "01100111010110000", -- t[52912] = 16
      "0010000" when "01100111010110001", -- t[52913] = 16
      "0010000" when "01100111010110010", -- t[52914] = 16
      "0010000" when "01100111010110011", -- t[52915] = 16
      "0010000" when "01100111010110100", -- t[52916] = 16
      "0010000" when "01100111010110101", -- t[52917] = 16
      "0010000" when "01100111010110110", -- t[52918] = 16
      "0010000" when "01100111010110111", -- t[52919] = 16
      "0010000" when "01100111010111000", -- t[52920] = 16
      "0010000" when "01100111010111001", -- t[52921] = 16
      "0010000" when "01100111010111010", -- t[52922] = 16
      "0010000" when "01100111010111011", -- t[52923] = 16
      "0010000" when "01100111010111100", -- t[52924] = 16
      "0010000" when "01100111010111101", -- t[52925] = 16
      "0010000" when "01100111010111110", -- t[52926] = 16
      "0010000" when "01100111010111111", -- t[52927] = 16
      "0010000" when "01100111011000000", -- t[52928] = 16
      "0010000" when "01100111011000001", -- t[52929] = 16
      "0010000" when "01100111011000010", -- t[52930] = 16
      "0010000" when "01100111011000011", -- t[52931] = 16
      "0010000" when "01100111011000100", -- t[52932] = 16
      "0010000" when "01100111011000101", -- t[52933] = 16
      "0010000" when "01100111011000110", -- t[52934] = 16
      "0010000" when "01100111011000111", -- t[52935] = 16
      "0010000" when "01100111011001000", -- t[52936] = 16
      "0010000" when "01100111011001001", -- t[52937] = 16
      "0010000" when "01100111011001010", -- t[52938] = 16
      "0010000" when "01100111011001011", -- t[52939] = 16
      "0010000" when "01100111011001100", -- t[52940] = 16
      "0010000" when "01100111011001101", -- t[52941] = 16
      "0010000" when "01100111011001110", -- t[52942] = 16
      "0010000" when "01100111011001111", -- t[52943] = 16
      "0010000" when "01100111011010000", -- t[52944] = 16
      "0010000" when "01100111011010001", -- t[52945] = 16
      "0010000" when "01100111011010010", -- t[52946] = 16
      "0010000" when "01100111011010011", -- t[52947] = 16
      "0010000" when "01100111011010100", -- t[52948] = 16
      "0010000" when "01100111011010101", -- t[52949] = 16
      "0010000" when "01100111011010110", -- t[52950] = 16
      "0010000" when "01100111011010111", -- t[52951] = 16
      "0010000" when "01100111011011000", -- t[52952] = 16
      "0010000" when "01100111011011001", -- t[52953] = 16
      "0010000" when "01100111011011010", -- t[52954] = 16
      "0010000" when "01100111011011011", -- t[52955] = 16
      "0010000" when "01100111011011100", -- t[52956] = 16
      "0010000" when "01100111011011101", -- t[52957] = 16
      "0010000" when "01100111011011110", -- t[52958] = 16
      "0010000" when "01100111011011111", -- t[52959] = 16
      "0010000" when "01100111011100000", -- t[52960] = 16
      "0010000" when "01100111011100001", -- t[52961] = 16
      "0010000" when "01100111011100010", -- t[52962] = 16
      "0010000" when "01100111011100011", -- t[52963] = 16
      "0010000" when "01100111011100100", -- t[52964] = 16
      "0010000" when "01100111011100101", -- t[52965] = 16
      "0010000" when "01100111011100110", -- t[52966] = 16
      "0010000" when "01100111011100111", -- t[52967] = 16
      "0010000" when "01100111011101000", -- t[52968] = 16
      "0010000" when "01100111011101001", -- t[52969] = 16
      "0010000" when "01100111011101010", -- t[52970] = 16
      "0010000" when "01100111011101011", -- t[52971] = 16
      "0010000" when "01100111011101100", -- t[52972] = 16
      "0010000" when "01100111011101101", -- t[52973] = 16
      "0010000" when "01100111011101110", -- t[52974] = 16
      "0010000" when "01100111011101111", -- t[52975] = 16
      "0010000" when "01100111011110000", -- t[52976] = 16
      "0010000" when "01100111011110001", -- t[52977] = 16
      "0010000" when "01100111011110010", -- t[52978] = 16
      "0010000" when "01100111011110011", -- t[52979] = 16
      "0010000" when "01100111011110100", -- t[52980] = 16
      "0010000" when "01100111011110101", -- t[52981] = 16
      "0010000" when "01100111011110110", -- t[52982] = 16
      "0010000" when "01100111011110111", -- t[52983] = 16
      "0010000" when "01100111011111000", -- t[52984] = 16
      "0010000" when "01100111011111001", -- t[52985] = 16
      "0010000" when "01100111011111010", -- t[52986] = 16
      "0010000" when "01100111011111011", -- t[52987] = 16
      "0010000" when "01100111011111100", -- t[52988] = 16
      "0010000" when "01100111011111101", -- t[52989] = 16
      "0010000" when "01100111011111110", -- t[52990] = 16
      "0010000" when "01100111011111111", -- t[52991] = 16
      "0010000" when "01100111100000000", -- t[52992] = 16
      "0010000" when "01100111100000001", -- t[52993] = 16
      "0010000" when "01100111100000010", -- t[52994] = 16
      "0010000" when "01100111100000011", -- t[52995] = 16
      "0010000" when "01100111100000100", -- t[52996] = 16
      "0010000" when "01100111100000101", -- t[52997] = 16
      "0010000" when "01100111100000110", -- t[52998] = 16
      "0010000" when "01100111100000111", -- t[52999] = 16
      "0010000" when "01100111100001000", -- t[53000] = 16
      "0010000" when "01100111100001001", -- t[53001] = 16
      "0010000" when "01100111100001010", -- t[53002] = 16
      "0010000" when "01100111100001011", -- t[53003] = 16
      "0010000" when "01100111100001100", -- t[53004] = 16
      "0010000" when "01100111100001101", -- t[53005] = 16
      "0010000" when "01100111100001110", -- t[53006] = 16
      "0010000" when "01100111100001111", -- t[53007] = 16
      "0010000" when "01100111100010000", -- t[53008] = 16
      "0010000" when "01100111100010001", -- t[53009] = 16
      "0010000" when "01100111100010010", -- t[53010] = 16
      "0010000" when "01100111100010011", -- t[53011] = 16
      "0010000" when "01100111100010100", -- t[53012] = 16
      "0010000" when "01100111100010101", -- t[53013] = 16
      "0010000" when "01100111100010110", -- t[53014] = 16
      "0010000" when "01100111100010111", -- t[53015] = 16
      "0010000" when "01100111100011000", -- t[53016] = 16
      "0010000" when "01100111100011001", -- t[53017] = 16
      "0010000" when "01100111100011010", -- t[53018] = 16
      "0010000" when "01100111100011011", -- t[53019] = 16
      "0010000" when "01100111100011100", -- t[53020] = 16
      "0010000" when "01100111100011101", -- t[53021] = 16
      "0010000" when "01100111100011110", -- t[53022] = 16
      "0010000" when "01100111100011111", -- t[53023] = 16
      "0010000" when "01100111100100000", -- t[53024] = 16
      "0010000" when "01100111100100001", -- t[53025] = 16
      "0010000" when "01100111100100010", -- t[53026] = 16
      "0010000" when "01100111100100011", -- t[53027] = 16
      "0010000" when "01100111100100100", -- t[53028] = 16
      "0010000" when "01100111100100101", -- t[53029] = 16
      "0010000" when "01100111100100110", -- t[53030] = 16
      "0010000" when "01100111100100111", -- t[53031] = 16
      "0010000" when "01100111100101000", -- t[53032] = 16
      "0010000" when "01100111100101001", -- t[53033] = 16
      "0010000" when "01100111100101010", -- t[53034] = 16
      "0010000" when "01100111100101011", -- t[53035] = 16
      "0010000" when "01100111100101100", -- t[53036] = 16
      "0010000" when "01100111100101101", -- t[53037] = 16
      "0010000" when "01100111100101110", -- t[53038] = 16
      "0010000" when "01100111100101111", -- t[53039] = 16
      "0010000" when "01100111100110000", -- t[53040] = 16
      "0010000" when "01100111100110001", -- t[53041] = 16
      "0010000" when "01100111100110010", -- t[53042] = 16
      "0010000" when "01100111100110011", -- t[53043] = 16
      "0010000" when "01100111100110100", -- t[53044] = 16
      "0010000" when "01100111100110101", -- t[53045] = 16
      "0010000" when "01100111100110110", -- t[53046] = 16
      "0010000" when "01100111100110111", -- t[53047] = 16
      "0010000" when "01100111100111000", -- t[53048] = 16
      "0010000" when "01100111100111001", -- t[53049] = 16
      "0010000" when "01100111100111010", -- t[53050] = 16
      "0010000" when "01100111100111011", -- t[53051] = 16
      "0010000" when "01100111100111100", -- t[53052] = 16
      "0010000" when "01100111100111101", -- t[53053] = 16
      "0010000" when "01100111100111110", -- t[53054] = 16
      "0010000" when "01100111100111111", -- t[53055] = 16
      "0010000" when "01100111101000000", -- t[53056] = 16
      "0010000" when "01100111101000001", -- t[53057] = 16
      "0010000" when "01100111101000010", -- t[53058] = 16
      "0010000" when "01100111101000011", -- t[53059] = 16
      "0010000" when "01100111101000100", -- t[53060] = 16
      "0010000" when "01100111101000101", -- t[53061] = 16
      "0010000" when "01100111101000110", -- t[53062] = 16
      "0010000" when "01100111101000111", -- t[53063] = 16
      "0010000" when "01100111101001000", -- t[53064] = 16
      "0010000" when "01100111101001001", -- t[53065] = 16
      "0010000" when "01100111101001010", -- t[53066] = 16
      "0010000" when "01100111101001011", -- t[53067] = 16
      "0010000" when "01100111101001100", -- t[53068] = 16
      "0010000" when "01100111101001101", -- t[53069] = 16
      "0010000" when "01100111101001110", -- t[53070] = 16
      "0010000" when "01100111101001111", -- t[53071] = 16
      "0010000" when "01100111101010000", -- t[53072] = 16
      "0010000" when "01100111101010001", -- t[53073] = 16
      "0010000" when "01100111101010010", -- t[53074] = 16
      "0010000" when "01100111101010011", -- t[53075] = 16
      "0010000" when "01100111101010100", -- t[53076] = 16
      "0010000" when "01100111101010101", -- t[53077] = 16
      "0010000" when "01100111101010110", -- t[53078] = 16
      "0010000" when "01100111101010111", -- t[53079] = 16
      "0010000" when "01100111101011000", -- t[53080] = 16
      "0010000" when "01100111101011001", -- t[53081] = 16
      "0010000" when "01100111101011010", -- t[53082] = 16
      "0010000" when "01100111101011011", -- t[53083] = 16
      "0010000" when "01100111101011100", -- t[53084] = 16
      "0010000" when "01100111101011101", -- t[53085] = 16
      "0010000" when "01100111101011110", -- t[53086] = 16
      "0010000" when "01100111101011111", -- t[53087] = 16
      "0010000" when "01100111101100000", -- t[53088] = 16
      "0010000" when "01100111101100001", -- t[53089] = 16
      "0010000" when "01100111101100010", -- t[53090] = 16
      "0010000" when "01100111101100011", -- t[53091] = 16
      "0010000" when "01100111101100100", -- t[53092] = 16
      "0010000" when "01100111101100101", -- t[53093] = 16
      "0010000" when "01100111101100110", -- t[53094] = 16
      "0010000" when "01100111101100111", -- t[53095] = 16
      "0010000" when "01100111101101000", -- t[53096] = 16
      "0010000" when "01100111101101001", -- t[53097] = 16
      "0010000" when "01100111101101010", -- t[53098] = 16
      "0010000" when "01100111101101011", -- t[53099] = 16
      "0010000" when "01100111101101100", -- t[53100] = 16
      "0010000" when "01100111101101101", -- t[53101] = 16
      "0010000" when "01100111101101110", -- t[53102] = 16
      "0010000" when "01100111101101111", -- t[53103] = 16
      "0010000" when "01100111101110000", -- t[53104] = 16
      "0010000" when "01100111101110001", -- t[53105] = 16
      "0010000" when "01100111101110010", -- t[53106] = 16
      "0010000" when "01100111101110011", -- t[53107] = 16
      "0010000" when "01100111101110100", -- t[53108] = 16
      "0010000" when "01100111101110101", -- t[53109] = 16
      "0010000" when "01100111101110110", -- t[53110] = 16
      "0010000" when "01100111101110111", -- t[53111] = 16
      "0010000" when "01100111101111000", -- t[53112] = 16
      "0010000" when "01100111101111001", -- t[53113] = 16
      "0010000" when "01100111101111010", -- t[53114] = 16
      "0010000" when "01100111101111011", -- t[53115] = 16
      "0010000" when "01100111101111100", -- t[53116] = 16
      "0010000" when "01100111101111101", -- t[53117] = 16
      "0010000" when "01100111101111110", -- t[53118] = 16
      "0010000" when "01100111101111111", -- t[53119] = 16
      "0010000" when "01100111110000000", -- t[53120] = 16
      "0010000" when "01100111110000001", -- t[53121] = 16
      "0010000" when "01100111110000010", -- t[53122] = 16
      "0010000" when "01100111110000011", -- t[53123] = 16
      "0010000" when "01100111110000100", -- t[53124] = 16
      "0010000" when "01100111110000101", -- t[53125] = 16
      "0010000" when "01100111110000110", -- t[53126] = 16
      "0010000" when "01100111110000111", -- t[53127] = 16
      "0010000" when "01100111110001000", -- t[53128] = 16
      "0010000" when "01100111110001001", -- t[53129] = 16
      "0010000" when "01100111110001010", -- t[53130] = 16
      "0010000" when "01100111110001011", -- t[53131] = 16
      "0010000" when "01100111110001100", -- t[53132] = 16
      "0010000" when "01100111110001101", -- t[53133] = 16
      "0010000" when "01100111110001110", -- t[53134] = 16
      "0010000" when "01100111110001111", -- t[53135] = 16
      "0010000" when "01100111110010000", -- t[53136] = 16
      "0010000" when "01100111110010001", -- t[53137] = 16
      "0010000" when "01100111110010010", -- t[53138] = 16
      "0010000" when "01100111110010011", -- t[53139] = 16
      "0010000" when "01100111110010100", -- t[53140] = 16
      "0010000" when "01100111110010101", -- t[53141] = 16
      "0010000" when "01100111110010110", -- t[53142] = 16
      "0010000" when "01100111110010111", -- t[53143] = 16
      "0010000" when "01100111110011000", -- t[53144] = 16
      "0010000" when "01100111110011001", -- t[53145] = 16
      "0010000" when "01100111110011010", -- t[53146] = 16
      "0010000" when "01100111110011011", -- t[53147] = 16
      "0010000" when "01100111110011100", -- t[53148] = 16
      "0010000" when "01100111110011101", -- t[53149] = 16
      "0010000" when "01100111110011110", -- t[53150] = 16
      "0010000" when "01100111110011111", -- t[53151] = 16
      "0010000" when "01100111110100000", -- t[53152] = 16
      "0010000" when "01100111110100001", -- t[53153] = 16
      "0010000" when "01100111110100010", -- t[53154] = 16
      "0010000" when "01100111110100011", -- t[53155] = 16
      "0010000" when "01100111110100100", -- t[53156] = 16
      "0010000" when "01100111110100101", -- t[53157] = 16
      "0010000" when "01100111110100110", -- t[53158] = 16
      "0010000" when "01100111110100111", -- t[53159] = 16
      "0010000" when "01100111110101000", -- t[53160] = 16
      "0010000" when "01100111110101001", -- t[53161] = 16
      "0010000" when "01100111110101010", -- t[53162] = 16
      "0010000" when "01100111110101011", -- t[53163] = 16
      "0010000" when "01100111110101100", -- t[53164] = 16
      "0010000" when "01100111110101101", -- t[53165] = 16
      "0010000" when "01100111110101110", -- t[53166] = 16
      "0010000" when "01100111110101111", -- t[53167] = 16
      "0010000" when "01100111110110000", -- t[53168] = 16
      "0010000" when "01100111110110001", -- t[53169] = 16
      "0010000" when "01100111110110010", -- t[53170] = 16
      "0010000" when "01100111110110011", -- t[53171] = 16
      "0010000" when "01100111110110100", -- t[53172] = 16
      "0010000" when "01100111110110101", -- t[53173] = 16
      "0010000" when "01100111110110110", -- t[53174] = 16
      "0010000" when "01100111110110111", -- t[53175] = 16
      "0010000" when "01100111110111000", -- t[53176] = 16
      "0010000" when "01100111110111001", -- t[53177] = 16
      "0010000" when "01100111110111010", -- t[53178] = 16
      "0010000" when "01100111110111011", -- t[53179] = 16
      "0010000" when "01100111110111100", -- t[53180] = 16
      "0010000" when "01100111110111101", -- t[53181] = 16
      "0010000" when "01100111110111110", -- t[53182] = 16
      "0010000" when "01100111110111111", -- t[53183] = 16
      "0010000" when "01100111111000000", -- t[53184] = 16
      "0010000" when "01100111111000001", -- t[53185] = 16
      "0010000" when "01100111111000010", -- t[53186] = 16
      "0010000" when "01100111111000011", -- t[53187] = 16
      "0010000" when "01100111111000100", -- t[53188] = 16
      "0010000" when "01100111111000101", -- t[53189] = 16
      "0010000" when "01100111111000110", -- t[53190] = 16
      "0010000" when "01100111111000111", -- t[53191] = 16
      "0010000" when "01100111111001000", -- t[53192] = 16
      "0010000" when "01100111111001001", -- t[53193] = 16
      "0010000" when "01100111111001010", -- t[53194] = 16
      "0010000" when "01100111111001011", -- t[53195] = 16
      "0010000" when "01100111111001100", -- t[53196] = 16
      "0010000" when "01100111111001101", -- t[53197] = 16
      "0010000" when "01100111111001110", -- t[53198] = 16
      "0010000" when "01100111111001111", -- t[53199] = 16
      "0010000" when "01100111111010000", -- t[53200] = 16
      "0010000" when "01100111111010001", -- t[53201] = 16
      "0010000" when "01100111111010010", -- t[53202] = 16
      "0010000" when "01100111111010011", -- t[53203] = 16
      "0010000" when "01100111111010100", -- t[53204] = 16
      "0010000" when "01100111111010101", -- t[53205] = 16
      "0010000" when "01100111111010110", -- t[53206] = 16
      "0010000" when "01100111111010111", -- t[53207] = 16
      "0010000" when "01100111111011000", -- t[53208] = 16
      "0010000" when "01100111111011001", -- t[53209] = 16
      "0010000" when "01100111111011010", -- t[53210] = 16
      "0010000" when "01100111111011011", -- t[53211] = 16
      "0010000" when "01100111111011100", -- t[53212] = 16
      "0010000" when "01100111111011101", -- t[53213] = 16
      "0010000" when "01100111111011110", -- t[53214] = 16
      "0010000" when "01100111111011111", -- t[53215] = 16
      "0010000" when "01100111111100000", -- t[53216] = 16
      "0010000" when "01100111111100001", -- t[53217] = 16
      "0010000" when "01100111111100010", -- t[53218] = 16
      "0010000" when "01100111111100011", -- t[53219] = 16
      "0010000" when "01100111111100100", -- t[53220] = 16
      "0010000" when "01100111111100101", -- t[53221] = 16
      "0010000" when "01100111111100110", -- t[53222] = 16
      "0010000" when "01100111111100111", -- t[53223] = 16
      "0010000" when "01100111111101000", -- t[53224] = 16
      "0010000" when "01100111111101001", -- t[53225] = 16
      "0010000" when "01100111111101010", -- t[53226] = 16
      "0010000" when "01100111111101011", -- t[53227] = 16
      "0010000" when "01100111111101100", -- t[53228] = 16
      "0010000" when "01100111111101101", -- t[53229] = 16
      "0010000" when "01100111111101110", -- t[53230] = 16
      "0010000" when "01100111111101111", -- t[53231] = 16
      "0010000" when "01100111111110000", -- t[53232] = 16
      "0010000" when "01100111111110001", -- t[53233] = 16
      "0010000" when "01100111111110010", -- t[53234] = 16
      "0010000" when "01100111111110011", -- t[53235] = 16
      "0010000" when "01100111111110100", -- t[53236] = 16
      "0010000" when "01100111111110101", -- t[53237] = 16
      "0010000" when "01100111111110110", -- t[53238] = 16
      "0010000" when "01100111111110111", -- t[53239] = 16
      "0010000" when "01100111111111000", -- t[53240] = 16
      "0010000" when "01100111111111001", -- t[53241] = 16
      "0010000" when "01100111111111010", -- t[53242] = 16
      "0010000" when "01100111111111011", -- t[53243] = 16
      "0010000" when "01100111111111100", -- t[53244] = 16
      "0010000" when "01100111111111101", -- t[53245] = 16
      "0010000" when "01100111111111110", -- t[53246] = 16
      "0010000" when "01100111111111111", -- t[53247] = 16
      "0010000" when "01101000000000000", -- t[53248] = 16
      "0010000" when "01101000000000001", -- t[53249] = 16
      "0010000" when "01101000000000010", -- t[53250] = 16
      "0010000" when "01101000000000011", -- t[53251] = 16
      "0010000" when "01101000000000100", -- t[53252] = 16
      "0010000" when "01101000000000101", -- t[53253] = 16
      "0010000" when "01101000000000110", -- t[53254] = 16
      "0010000" when "01101000000000111", -- t[53255] = 16
      "0010000" when "01101000000001000", -- t[53256] = 16
      "0010000" when "01101000000001001", -- t[53257] = 16
      "0010000" when "01101000000001010", -- t[53258] = 16
      "0010000" when "01101000000001011", -- t[53259] = 16
      "0010000" when "01101000000001100", -- t[53260] = 16
      "0010000" when "01101000000001101", -- t[53261] = 16
      "0010000" when "01101000000001110", -- t[53262] = 16
      "0010000" when "01101000000001111", -- t[53263] = 16
      "0010000" when "01101000000010000", -- t[53264] = 16
      "0010000" when "01101000000010001", -- t[53265] = 16
      "0010000" when "01101000000010010", -- t[53266] = 16
      "0010000" when "01101000000010011", -- t[53267] = 16
      "0010000" when "01101000000010100", -- t[53268] = 16
      "0010000" when "01101000000010101", -- t[53269] = 16
      "0010000" when "01101000000010110", -- t[53270] = 16
      "0010000" when "01101000000010111", -- t[53271] = 16
      "0010000" when "01101000000011000", -- t[53272] = 16
      "0010000" when "01101000000011001", -- t[53273] = 16
      "0010000" when "01101000000011010", -- t[53274] = 16
      "0010000" when "01101000000011011", -- t[53275] = 16
      "0010000" when "01101000000011100", -- t[53276] = 16
      "0010000" when "01101000000011101", -- t[53277] = 16
      "0010000" when "01101000000011110", -- t[53278] = 16
      "0010000" when "01101000000011111", -- t[53279] = 16
      "0010000" when "01101000000100000", -- t[53280] = 16
      "0010000" when "01101000000100001", -- t[53281] = 16
      "0010000" when "01101000000100010", -- t[53282] = 16
      "0010000" when "01101000000100011", -- t[53283] = 16
      "0010000" when "01101000000100100", -- t[53284] = 16
      "0010000" when "01101000000100101", -- t[53285] = 16
      "0010000" when "01101000000100110", -- t[53286] = 16
      "0010000" when "01101000000100111", -- t[53287] = 16
      "0010000" when "01101000000101000", -- t[53288] = 16
      "0010000" when "01101000000101001", -- t[53289] = 16
      "0010000" when "01101000000101010", -- t[53290] = 16
      "0010000" when "01101000000101011", -- t[53291] = 16
      "0010000" when "01101000000101100", -- t[53292] = 16
      "0010000" when "01101000000101101", -- t[53293] = 16
      "0010000" when "01101000000101110", -- t[53294] = 16
      "0010000" when "01101000000101111", -- t[53295] = 16
      "0010000" when "01101000000110000", -- t[53296] = 16
      "0010000" when "01101000000110001", -- t[53297] = 16
      "0010000" when "01101000000110010", -- t[53298] = 16
      "0010000" when "01101000000110011", -- t[53299] = 16
      "0010000" when "01101000000110100", -- t[53300] = 16
      "0010000" when "01101000000110101", -- t[53301] = 16
      "0010000" when "01101000000110110", -- t[53302] = 16
      "0010000" when "01101000000110111", -- t[53303] = 16
      "0010000" when "01101000000111000", -- t[53304] = 16
      "0010000" when "01101000000111001", -- t[53305] = 16
      "0010000" when "01101000000111010", -- t[53306] = 16
      "0010000" when "01101000000111011", -- t[53307] = 16
      "0010000" when "01101000000111100", -- t[53308] = 16
      "0010000" when "01101000000111101", -- t[53309] = 16
      "0010000" when "01101000000111110", -- t[53310] = 16
      "0010000" when "01101000000111111", -- t[53311] = 16
      "0010000" when "01101000001000000", -- t[53312] = 16
      "0010000" when "01101000001000001", -- t[53313] = 16
      "0010000" when "01101000001000010", -- t[53314] = 16
      "0010000" when "01101000001000011", -- t[53315] = 16
      "0010000" when "01101000001000100", -- t[53316] = 16
      "0010000" when "01101000001000101", -- t[53317] = 16
      "0010000" when "01101000001000110", -- t[53318] = 16
      "0010000" when "01101000001000111", -- t[53319] = 16
      "0010000" when "01101000001001000", -- t[53320] = 16
      "0010000" when "01101000001001001", -- t[53321] = 16
      "0010000" when "01101000001001010", -- t[53322] = 16
      "0010000" when "01101000001001011", -- t[53323] = 16
      "0010000" when "01101000001001100", -- t[53324] = 16
      "0010000" when "01101000001001101", -- t[53325] = 16
      "0010000" when "01101000001001110", -- t[53326] = 16
      "0010000" when "01101000001001111", -- t[53327] = 16
      "0010000" when "01101000001010000", -- t[53328] = 16
      "0010000" when "01101000001010001", -- t[53329] = 16
      "0010000" when "01101000001010010", -- t[53330] = 16
      "0010000" when "01101000001010011", -- t[53331] = 16
      "0010000" when "01101000001010100", -- t[53332] = 16
      "0010000" when "01101000001010101", -- t[53333] = 16
      "0010000" when "01101000001010110", -- t[53334] = 16
      "0010000" when "01101000001010111", -- t[53335] = 16
      "0010000" when "01101000001011000", -- t[53336] = 16
      "0010000" when "01101000001011001", -- t[53337] = 16
      "0010000" when "01101000001011010", -- t[53338] = 16
      "0010000" when "01101000001011011", -- t[53339] = 16
      "0010000" when "01101000001011100", -- t[53340] = 16
      "0010000" when "01101000001011101", -- t[53341] = 16
      "0010000" when "01101000001011110", -- t[53342] = 16
      "0010000" when "01101000001011111", -- t[53343] = 16
      "0010000" when "01101000001100000", -- t[53344] = 16
      "0010000" when "01101000001100001", -- t[53345] = 16
      "0010000" when "01101000001100010", -- t[53346] = 16
      "0010000" when "01101000001100011", -- t[53347] = 16
      "0010000" when "01101000001100100", -- t[53348] = 16
      "0010000" when "01101000001100101", -- t[53349] = 16
      "0010000" when "01101000001100110", -- t[53350] = 16
      "0010000" when "01101000001100111", -- t[53351] = 16
      "0010000" when "01101000001101000", -- t[53352] = 16
      "0010000" when "01101000001101001", -- t[53353] = 16
      "0010000" when "01101000001101010", -- t[53354] = 16
      "0010000" when "01101000001101011", -- t[53355] = 16
      "0010000" when "01101000001101100", -- t[53356] = 16
      "0010000" when "01101000001101101", -- t[53357] = 16
      "0010000" when "01101000001101110", -- t[53358] = 16
      "0010000" when "01101000001101111", -- t[53359] = 16
      "0010000" when "01101000001110000", -- t[53360] = 16
      "0010000" when "01101000001110001", -- t[53361] = 16
      "0010000" when "01101000001110010", -- t[53362] = 16
      "0010000" when "01101000001110011", -- t[53363] = 16
      "0010000" when "01101000001110100", -- t[53364] = 16
      "0010000" when "01101000001110101", -- t[53365] = 16
      "0010000" when "01101000001110110", -- t[53366] = 16
      "0010000" when "01101000001110111", -- t[53367] = 16
      "0010001" when "01101000001111000", -- t[53368] = 17
      "0010001" when "01101000001111001", -- t[53369] = 17
      "0010001" when "01101000001111010", -- t[53370] = 17
      "0010001" when "01101000001111011", -- t[53371] = 17
      "0010001" when "01101000001111100", -- t[53372] = 17
      "0010001" when "01101000001111101", -- t[53373] = 17
      "0010001" when "01101000001111110", -- t[53374] = 17
      "0010001" when "01101000001111111", -- t[53375] = 17
      "0010001" when "01101000010000000", -- t[53376] = 17
      "0010001" when "01101000010000001", -- t[53377] = 17
      "0010001" when "01101000010000010", -- t[53378] = 17
      "0010001" when "01101000010000011", -- t[53379] = 17
      "0010001" when "01101000010000100", -- t[53380] = 17
      "0010001" when "01101000010000101", -- t[53381] = 17
      "0010001" when "01101000010000110", -- t[53382] = 17
      "0010001" when "01101000010000111", -- t[53383] = 17
      "0010001" when "01101000010001000", -- t[53384] = 17
      "0010001" when "01101000010001001", -- t[53385] = 17
      "0010001" when "01101000010001010", -- t[53386] = 17
      "0010001" when "01101000010001011", -- t[53387] = 17
      "0010001" when "01101000010001100", -- t[53388] = 17
      "0010001" when "01101000010001101", -- t[53389] = 17
      "0010001" when "01101000010001110", -- t[53390] = 17
      "0010001" when "01101000010001111", -- t[53391] = 17
      "0010001" when "01101000010010000", -- t[53392] = 17
      "0010001" when "01101000010010001", -- t[53393] = 17
      "0010001" when "01101000010010010", -- t[53394] = 17
      "0010001" when "01101000010010011", -- t[53395] = 17
      "0010001" when "01101000010010100", -- t[53396] = 17
      "0010001" when "01101000010010101", -- t[53397] = 17
      "0010001" when "01101000010010110", -- t[53398] = 17
      "0010001" when "01101000010010111", -- t[53399] = 17
      "0010001" when "01101000010011000", -- t[53400] = 17
      "0010001" when "01101000010011001", -- t[53401] = 17
      "0010001" when "01101000010011010", -- t[53402] = 17
      "0010001" when "01101000010011011", -- t[53403] = 17
      "0010001" when "01101000010011100", -- t[53404] = 17
      "0010001" when "01101000010011101", -- t[53405] = 17
      "0010001" when "01101000010011110", -- t[53406] = 17
      "0010001" when "01101000010011111", -- t[53407] = 17
      "0010001" when "01101000010100000", -- t[53408] = 17
      "0010001" when "01101000010100001", -- t[53409] = 17
      "0010001" when "01101000010100010", -- t[53410] = 17
      "0010001" when "01101000010100011", -- t[53411] = 17
      "0010001" when "01101000010100100", -- t[53412] = 17
      "0010001" when "01101000010100101", -- t[53413] = 17
      "0010001" when "01101000010100110", -- t[53414] = 17
      "0010001" when "01101000010100111", -- t[53415] = 17
      "0010001" when "01101000010101000", -- t[53416] = 17
      "0010001" when "01101000010101001", -- t[53417] = 17
      "0010001" when "01101000010101010", -- t[53418] = 17
      "0010001" when "01101000010101011", -- t[53419] = 17
      "0010001" when "01101000010101100", -- t[53420] = 17
      "0010001" when "01101000010101101", -- t[53421] = 17
      "0010001" when "01101000010101110", -- t[53422] = 17
      "0010001" when "01101000010101111", -- t[53423] = 17
      "0010001" when "01101000010110000", -- t[53424] = 17
      "0010001" when "01101000010110001", -- t[53425] = 17
      "0010001" when "01101000010110010", -- t[53426] = 17
      "0010001" when "01101000010110011", -- t[53427] = 17
      "0010001" when "01101000010110100", -- t[53428] = 17
      "0010001" when "01101000010110101", -- t[53429] = 17
      "0010001" when "01101000010110110", -- t[53430] = 17
      "0010001" when "01101000010110111", -- t[53431] = 17
      "0010001" when "01101000010111000", -- t[53432] = 17
      "0010001" when "01101000010111001", -- t[53433] = 17
      "0010001" when "01101000010111010", -- t[53434] = 17
      "0010001" when "01101000010111011", -- t[53435] = 17
      "0010001" when "01101000010111100", -- t[53436] = 17
      "0010001" when "01101000010111101", -- t[53437] = 17
      "0010001" when "01101000010111110", -- t[53438] = 17
      "0010001" when "01101000010111111", -- t[53439] = 17
      "0010001" when "01101000011000000", -- t[53440] = 17
      "0010001" when "01101000011000001", -- t[53441] = 17
      "0010001" when "01101000011000010", -- t[53442] = 17
      "0010001" when "01101000011000011", -- t[53443] = 17
      "0010001" when "01101000011000100", -- t[53444] = 17
      "0010001" when "01101000011000101", -- t[53445] = 17
      "0010001" when "01101000011000110", -- t[53446] = 17
      "0010001" when "01101000011000111", -- t[53447] = 17
      "0010001" when "01101000011001000", -- t[53448] = 17
      "0010001" when "01101000011001001", -- t[53449] = 17
      "0010001" when "01101000011001010", -- t[53450] = 17
      "0010001" when "01101000011001011", -- t[53451] = 17
      "0010001" when "01101000011001100", -- t[53452] = 17
      "0010001" when "01101000011001101", -- t[53453] = 17
      "0010001" when "01101000011001110", -- t[53454] = 17
      "0010001" when "01101000011001111", -- t[53455] = 17
      "0010001" when "01101000011010000", -- t[53456] = 17
      "0010001" when "01101000011010001", -- t[53457] = 17
      "0010001" when "01101000011010010", -- t[53458] = 17
      "0010001" when "01101000011010011", -- t[53459] = 17
      "0010001" when "01101000011010100", -- t[53460] = 17
      "0010001" when "01101000011010101", -- t[53461] = 17
      "0010001" when "01101000011010110", -- t[53462] = 17
      "0010001" when "01101000011010111", -- t[53463] = 17
      "0010001" when "01101000011011000", -- t[53464] = 17
      "0010001" when "01101000011011001", -- t[53465] = 17
      "0010001" when "01101000011011010", -- t[53466] = 17
      "0010001" when "01101000011011011", -- t[53467] = 17
      "0010001" when "01101000011011100", -- t[53468] = 17
      "0010001" when "01101000011011101", -- t[53469] = 17
      "0010001" when "01101000011011110", -- t[53470] = 17
      "0010001" when "01101000011011111", -- t[53471] = 17
      "0010001" when "01101000011100000", -- t[53472] = 17
      "0010001" when "01101000011100001", -- t[53473] = 17
      "0010001" when "01101000011100010", -- t[53474] = 17
      "0010001" when "01101000011100011", -- t[53475] = 17
      "0010001" when "01101000011100100", -- t[53476] = 17
      "0010001" when "01101000011100101", -- t[53477] = 17
      "0010001" when "01101000011100110", -- t[53478] = 17
      "0010001" when "01101000011100111", -- t[53479] = 17
      "0010001" when "01101000011101000", -- t[53480] = 17
      "0010001" when "01101000011101001", -- t[53481] = 17
      "0010001" when "01101000011101010", -- t[53482] = 17
      "0010001" when "01101000011101011", -- t[53483] = 17
      "0010001" when "01101000011101100", -- t[53484] = 17
      "0010001" when "01101000011101101", -- t[53485] = 17
      "0010001" when "01101000011101110", -- t[53486] = 17
      "0010001" when "01101000011101111", -- t[53487] = 17
      "0010001" when "01101000011110000", -- t[53488] = 17
      "0010001" when "01101000011110001", -- t[53489] = 17
      "0010001" when "01101000011110010", -- t[53490] = 17
      "0010001" when "01101000011110011", -- t[53491] = 17
      "0010001" when "01101000011110100", -- t[53492] = 17
      "0010001" when "01101000011110101", -- t[53493] = 17
      "0010001" when "01101000011110110", -- t[53494] = 17
      "0010001" when "01101000011110111", -- t[53495] = 17
      "0010001" when "01101000011111000", -- t[53496] = 17
      "0010001" when "01101000011111001", -- t[53497] = 17
      "0010001" when "01101000011111010", -- t[53498] = 17
      "0010001" when "01101000011111011", -- t[53499] = 17
      "0010001" when "01101000011111100", -- t[53500] = 17
      "0010001" when "01101000011111101", -- t[53501] = 17
      "0010001" when "01101000011111110", -- t[53502] = 17
      "0010001" when "01101000011111111", -- t[53503] = 17
      "0010001" when "01101000100000000", -- t[53504] = 17
      "0010001" when "01101000100000001", -- t[53505] = 17
      "0010001" when "01101000100000010", -- t[53506] = 17
      "0010001" when "01101000100000011", -- t[53507] = 17
      "0010001" when "01101000100000100", -- t[53508] = 17
      "0010001" when "01101000100000101", -- t[53509] = 17
      "0010001" when "01101000100000110", -- t[53510] = 17
      "0010001" when "01101000100000111", -- t[53511] = 17
      "0010001" when "01101000100001000", -- t[53512] = 17
      "0010001" when "01101000100001001", -- t[53513] = 17
      "0010001" when "01101000100001010", -- t[53514] = 17
      "0010001" when "01101000100001011", -- t[53515] = 17
      "0010001" when "01101000100001100", -- t[53516] = 17
      "0010001" when "01101000100001101", -- t[53517] = 17
      "0010001" when "01101000100001110", -- t[53518] = 17
      "0010001" when "01101000100001111", -- t[53519] = 17
      "0010001" when "01101000100010000", -- t[53520] = 17
      "0010001" when "01101000100010001", -- t[53521] = 17
      "0010001" when "01101000100010010", -- t[53522] = 17
      "0010001" when "01101000100010011", -- t[53523] = 17
      "0010001" when "01101000100010100", -- t[53524] = 17
      "0010001" when "01101000100010101", -- t[53525] = 17
      "0010001" when "01101000100010110", -- t[53526] = 17
      "0010001" when "01101000100010111", -- t[53527] = 17
      "0010001" when "01101000100011000", -- t[53528] = 17
      "0010001" when "01101000100011001", -- t[53529] = 17
      "0010001" when "01101000100011010", -- t[53530] = 17
      "0010001" when "01101000100011011", -- t[53531] = 17
      "0010001" when "01101000100011100", -- t[53532] = 17
      "0010001" when "01101000100011101", -- t[53533] = 17
      "0010001" when "01101000100011110", -- t[53534] = 17
      "0010001" when "01101000100011111", -- t[53535] = 17
      "0010001" when "01101000100100000", -- t[53536] = 17
      "0010001" when "01101000100100001", -- t[53537] = 17
      "0010001" when "01101000100100010", -- t[53538] = 17
      "0010001" when "01101000100100011", -- t[53539] = 17
      "0010001" when "01101000100100100", -- t[53540] = 17
      "0010001" when "01101000100100101", -- t[53541] = 17
      "0010001" when "01101000100100110", -- t[53542] = 17
      "0010001" when "01101000100100111", -- t[53543] = 17
      "0010001" when "01101000100101000", -- t[53544] = 17
      "0010001" when "01101000100101001", -- t[53545] = 17
      "0010001" when "01101000100101010", -- t[53546] = 17
      "0010001" when "01101000100101011", -- t[53547] = 17
      "0010001" when "01101000100101100", -- t[53548] = 17
      "0010001" when "01101000100101101", -- t[53549] = 17
      "0010001" when "01101000100101110", -- t[53550] = 17
      "0010001" when "01101000100101111", -- t[53551] = 17
      "0010001" when "01101000100110000", -- t[53552] = 17
      "0010001" when "01101000100110001", -- t[53553] = 17
      "0010001" when "01101000100110010", -- t[53554] = 17
      "0010001" when "01101000100110011", -- t[53555] = 17
      "0010001" when "01101000100110100", -- t[53556] = 17
      "0010001" when "01101000100110101", -- t[53557] = 17
      "0010001" when "01101000100110110", -- t[53558] = 17
      "0010001" when "01101000100110111", -- t[53559] = 17
      "0010001" when "01101000100111000", -- t[53560] = 17
      "0010001" when "01101000100111001", -- t[53561] = 17
      "0010001" when "01101000100111010", -- t[53562] = 17
      "0010001" when "01101000100111011", -- t[53563] = 17
      "0010001" when "01101000100111100", -- t[53564] = 17
      "0010001" when "01101000100111101", -- t[53565] = 17
      "0010001" when "01101000100111110", -- t[53566] = 17
      "0010001" when "01101000100111111", -- t[53567] = 17
      "0010001" when "01101000101000000", -- t[53568] = 17
      "0010001" when "01101000101000001", -- t[53569] = 17
      "0010001" when "01101000101000010", -- t[53570] = 17
      "0010001" when "01101000101000011", -- t[53571] = 17
      "0010001" when "01101000101000100", -- t[53572] = 17
      "0010001" when "01101000101000101", -- t[53573] = 17
      "0010001" when "01101000101000110", -- t[53574] = 17
      "0010001" when "01101000101000111", -- t[53575] = 17
      "0010001" when "01101000101001000", -- t[53576] = 17
      "0010001" when "01101000101001001", -- t[53577] = 17
      "0010001" when "01101000101001010", -- t[53578] = 17
      "0010001" when "01101000101001011", -- t[53579] = 17
      "0010001" when "01101000101001100", -- t[53580] = 17
      "0010001" when "01101000101001101", -- t[53581] = 17
      "0010001" when "01101000101001110", -- t[53582] = 17
      "0010001" when "01101000101001111", -- t[53583] = 17
      "0010001" when "01101000101010000", -- t[53584] = 17
      "0010001" when "01101000101010001", -- t[53585] = 17
      "0010001" when "01101000101010010", -- t[53586] = 17
      "0010001" when "01101000101010011", -- t[53587] = 17
      "0010001" when "01101000101010100", -- t[53588] = 17
      "0010001" when "01101000101010101", -- t[53589] = 17
      "0010001" when "01101000101010110", -- t[53590] = 17
      "0010001" when "01101000101010111", -- t[53591] = 17
      "0010001" when "01101000101011000", -- t[53592] = 17
      "0010001" when "01101000101011001", -- t[53593] = 17
      "0010001" when "01101000101011010", -- t[53594] = 17
      "0010001" when "01101000101011011", -- t[53595] = 17
      "0010001" when "01101000101011100", -- t[53596] = 17
      "0010001" when "01101000101011101", -- t[53597] = 17
      "0010001" when "01101000101011110", -- t[53598] = 17
      "0010001" when "01101000101011111", -- t[53599] = 17
      "0010001" when "01101000101100000", -- t[53600] = 17
      "0010001" when "01101000101100001", -- t[53601] = 17
      "0010001" when "01101000101100010", -- t[53602] = 17
      "0010001" when "01101000101100011", -- t[53603] = 17
      "0010001" when "01101000101100100", -- t[53604] = 17
      "0010001" when "01101000101100101", -- t[53605] = 17
      "0010001" when "01101000101100110", -- t[53606] = 17
      "0010001" when "01101000101100111", -- t[53607] = 17
      "0010001" when "01101000101101000", -- t[53608] = 17
      "0010001" when "01101000101101001", -- t[53609] = 17
      "0010001" when "01101000101101010", -- t[53610] = 17
      "0010001" when "01101000101101011", -- t[53611] = 17
      "0010001" when "01101000101101100", -- t[53612] = 17
      "0010001" when "01101000101101101", -- t[53613] = 17
      "0010001" when "01101000101101110", -- t[53614] = 17
      "0010001" when "01101000101101111", -- t[53615] = 17
      "0010001" when "01101000101110000", -- t[53616] = 17
      "0010001" when "01101000101110001", -- t[53617] = 17
      "0010001" when "01101000101110010", -- t[53618] = 17
      "0010001" when "01101000101110011", -- t[53619] = 17
      "0010001" when "01101000101110100", -- t[53620] = 17
      "0010001" when "01101000101110101", -- t[53621] = 17
      "0010001" when "01101000101110110", -- t[53622] = 17
      "0010001" when "01101000101110111", -- t[53623] = 17
      "0010001" when "01101000101111000", -- t[53624] = 17
      "0010001" when "01101000101111001", -- t[53625] = 17
      "0010001" when "01101000101111010", -- t[53626] = 17
      "0010001" when "01101000101111011", -- t[53627] = 17
      "0010001" when "01101000101111100", -- t[53628] = 17
      "0010001" when "01101000101111101", -- t[53629] = 17
      "0010001" when "01101000101111110", -- t[53630] = 17
      "0010001" when "01101000101111111", -- t[53631] = 17
      "0010001" when "01101000110000000", -- t[53632] = 17
      "0010001" when "01101000110000001", -- t[53633] = 17
      "0010001" when "01101000110000010", -- t[53634] = 17
      "0010001" when "01101000110000011", -- t[53635] = 17
      "0010001" when "01101000110000100", -- t[53636] = 17
      "0010001" when "01101000110000101", -- t[53637] = 17
      "0010001" when "01101000110000110", -- t[53638] = 17
      "0010001" when "01101000110000111", -- t[53639] = 17
      "0010001" when "01101000110001000", -- t[53640] = 17
      "0010001" when "01101000110001001", -- t[53641] = 17
      "0010001" when "01101000110001010", -- t[53642] = 17
      "0010001" when "01101000110001011", -- t[53643] = 17
      "0010001" when "01101000110001100", -- t[53644] = 17
      "0010001" when "01101000110001101", -- t[53645] = 17
      "0010001" when "01101000110001110", -- t[53646] = 17
      "0010001" when "01101000110001111", -- t[53647] = 17
      "0010001" when "01101000110010000", -- t[53648] = 17
      "0010001" when "01101000110010001", -- t[53649] = 17
      "0010001" when "01101000110010010", -- t[53650] = 17
      "0010001" when "01101000110010011", -- t[53651] = 17
      "0010001" when "01101000110010100", -- t[53652] = 17
      "0010001" when "01101000110010101", -- t[53653] = 17
      "0010001" when "01101000110010110", -- t[53654] = 17
      "0010001" when "01101000110010111", -- t[53655] = 17
      "0010001" when "01101000110011000", -- t[53656] = 17
      "0010001" when "01101000110011001", -- t[53657] = 17
      "0010001" when "01101000110011010", -- t[53658] = 17
      "0010001" when "01101000110011011", -- t[53659] = 17
      "0010001" when "01101000110011100", -- t[53660] = 17
      "0010001" when "01101000110011101", -- t[53661] = 17
      "0010001" when "01101000110011110", -- t[53662] = 17
      "0010001" when "01101000110011111", -- t[53663] = 17
      "0010001" when "01101000110100000", -- t[53664] = 17
      "0010001" when "01101000110100001", -- t[53665] = 17
      "0010001" when "01101000110100010", -- t[53666] = 17
      "0010001" when "01101000110100011", -- t[53667] = 17
      "0010001" when "01101000110100100", -- t[53668] = 17
      "0010001" when "01101000110100101", -- t[53669] = 17
      "0010001" when "01101000110100110", -- t[53670] = 17
      "0010001" when "01101000110100111", -- t[53671] = 17
      "0010001" when "01101000110101000", -- t[53672] = 17
      "0010001" when "01101000110101001", -- t[53673] = 17
      "0010001" when "01101000110101010", -- t[53674] = 17
      "0010001" when "01101000110101011", -- t[53675] = 17
      "0010001" when "01101000110101100", -- t[53676] = 17
      "0010001" when "01101000110101101", -- t[53677] = 17
      "0010001" when "01101000110101110", -- t[53678] = 17
      "0010001" when "01101000110101111", -- t[53679] = 17
      "0010001" when "01101000110110000", -- t[53680] = 17
      "0010001" when "01101000110110001", -- t[53681] = 17
      "0010001" when "01101000110110010", -- t[53682] = 17
      "0010001" when "01101000110110011", -- t[53683] = 17
      "0010001" when "01101000110110100", -- t[53684] = 17
      "0010001" when "01101000110110101", -- t[53685] = 17
      "0010001" when "01101000110110110", -- t[53686] = 17
      "0010001" when "01101000110110111", -- t[53687] = 17
      "0010001" when "01101000110111000", -- t[53688] = 17
      "0010001" when "01101000110111001", -- t[53689] = 17
      "0010001" when "01101000110111010", -- t[53690] = 17
      "0010001" when "01101000110111011", -- t[53691] = 17
      "0010001" when "01101000110111100", -- t[53692] = 17
      "0010001" when "01101000110111101", -- t[53693] = 17
      "0010001" when "01101000110111110", -- t[53694] = 17
      "0010001" when "01101000110111111", -- t[53695] = 17
      "0010001" when "01101000111000000", -- t[53696] = 17
      "0010001" when "01101000111000001", -- t[53697] = 17
      "0010001" when "01101000111000010", -- t[53698] = 17
      "0010001" when "01101000111000011", -- t[53699] = 17
      "0010001" when "01101000111000100", -- t[53700] = 17
      "0010001" when "01101000111000101", -- t[53701] = 17
      "0010001" when "01101000111000110", -- t[53702] = 17
      "0010001" when "01101000111000111", -- t[53703] = 17
      "0010001" when "01101000111001000", -- t[53704] = 17
      "0010001" when "01101000111001001", -- t[53705] = 17
      "0010001" when "01101000111001010", -- t[53706] = 17
      "0010001" when "01101000111001011", -- t[53707] = 17
      "0010001" when "01101000111001100", -- t[53708] = 17
      "0010001" when "01101000111001101", -- t[53709] = 17
      "0010001" when "01101000111001110", -- t[53710] = 17
      "0010001" when "01101000111001111", -- t[53711] = 17
      "0010001" when "01101000111010000", -- t[53712] = 17
      "0010001" when "01101000111010001", -- t[53713] = 17
      "0010001" when "01101000111010010", -- t[53714] = 17
      "0010001" when "01101000111010011", -- t[53715] = 17
      "0010001" when "01101000111010100", -- t[53716] = 17
      "0010001" when "01101000111010101", -- t[53717] = 17
      "0010001" when "01101000111010110", -- t[53718] = 17
      "0010001" when "01101000111010111", -- t[53719] = 17
      "0010001" when "01101000111011000", -- t[53720] = 17
      "0010001" when "01101000111011001", -- t[53721] = 17
      "0010001" when "01101000111011010", -- t[53722] = 17
      "0010001" when "01101000111011011", -- t[53723] = 17
      "0010001" when "01101000111011100", -- t[53724] = 17
      "0010001" when "01101000111011101", -- t[53725] = 17
      "0010001" when "01101000111011110", -- t[53726] = 17
      "0010001" when "01101000111011111", -- t[53727] = 17
      "0010001" when "01101000111100000", -- t[53728] = 17
      "0010001" when "01101000111100001", -- t[53729] = 17
      "0010001" when "01101000111100010", -- t[53730] = 17
      "0010001" when "01101000111100011", -- t[53731] = 17
      "0010001" when "01101000111100100", -- t[53732] = 17
      "0010001" when "01101000111100101", -- t[53733] = 17
      "0010001" when "01101000111100110", -- t[53734] = 17
      "0010001" when "01101000111100111", -- t[53735] = 17
      "0010001" when "01101000111101000", -- t[53736] = 17
      "0010001" when "01101000111101001", -- t[53737] = 17
      "0010001" when "01101000111101010", -- t[53738] = 17
      "0010001" when "01101000111101011", -- t[53739] = 17
      "0010001" when "01101000111101100", -- t[53740] = 17
      "0010001" when "01101000111101101", -- t[53741] = 17
      "0010001" when "01101000111101110", -- t[53742] = 17
      "0010001" when "01101000111101111", -- t[53743] = 17
      "0010001" when "01101000111110000", -- t[53744] = 17
      "0010001" when "01101000111110001", -- t[53745] = 17
      "0010001" when "01101000111110010", -- t[53746] = 17
      "0010001" when "01101000111110011", -- t[53747] = 17
      "0010001" when "01101000111110100", -- t[53748] = 17
      "0010001" when "01101000111110101", -- t[53749] = 17
      "0010001" when "01101000111110110", -- t[53750] = 17
      "0010001" when "01101000111110111", -- t[53751] = 17
      "0010001" when "01101000111111000", -- t[53752] = 17
      "0010001" when "01101000111111001", -- t[53753] = 17
      "0010001" when "01101000111111010", -- t[53754] = 17
      "0010001" when "01101000111111011", -- t[53755] = 17
      "0010001" when "01101000111111100", -- t[53756] = 17
      "0010001" when "01101000111111101", -- t[53757] = 17
      "0010001" when "01101000111111110", -- t[53758] = 17
      "0010001" when "01101000111111111", -- t[53759] = 17
      "0010001" when "01101001000000000", -- t[53760] = 17
      "0010001" when "01101001000000001", -- t[53761] = 17
      "0010001" when "01101001000000010", -- t[53762] = 17
      "0010001" when "01101001000000011", -- t[53763] = 17
      "0010001" when "01101001000000100", -- t[53764] = 17
      "0010001" when "01101001000000101", -- t[53765] = 17
      "0010001" when "01101001000000110", -- t[53766] = 17
      "0010001" when "01101001000000111", -- t[53767] = 17
      "0010001" when "01101001000001000", -- t[53768] = 17
      "0010001" when "01101001000001001", -- t[53769] = 17
      "0010001" when "01101001000001010", -- t[53770] = 17
      "0010001" when "01101001000001011", -- t[53771] = 17
      "0010001" when "01101001000001100", -- t[53772] = 17
      "0010001" when "01101001000001101", -- t[53773] = 17
      "0010001" when "01101001000001110", -- t[53774] = 17
      "0010001" when "01101001000001111", -- t[53775] = 17
      "0010001" when "01101001000010000", -- t[53776] = 17
      "0010001" when "01101001000010001", -- t[53777] = 17
      "0010001" when "01101001000010010", -- t[53778] = 17
      "0010001" when "01101001000010011", -- t[53779] = 17
      "0010001" when "01101001000010100", -- t[53780] = 17
      "0010001" when "01101001000010101", -- t[53781] = 17
      "0010001" when "01101001000010110", -- t[53782] = 17
      "0010001" when "01101001000010111", -- t[53783] = 17
      "0010001" when "01101001000011000", -- t[53784] = 17
      "0010001" when "01101001000011001", -- t[53785] = 17
      "0010001" when "01101001000011010", -- t[53786] = 17
      "0010001" when "01101001000011011", -- t[53787] = 17
      "0010001" when "01101001000011100", -- t[53788] = 17
      "0010001" when "01101001000011101", -- t[53789] = 17
      "0010001" when "01101001000011110", -- t[53790] = 17
      "0010001" when "01101001000011111", -- t[53791] = 17
      "0010001" when "01101001000100000", -- t[53792] = 17
      "0010001" when "01101001000100001", -- t[53793] = 17
      "0010001" when "01101001000100010", -- t[53794] = 17
      "0010001" when "01101001000100011", -- t[53795] = 17
      "0010001" when "01101001000100100", -- t[53796] = 17
      "0010001" when "01101001000100101", -- t[53797] = 17
      "0010001" when "01101001000100110", -- t[53798] = 17
      "0010001" when "01101001000100111", -- t[53799] = 17
      "0010001" when "01101001000101000", -- t[53800] = 17
      "0010001" when "01101001000101001", -- t[53801] = 17
      "0010001" when "01101001000101010", -- t[53802] = 17
      "0010001" when "01101001000101011", -- t[53803] = 17
      "0010001" when "01101001000101100", -- t[53804] = 17
      "0010001" when "01101001000101101", -- t[53805] = 17
      "0010001" when "01101001000101110", -- t[53806] = 17
      "0010001" when "01101001000101111", -- t[53807] = 17
      "0010001" when "01101001000110000", -- t[53808] = 17
      "0010001" when "01101001000110001", -- t[53809] = 17
      "0010001" when "01101001000110010", -- t[53810] = 17
      "0010001" when "01101001000110011", -- t[53811] = 17
      "0010001" when "01101001000110100", -- t[53812] = 17
      "0010001" when "01101001000110101", -- t[53813] = 17
      "0010001" when "01101001000110110", -- t[53814] = 17
      "0010001" when "01101001000110111", -- t[53815] = 17
      "0010001" when "01101001000111000", -- t[53816] = 17
      "0010001" when "01101001000111001", -- t[53817] = 17
      "0010001" when "01101001000111010", -- t[53818] = 17
      "0010001" when "01101001000111011", -- t[53819] = 17
      "0010001" when "01101001000111100", -- t[53820] = 17
      "0010001" when "01101001000111101", -- t[53821] = 17
      "0010001" when "01101001000111110", -- t[53822] = 17
      "0010001" when "01101001000111111", -- t[53823] = 17
      "0010001" when "01101001001000000", -- t[53824] = 17
      "0010001" when "01101001001000001", -- t[53825] = 17
      "0010001" when "01101001001000010", -- t[53826] = 17
      "0010001" when "01101001001000011", -- t[53827] = 17
      "0010001" when "01101001001000100", -- t[53828] = 17
      "0010001" when "01101001001000101", -- t[53829] = 17
      "0010001" when "01101001001000110", -- t[53830] = 17
      "0010001" when "01101001001000111", -- t[53831] = 17
      "0010001" when "01101001001001000", -- t[53832] = 17
      "0010001" when "01101001001001001", -- t[53833] = 17
      "0010001" when "01101001001001010", -- t[53834] = 17
      "0010001" when "01101001001001011", -- t[53835] = 17
      "0010001" when "01101001001001100", -- t[53836] = 17
      "0010001" when "01101001001001101", -- t[53837] = 17
      "0010001" when "01101001001001110", -- t[53838] = 17
      "0010001" when "01101001001001111", -- t[53839] = 17
      "0010001" when "01101001001010000", -- t[53840] = 17
      "0010001" when "01101001001010001", -- t[53841] = 17
      "0010001" when "01101001001010010", -- t[53842] = 17
      "0010001" when "01101001001010011", -- t[53843] = 17
      "0010001" when "01101001001010100", -- t[53844] = 17
      "0010001" when "01101001001010101", -- t[53845] = 17
      "0010001" when "01101001001010110", -- t[53846] = 17
      "0010001" when "01101001001010111", -- t[53847] = 17
      "0010001" when "01101001001011000", -- t[53848] = 17
      "0010001" when "01101001001011001", -- t[53849] = 17
      "0010001" when "01101001001011010", -- t[53850] = 17
      "0010001" when "01101001001011011", -- t[53851] = 17
      "0010001" when "01101001001011100", -- t[53852] = 17
      "0010001" when "01101001001011101", -- t[53853] = 17
      "0010001" when "01101001001011110", -- t[53854] = 17
      "0010001" when "01101001001011111", -- t[53855] = 17
      "0010001" when "01101001001100000", -- t[53856] = 17
      "0010001" when "01101001001100001", -- t[53857] = 17
      "0010001" when "01101001001100010", -- t[53858] = 17
      "0010001" when "01101001001100011", -- t[53859] = 17
      "0010001" when "01101001001100100", -- t[53860] = 17
      "0010001" when "01101001001100101", -- t[53861] = 17
      "0010001" when "01101001001100110", -- t[53862] = 17
      "0010001" when "01101001001100111", -- t[53863] = 17
      "0010001" when "01101001001101000", -- t[53864] = 17
      "0010001" when "01101001001101001", -- t[53865] = 17
      "0010001" when "01101001001101010", -- t[53866] = 17
      "0010001" when "01101001001101011", -- t[53867] = 17
      "0010001" when "01101001001101100", -- t[53868] = 17
      "0010001" when "01101001001101101", -- t[53869] = 17
      "0010001" when "01101001001101110", -- t[53870] = 17
      "0010001" when "01101001001101111", -- t[53871] = 17
      "0010001" when "01101001001110000", -- t[53872] = 17
      "0010001" when "01101001001110001", -- t[53873] = 17
      "0010001" when "01101001001110010", -- t[53874] = 17
      "0010001" when "01101001001110011", -- t[53875] = 17
      "0010001" when "01101001001110100", -- t[53876] = 17
      "0010001" when "01101001001110101", -- t[53877] = 17
      "0010001" when "01101001001110110", -- t[53878] = 17
      "0010001" when "01101001001110111", -- t[53879] = 17
      "0010001" when "01101001001111000", -- t[53880] = 17
      "0010001" when "01101001001111001", -- t[53881] = 17
      "0010001" when "01101001001111010", -- t[53882] = 17
      "0010001" when "01101001001111011", -- t[53883] = 17
      "0010001" when "01101001001111100", -- t[53884] = 17
      "0010001" when "01101001001111101", -- t[53885] = 17
      "0010001" when "01101001001111110", -- t[53886] = 17
      "0010001" when "01101001001111111", -- t[53887] = 17
      "0010001" when "01101001010000000", -- t[53888] = 17
      "0010001" when "01101001010000001", -- t[53889] = 17
      "0010001" when "01101001010000010", -- t[53890] = 17
      "0010001" when "01101001010000011", -- t[53891] = 17
      "0010001" when "01101001010000100", -- t[53892] = 17
      "0010001" when "01101001010000101", -- t[53893] = 17
      "0010001" when "01101001010000110", -- t[53894] = 17
      "0010001" when "01101001010000111", -- t[53895] = 17
      "0010001" when "01101001010001000", -- t[53896] = 17
      "0010001" when "01101001010001001", -- t[53897] = 17
      "0010001" when "01101001010001010", -- t[53898] = 17
      "0010001" when "01101001010001011", -- t[53899] = 17
      "0010001" when "01101001010001100", -- t[53900] = 17
      "0010001" when "01101001010001101", -- t[53901] = 17
      "0010001" when "01101001010001110", -- t[53902] = 17
      "0010001" when "01101001010001111", -- t[53903] = 17
      "0010001" when "01101001010010000", -- t[53904] = 17
      "0010001" when "01101001010010001", -- t[53905] = 17
      "0010001" when "01101001010010010", -- t[53906] = 17
      "0010001" when "01101001010010011", -- t[53907] = 17
      "0010001" when "01101001010010100", -- t[53908] = 17
      "0010001" when "01101001010010101", -- t[53909] = 17
      "0010001" when "01101001010010110", -- t[53910] = 17
      "0010001" when "01101001010010111", -- t[53911] = 17
      "0010001" when "01101001010011000", -- t[53912] = 17
      "0010001" when "01101001010011001", -- t[53913] = 17
      "0010001" when "01101001010011010", -- t[53914] = 17
      "0010001" when "01101001010011011", -- t[53915] = 17
      "0010001" when "01101001010011100", -- t[53916] = 17
      "0010001" when "01101001010011101", -- t[53917] = 17
      "0010001" when "01101001010011110", -- t[53918] = 17
      "0010001" when "01101001010011111", -- t[53919] = 17
      "0010001" when "01101001010100000", -- t[53920] = 17
      "0010001" when "01101001010100001", -- t[53921] = 17
      "0010001" when "01101001010100010", -- t[53922] = 17
      "0010001" when "01101001010100011", -- t[53923] = 17
      "0010001" when "01101001010100100", -- t[53924] = 17
      "0010001" when "01101001010100101", -- t[53925] = 17
      "0010001" when "01101001010100110", -- t[53926] = 17
      "0010001" when "01101001010100111", -- t[53927] = 17
      "0010001" when "01101001010101000", -- t[53928] = 17
      "0010001" when "01101001010101001", -- t[53929] = 17
      "0010001" when "01101001010101010", -- t[53930] = 17
      "0010001" when "01101001010101011", -- t[53931] = 17
      "0010001" when "01101001010101100", -- t[53932] = 17
      "0010001" when "01101001010101101", -- t[53933] = 17
      "0010001" when "01101001010101110", -- t[53934] = 17
      "0010001" when "01101001010101111", -- t[53935] = 17
      "0010001" when "01101001010110000", -- t[53936] = 17
      "0010001" when "01101001010110001", -- t[53937] = 17
      "0010001" when "01101001010110010", -- t[53938] = 17
      "0010001" when "01101001010110011", -- t[53939] = 17
      "0010001" when "01101001010110100", -- t[53940] = 17
      "0010001" when "01101001010110101", -- t[53941] = 17
      "0010001" when "01101001010110110", -- t[53942] = 17
      "0010001" when "01101001010110111", -- t[53943] = 17
      "0010001" when "01101001010111000", -- t[53944] = 17
      "0010001" when "01101001010111001", -- t[53945] = 17
      "0010001" when "01101001010111010", -- t[53946] = 17
      "0010001" when "01101001010111011", -- t[53947] = 17
      "0010001" when "01101001010111100", -- t[53948] = 17
      "0010001" when "01101001010111101", -- t[53949] = 17
      "0010001" when "01101001010111110", -- t[53950] = 17
      "0010001" when "01101001010111111", -- t[53951] = 17
      "0010001" when "01101001011000000", -- t[53952] = 17
      "0010001" when "01101001011000001", -- t[53953] = 17
      "0010001" when "01101001011000010", -- t[53954] = 17
      "0010001" when "01101001011000011", -- t[53955] = 17
      "0010001" when "01101001011000100", -- t[53956] = 17
      "0010001" when "01101001011000101", -- t[53957] = 17
      "0010001" when "01101001011000110", -- t[53958] = 17
      "0010001" when "01101001011000111", -- t[53959] = 17
      "0010001" when "01101001011001000", -- t[53960] = 17
      "0010001" when "01101001011001001", -- t[53961] = 17
      "0010001" when "01101001011001010", -- t[53962] = 17
      "0010001" when "01101001011001011", -- t[53963] = 17
      "0010001" when "01101001011001100", -- t[53964] = 17
      "0010001" when "01101001011001101", -- t[53965] = 17
      "0010001" when "01101001011001110", -- t[53966] = 17
      "0010001" when "01101001011001111", -- t[53967] = 17
      "0010001" when "01101001011010000", -- t[53968] = 17
      "0010001" when "01101001011010001", -- t[53969] = 17
      "0010001" when "01101001011010010", -- t[53970] = 17
      "0010001" when "01101001011010011", -- t[53971] = 17
      "0010001" when "01101001011010100", -- t[53972] = 17
      "0010001" when "01101001011010101", -- t[53973] = 17
      "0010001" when "01101001011010110", -- t[53974] = 17
      "0010001" when "01101001011010111", -- t[53975] = 17
      "0010001" when "01101001011011000", -- t[53976] = 17
      "0010001" when "01101001011011001", -- t[53977] = 17
      "0010001" when "01101001011011010", -- t[53978] = 17
      "0010001" when "01101001011011011", -- t[53979] = 17
      "0010001" when "01101001011011100", -- t[53980] = 17
      "0010001" when "01101001011011101", -- t[53981] = 17
      "0010001" when "01101001011011110", -- t[53982] = 17
      "0010001" when "01101001011011111", -- t[53983] = 17
      "0010001" when "01101001011100000", -- t[53984] = 17
      "0010001" when "01101001011100001", -- t[53985] = 17
      "0010001" when "01101001011100010", -- t[53986] = 17
      "0010001" when "01101001011100011", -- t[53987] = 17
      "0010001" when "01101001011100100", -- t[53988] = 17
      "0010001" when "01101001011100101", -- t[53989] = 17
      "0010001" when "01101001011100110", -- t[53990] = 17
      "0010001" when "01101001011100111", -- t[53991] = 17
      "0010001" when "01101001011101000", -- t[53992] = 17
      "0010001" when "01101001011101001", -- t[53993] = 17
      "0010001" when "01101001011101010", -- t[53994] = 17
      "0010001" when "01101001011101011", -- t[53995] = 17
      "0010001" when "01101001011101100", -- t[53996] = 17
      "0010001" when "01101001011101101", -- t[53997] = 17
      "0010001" when "01101001011101110", -- t[53998] = 17
      "0010001" when "01101001011101111", -- t[53999] = 17
      "0010001" when "01101001011110000", -- t[54000] = 17
      "0010001" when "01101001011110001", -- t[54001] = 17
      "0010001" when "01101001011110010", -- t[54002] = 17
      "0010001" when "01101001011110011", -- t[54003] = 17
      "0010001" when "01101001011110100", -- t[54004] = 17
      "0010001" when "01101001011110101", -- t[54005] = 17
      "0010001" when "01101001011110110", -- t[54006] = 17
      "0010001" when "01101001011110111", -- t[54007] = 17
      "0010001" when "01101001011111000", -- t[54008] = 17
      "0010001" when "01101001011111001", -- t[54009] = 17
      "0010001" when "01101001011111010", -- t[54010] = 17
      "0010001" when "01101001011111011", -- t[54011] = 17
      "0010001" when "01101001011111100", -- t[54012] = 17
      "0010001" when "01101001011111101", -- t[54013] = 17
      "0010001" when "01101001011111110", -- t[54014] = 17
      "0010001" when "01101001011111111", -- t[54015] = 17
      "0010001" when "01101001100000000", -- t[54016] = 17
      "0010001" when "01101001100000001", -- t[54017] = 17
      "0010001" when "01101001100000010", -- t[54018] = 17
      "0010001" when "01101001100000011", -- t[54019] = 17
      "0010001" when "01101001100000100", -- t[54020] = 17
      "0010001" when "01101001100000101", -- t[54021] = 17
      "0010001" when "01101001100000110", -- t[54022] = 17
      "0010001" when "01101001100000111", -- t[54023] = 17
      "0010001" when "01101001100001000", -- t[54024] = 17
      "0010001" when "01101001100001001", -- t[54025] = 17
      "0010001" when "01101001100001010", -- t[54026] = 17
      "0010001" when "01101001100001011", -- t[54027] = 17
      "0010001" when "01101001100001100", -- t[54028] = 17
      "0010001" when "01101001100001101", -- t[54029] = 17
      "0010001" when "01101001100001110", -- t[54030] = 17
      "0010001" when "01101001100001111", -- t[54031] = 17
      "0010001" when "01101001100010000", -- t[54032] = 17
      "0010001" when "01101001100010001", -- t[54033] = 17
      "0010001" when "01101001100010010", -- t[54034] = 17
      "0010001" when "01101001100010011", -- t[54035] = 17
      "0010001" when "01101001100010100", -- t[54036] = 17
      "0010001" when "01101001100010101", -- t[54037] = 17
      "0010001" when "01101001100010110", -- t[54038] = 17
      "0010001" when "01101001100010111", -- t[54039] = 17
      "0010001" when "01101001100011000", -- t[54040] = 17
      "0010001" when "01101001100011001", -- t[54041] = 17
      "0010001" when "01101001100011010", -- t[54042] = 17
      "0010001" when "01101001100011011", -- t[54043] = 17
      "0010001" when "01101001100011100", -- t[54044] = 17
      "0010001" when "01101001100011101", -- t[54045] = 17
      "0010001" when "01101001100011110", -- t[54046] = 17
      "0010001" when "01101001100011111", -- t[54047] = 17
      "0010001" when "01101001100100000", -- t[54048] = 17
      "0010001" when "01101001100100001", -- t[54049] = 17
      "0010001" when "01101001100100010", -- t[54050] = 17
      "0010001" when "01101001100100011", -- t[54051] = 17
      "0010001" when "01101001100100100", -- t[54052] = 17
      "0010001" when "01101001100100101", -- t[54053] = 17
      "0010001" when "01101001100100110", -- t[54054] = 17
      "0010001" when "01101001100100111", -- t[54055] = 17
      "0010001" when "01101001100101000", -- t[54056] = 17
      "0010001" when "01101001100101001", -- t[54057] = 17
      "0010001" when "01101001100101010", -- t[54058] = 17
      "0010001" when "01101001100101011", -- t[54059] = 17
      "0010001" when "01101001100101100", -- t[54060] = 17
      "0010001" when "01101001100101101", -- t[54061] = 17
      "0010001" when "01101001100101110", -- t[54062] = 17
      "0010010" when "01101001100101111", -- t[54063] = 18
      "0010010" when "01101001100110000", -- t[54064] = 18
      "0010010" when "01101001100110001", -- t[54065] = 18
      "0010010" when "01101001100110010", -- t[54066] = 18
      "0010010" when "01101001100110011", -- t[54067] = 18
      "0010010" when "01101001100110100", -- t[54068] = 18
      "0010010" when "01101001100110101", -- t[54069] = 18
      "0010010" when "01101001100110110", -- t[54070] = 18
      "0010010" when "01101001100110111", -- t[54071] = 18
      "0010010" when "01101001100111000", -- t[54072] = 18
      "0010010" when "01101001100111001", -- t[54073] = 18
      "0010010" when "01101001100111010", -- t[54074] = 18
      "0010010" when "01101001100111011", -- t[54075] = 18
      "0010010" when "01101001100111100", -- t[54076] = 18
      "0010010" when "01101001100111101", -- t[54077] = 18
      "0010010" when "01101001100111110", -- t[54078] = 18
      "0010010" when "01101001100111111", -- t[54079] = 18
      "0010010" when "01101001101000000", -- t[54080] = 18
      "0010010" when "01101001101000001", -- t[54081] = 18
      "0010010" when "01101001101000010", -- t[54082] = 18
      "0010010" when "01101001101000011", -- t[54083] = 18
      "0010010" when "01101001101000100", -- t[54084] = 18
      "0010010" when "01101001101000101", -- t[54085] = 18
      "0010010" when "01101001101000110", -- t[54086] = 18
      "0010010" when "01101001101000111", -- t[54087] = 18
      "0010010" when "01101001101001000", -- t[54088] = 18
      "0010010" when "01101001101001001", -- t[54089] = 18
      "0010010" when "01101001101001010", -- t[54090] = 18
      "0010010" when "01101001101001011", -- t[54091] = 18
      "0010010" when "01101001101001100", -- t[54092] = 18
      "0010010" when "01101001101001101", -- t[54093] = 18
      "0010010" when "01101001101001110", -- t[54094] = 18
      "0010010" when "01101001101001111", -- t[54095] = 18
      "0010010" when "01101001101010000", -- t[54096] = 18
      "0010010" when "01101001101010001", -- t[54097] = 18
      "0010010" when "01101001101010010", -- t[54098] = 18
      "0010010" when "01101001101010011", -- t[54099] = 18
      "0010010" when "01101001101010100", -- t[54100] = 18
      "0010010" when "01101001101010101", -- t[54101] = 18
      "0010010" when "01101001101010110", -- t[54102] = 18
      "0010010" when "01101001101010111", -- t[54103] = 18
      "0010010" when "01101001101011000", -- t[54104] = 18
      "0010010" when "01101001101011001", -- t[54105] = 18
      "0010010" when "01101001101011010", -- t[54106] = 18
      "0010010" when "01101001101011011", -- t[54107] = 18
      "0010010" when "01101001101011100", -- t[54108] = 18
      "0010010" when "01101001101011101", -- t[54109] = 18
      "0010010" when "01101001101011110", -- t[54110] = 18
      "0010010" when "01101001101011111", -- t[54111] = 18
      "0010010" when "01101001101100000", -- t[54112] = 18
      "0010010" when "01101001101100001", -- t[54113] = 18
      "0010010" when "01101001101100010", -- t[54114] = 18
      "0010010" when "01101001101100011", -- t[54115] = 18
      "0010010" when "01101001101100100", -- t[54116] = 18
      "0010010" when "01101001101100101", -- t[54117] = 18
      "0010010" when "01101001101100110", -- t[54118] = 18
      "0010010" when "01101001101100111", -- t[54119] = 18
      "0010010" when "01101001101101000", -- t[54120] = 18
      "0010010" when "01101001101101001", -- t[54121] = 18
      "0010010" when "01101001101101010", -- t[54122] = 18
      "0010010" when "01101001101101011", -- t[54123] = 18
      "0010010" when "01101001101101100", -- t[54124] = 18
      "0010010" when "01101001101101101", -- t[54125] = 18
      "0010010" when "01101001101101110", -- t[54126] = 18
      "0010010" when "01101001101101111", -- t[54127] = 18
      "0010010" when "01101001101110000", -- t[54128] = 18
      "0010010" when "01101001101110001", -- t[54129] = 18
      "0010010" when "01101001101110010", -- t[54130] = 18
      "0010010" when "01101001101110011", -- t[54131] = 18
      "0010010" when "01101001101110100", -- t[54132] = 18
      "0010010" when "01101001101110101", -- t[54133] = 18
      "0010010" when "01101001101110110", -- t[54134] = 18
      "0010010" when "01101001101110111", -- t[54135] = 18
      "0010010" when "01101001101111000", -- t[54136] = 18
      "0010010" when "01101001101111001", -- t[54137] = 18
      "0010010" when "01101001101111010", -- t[54138] = 18
      "0010010" when "01101001101111011", -- t[54139] = 18
      "0010010" when "01101001101111100", -- t[54140] = 18
      "0010010" when "01101001101111101", -- t[54141] = 18
      "0010010" when "01101001101111110", -- t[54142] = 18
      "0010010" when "01101001101111111", -- t[54143] = 18
      "0010010" when "01101001110000000", -- t[54144] = 18
      "0010010" when "01101001110000001", -- t[54145] = 18
      "0010010" when "01101001110000010", -- t[54146] = 18
      "0010010" when "01101001110000011", -- t[54147] = 18
      "0010010" when "01101001110000100", -- t[54148] = 18
      "0010010" when "01101001110000101", -- t[54149] = 18
      "0010010" when "01101001110000110", -- t[54150] = 18
      "0010010" when "01101001110000111", -- t[54151] = 18
      "0010010" when "01101001110001000", -- t[54152] = 18
      "0010010" when "01101001110001001", -- t[54153] = 18
      "0010010" when "01101001110001010", -- t[54154] = 18
      "0010010" when "01101001110001011", -- t[54155] = 18
      "0010010" when "01101001110001100", -- t[54156] = 18
      "0010010" when "01101001110001101", -- t[54157] = 18
      "0010010" when "01101001110001110", -- t[54158] = 18
      "0010010" when "01101001110001111", -- t[54159] = 18
      "0010010" when "01101001110010000", -- t[54160] = 18
      "0010010" when "01101001110010001", -- t[54161] = 18
      "0010010" when "01101001110010010", -- t[54162] = 18
      "0010010" when "01101001110010011", -- t[54163] = 18
      "0010010" when "01101001110010100", -- t[54164] = 18
      "0010010" when "01101001110010101", -- t[54165] = 18
      "0010010" when "01101001110010110", -- t[54166] = 18
      "0010010" when "01101001110010111", -- t[54167] = 18
      "0010010" when "01101001110011000", -- t[54168] = 18
      "0010010" when "01101001110011001", -- t[54169] = 18
      "0010010" when "01101001110011010", -- t[54170] = 18
      "0010010" when "01101001110011011", -- t[54171] = 18
      "0010010" when "01101001110011100", -- t[54172] = 18
      "0010010" when "01101001110011101", -- t[54173] = 18
      "0010010" when "01101001110011110", -- t[54174] = 18
      "0010010" when "01101001110011111", -- t[54175] = 18
      "0010010" when "01101001110100000", -- t[54176] = 18
      "0010010" when "01101001110100001", -- t[54177] = 18
      "0010010" when "01101001110100010", -- t[54178] = 18
      "0010010" when "01101001110100011", -- t[54179] = 18
      "0010010" when "01101001110100100", -- t[54180] = 18
      "0010010" when "01101001110100101", -- t[54181] = 18
      "0010010" when "01101001110100110", -- t[54182] = 18
      "0010010" when "01101001110100111", -- t[54183] = 18
      "0010010" when "01101001110101000", -- t[54184] = 18
      "0010010" when "01101001110101001", -- t[54185] = 18
      "0010010" when "01101001110101010", -- t[54186] = 18
      "0010010" when "01101001110101011", -- t[54187] = 18
      "0010010" when "01101001110101100", -- t[54188] = 18
      "0010010" when "01101001110101101", -- t[54189] = 18
      "0010010" when "01101001110101110", -- t[54190] = 18
      "0010010" when "01101001110101111", -- t[54191] = 18
      "0010010" when "01101001110110000", -- t[54192] = 18
      "0010010" when "01101001110110001", -- t[54193] = 18
      "0010010" when "01101001110110010", -- t[54194] = 18
      "0010010" when "01101001110110011", -- t[54195] = 18
      "0010010" when "01101001110110100", -- t[54196] = 18
      "0010010" when "01101001110110101", -- t[54197] = 18
      "0010010" when "01101001110110110", -- t[54198] = 18
      "0010010" when "01101001110110111", -- t[54199] = 18
      "0010010" when "01101001110111000", -- t[54200] = 18
      "0010010" when "01101001110111001", -- t[54201] = 18
      "0010010" when "01101001110111010", -- t[54202] = 18
      "0010010" when "01101001110111011", -- t[54203] = 18
      "0010010" when "01101001110111100", -- t[54204] = 18
      "0010010" when "01101001110111101", -- t[54205] = 18
      "0010010" when "01101001110111110", -- t[54206] = 18
      "0010010" when "01101001110111111", -- t[54207] = 18
      "0010010" when "01101001111000000", -- t[54208] = 18
      "0010010" when "01101001111000001", -- t[54209] = 18
      "0010010" when "01101001111000010", -- t[54210] = 18
      "0010010" when "01101001111000011", -- t[54211] = 18
      "0010010" when "01101001111000100", -- t[54212] = 18
      "0010010" when "01101001111000101", -- t[54213] = 18
      "0010010" when "01101001111000110", -- t[54214] = 18
      "0010010" when "01101001111000111", -- t[54215] = 18
      "0010010" when "01101001111001000", -- t[54216] = 18
      "0010010" when "01101001111001001", -- t[54217] = 18
      "0010010" when "01101001111001010", -- t[54218] = 18
      "0010010" when "01101001111001011", -- t[54219] = 18
      "0010010" when "01101001111001100", -- t[54220] = 18
      "0010010" when "01101001111001101", -- t[54221] = 18
      "0010010" when "01101001111001110", -- t[54222] = 18
      "0010010" when "01101001111001111", -- t[54223] = 18
      "0010010" when "01101001111010000", -- t[54224] = 18
      "0010010" when "01101001111010001", -- t[54225] = 18
      "0010010" when "01101001111010010", -- t[54226] = 18
      "0010010" when "01101001111010011", -- t[54227] = 18
      "0010010" when "01101001111010100", -- t[54228] = 18
      "0010010" when "01101001111010101", -- t[54229] = 18
      "0010010" when "01101001111010110", -- t[54230] = 18
      "0010010" when "01101001111010111", -- t[54231] = 18
      "0010010" when "01101001111011000", -- t[54232] = 18
      "0010010" when "01101001111011001", -- t[54233] = 18
      "0010010" when "01101001111011010", -- t[54234] = 18
      "0010010" when "01101001111011011", -- t[54235] = 18
      "0010010" when "01101001111011100", -- t[54236] = 18
      "0010010" when "01101001111011101", -- t[54237] = 18
      "0010010" when "01101001111011110", -- t[54238] = 18
      "0010010" when "01101001111011111", -- t[54239] = 18
      "0010010" when "01101001111100000", -- t[54240] = 18
      "0010010" when "01101001111100001", -- t[54241] = 18
      "0010010" when "01101001111100010", -- t[54242] = 18
      "0010010" when "01101001111100011", -- t[54243] = 18
      "0010010" when "01101001111100100", -- t[54244] = 18
      "0010010" when "01101001111100101", -- t[54245] = 18
      "0010010" when "01101001111100110", -- t[54246] = 18
      "0010010" when "01101001111100111", -- t[54247] = 18
      "0010010" when "01101001111101000", -- t[54248] = 18
      "0010010" when "01101001111101001", -- t[54249] = 18
      "0010010" when "01101001111101010", -- t[54250] = 18
      "0010010" when "01101001111101011", -- t[54251] = 18
      "0010010" when "01101001111101100", -- t[54252] = 18
      "0010010" when "01101001111101101", -- t[54253] = 18
      "0010010" when "01101001111101110", -- t[54254] = 18
      "0010010" when "01101001111101111", -- t[54255] = 18
      "0010010" when "01101001111110000", -- t[54256] = 18
      "0010010" when "01101001111110001", -- t[54257] = 18
      "0010010" when "01101001111110010", -- t[54258] = 18
      "0010010" when "01101001111110011", -- t[54259] = 18
      "0010010" when "01101001111110100", -- t[54260] = 18
      "0010010" when "01101001111110101", -- t[54261] = 18
      "0010010" when "01101001111110110", -- t[54262] = 18
      "0010010" when "01101001111110111", -- t[54263] = 18
      "0010010" when "01101001111111000", -- t[54264] = 18
      "0010010" when "01101001111111001", -- t[54265] = 18
      "0010010" when "01101001111111010", -- t[54266] = 18
      "0010010" when "01101001111111011", -- t[54267] = 18
      "0010010" when "01101001111111100", -- t[54268] = 18
      "0010010" when "01101001111111101", -- t[54269] = 18
      "0010010" when "01101001111111110", -- t[54270] = 18
      "0010010" when "01101001111111111", -- t[54271] = 18
      "0010010" when "01101010000000000", -- t[54272] = 18
      "0010010" when "01101010000000001", -- t[54273] = 18
      "0010010" when "01101010000000010", -- t[54274] = 18
      "0010010" when "01101010000000011", -- t[54275] = 18
      "0010010" when "01101010000000100", -- t[54276] = 18
      "0010010" when "01101010000000101", -- t[54277] = 18
      "0010010" when "01101010000000110", -- t[54278] = 18
      "0010010" when "01101010000000111", -- t[54279] = 18
      "0010010" when "01101010000001000", -- t[54280] = 18
      "0010010" when "01101010000001001", -- t[54281] = 18
      "0010010" when "01101010000001010", -- t[54282] = 18
      "0010010" when "01101010000001011", -- t[54283] = 18
      "0010010" when "01101010000001100", -- t[54284] = 18
      "0010010" when "01101010000001101", -- t[54285] = 18
      "0010010" when "01101010000001110", -- t[54286] = 18
      "0010010" when "01101010000001111", -- t[54287] = 18
      "0010010" when "01101010000010000", -- t[54288] = 18
      "0010010" when "01101010000010001", -- t[54289] = 18
      "0010010" when "01101010000010010", -- t[54290] = 18
      "0010010" when "01101010000010011", -- t[54291] = 18
      "0010010" when "01101010000010100", -- t[54292] = 18
      "0010010" when "01101010000010101", -- t[54293] = 18
      "0010010" when "01101010000010110", -- t[54294] = 18
      "0010010" when "01101010000010111", -- t[54295] = 18
      "0010010" when "01101010000011000", -- t[54296] = 18
      "0010010" when "01101010000011001", -- t[54297] = 18
      "0010010" when "01101010000011010", -- t[54298] = 18
      "0010010" when "01101010000011011", -- t[54299] = 18
      "0010010" when "01101010000011100", -- t[54300] = 18
      "0010010" when "01101010000011101", -- t[54301] = 18
      "0010010" when "01101010000011110", -- t[54302] = 18
      "0010010" when "01101010000011111", -- t[54303] = 18
      "0010010" when "01101010000100000", -- t[54304] = 18
      "0010010" when "01101010000100001", -- t[54305] = 18
      "0010010" when "01101010000100010", -- t[54306] = 18
      "0010010" when "01101010000100011", -- t[54307] = 18
      "0010010" when "01101010000100100", -- t[54308] = 18
      "0010010" when "01101010000100101", -- t[54309] = 18
      "0010010" when "01101010000100110", -- t[54310] = 18
      "0010010" when "01101010000100111", -- t[54311] = 18
      "0010010" when "01101010000101000", -- t[54312] = 18
      "0010010" when "01101010000101001", -- t[54313] = 18
      "0010010" when "01101010000101010", -- t[54314] = 18
      "0010010" when "01101010000101011", -- t[54315] = 18
      "0010010" when "01101010000101100", -- t[54316] = 18
      "0010010" when "01101010000101101", -- t[54317] = 18
      "0010010" when "01101010000101110", -- t[54318] = 18
      "0010010" when "01101010000101111", -- t[54319] = 18
      "0010010" when "01101010000110000", -- t[54320] = 18
      "0010010" when "01101010000110001", -- t[54321] = 18
      "0010010" when "01101010000110010", -- t[54322] = 18
      "0010010" when "01101010000110011", -- t[54323] = 18
      "0010010" when "01101010000110100", -- t[54324] = 18
      "0010010" when "01101010000110101", -- t[54325] = 18
      "0010010" when "01101010000110110", -- t[54326] = 18
      "0010010" when "01101010000110111", -- t[54327] = 18
      "0010010" when "01101010000111000", -- t[54328] = 18
      "0010010" when "01101010000111001", -- t[54329] = 18
      "0010010" when "01101010000111010", -- t[54330] = 18
      "0010010" when "01101010000111011", -- t[54331] = 18
      "0010010" when "01101010000111100", -- t[54332] = 18
      "0010010" when "01101010000111101", -- t[54333] = 18
      "0010010" when "01101010000111110", -- t[54334] = 18
      "0010010" when "01101010000111111", -- t[54335] = 18
      "0010010" when "01101010001000000", -- t[54336] = 18
      "0010010" when "01101010001000001", -- t[54337] = 18
      "0010010" when "01101010001000010", -- t[54338] = 18
      "0010010" when "01101010001000011", -- t[54339] = 18
      "0010010" when "01101010001000100", -- t[54340] = 18
      "0010010" when "01101010001000101", -- t[54341] = 18
      "0010010" when "01101010001000110", -- t[54342] = 18
      "0010010" when "01101010001000111", -- t[54343] = 18
      "0010010" when "01101010001001000", -- t[54344] = 18
      "0010010" when "01101010001001001", -- t[54345] = 18
      "0010010" when "01101010001001010", -- t[54346] = 18
      "0010010" when "01101010001001011", -- t[54347] = 18
      "0010010" when "01101010001001100", -- t[54348] = 18
      "0010010" when "01101010001001101", -- t[54349] = 18
      "0010010" when "01101010001001110", -- t[54350] = 18
      "0010010" when "01101010001001111", -- t[54351] = 18
      "0010010" when "01101010001010000", -- t[54352] = 18
      "0010010" when "01101010001010001", -- t[54353] = 18
      "0010010" when "01101010001010010", -- t[54354] = 18
      "0010010" when "01101010001010011", -- t[54355] = 18
      "0010010" when "01101010001010100", -- t[54356] = 18
      "0010010" when "01101010001010101", -- t[54357] = 18
      "0010010" when "01101010001010110", -- t[54358] = 18
      "0010010" when "01101010001010111", -- t[54359] = 18
      "0010010" when "01101010001011000", -- t[54360] = 18
      "0010010" when "01101010001011001", -- t[54361] = 18
      "0010010" when "01101010001011010", -- t[54362] = 18
      "0010010" when "01101010001011011", -- t[54363] = 18
      "0010010" when "01101010001011100", -- t[54364] = 18
      "0010010" when "01101010001011101", -- t[54365] = 18
      "0010010" when "01101010001011110", -- t[54366] = 18
      "0010010" when "01101010001011111", -- t[54367] = 18
      "0010010" when "01101010001100000", -- t[54368] = 18
      "0010010" when "01101010001100001", -- t[54369] = 18
      "0010010" when "01101010001100010", -- t[54370] = 18
      "0010010" when "01101010001100011", -- t[54371] = 18
      "0010010" when "01101010001100100", -- t[54372] = 18
      "0010010" when "01101010001100101", -- t[54373] = 18
      "0010010" when "01101010001100110", -- t[54374] = 18
      "0010010" when "01101010001100111", -- t[54375] = 18
      "0010010" when "01101010001101000", -- t[54376] = 18
      "0010010" when "01101010001101001", -- t[54377] = 18
      "0010010" when "01101010001101010", -- t[54378] = 18
      "0010010" when "01101010001101011", -- t[54379] = 18
      "0010010" when "01101010001101100", -- t[54380] = 18
      "0010010" when "01101010001101101", -- t[54381] = 18
      "0010010" when "01101010001101110", -- t[54382] = 18
      "0010010" when "01101010001101111", -- t[54383] = 18
      "0010010" when "01101010001110000", -- t[54384] = 18
      "0010010" when "01101010001110001", -- t[54385] = 18
      "0010010" when "01101010001110010", -- t[54386] = 18
      "0010010" when "01101010001110011", -- t[54387] = 18
      "0010010" when "01101010001110100", -- t[54388] = 18
      "0010010" when "01101010001110101", -- t[54389] = 18
      "0010010" when "01101010001110110", -- t[54390] = 18
      "0010010" when "01101010001110111", -- t[54391] = 18
      "0010010" when "01101010001111000", -- t[54392] = 18
      "0010010" when "01101010001111001", -- t[54393] = 18
      "0010010" when "01101010001111010", -- t[54394] = 18
      "0010010" when "01101010001111011", -- t[54395] = 18
      "0010010" when "01101010001111100", -- t[54396] = 18
      "0010010" when "01101010001111101", -- t[54397] = 18
      "0010010" when "01101010001111110", -- t[54398] = 18
      "0010010" when "01101010001111111", -- t[54399] = 18
      "0010010" when "01101010010000000", -- t[54400] = 18
      "0010010" when "01101010010000001", -- t[54401] = 18
      "0010010" when "01101010010000010", -- t[54402] = 18
      "0010010" when "01101010010000011", -- t[54403] = 18
      "0010010" when "01101010010000100", -- t[54404] = 18
      "0010010" when "01101010010000101", -- t[54405] = 18
      "0010010" when "01101010010000110", -- t[54406] = 18
      "0010010" when "01101010010000111", -- t[54407] = 18
      "0010010" when "01101010010001000", -- t[54408] = 18
      "0010010" when "01101010010001001", -- t[54409] = 18
      "0010010" when "01101010010001010", -- t[54410] = 18
      "0010010" when "01101010010001011", -- t[54411] = 18
      "0010010" when "01101010010001100", -- t[54412] = 18
      "0010010" when "01101010010001101", -- t[54413] = 18
      "0010010" when "01101010010001110", -- t[54414] = 18
      "0010010" when "01101010010001111", -- t[54415] = 18
      "0010010" when "01101010010010000", -- t[54416] = 18
      "0010010" when "01101010010010001", -- t[54417] = 18
      "0010010" when "01101010010010010", -- t[54418] = 18
      "0010010" when "01101010010010011", -- t[54419] = 18
      "0010010" when "01101010010010100", -- t[54420] = 18
      "0010010" when "01101010010010101", -- t[54421] = 18
      "0010010" when "01101010010010110", -- t[54422] = 18
      "0010010" when "01101010010010111", -- t[54423] = 18
      "0010010" when "01101010010011000", -- t[54424] = 18
      "0010010" when "01101010010011001", -- t[54425] = 18
      "0010010" when "01101010010011010", -- t[54426] = 18
      "0010010" when "01101010010011011", -- t[54427] = 18
      "0010010" when "01101010010011100", -- t[54428] = 18
      "0010010" when "01101010010011101", -- t[54429] = 18
      "0010010" when "01101010010011110", -- t[54430] = 18
      "0010010" when "01101010010011111", -- t[54431] = 18
      "0010010" when "01101010010100000", -- t[54432] = 18
      "0010010" when "01101010010100001", -- t[54433] = 18
      "0010010" when "01101010010100010", -- t[54434] = 18
      "0010010" when "01101010010100011", -- t[54435] = 18
      "0010010" when "01101010010100100", -- t[54436] = 18
      "0010010" when "01101010010100101", -- t[54437] = 18
      "0010010" when "01101010010100110", -- t[54438] = 18
      "0010010" when "01101010010100111", -- t[54439] = 18
      "0010010" when "01101010010101000", -- t[54440] = 18
      "0010010" when "01101010010101001", -- t[54441] = 18
      "0010010" when "01101010010101010", -- t[54442] = 18
      "0010010" when "01101010010101011", -- t[54443] = 18
      "0010010" when "01101010010101100", -- t[54444] = 18
      "0010010" when "01101010010101101", -- t[54445] = 18
      "0010010" when "01101010010101110", -- t[54446] = 18
      "0010010" when "01101010010101111", -- t[54447] = 18
      "0010010" when "01101010010110000", -- t[54448] = 18
      "0010010" when "01101010010110001", -- t[54449] = 18
      "0010010" when "01101010010110010", -- t[54450] = 18
      "0010010" when "01101010010110011", -- t[54451] = 18
      "0010010" when "01101010010110100", -- t[54452] = 18
      "0010010" when "01101010010110101", -- t[54453] = 18
      "0010010" when "01101010010110110", -- t[54454] = 18
      "0010010" when "01101010010110111", -- t[54455] = 18
      "0010010" when "01101010010111000", -- t[54456] = 18
      "0010010" when "01101010010111001", -- t[54457] = 18
      "0010010" when "01101010010111010", -- t[54458] = 18
      "0010010" when "01101010010111011", -- t[54459] = 18
      "0010010" when "01101010010111100", -- t[54460] = 18
      "0010010" when "01101010010111101", -- t[54461] = 18
      "0010010" when "01101010010111110", -- t[54462] = 18
      "0010010" when "01101010010111111", -- t[54463] = 18
      "0010010" when "01101010011000000", -- t[54464] = 18
      "0010010" when "01101010011000001", -- t[54465] = 18
      "0010010" when "01101010011000010", -- t[54466] = 18
      "0010010" when "01101010011000011", -- t[54467] = 18
      "0010010" when "01101010011000100", -- t[54468] = 18
      "0010010" when "01101010011000101", -- t[54469] = 18
      "0010010" when "01101010011000110", -- t[54470] = 18
      "0010010" when "01101010011000111", -- t[54471] = 18
      "0010010" when "01101010011001000", -- t[54472] = 18
      "0010010" when "01101010011001001", -- t[54473] = 18
      "0010010" when "01101010011001010", -- t[54474] = 18
      "0010010" when "01101010011001011", -- t[54475] = 18
      "0010010" when "01101010011001100", -- t[54476] = 18
      "0010010" when "01101010011001101", -- t[54477] = 18
      "0010010" when "01101010011001110", -- t[54478] = 18
      "0010010" when "01101010011001111", -- t[54479] = 18
      "0010010" when "01101010011010000", -- t[54480] = 18
      "0010010" when "01101010011010001", -- t[54481] = 18
      "0010010" when "01101010011010010", -- t[54482] = 18
      "0010010" when "01101010011010011", -- t[54483] = 18
      "0010010" when "01101010011010100", -- t[54484] = 18
      "0010010" when "01101010011010101", -- t[54485] = 18
      "0010010" when "01101010011010110", -- t[54486] = 18
      "0010010" when "01101010011010111", -- t[54487] = 18
      "0010010" when "01101010011011000", -- t[54488] = 18
      "0010010" when "01101010011011001", -- t[54489] = 18
      "0010010" when "01101010011011010", -- t[54490] = 18
      "0010010" when "01101010011011011", -- t[54491] = 18
      "0010010" when "01101010011011100", -- t[54492] = 18
      "0010010" when "01101010011011101", -- t[54493] = 18
      "0010010" when "01101010011011110", -- t[54494] = 18
      "0010010" when "01101010011011111", -- t[54495] = 18
      "0010010" when "01101010011100000", -- t[54496] = 18
      "0010010" when "01101010011100001", -- t[54497] = 18
      "0010010" when "01101010011100010", -- t[54498] = 18
      "0010010" when "01101010011100011", -- t[54499] = 18
      "0010010" when "01101010011100100", -- t[54500] = 18
      "0010010" when "01101010011100101", -- t[54501] = 18
      "0010010" when "01101010011100110", -- t[54502] = 18
      "0010010" when "01101010011100111", -- t[54503] = 18
      "0010010" when "01101010011101000", -- t[54504] = 18
      "0010010" when "01101010011101001", -- t[54505] = 18
      "0010010" when "01101010011101010", -- t[54506] = 18
      "0010010" when "01101010011101011", -- t[54507] = 18
      "0010010" when "01101010011101100", -- t[54508] = 18
      "0010010" when "01101010011101101", -- t[54509] = 18
      "0010010" when "01101010011101110", -- t[54510] = 18
      "0010010" when "01101010011101111", -- t[54511] = 18
      "0010010" when "01101010011110000", -- t[54512] = 18
      "0010010" when "01101010011110001", -- t[54513] = 18
      "0010010" when "01101010011110010", -- t[54514] = 18
      "0010010" when "01101010011110011", -- t[54515] = 18
      "0010010" when "01101010011110100", -- t[54516] = 18
      "0010010" when "01101010011110101", -- t[54517] = 18
      "0010010" when "01101010011110110", -- t[54518] = 18
      "0010010" when "01101010011110111", -- t[54519] = 18
      "0010010" when "01101010011111000", -- t[54520] = 18
      "0010010" when "01101010011111001", -- t[54521] = 18
      "0010010" when "01101010011111010", -- t[54522] = 18
      "0010010" when "01101010011111011", -- t[54523] = 18
      "0010010" when "01101010011111100", -- t[54524] = 18
      "0010010" when "01101010011111101", -- t[54525] = 18
      "0010010" when "01101010011111110", -- t[54526] = 18
      "0010010" when "01101010011111111", -- t[54527] = 18
      "0010010" when "01101010100000000", -- t[54528] = 18
      "0010010" when "01101010100000001", -- t[54529] = 18
      "0010010" when "01101010100000010", -- t[54530] = 18
      "0010010" when "01101010100000011", -- t[54531] = 18
      "0010010" when "01101010100000100", -- t[54532] = 18
      "0010010" when "01101010100000101", -- t[54533] = 18
      "0010010" when "01101010100000110", -- t[54534] = 18
      "0010010" when "01101010100000111", -- t[54535] = 18
      "0010010" when "01101010100001000", -- t[54536] = 18
      "0010010" when "01101010100001001", -- t[54537] = 18
      "0010010" when "01101010100001010", -- t[54538] = 18
      "0010010" when "01101010100001011", -- t[54539] = 18
      "0010010" when "01101010100001100", -- t[54540] = 18
      "0010010" when "01101010100001101", -- t[54541] = 18
      "0010010" when "01101010100001110", -- t[54542] = 18
      "0010010" when "01101010100001111", -- t[54543] = 18
      "0010010" when "01101010100010000", -- t[54544] = 18
      "0010010" when "01101010100010001", -- t[54545] = 18
      "0010010" when "01101010100010010", -- t[54546] = 18
      "0010010" when "01101010100010011", -- t[54547] = 18
      "0010010" when "01101010100010100", -- t[54548] = 18
      "0010010" when "01101010100010101", -- t[54549] = 18
      "0010010" when "01101010100010110", -- t[54550] = 18
      "0010010" when "01101010100010111", -- t[54551] = 18
      "0010010" when "01101010100011000", -- t[54552] = 18
      "0010010" when "01101010100011001", -- t[54553] = 18
      "0010010" when "01101010100011010", -- t[54554] = 18
      "0010010" when "01101010100011011", -- t[54555] = 18
      "0010010" when "01101010100011100", -- t[54556] = 18
      "0010010" when "01101010100011101", -- t[54557] = 18
      "0010010" when "01101010100011110", -- t[54558] = 18
      "0010010" when "01101010100011111", -- t[54559] = 18
      "0010010" when "01101010100100000", -- t[54560] = 18
      "0010010" when "01101010100100001", -- t[54561] = 18
      "0010010" when "01101010100100010", -- t[54562] = 18
      "0010010" when "01101010100100011", -- t[54563] = 18
      "0010010" when "01101010100100100", -- t[54564] = 18
      "0010010" when "01101010100100101", -- t[54565] = 18
      "0010010" when "01101010100100110", -- t[54566] = 18
      "0010010" when "01101010100100111", -- t[54567] = 18
      "0010010" when "01101010100101000", -- t[54568] = 18
      "0010010" when "01101010100101001", -- t[54569] = 18
      "0010010" when "01101010100101010", -- t[54570] = 18
      "0010010" when "01101010100101011", -- t[54571] = 18
      "0010010" when "01101010100101100", -- t[54572] = 18
      "0010010" when "01101010100101101", -- t[54573] = 18
      "0010010" when "01101010100101110", -- t[54574] = 18
      "0010010" when "01101010100101111", -- t[54575] = 18
      "0010010" when "01101010100110000", -- t[54576] = 18
      "0010010" when "01101010100110001", -- t[54577] = 18
      "0010010" when "01101010100110010", -- t[54578] = 18
      "0010010" when "01101010100110011", -- t[54579] = 18
      "0010010" when "01101010100110100", -- t[54580] = 18
      "0010010" when "01101010100110101", -- t[54581] = 18
      "0010010" when "01101010100110110", -- t[54582] = 18
      "0010010" when "01101010100110111", -- t[54583] = 18
      "0010010" when "01101010100111000", -- t[54584] = 18
      "0010010" when "01101010100111001", -- t[54585] = 18
      "0010010" when "01101010100111010", -- t[54586] = 18
      "0010010" when "01101010100111011", -- t[54587] = 18
      "0010010" when "01101010100111100", -- t[54588] = 18
      "0010010" when "01101010100111101", -- t[54589] = 18
      "0010010" when "01101010100111110", -- t[54590] = 18
      "0010010" when "01101010100111111", -- t[54591] = 18
      "0010010" when "01101010101000000", -- t[54592] = 18
      "0010010" when "01101010101000001", -- t[54593] = 18
      "0010010" when "01101010101000010", -- t[54594] = 18
      "0010010" when "01101010101000011", -- t[54595] = 18
      "0010010" when "01101010101000100", -- t[54596] = 18
      "0010010" when "01101010101000101", -- t[54597] = 18
      "0010010" when "01101010101000110", -- t[54598] = 18
      "0010010" when "01101010101000111", -- t[54599] = 18
      "0010010" when "01101010101001000", -- t[54600] = 18
      "0010010" when "01101010101001001", -- t[54601] = 18
      "0010010" when "01101010101001010", -- t[54602] = 18
      "0010010" when "01101010101001011", -- t[54603] = 18
      "0010010" when "01101010101001100", -- t[54604] = 18
      "0010010" when "01101010101001101", -- t[54605] = 18
      "0010010" when "01101010101001110", -- t[54606] = 18
      "0010010" when "01101010101001111", -- t[54607] = 18
      "0010010" when "01101010101010000", -- t[54608] = 18
      "0010010" when "01101010101010001", -- t[54609] = 18
      "0010010" when "01101010101010010", -- t[54610] = 18
      "0010010" when "01101010101010011", -- t[54611] = 18
      "0010010" when "01101010101010100", -- t[54612] = 18
      "0010010" when "01101010101010101", -- t[54613] = 18
      "0010010" when "01101010101010110", -- t[54614] = 18
      "0010010" when "01101010101010111", -- t[54615] = 18
      "0010010" when "01101010101011000", -- t[54616] = 18
      "0010010" when "01101010101011001", -- t[54617] = 18
      "0010010" when "01101010101011010", -- t[54618] = 18
      "0010010" when "01101010101011011", -- t[54619] = 18
      "0010010" when "01101010101011100", -- t[54620] = 18
      "0010010" when "01101010101011101", -- t[54621] = 18
      "0010010" when "01101010101011110", -- t[54622] = 18
      "0010010" when "01101010101011111", -- t[54623] = 18
      "0010010" when "01101010101100000", -- t[54624] = 18
      "0010010" when "01101010101100001", -- t[54625] = 18
      "0010010" when "01101010101100010", -- t[54626] = 18
      "0010010" when "01101010101100011", -- t[54627] = 18
      "0010010" when "01101010101100100", -- t[54628] = 18
      "0010010" when "01101010101100101", -- t[54629] = 18
      "0010010" when "01101010101100110", -- t[54630] = 18
      "0010010" when "01101010101100111", -- t[54631] = 18
      "0010010" when "01101010101101000", -- t[54632] = 18
      "0010010" when "01101010101101001", -- t[54633] = 18
      "0010010" when "01101010101101010", -- t[54634] = 18
      "0010010" when "01101010101101011", -- t[54635] = 18
      "0010010" when "01101010101101100", -- t[54636] = 18
      "0010010" when "01101010101101101", -- t[54637] = 18
      "0010010" when "01101010101101110", -- t[54638] = 18
      "0010010" when "01101010101101111", -- t[54639] = 18
      "0010010" when "01101010101110000", -- t[54640] = 18
      "0010010" when "01101010101110001", -- t[54641] = 18
      "0010010" when "01101010101110010", -- t[54642] = 18
      "0010010" when "01101010101110011", -- t[54643] = 18
      "0010010" when "01101010101110100", -- t[54644] = 18
      "0010010" when "01101010101110101", -- t[54645] = 18
      "0010010" when "01101010101110110", -- t[54646] = 18
      "0010010" when "01101010101110111", -- t[54647] = 18
      "0010010" when "01101010101111000", -- t[54648] = 18
      "0010010" when "01101010101111001", -- t[54649] = 18
      "0010010" when "01101010101111010", -- t[54650] = 18
      "0010010" when "01101010101111011", -- t[54651] = 18
      "0010010" when "01101010101111100", -- t[54652] = 18
      "0010010" when "01101010101111101", -- t[54653] = 18
      "0010010" when "01101010101111110", -- t[54654] = 18
      "0010010" when "01101010101111111", -- t[54655] = 18
      "0010010" when "01101010110000000", -- t[54656] = 18
      "0010010" when "01101010110000001", -- t[54657] = 18
      "0010010" when "01101010110000010", -- t[54658] = 18
      "0010010" when "01101010110000011", -- t[54659] = 18
      "0010010" when "01101010110000100", -- t[54660] = 18
      "0010010" when "01101010110000101", -- t[54661] = 18
      "0010010" when "01101010110000110", -- t[54662] = 18
      "0010010" when "01101010110000111", -- t[54663] = 18
      "0010010" when "01101010110001000", -- t[54664] = 18
      "0010010" when "01101010110001001", -- t[54665] = 18
      "0010010" when "01101010110001010", -- t[54666] = 18
      "0010010" when "01101010110001011", -- t[54667] = 18
      "0010010" when "01101010110001100", -- t[54668] = 18
      "0010010" when "01101010110001101", -- t[54669] = 18
      "0010010" when "01101010110001110", -- t[54670] = 18
      "0010010" when "01101010110001111", -- t[54671] = 18
      "0010010" when "01101010110010000", -- t[54672] = 18
      "0010010" when "01101010110010001", -- t[54673] = 18
      "0010010" when "01101010110010010", -- t[54674] = 18
      "0010010" when "01101010110010011", -- t[54675] = 18
      "0010010" when "01101010110010100", -- t[54676] = 18
      "0010010" when "01101010110010101", -- t[54677] = 18
      "0010010" when "01101010110010110", -- t[54678] = 18
      "0010010" when "01101010110010111", -- t[54679] = 18
      "0010010" when "01101010110011000", -- t[54680] = 18
      "0010010" when "01101010110011001", -- t[54681] = 18
      "0010010" when "01101010110011010", -- t[54682] = 18
      "0010010" when "01101010110011011", -- t[54683] = 18
      "0010010" when "01101010110011100", -- t[54684] = 18
      "0010010" when "01101010110011101", -- t[54685] = 18
      "0010010" when "01101010110011110", -- t[54686] = 18
      "0010010" when "01101010110011111", -- t[54687] = 18
      "0010010" when "01101010110100000", -- t[54688] = 18
      "0010010" when "01101010110100001", -- t[54689] = 18
      "0010010" when "01101010110100010", -- t[54690] = 18
      "0010010" when "01101010110100011", -- t[54691] = 18
      "0010010" when "01101010110100100", -- t[54692] = 18
      "0010010" when "01101010110100101", -- t[54693] = 18
      "0010010" when "01101010110100110", -- t[54694] = 18
      "0010010" when "01101010110100111", -- t[54695] = 18
      "0010010" when "01101010110101000", -- t[54696] = 18
      "0010010" when "01101010110101001", -- t[54697] = 18
      "0010010" when "01101010110101010", -- t[54698] = 18
      "0010010" when "01101010110101011", -- t[54699] = 18
      "0010010" when "01101010110101100", -- t[54700] = 18
      "0010010" when "01101010110101101", -- t[54701] = 18
      "0010010" when "01101010110101110", -- t[54702] = 18
      "0010010" when "01101010110101111", -- t[54703] = 18
      "0010010" when "01101010110110000", -- t[54704] = 18
      "0010010" when "01101010110110001", -- t[54705] = 18
      "0010010" when "01101010110110010", -- t[54706] = 18
      "0010010" when "01101010110110011", -- t[54707] = 18
      "0010010" when "01101010110110100", -- t[54708] = 18
      "0010010" when "01101010110110101", -- t[54709] = 18
      "0010010" when "01101010110110110", -- t[54710] = 18
      "0010010" when "01101010110110111", -- t[54711] = 18
      "0010010" when "01101010110111000", -- t[54712] = 18
      "0010010" when "01101010110111001", -- t[54713] = 18
      "0010010" when "01101010110111010", -- t[54714] = 18
      "0010010" when "01101010110111011", -- t[54715] = 18
      "0010010" when "01101010110111100", -- t[54716] = 18
      "0010010" when "01101010110111101", -- t[54717] = 18
      "0010010" when "01101010110111110", -- t[54718] = 18
      "0010011" when "01101010110111111", -- t[54719] = 19
      "0010011" when "01101010111000000", -- t[54720] = 19
      "0010011" when "01101010111000001", -- t[54721] = 19
      "0010011" when "01101010111000010", -- t[54722] = 19
      "0010011" when "01101010111000011", -- t[54723] = 19
      "0010011" when "01101010111000100", -- t[54724] = 19
      "0010011" when "01101010111000101", -- t[54725] = 19
      "0010011" when "01101010111000110", -- t[54726] = 19
      "0010011" when "01101010111000111", -- t[54727] = 19
      "0010011" when "01101010111001000", -- t[54728] = 19
      "0010011" when "01101010111001001", -- t[54729] = 19
      "0010011" when "01101010111001010", -- t[54730] = 19
      "0010011" when "01101010111001011", -- t[54731] = 19
      "0010011" when "01101010111001100", -- t[54732] = 19
      "0010011" when "01101010111001101", -- t[54733] = 19
      "0010011" when "01101010111001110", -- t[54734] = 19
      "0010011" when "01101010111001111", -- t[54735] = 19
      "0010011" when "01101010111010000", -- t[54736] = 19
      "0010011" when "01101010111010001", -- t[54737] = 19
      "0010011" when "01101010111010010", -- t[54738] = 19
      "0010011" when "01101010111010011", -- t[54739] = 19
      "0010011" when "01101010111010100", -- t[54740] = 19
      "0010011" when "01101010111010101", -- t[54741] = 19
      "0010011" when "01101010111010110", -- t[54742] = 19
      "0010011" when "01101010111010111", -- t[54743] = 19
      "0010011" when "01101010111011000", -- t[54744] = 19
      "0010011" when "01101010111011001", -- t[54745] = 19
      "0010011" when "01101010111011010", -- t[54746] = 19
      "0010011" when "01101010111011011", -- t[54747] = 19
      "0010011" when "01101010111011100", -- t[54748] = 19
      "0010011" when "01101010111011101", -- t[54749] = 19
      "0010011" when "01101010111011110", -- t[54750] = 19
      "0010011" when "01101010111011111", -- t[54751] = 19
      "0010011" when "01101010111100000", -- t[54752] = 19
      "0010011" when "01101010111100001", -- t[54753] = 19
      "0010011" when "01101010111100010", -- t[54754] = 19
      "0010011" when "01101010111100011", -- t[54755] = 19
      "0010011" when "01101010111100100", -- t[54756] = 19
      "0010011" when "01101010111100101", -- t[54757] = 19
      "0010011" when "01101010111100110", -- t[54758] = 19
      "0010011" when "01101010111100111", -- t[54759] = 19
      "0010011" when "01101010111101000", -- t[54760] = 19
      "0010011" when "01101010111101001", -- t[54761] = 19
      "0010011" when "01101010111101010", -- t[54762] = 19
      "0010011" when "01101010111101011", -- t[54763] = 19
      "0010011" when "01101010111101100", -- t[54764] = 19
      "0010011" when "01101010111101101", -- t[54765] = 19
      "0010011" when "01101010111101110", -- t[54766] = 19
      "0010011" when "01101010111101111", -- t[54767] = 19
      "0010011" when "01101010111110000", -- t[54768] = 19
      "0010011" when "01101010111110001", -- t[54769] = 19
      "0010011" when "01101010111110010", -- t[54770] = 19
      "0010011" when "01101010111110011", -- t[54771] = 19
      "0010011" when "01101010111110100", -- t[54772] = 19
      "0010011" when "01101010111110101", -- t[54773] = 19
      "0010011" when "01101010111110110", -- t[54774] = 19
      "0010011" when "01101010111110111", -- t[54775] = 19
      "0010011" when "01101010111111000", -- t[54776] = 19
      "0010011" when "01101010111111001", -- t[54777] = 19
      "0010011" when "01101010111111010", -- t[54778] = 19
      "0010011" when "01101010111111011", -- t[54779] = 19
      "0010011" when "01101010111111100", -- t[54780] = 19
      "0010011" when "01101010111111101", -- t[54781] = 19
      "0010011" when "01101010111111110", -- t[54782] = 19
      "0010011" when "01101010111111111", -- t[54783] = 19
      "0010011" when "01101011000000000", -- t[54784] = 19
      "0010011" when "01101011000000001", -- t[54785] = 19
      "0010011" when "01101011000000010", -- t[54786] = 19
      "0010011" when "01101011000000011", -- t[54787] = 19
      "0010011" when "01101011000000100", -- t[54788] = 19
      "0010011" when "01101011000000101", -- t[54789] = 19
      "0010011" when "01101011000000110", -- t[54790] = 19
      "0010011" when "01101011000000111", -- t[54791] = 19
      "0010011" when "01101011000001000", -- t[54792] = 19
      "0010011" when "01101011000001001", -- t[54793] = 19
      "0010011" when "01101011000001010", -- t[54794] = 19
      "0010011" when "01101011000001011", -- t[54795] = 19
      "0010011" when "01101011000001100", -- t[54796] = 19
      "0010011" when "01101011000001101", -- t[54797] = 19
      "0010011" when "01101011000001110", -- t[54798] = 19
      "0010011" when "01101011000001111", -- t[54799] = 19
      "0010011" when "01101011000010000", -- t[54800] = 19
      "0010011" when "01101011000010001", -- t[54801] = 19
      "0010011" when "01101011000010010", -- t[54802] = 19
      "0010011" when "01101011000010011", -- t[54803] = 19
      "0010011" when "01101011000010100", -- t[54804] = 19
      "0010011" when "01101011000010101", -- t[54805] = 19
      "0010011" when "01101011000010110", -- t[54806] = 19
      "0010011" when "01101011000010111", -- t[54807] = 19
      "0010011" when "01101011000011000", -- t[54808] = 19
      "0010011" when "01101011000011001", -- t[54809] = 19
      "0010011" when "01101011000011010", -- t[54810] = 19
      "0010011" when "01101011000011011", -- t[54811] = 19
      "0010011" when "01101011000011100", -- t[54812] = 19
      "0010011" when "01101011000011101", -- t[54813] = 19
      "0010011" when "01101011000011110", -- t[54814] = 19
      "0010011" when "01101011000011111", -- t[54815] = 19
      "0010011" when "01101011000100000", -- t[54816] = 19
      "0010011" when "01101011000100001", -- t[54817] = 19
      "0010011" when "01101011000100010", -- t[54818] = 19
      "0010011" when "01101011000100011", -- t[54819] = 19
      "0010011" when "01101011000100100", -- t[54820] = 19
      "0010011" when "01101011000100101", -- t[54821] = 19
      "0010011" when "01101011000100110", -- t[54822] = 19
      "0010011" when "01101011000100111", -- t[54823] = 19
      "0010011" when "01101011000101000", -- t[54824] = 19
      "0010011" when "01101011000101001", -- t[54825] = 19
      "0010011" when "01101011000101010", -- t[54826] = 19
      "0010011" when "01101011000101011", -- t[54827] = 19
      "0010011" when "01101011000101100", -- t[54828] = 19
      "0010011" when "01101011000101101", -- t[54829] = 19
      "0010011" when "01101011000101110", -- t[54830] = 19
      "0010011" when "01101011000101111", -- t[54831] = 19
      "0010011" when "01101011000110000", -- t[54832] = 19
      "0010011" when "01101011000110001", -- t[54833] = 19
      "0010011" when "01101011000110010", -- t[54834] = 19
      "0010011" when "01101011000110011", -- t[54835] = 19
      "0010011" when "01101011000110100", -- t[54836] = 19
      "0010011" when "01101011000110101", -- t[54837] = 19
      "0010011" when "01101011000110110", -- t[54838] = 19
      "0010011" when "01101011000110111", -- t[54839] = 19
      "0010011" when "01101011000111000", -- t[54840] = 19
      "0010011" when "01101011000111001", -- t[54841] = 19
      "0010011" when "01101011000111010", -- t[54842] = 19
      "0010011" when "01101011000111011", -- t[54843] = 19
      "0010011" when "01101011000111100", -- t[54844] = 19
      "0010011" when "01101011000111101", -- t[54845] = 19
      "0010011" when "01101011000111110", -- t[54846] = 19
      "0010011" when "01101011000111111", -- t[54847] = 19
      "0010011" when "01101011001000000", -- t[54848] = 19
      "0010011" when "01101011001000001", -- t[54849] = 19
      "0010011" when "01101011001000010", -- t[54850] = 19
      "0010011" when "01101011001000011", -- t[54851] = 19
      "0010011" when "01101011001000100", -- t[54852] = 19
      "0010011" when "01101011001000101", -- t[54853] = 19
      "0010011" when "01101011001000110", -- t[54854] = 19
      "0010011" when "01101011001000111", -- t[54855] = 19
      "0010011" when "01101011001001000", -- t[54856] = 19
      "0010011" when "01101011001001001", -- t[54857] = 19
      "0010011" when "01101011001001010", -- t[54858] = 19
      "0010011" when "01101011001001011", -- t[54859] = 19
      "0010011" when "01101011001001100", -- t[54860] = 19
      "0010011" when "01101011001001101", -- t[54861] = 19
      "0010011" when "01101011001001110", -- t[54862] = 19
      "0010011" when "01101011001001111", -- t[54863] = 19
      "0010011" when "01101011001010000", -- t[54864] = 19
      "0010011" when "01101011001010001", -- t[54865] = 19
      "0010011" when "01101011001010010", -- t[54866] = 19
      "0010011" when "01101011001010011", -- t[54867] = 19
      "0010011" when "01101011001010100", -- t[54868] = 19
      "0010011" when "01101011001010101", -- t[54869] = 19
      "0010011" when "01101011001010110", -- t[54870] = 19
      "0010011" when "01101011001010111", -- t[54871] = 19
      "0010011" when "01101011001011000", -- t[54872] = 19
      "0010011" when "01101011001011001", -- t[54873] = 19
      "0010011" when "01101011001011010", -- t[54874] = 19
      "0010011" when "01101011001011011", -- t[54875] = 19
      "0010011" when "01101011001011100", -- t[54876] = 19
      "0010011" when "01101011001011101", -- t[54877] = 19
      "0010011" when "01101011001011110", -- t[54878] = 19
      "0010011" when "01101011001011111", -- t[54879] = 19
      "0010011" when "01101011001100000", -- t[54880] = 19
      "0010011" when "01101011001100001", -- t[54881] = 19
      "0010011" when "01101011001100010", -- t[54882] = 19
      "0010011" when "01101011001100011", -- t[54883] = 19
      "0010011" when "01101011001100100", -- t[54884] = 19
      "0010011" when "01101011001100101", -- t[54885] = 19
      "0010011" when "01101011001100110", -- t[54886] = 19
      "0010011" when "01101011001100111", -- t[54887] = 19
      "0010011" when "01101011001101000", -- t[54888] = 19
      "0010011" when "01101011001101001", -- t[54889] = 19
      "0010011" when "01101011001101010", -- t[54890] = 19
      "0010011" when "01101011001101011", -- t[54891] = 19
      "0010011" when "01101011001101100", -- t[54892] = 19
      "0010011" when "01101011001101101", -- t[54893] = 19
      "0010011" when "01101011001101110", -- t[54894] = 19
      "0010011" when "01101011001101111", -- t[54895] = 19
      "0010011" when "01101011001110000", -- t[54896] = 19
      "0010011" when "01101011001110001", -- t[54897] = 19
      "0010011" when "01101011001110010", -- t[54898] = 19
      "0010011" when "01101011001110011", -- t[54899] = 19
      "0010011" when "01101011001110100", -- t[54900] = 19
      "0010011" when "01101011001110101", -- t[54901] = 19
      "0010011" when "01101011001110110", -- t[54902] = 19
      "0010011" when "01101011001110111", -- t[54903] = 19
      "0010011" when "01101011001111000", -- t[54904] = 19
      "0010011" when "01101011001111001", -- t[54905] = 19
      "0010011" when "01101011001111010", -- t[54906] = 19
      "0010011" when "01101011001111011", -- t[54907] = 19
      "0010011" when "01101011001111100", -- t[54908] = 19
      "0010011" when "01101011001111101", -- t[54909] = 19
      "0010011" when "01101011001111110", -- t[54910] = 19
      "0010011" when "01101011001111111", -- t[54911] = 19
      "0010011" when "01101011010000000", -- t[54912] = 19
      "0010011" when "01101011010000001", -- t[54913] = 19
      "0010011" when "01101011010000010", -- t[54914] = 19
      "0010011" when "01101011010000011", -- t[54915] = 19
      "0010011" when "01101011010000100", -- t[54916] = 19
      "0010011" when "01101011010000101", -- t[54917] = 19
      "0010011" when "01101011010000110", -- t[54918] = 19
      "0010011" when "01101011010000111", -- t[54919] = 19
      "0010011" when "01101011010001000", -- t[54920] = 19
      "0010011" when "01101011010001001", -- t[54921] = 19
      "0010011" when "01101011010001010", -- t[54922] = 19
      "0010011" when "01101011010001011", -- t[54923] = 19
      "0010011" when "01101011010001100", -- t[54924] = 19
      "0010011" when "01101011010001101", -- t[54925] = 19
      "0010011" when "01101011010001110", -- t[54926] = 19
      "0010011" when "01101011010001111", -- t[54927] = 19
      "0010011" when "01101011010010000", -- t[54928] = 19
      "0010011" when "01101011010010001", -- t[54929] = 19
      "0010011" when "01101011010010010", -- t[54930] = 19
      "0010011" when "01101011010010011", -- t[54931] = 19
      "0010011" when "01101011010010100", -- t[54932] = 19
      "0010011" when "01101011010010101", -- t[54933] = 19
      "0010011" when "01101011010010110", -- t[54934] = 19
      "0010011" when "01101011010010111", -- t[54935] = 19
      "0010011" when "01101011010011000", -- t[54936] = 19
      "0010011" when "01101011010011001", -- t[54937] = 19
      "0010011" when "01101011010011010", -- t[54938] = 19
      "0010011" when "01101011010011011", -- t[54939] = 19
      "0010011" when "01101011010011100", -- t[54940] = 19
      "0010011" when "01101011010011101", -- t[54941] = 19
      "0010011" when "01101011010011110", -- t[54942] = 19
      "0010011" when "01101011010011111", -- t[54943] = 19
      "0010011" when "01101011010100000", -- t[54944] = 19
      "0010011" when "01101011010100001", -- t[54945] = 19
      "0010011" when "01101011010100010", -- t[54946] = 19
      "0010011" when "01101011010100011", -- t[54947] = 19
      "0010011" when "01101011010100100", -- t[54948] = 19
      "0010011" when "01101011010100101", -- t[54949] = 19
      "0010011" when "01101011010100110", -- t[54950] = 19
      "0010011" when "01101011010100111", -- t[54951] = 19
      "0010011" when "01101011010101000", -- t[54952] = 19
      "0010011" when "01101011010101001", -- t[54953] = 19
      "0010011" when "01101011010101010", -- t[54954] = 19
      "0010011" when "01101011010101011", -- t[54955] = 19
      "0010011" when "01101011010101100", -- t[54956] = 19
      "0010011" when "01101011010101101", -- t[54957] = 19
      "0010011" when "01101011010101110", -- t[54958] = 19
      "0010011" when "01101011010101111", -- t[54959] = 19
      "0010011" when "01101011010110000", -- t[54960] = 19
      "0010011" when "01101011010110001", -- t[54961] = 19
      "0010011" when "01101011010110010", -- t[54962] = 19
      "0010011" when "01101011010110011", -- t[54963] = 19
      "0010011" when "01101011010110100", -- t[54964] = 19
      "0010011" when "01101011010110101", -- t[54965] = 19
      "0010011" when "01101011010110110", -- t[54966] = 19
      "0010011" when "01101011010110111", -- t[54967] = 19
      "0010011" when "01101011010111000", -- t[54968] = 19
      "0010011" when "01101011010111001", -- t[54969] = 19
      "0010011" when "01101011010111010", -- t[54970] = 19
      "0010011" when "01101011010111011", -- t[54971] = 19
      "0010011" when "01101011010111100", -- t[54972] = 19
      "0010011" when "01101011010111101", -- t[54973] = 19
      "0010011" when "01101011010111110", -- t[54974] = 19
      "0010011" when "01101011010111111", -- t[54975] = 19
      "0010011" when "01101011011000000", -- t[54976] = 19
      "0010011" when "01101011011000001", -- t[54977] = 19
      "0010011" when "01101011011000010", -- t[54978] = 19
      "0010011" when "01101011011000011", -- t[54979] = 19
      "0010011" when "01101011011000100", -- t[54980] = 19
      "0010011" when "01101011011000101", -- t[54981] = 19
      "0010011" when "01101011011000110", -- t[54982] = 19
      "0010011" when "01101011011000111", -- t[54983] = 19
      "0010011" when "01101011011001000", -- t[54984] = 19
      "0010011" when "01101011011001001", -- t[54985] = 19
      "0010011" when "01101011011001010", -- t[54986] = 19
      "0010011" when "01101011011001011", -- t[54987] = 19
      "0010011" when "01101011011001100", -- t[54988] = 19
      "0010011" when "01101011011001101", -- t[54989] = 19
      "0010011" when "01101011011001110", -- t[54990] = 19
      "0010011" when "01101011011001111", -- t[54991] = 19
      "0010011" when "01101011011010000", -- t[54992] = 19
      "0010011" when "01101011011010001", -- t[54993] = 19
      "0010011" when "01101011011010010", -- t[54994] = 19
      "0010011" when "01101011011010011", -- t[54995] = 19
      "0010011" when "01101011011010100", -- t[54996] = 19
      "0010011" when "01101011011010101", -- t[54997] = 19
      "0010011" when "01101011011010110", -- t[54998] = 19
      "0010011" when "01101011011010111", -- t[54999] = 19
      "0010011" when "01101011011011000", -- t[55000] = 19
      "0010011" when "01101011011011001", -- t[55001] = 19
      "0010011" when "01101011011011010", -- t[55002] = 19
      "0010011" when "01101011011011011", -- t[55003] = 19
      "0010011" when "01101011011011100", -- t[55004] = 19
      "0010011" when "01101011011011101", -- t[55005] = 19
      "0010011" when "01101011011011110", -- t[55006] = 19
      "0010011" when "01101011011011111", -- t[55007] = 19
      "0010011" when "01101011011100000", -- t[55008] = 19
      "0010011" when "01101011011100001", -- t[55009] = 19
      "0010011" when "01101011011100010", -- t[55010] = 19
      "0010011" when "01101011011100011", -- t[55011] = 19
      "0010011" when "01101011011100100", -- t[55012] = 19
      "0010011" when "01101011011100101", -- t[55013] = 19
      "0010011" when "01101011011100110", -- t[55014] = 19
      "0010011" when "01101011011100111", -- t[55015] = 19
      "0010011" when "01101011011101000", -- t[55016] = 19
      "0010011" when "01101011011101001", -- t[55017] = 19
      "0010011" when "01101011011101010", -- t[55018] = 19
      "0010011" when "01101011011101011", -- t[55019] = 19
      "0010011" when "01101011011101100", -- t[55020] = 19
      "0010011" when "01101011011101101", -- t[55021] = 19
      "0010011" when "01101011011101110", -- t[55022] = 19
      "0010011" when "01101011011101111", -- t[55023] = 19
      "0010011" when "01101011011110000", -- t[55024] = 19
      "0010011" when "01101011011110001", -- t[55025] = 19
      "0010011" when "01101011011110010", -- t[55026] = 19
      "0010011" when "01101011011110011", -- t[55027] = 19
      "0010011" when "01101011011110100", -- t[55028] = 19
      "0010011" when "01101011011110101", -- t[55029] = 19
      "0010011" when "01101011011110110", -- t[55030] = 19
      "0010011" when "01101011011110111", -- t[55031] = 19
      "0010011" when "01101011011111000", -- t[55032] = 19
      "0010011" when "01101011011111001", -- t[55033] = 19
      "0010011" when "01101011011111010", -- t[55034] = 19
      "0010011" when "01101011011111011", -- t[55035] = 19
      "0010011" when "01101011011111100", -- t[55036] = 19
      "0010011" when "01101011011111101", -- t[55037] = 19
      "0010011" when "01101011011111110", -- t[55038] = 19
      "0010011" when "01101011011111111", -- t[55039] = 19
      "0010011" when "01101011100000000", -- t[55040] = 19
      "0010011" when "01101011100000001", -- t[55041] = 19
      "0010011" when "01101011100000010", -- t[55042] = 19
      "0010011" when "01101011100000011", -- t[55043] = 19
      "0010011" when "01101011100000100", -- t[55044] = 19
      "0010011" when "01101011100000101", -- t[55045] = 19
      "0010011" when "01101011100000110", -- t[55046] = 19
      "0010011" when "01101011100000111", -- t[55047] = 19
      "0010011" when "01101011100001000", -- t[55048] = 19
      "0010011" when "01101011100001001", -- t[55049] = 19
      "0010011" when "01101011100001010", -- t[55050] = 19
      "0010011" when "01101011100001011", -- t[55051] = 19
      "0010011" when "01101011100001100", -- t[55052] = 19
      "0010011" when "01101011100001101", -- t[55053] = 19
      "0010011" when "01101011100001110", -- t[55054] = 19
      "0010011" when "01101011100001111", -- t[55055] = 19
      "0010011" when "01101011100010000", -- t[55056] = 19
      "0010011" when "01101011100010001", -- t[55057] = 19
      "0010011" when "01101011100010010", -- t[55058] = 19
      "0010011" when "01101011100010011", -- t[55059] = 19
      "0010011" when "01101011100010100", -- t[55060] = 19
      "0010011" when "01101011100010101", -- t[55061] = 19
      "0010011" when "01101011100010110", -- t[55062] = 19
      "0010011" when "01101011100010111", -- t[55063] = 19
      "0010011" when "01101011100011000", -- t[55064] = 19
      "0010011" when "01101011100011001", -- t[55065] = 19
      "0010011" when "01101011100011010", -- t[55066] = 19
      "0010011" when "01101011100011011", -- t[55067] = 19
      "0010011" when "01101011100011100", -- t[55068] = 19
      "0010011" when "01101011100011101", -- t[55069] = 19
      "0010011" when "01101011100011110", -- t[55070] = 19
      "0010011" when "01101011100011111", -- t[55071] = 19
      "0010011" when "01101011100100000", -- t[55072] = 19
      "0010011" when "01101011100100001", -- t[55073] = 19
      "0010011" when "01101011100100010", -- t[55074] = 19
      "0010011" when "01101011100100011", -- t[55075] = 19
      "0010011" when "01101011100100100", -- t[55076] = 19
      "0010011" when "01101011100100101", -- t[55077] = 19
      "0010011" when "01101011100100110", -- t[55078] = 19
      "0010011" when "01101011100100111", -- t[55079] = 19
      "0010011" when "01101011100101000", -- t[55080] = 19
      "0010011" when "01101011100101001", -- t[55081] = 19
      "0010011" when "01101011100101010", -- t[55082] = 19
      "0010011" when "01101011100101011", -- t[55083] = 19
      "0010011" when "01101011100101100", -- t[55084] = 19
      "0010011" when "01101011100101101", -- t[55085] = 19
      "0010011" when "01101011100101110", -- t[55086] = 19
      "0010011" when "01101011100101111", -- t[55087] = 19
      "0010011" when "01101011100110000", -- t[55088] = 19
      "0010011" when "01101011100110001", -- t[55089] = 19
      "0010011" when "01101011100110010", -- t[55090] = 19
      "0010011" when "01101011100110011", -- t[55091] = 19
      "0010011" when "01101011100110100", -- t[55092] = 19
      "0010011" when "01101011100110101", -- t[55093] = 19
      "0010011" when "01101011100110110", -- t[55094] = 19
      "0010011" when "01101011100110111", -- t[55095] = 19
      "0010011" when "01101011100111000", -- t[55096] = 19
      "0010011" when "01101011100111001", -- t[55097] = 19
      "0010011" when "01101011100111010", -- t[55098] = 19
      "0010011" when "01101011100111011", -- t[55099] = 19
      "0010011" when "01101011100111100", -- t[55100] = 19
      "0010011" when "01101011100111101", -- t[55101] = 19
      "0010011" when "01101011100111110", -- t[55102] = 19
      "0010011" when "01101011100111111", -- t[55103] = 19
      "0010011" when "01101011101000000", -- t[55104] = 19
      "0010011" when "01101011101000001", -- t[55105] = 19
      "0010011" when "01101011101000010", -- t[55106] = 19
      "0010011" when "01101011101000011", -- t[55107] = 19
      "0010011" when "01101011101000100", -- t[55108] = 19
      "0010011" when "01101011101000101", -- t[55109] = 19
      "0010011" when "01101011101000110", -- t[55110] = 19
      "0010011" when "01101011101000111", -- t[55111] = 19
      "0010011" when "01101011101001000", -- t[55112] = 19
      "0010011" when "01101011101001001", -- t[55113] = 19
      "0010011" when "01101011101001010", -- t[55114] = 19
      "0010011" when "01101011101001011", -- t[55115] = 19
      "0010011" when "01101011101001100", -- t[55116] = 19
      "0010011" when "01101011101001101", -- t[55117] = 19
      "0010011" when "01101011101001110", -- t[55118] = 19
      "0010011" when "01101011101001111", -- t[55119] = 19
      "0010011" when "01101011101010000", -- t[55120] = 19
      "0010011" when "01101011101010001", -- t[55121] = 19
      "0010011" when "01101011101010010", -- t[55122] = 19
      "0010011" when "01101011101010011", -- t[55123] = 19
      "0010011" when "01101011101010100", -- t[55124] = 19
      "0010011" when "01101011101010101", -- t[55125] = 19
      "0010011" when "01101011101010110", -- t[55126] = 19
      "0010011" when "01101011101010111", -- t[55127] = 19
      "0010011" when "01101011101011000", -- t[55128] = 19
      "0010011" when "01101011101011001", -- t[55129] = 19
      "0010011" when "01101011101011010", -- t[55130] = 19
      "0010011" when "01101011101011011", -- t[55131] = 19
      "0010011" when "01101011101011100", -- t[55132] = 19
      "0010011" when "01101011101011101", -- t[55133] = 19
      "0010011" when "01101011101011110", -- t[55134] = 19
      "0010011" when "01101011101011111", -- t[55135] = 19
      "0010011" when "01101011101100000", -- t[55136] = 19
      "0010011" when "01101011101100001", -- t[55137] = 19
      "0010011" when "01101011101100010", -- t[55138] = 19
      "0010011" when "01101011101100011", -- t[55139] = 19
      "0010011" when "01101011101100100", -- t[55140] = 19
      "0010011" when "01101011101100101", -- t[55141] = 19
      "0010011" when "01101011101100110", -- t[55142] = 19
      "0010011" when "01101011101100111", -- t[55143] = 19
      "0010011" when "01101011101101000", -- t[55144] = 19
      "0010011" when "01101011101101001", -- t[55145] = 19
      "0010011" when "01101011101101010", -- t[55146] = 19
      "0010011" when "01101011101101011", -- t[55147] = 19
      "0010011" when "01101011101101100", -- t[55148] = 19
      "0010011" when "01101011101101101", -- t[55149] = 19
      "0010011" when "01101011101101110", -- t[55150] = 19
      "0010011" when "01101011101101111", -- t[55151] = 19
      "0010011" when "01101011101110000", -- t[55152] = 19
      "0010011" when "01101011101110001", -- t[55153] = 19
      "0010011" when "01101011101110010", -- t[55154] = 19
      "0010011" when "01101011101110011", -- t[55155] = 19
      "0010011" when "01101011101110100", -- t[55156] = 19
      "0010011" when "01101011101110101", -- t[55157] = 19
      "0010011" when "01101011101110110", -- t[55158] = 19
      "0010011" when "01101011101110111", -- t[55159] = 19
      "0010011" when "01101011101111000", -- t[55160] = 19
      "0010011" when "01101011101111001", -- t[55161] = 19
      "0010011" when "01101011101111010", -- t[55162] = 19
      "0010011" when "01101011101111011", -- t[55163] = 19
      "0010011" when "01101011101111100", -- t[55164] = 19
      "0010011" when "01101011101111101", -- t[55165] = 19
      "0010011" when "01101011101111110", -- t[55166] = 19
      "0010011" when "01101011101111111", -- t[55167] = 19
      "0010011" when "01101011110000000", -- t[55168] = 19
      "0010011" when "01101011110000001", -- t[55169] = 19
      "0010011" when "01101011110000010", -- t[55170] = 19
      "0010011" when "01101011110000011", -- t[55171] = 19
      "0010011" when "01101011110000100", -- t[55172] = 19
      "0010011" when "01101011110000101", -- t[55173] = 19
      "0010011" when "01101011110000110", -- t[55174] = 19
      "0010011" when "01101011110000111", -- t[55175] = 19
      "0010011" when "01101011110001000", -- t[55176] = 19
      "0010011" when "01101011110001001", -- t[55177] = 19
      "0010011" when "01101011110001010", -- t[55178] = 19
      "0010011" when "01101011110001011", -- t[55179] = 19
      "0010011" when "01101011110001100", -- t[55180] = 19
      "0010011" when "01101011110001101", -- t[55181] = 19
      "0010011" when "01101011110001110", -- t[55182] = 19
      "0010011" when "01101011110001111", -- t[55183] = 19
      "0010011" when "01101011110010000", -- t[55184] = 19
      "0010011" when "01101011110010001", -- t[55185] = 19
      "0010011" when "01101011110010010", -- t[55186] = 19
      "0010011" when "01101011110010011", -- t[55187] = 19
      "0010011" when "01101011110010100", -- t[55188] = 19
      "0010011" when "01101011110010101", -- t[55189] = 19
      "0010011" when "01101011110010110", -- t[55190] = 19
      "0010011" when "01101011110010111", -- t[55191] = 19
      "0010011" when "01101011110011000", -- t[55192] = 19
      "0010011" when "01101011110011001", -- t[55193] = 19
      "0010011" when "01101011110011010", -- t[55194] = 19
      "0010011" when "01101011110011011", -- t[55195] = 19
      "0010011" when "01101011110011100", -- t[55196] = 19
      "0010011" when "01101011110011101", -- t[55197] = 19
      "0010011" when "01101011110011110", -- t[55198] = 19
      "0010011" when "01101011110011111", -- t[55199] = 19
      "0010011" when "01101011110100000", -- t[55200] = 19
      "0010011" when "01101011110100001", -- t[55201] = 19
      "0010011" when "01101011110100010", -- t[55202] = 19
      "0010011" when "01101011110100011", -- t[55203] = 19
      "0010011" when "01101011110100100", -- t[55204] = 19
      "0010011" when "01101011110100101", -- t[55205] = 19
      "0010011" when "01101011110100110", -- t[55206] = 19
      "0010011" when "01101011110100111", -- t[55207] = 19
      "0010011" when "01101011110101000", -- t[55208] = 19
      "0010011" when "01101011110101001", -- t[55209] = 19
      "0010011" when "01101011110101010", -- t[55210] = 19
      "0010011" when "01101011110101011", -- t[55211] = 19
      "0010011" when "01101011110101100", -- t[55212] = 19
      "0010011" when "01101011110101101", -- t[55213] = 19
      "0010011" when "01101011110101110", -- t[55214] = 19
      "0010011" when "01101011110101111", -- t[55215] = 19
      "0010011" when "01101011110110000", -- t[55216] = 19
      "0010011" when "01101011110110001", -- t[55217] = 19
      "0010011" when "01101011110110010", -- t[55218] = 19
      "0010011" when "01101011110110011", -- t[55219] = 19
      "0010011" when "01101011110110100", -- t[55220] = 19
      "0010011" when "01101011110110101", -- t[55221] = 19
      "0010011" when "01101011110110110", -- t[55222] = 19
      "0010011" when "01101011110110111", -- t[55223] = 19
      "0010011" when "01101011110111000", -- t[55224] = 19
      "0010011" when "01101011110111001", -- t[55225] = 19
      "0010011" when "01101011110111010", -- t[55226] = 19
      "0010011" when "01101011110111011", -- t[55227] = 19
      "0010011" when "01101011110111100", -- t[55228] = 19
      "0010011" when "01101011110111101", -- t[55229] = 19
      "0010011" when "01101011110111110", -- t[55230] = 19
      "0010011" when "01101011110111111", -- t[55231] = 19
      "0010011" when "01101011111000000", -- t[55232] = 19
      "0010011" when "01101011111000001", -- t[55233] = 19
      "0010011" when "01101011111000010", -- t[55234] = 19
      "0010011" when "01101011111000011", -- t[55235] = 19
      "0010011" when "01101011111000100", -- t[55236] = 19
      "0010011" when "01101011111000101", -- t[55237] = 19
      "0010011" when "01101011111000110", -- t[55238] = 19
      "0010011" when "01101011111000111", -- t[55239] = 19
      "0010011" when "01101011111001000", -- t[55240] = 19
      "0010011" when "01101011111001001", -- t[55241] = 19
      "0010011" when "01101011111001010", -- t[55242] = 19
      "0010011" when "01101011111001011", -- t[55243] = 19
      "0010011" when "01101011111001100", -- t[55244] = 19
      "0010011" when "01101011111001101", -- t[55245] = 19
      "0010011" when "01101011111001110", -- t[55246] = 19
      "0010011" when "01101011111001111", -- t[55247] = 19
      "0010011" when "01101011111010000", -- t[55248] = 19
      "0010011" when "01101011111010001", -- t[55249] = 19
      "0010011" when "01101011111010010", -- t[55250] = 19
      "0010011" when "01101011111010011", -- t[55251] = 19
      "0010011" when "01101011111010100", -- t[55252] = 19
      "0010011" when "01101011111010101", -- t[55253] = 19
      "0010011" when "01101011111010110", -- t[55254] = 19
      "0010011" when "01101011111010111", -- t[55255] = 19
      "0010011" when "01101011111011000", -- t[55256] = 19
      "0010011" when "01101011111011001", -- t[55257] = 19
      "0010011" when "01101011111011010", -- t[55258] = 19
      "0010011" when "01101011111011011", -- t[55259] = 19
      "0010011" when "01101011111011100", -- t[55260] = 19
      "0010011" when "01101011111011101", -- t[55261] = 19
      "0010011" when "01101011111011110", -- t[55262] = 19
      "0010011" when "01101011111011111", -- t[55263] = 19
      "0010011" when "01101011111100000", -- t[55264] = 19
      "0010011" when "01101011111100001", -- t[55265] = 19
      "0010011" when "01101011111100010", -- t[55266] = 19
      "0010011" when "01101011111100011", -- t[55267] = 19
      "0010011" when "01101011111100100", -- t[55268] = 19
      "0010011" when "01101011111100101", -- t[55269] = 19
      "0010011" when "01101011111100110", -- t[55270] = 19
      "0010011" when "01101011111100111", -- t[55271] = 19
      "0010011" when "01101011111101000", -- t[55272] = 19
      "0010011" when "01101011111101001", -- t[55273] = 19
      "0010011" when "01101011111101010", -- t[55274] = 19
      "0010011" when "01101011111101011", -- t[55275] = 19
      "0010011" when "01101011111101100", -- t[55276] = 19
      "0010011" when "01101011111101101", -- t[55277] = 19
      "0010011" when "01101011111101110", -- t[55278] = 19
      "0010011" when "01101011111101111", -- t[55279] = 19
      "0010011" when "01101011111110000", -- t[55280] = 19
      "0010011" when "01101011111110001", -- t[55281] = 19
      "0010011" when "01101011111110010", -- t[55282] = 19
      "0010011" when "01101011111110011", -- t[55283] = 19
      "0010011" when "01101011111110100", -- t[55284] = 19
      "0010011" when "01101011111110101", -- t[55285] = 19
      "0010011" when "01101011111110110", -- t[55286] = 19
      "0010011" when "01101011111110111", -- t[55287] = 19
      "0010011" when "01101011111111000", -- t[55288] = 19
      "0010011" when "01101011111111001", -- t[55289] = 19
      "0010011" when "01101011111111010", -- t[55290] = 19
      "0010011" when "01101011111111011", -- t[55291] = 19
      "0010011" when "01101011111111100", -- t[55292] = 19
      "0010011" when "01101011111111101", -- t[55293] = 19
      "0010011" when "01101011111111110", -- t[55294] = 19
      "0010011" when "01101011111111111", -- t[55295] = 19
      "0010011" when "01101100000000000", -- t[55296] = 19
      "0010011" when "01101100000000001", -- t[55297] = 19
      "0010011" when "01101100000000010", -- t[55298] = 19
      "0010011" when "01101100000000011", -- t[55299] = 19
      "0010011" when "01101100000000100", -- t[55300] = 19
      "0010011" when "01101100000000101", -- t[55301] = 19
      "0010011" when "01101100000000110", -- t[55302] = 19
      "0010011" when "01101100000000111", -- t[55303] = 19
      "0010011" when "01101100000001000", -- t[55304] = 19
      "0010011" when "01101100000001001", -- t[55305] = 19
      "0010011" when "01101100000001010", -- t[55306] = 19
      "0010011" when "01101100000001011", -- t[55307] = 19
      "0010011" when "01101100000001100", -- t[55308] = 19
      "0010011" when "01101100000001101", -- t[55309] = 19
      "0010011" when "01101100000001110", -- t[55310] = 19
      "0010011" when "01101100000001111", -- t[55311] = 19
      "0010011" when "01101100000010000", -- t[55312] = 19
      "0010011" when "01101100000010001", -- t[55313] = 19
      "0010011" when "01101100000010010", -- t[55314] = 19
      "0010011" when "01101100000010011", -- t[55315] = 19
      "0010011" when "01101100000010100", -- t[55316] = 19
      "0010011" when "01101100000010101", -- t[55317] = 19
      "0010011" when "01101100000010110", -- t[55318] = 19
      "0010011" when "01101100000010111", -- t[55319] = 19
      "0010011" when "01101100000011000", -- t[55320] = 19
      "0010011" when "01101100000011001", -- t[55321] = 19
      "0010011" when "01101100000011010", -- t[55322] = 19
      "0010011" when "01101100000011011", -- t[55323] = 19
      "0010011" when "01101100000011100", -- t[55324] = 19
      "0010011" when "01101100000011101", -- t[55325] = 19
      "0010011" when "01101100000011110", -- t[55326] = 19
      "0010011" when "01101100000011111", -- t[55327] = 19
      "0010011" when "01101100000100000", -- t[55328] = 19
      "0010011" when "01101100000100001", -- t[55329] = 19
      "0010011" when "01101100000100010", -- t[55330] = 19
      "0010011" when "01101100000100011", -- t[55331] = 19
      "0010011" when "01101100000100100", -- t[55332] = 19
      "0010011" when "01101100000100101", -- t[55333] = 19
      "0010011" when "01101100000100110", -- t[55334] = 19
      "0010011" when "01101100000100111", -- t[55335] = 19
      "0010011" when "01101100000101000", -- t[55336] = 19
      "0010011" when "01101100000101001", -- t[55337] = 19
      "0010011" when "01101100000101010", -- t[55338] = 19
      "0010011" when "01101100000101011", -- t[55339] = 19
      "0010011" when "01101100000101100", -- t[55340] = 19
      "0010100" when "01101100000101101", -- t[55341] = 20
      "0010100" when "01101100000101110", -- t[55342] = 20
      "0010100" when "01101100000101111", -- t[55343] = 20
      "0010100" when "01101100000110000", -- t[55344] = 20
      "0010100" when "01101100000110001", -- t[55345] = 20
      "0010100" when "01101100000110010", -- t[55346] = 20
      "0010100" when "01101100000110011", -- t[55347] = 20
      "0010100" when "01101100000110100", -- t[55348] = 20
      "0010100" when "01101100000110101", -- t[55349] = 20
      "0010100" when "01101100000110110", -- t[55350] = 20
      "0010100" when "01101100000110111", -- t[55351] = 20
      "0010100" when "01101100000111000", -- t[55352] = 20
      "0010100" when "01101100000111001", -- t[55353] = 20
      "0010100" when "01101100000111010", -- t[55354] = 20
      "0010100" when "01101100000111011", -- t[55355] = 20
      "0010100" when "01101100000111100", -- t[55356] = 20
      "0010100" when "01101100000111101", -- t[55357] = 20
      "0010100" when "01101100000111110", -- t[55358] = 20
      "0010100" when "01101100000111111", -- t[55359] = 20
      "0010100" when "01101100001000000", -- t[55360] = 20
      "0010100" when "01101100001000001", -- t[55361] = 20
      "0010100" when "01101100001000010", -- t[55362] = 20
      "0010100" when "01101100001000011", -- t[55363] = 20
      "0010100" when "01101100001000100", -- t[55364] = 20
      "0010100" when "01101100001000101", -- t[55365] = 20
      "0010100" when "01101100001000110", -- t[55366] = 20
      "0010100" when "01101100001000111", -- t[55367] = 20
      "0010100" when "01101100001001000", -- t[55368] = 20
      "0010100" when "01101100001001001", -- t[55369] = 20
      "0010100" when "01101100001001010", -- t[55370] = 20
      "0010100" when "01101100001001011", -- t[55371] = 20
      "0010100" when "01101100001001100", -- t[55372] = 20
      "0010100" when "01101100001001101", -- t[55373] = 20
      "0010100" when "01101100001001110", -- t[55374] = 20
      "0010100" when "01101100001001111", -- t[55375] = 20
      "0010100" when "01101100001010000", -- t[55376] = 20
      "0010100" when "01101100001010001", -- t[55377] = 20
      "0010100" when "01101100001010010", -- t[55378] = 20
      "0010100" when "01101100001010011", -- t[55379] = 20
      "0010100" when "01101100001010100", -- t[55380] = 20
      "0010100" when "01101100001010101", -- t[55381] = 20
      "0010100" when "01101100001010110", -- t[55382] = 20
      "0010100" when "01101100001010111", -- t[55383] = 20
      "0010100" when "01101100001011000", -- t[55384] = 20
      "0010100" when "01101100001011001", -- t[55385] = 20
      "0010100" when "01101100001011010", -- t[55386] = 20
      "0010100" when "01101100001011011", -- t[55387] = 20
      "0010100" when "01101100001011100", -- t[55388] = 20
      "0010100" when "01101100001011101", -- t[55389] = 20
      "0010100" when "01101100001011110", -- t[55390] = 20
      "0010100" when "01101100001011111", -- t[55391] = 20
      "0010100" when "01101100001100000", -- t[55392] = 20
      "0010100" when "01101100001100001", -- t[55393] = 20
      "0010100" when "01101100001100010", -- t[55394] = 20
      "0010100" when "01101100001100011", -- t[55395] = 20
      "0010100" when "01101100001100100", -- t[55396] = 20
      "0010100" when "01101100001100101", -- t[55397] = 20
      "0010100" when "01101100001100110", -- t[55398] = 20
      "0010100" when "01101100001100111", -- t[55399] = 20
      "0010100" when "01101100001101000", -- t[55400] = 20
      "0010100" when "01101100001101001", -- t[55401] = 20
      "0010100" when "01101100001101010", -- t[55402] = 20
      "0010100" when "01101100001101011", -- t[55403] = 20
      "0010100" when "01101100001101100", -- t[55404] = 20
      "0010100" when "01101100001101101", -- t[55405] = 20
      "0010100" when "01101100001101110", -- t[55406] = 20
      "0010100" when "01101100001101111", -- t[55407] = 20
      "0010100" when "01101100001110000", -- t[55408] = 20
      "0010100" when "01101100001110001", -- t[55409] = 20
      "0010100" when "01101100001110010", -- t[55410] = 20
      "0010100" when "01101100001110011", -- t[55411] = 20
      "0010100" when "01101100001110100", -- t[55412] = 20
      "0010100" when "01101100001110101", -- t[55413] = 20
      "0010100" when "01101100001110110", -- t[55414] = 20
      "0010100" when "01101100001110111", -- t[55415] = 20
      "0010100" when "01101100001111000", -- t[55416] = 20
      "0010100" when "01101100001111001", -- t[55417] = 20
      "0010100" when "01101100001111010", -- t[55418] = 20
      "0010100" when "01101100001111011", -- t[55419] = 20
      "0010100" when "01101100001111100", -- t[55420] = 20
      "0010100" when "01101100001111101", -- t[55421] = 20
      "0010100" when "01101100001111110", -- t[55422] = 20
      "0010100" when "01101100001111111", -- t[55423] = 20
      "0010100" when "01101100010000000", -- t[55424] = 20
      "0010100" when "01101100010000001", -- t[55425] = 20
      "0010100" when "01101100010000010", -- t[55426] = 20
      "0010100" when "01101100010000011", -- t[55427] = 20
      "0010100" when "01101100010000100", -- t[55428] = 20
      "0010100" when "01101100010000101", -- t[55429] = 20
      "0010100" when "01101100010000110", -- t[55430] = 20
      "0010100" when "01101100010000111", -- t[55431] = 20
      "0010100" when "01101100010001000", -- t[55432] = 20
      "0010100" when "01101100010001001", -- t[55433] = 20
      "0010100" when "01101100010001010", -- t[55434] = 20
      "0010100" when "01101100010001011", -- t[55435] = 20
      "0010100" when "01101100010001100", -- t[55436] = 20
      "0010100" when "01101100010001101", -- t[55437] = 20
      "0010100" when "01101100010001110", -- t[55438] = 20
      "0010100" when "01101100010001111", -- t[55439] = 20
      "0010100" when "01101100010010000", -- t[55440] = 20
      "0010100" when "01101100010010001", -- t[55441] = 20
      "0010100" when "01101100010010010", -- t[55442] = 20
      "0010100" when "01101100010010011", -- t[55443] = 20
      "0010100" when "01101100010010100", -- t[55444] = 20
      "0010100" when "01101100010010101", -- t[55445] = 20
      "0010100" when "01101100010010110", -- t[55446] = 20
      "0010100" when "01101100010010111", -- t[55447] = 20
      "0010100" when "01101100010011000", -- t[55448] = 20
      "0010100" when "01101100010011001", -- t[55449] = 20
      "0010100" when "01101100010011010", -- t[55450] = 20
      "0010100" when "01101100010011011", -- t[55451] = 20
      "0010100" when "01101100010011100", -- t[55452] = 20
      "0010100" when "01101100010011101", -- t[55453] = 20
      "0010100" when "01101100010011110", -- t[55454] = 20
      "0010100" when "01101100010011111", -- t[55455] = 20
      "0010100" when "01101100010100000", -- t[55456] = 20
      "0010100" when "01101100010100001", -- t[55457] = 20
      "0010100" when "01101100010100010", -- t[55458] = 20
      "0010100" when "01101100010100011", -- t[55459] = 20
      "0010100" when "01101100010100100", -- t[55460] = 20
      "0010100" when "01101100010100101", -- t[55461] = 20
      "0010100" when "01101100010100110", -- t[55462] = 20
      "0010100" when "01101100010100111", -- t[55463] = 20
      "0010100" when "01101100010101000", -- t[55464] = 20
      "0010100" when "01101100010101001", -- t[55465] = 20
      "0010100" when "01101100010101010", -- t[55466] = 20
      "0010100" when "01101100010101011", -- t[55467] = 20
      "0010100" when "01101100010101100", -- t[55468] = 20
      "0010100" when "01101100010101101", -- t[55469] = 20
      "0010100" when "01101100010101110", -- t[55470] = 20
      "0010100" when "01101100010101111", -- t[55471] = 20
      "0010100" when "01101100010110000", -- t[55472] = 20
      "0010100" when "01101100010110001", -- t[55473] = 20
      "0010100" when "01101100010110010", -- t[55474] = 20
      "0010100" when "01101100010110011", -- t[55475] = 20
      "0010100" when "01101100010110100", -- t[55476] = 20
      "0010100" when "01101100010110101", -- t[55477] = 20
      "0010100" when "01101100010110110", -- t[55478] = 20
      "0010100" when "01101100010110111", -- t[55479] = 20
      "0010100" when "01101100010111000", -- t[55480] = 20
      "0010100" when "01101100010111001", -- t[55481] = 20
      "0010100" when "01101100010111010", -- t[55482] = 20
      "0010100" when "01101100010111011", -- t[55483] = 20
      "0010100" when "01101100010111100", -- t[55484] = 20
      "0010100" when "01101100010111101", -- t[55485] = 20
      "0010100" when "01101100010111110", -- t[55486] = 20
      "0010100" when "01101100010111111", -- t[55487] = 20
      "0010100" when "01101100011000000", -- t[55488] = 20
      "0010100" when "01101100011000001", -- t[55489] = 20
      "0010100" when "01101100011000010", -- t[55490] = 20
      "0010100" when "01101100011000011", -- t[55491] = 20
      "0010100" when "01101100011000100", -- t[55492] = 20
      "0010100" when "01101100011000101", -- t[55493] = 20
      "0010100" when "01101100011000110", -- t[55494] = 20
      "0010100" when "01101100011000111", -- t[55495] = 20
      "0010100" when "01101100011001000", -- t[55496] = 20
      "0010100" when "01101100011001001", -- t[55497] = 20
      "0010100" when "01101100011001010", -- t[55498] = 20
      "0010100" when "01101100011001011", -- t[55499] = 20
      "0010100" when "01101100011001100", -- t[55500] = 20
      "0010100" when "01101100011001101", -- t[55501] = 20
      "0010100" when "01101100011001110", -- t[55502] = 20
      "0010100" when "01101100011001111", -- t[55503] = 20
      "0010100" when "01101100011010000", -- t[55504] = 20
      "0010100" when "01101100011010001", -- t[55505] = 20
      "0010100" when "01101100011010010", -- t[55506] = 20
      "0010100" when "01101100011010011", -- t[55507] = 20
      "0010100" when "01101100011010100", -- t[55508] = 20
      "0010100" when "01101100011010101", -- t[55509] = 20
      "0010100" when "01101100011010110", -- t[55510] = 20
      "0010100" when "01101100011010111", -- t[55511] = 20
      "0010100" when "01101100011011000", -- t[55512] = 20
      "0010100" when "01101100011011001", -- t[55513] = 20
      "0010100" when "01101100011011010", -- t[55514] = 20
      "0010100" when "01101100011011011", -- t[55515] = 20
      "0010100" when "01101100011011100", -- t[55516] = 20
      "0010100" when "01101100011011101", -- t[55517] = 20
      "0010100" when "01101100011011110", -- t[55518] = 20
      "0010100" when "01101100011011111", -- t[55519] = 20
      "0010100" when "01101100011100000", -- t[55520] = 20
      "0010100" when "01101100011100001", -- t[55521] = 20
      "0010100" when "01101100011100010", -- t[55522] = 20
      "0010100" when "01101100011100011", -- t[55523] = 20
      "0010100" when "01101100011100100", -- t[55524] = 20
      "0010100" when "01101100011100101", -- t[55525] = 20
      "0010100" when "01101100011100110", -- t[55526] = 20
      "0010100" when "01101100011100111", -- t[55527] = 20
      "0010100" when "01101100011101000", -- t[55528] = 20
      "0010100" when "01101100011101001", -- t[55529] = 20
      "0010100" when "01101100011101010", -- t[55530] = 20
      "0010100" when "01101100011101011", -- t[55531] = 20
      "0010100" when "01101100011101100", -- t[55532] = 20
      "0010100" when "01101100011101101", -- t[55533] = 20
      "0010100" when "01101100011101110", -- t[55534] = 20
      "0010100" when "01101100011101111", -- t[55535] = 20
      "0010100" when "01101100011110000", -- t[55536] = 20
      "0010100" when "01101100011110001", -- t[55537] = 20
      "0010100" when "01101100011110010", -- t[55538] = 20
      "0010100" when "01101100011110011", -- t[55539] = 20
      "0010100" when "01101100011110100", -- t[55540] = 20
      "0010100" when "01101100011110101", -- t[55541] = 20
      "0010100" when "01101100011110110", -- t[55542] = 20
      "0010100" when "01101100011110111", -- t[55543] = 20
      "0010100" when "01101100011111000", -- t[55544] = 20
      "0010100" when "01101100011111001", -- t[55545] = 20
      "0010100" when "01101100011111010", -- t[55546] = 20
      "0010100" when "01101100011111011", -- t[55547] = 20
      "0010100" when "01101100011111100", -- t[55548] = 20
      "0010100" when "01101100011111101", -- t[55549] = 20
      "0010100" when "01101100011111110", -- t[55550] = 20
      "0010100" when "01101100011111111", -- t[55551] = 20
      "0010100" when "01101100100000000", -- t[55552] = 20
      "0010100" when "01101100100000001", -- t[55553] = 20
      "0010100" when "01101100100000010", -- t[55554] = 20
      "0010100" when "01101100100000011", -- t[55555] = 20
      "0010100" when "01101100100000100", -- t[55556] = 20
      "0010100" when "01101100100000101", -- t[55557] = 20
      "0010100" when "01101100100000110", -- t[55558] = 20
      "0010100" when "01101100100000111", -- t[55559] = 20
      "0010100" when "01101100100001000", -- t[55560] = 20
      "0010100" when "01101100100001001", -- t[55561] = 20
      "0010100" when "01101100100001010", -- t[55562] = 20
      "0010100" when "01101100100001011", -- t[55563] = 20
      "0010100" when "01101100100001100", -- t[55564] = 20
      "0010100" when "01101100100001101", -- t[55565] = 20
      "0010100" when "01101100100001110", -- t[55566] = 20
      "0010100" when "01101100100001111", -- t[55567] = 20
      "0010100" when "01101100100010000", -- t[55568] = 20
      "0010100" when "01101100100010001", -- t[55569] = 20
      "0010100" when "01101100100010010", -- t[55570] = 20
      "0010100" when "01101100100010011", -- t[55571] = 20
      "0010100" when "01101100100010100", -- t[55572] = 20
      "0010100" when "01101100100010101", -- t[55573] = 20
      "0010100" when "01101100100010110", -- t[55574] = 20
      "0010100" when "01101100100010111", -- t[55575] = 20
      "0010100" when "01101100100011000", -- t[55576] = 20
      "0010100" when "01101100100011001", -- t[55577] = 20
      "0010100" when "01101100100011010", -- t[55578] = 20
      "0010100" when "01101100100011011", -- t[55579] = 20
      "0010100" when "01101100100011100", -- t[55580] = 20
      "0010100" when "01101100100011101", -- t[55581] = 20
      "0010100" when "01101100100011110", -- t[55582] = 20
      "0010100" when "01101100100011111", -- t[55583] = 20
      "0010100" when "01101100100100000", -- t[55584] = 20
      "0010100" when "01101100100100001", -- t[55585] = 20
      "0010100" when "01101100100100010", -- t[55586] = 20
      "0010100" when "01101100100100011", -- t[55587] = 20
      "0010100" when "01101100100100100", -- t[55588] = 20
      "0010100" when "01101100100100101", -- t[55589] = 20
      "0010100" when "01101100100100110", -- t[55590] = 20
      "0010100" when "01101100100100111", -- t[55591] = 20
      "0010100" when "01101100100101000", -- t[55592] = 20
      "0010100" when "01101100100101001", -- t[55593] = 20
      "0010100" when "01101100100101010", -- t[55594] = 20
      "0010100" when "01101100100101011", -- t[55595] = 20
      "0010100" when "01101100100101100", -- t[55596] = 20
      "0010100" when "01101100100101101", -- t[55597] = 20
      "0010100" when "01101100100101110", -- t[55598] = 20
      "0010100" when "01101100100101111", -- t[55599] = 20
      "0010100" when "01101100100110000", -- t[55600] = 20
      "0010100" when "01101100100110001", -- t[55601] = 20
      "0010100" when "01101100100110010", -- t[55602] = 20
      "0010100" when "01101100100110011", -- t[55603] = 20
      "0010100" when "01101100100110100", -- t[55604] = 20
      "0010100" when "01101100100110101", -- t[55605] = 20
      "0010100" when "01101100100110110", -- t[55606] = 20
      "0010100" when "01101100100110111", -- t[55607] = 20
      "0010100" when "01101100100111000", -- t[55608] = 20
      "0010100" when "01101100100111001", -- t[55609] = 20
      "0010100" when "01101100100111010", -- t[55610] = 20
      "0010100" when "01101100100111011", -- t[55611] = 20
      "0010100" when "01101100100111100", -- t[55612] = 20
      "0010100" when "01101100100111101", -- t[55613] = 20
      "0010100" when "01101100100111110", -- t[55614] = 20
      "0010100" when "01101100100111111", -- t[55615] = 20
      "0010100" when "01101100101000000", -- t[55616] = 20
      "0010100" when "01101100101000001", -- t[55617] = 20
      "0010100" when "01101100101000010", -- t[55618] = 20
      "0010100" when "01101100101000011", -- t[55619] = 20
      "0010100" when "01101100101000100", -- t[55620] = 20
      "0010100" when "01101100101000101", -- t[55621] = 20
      "0010100" when "01101100101000110", -- t[55622] = 20
      "0010100" when "01101100101000111", -- t[55623] = 20
      "0010100" when "01101100101001000", -- t[55624] = 20
      "0010100" when "01101100101001001", -- t[55625] = 20
      "0010100" when "01101100101001010", -- t[55626] = 20
      "0010100" when "01101100101001011", -- t[55627] = 20
      "0010100" when "01101100101001100", -- t[55628] = 20
      "0010100" when "01101100101001101", -- t[55629] = 20
      "0010100" when "01101100101001110", -- t[55630] = 20
      "0010100" when "01101100101001111", -- t[55631] = 20
      "0010100" when "01101100101010000", -- t[55632] = 20
      "0010100" when "01101100101010001", -- t[55633] = 20
      "0010100" when "01101100101010010", -- t[55634] = 20
      "0010100" when "01101100101010011", -- t[55635] = 20
      "0010100" when "01101100101010100", -- t[55636] = 20
      "0010100" when "01101100101010101", -- t[55637] = 20
      "0010100" when "01101100101010110", -- t[55638] = 20
      "0010100" when "01101100101010111", -- t[55639] = 20
      "0010100" when "01101100101011000", -- t[55640] = 20
      "0010100" when "01101100101011001", -- t[55641] = 20
      "0010100" when "01101100101011010", -- t[55642] = 20
      "0010100" when "01101100101011011", -- t[55643] = 20
      "0010100" when "01101100101011100", -- t[55644] = 20
      "0010100" when "01101100101011101", -- t[55645] = 20
      "0010100" when "01101100101011110", -- t[55646] = 20
      "0010100" when "01101100101011111", -- t[55647] = 20
      "0010100" when "01101100101100000", -- t[55648] = 20
      "0010100" when "01101100101100001", -- t[55649] = 20
      "0010100" when "01101100101100010", -- t[55650] = 20
      "0010100" when "01101100101100011", -- t[55651] = 20
      "0010100" when "01101100101100100", -- t[55652] = 20
      "0010100" when "01101100101100101", -- t[55653] = 20
      "0010100" when "01101100101100110", -- t[55654] = 20
      "0010100" when "01101100101100111", -- t[55655] = 20
      "0010100" when "01101100101101000", -- t[55656] = 20
      "0010100" when "01101100101101001", -- t[55657] = 20
      "0010100" when "01101100101101010", -- t[55658] = 20
      "0010100" when "01101100101101011", -- t[55659] = 20
      "0010100" when "01101100101101100", -- t[55660] = 20
      "0010100" when "01101100101101101", -- t[55661] = 20
      "0010100" when "01101100101101110", -- t[55662] = 20
      "0010100" when "01101100101101111", -- t[55663] = 20
      "0010100" when "01101100101110000", -- t[55664] = 20
      "0010100" when "01101100101110001", -- t[55665] = 20
      "0010100" when "01101100101110010", -- t[55666] = 20
      "0010100" when "01101100101110011", -- t[55667] = 20
      "0010100" when "01101100101110100", -- t[55668] = 20
      "0010100" when "01101100101110101", -- t[55669] = 20
      "0010100" when "01101100101110110", -- t[55670] = 20
      "0010100" when "01101100101110111", -- t[55671] = 20
      "0010100" when "01101100101111000", -- t[55672] = 20
      "0010100" when "01101100101111001", -- t[55673] = 20
      "0010100" when "01101100101111010", -- t[55674] = 20
      "0010100" when "01101100101111011", -- t[55675] = 20
      "0010100" when "01101100101111100", -- t[55676] = 20
      "0010100" when "01101100101111101", -- t[55677] = 20
      "0010100" when "01101100101111110", -- t[55678] = 20
      "0010100" when "01101100101111111", -- t[55679] = 20
      "0010100" when "01101100110000000", -- t[55680] = 20
      "0010100" when "01101100110000001", -- t[55681] = 20
      "0010100" when "01101100110000010", -- t[55682] = 20
      "0010100" when "01101100110000011", -- t[55683] = 20
      "0010100" when "01101100110000100", -- t[55684] = 20
      "0010100" when "01101100110000101", -- t[55685] = 20
      "0010100" when "01101100110000110", -- t[55686] = 20
      "0010100" when "01101100110000111", -- t[55687] = 20
      "0010100" when "01101100110001000", -- t[55688] = 20
      "0010100" when "01101100110001001", -- t[55689] = 20
      "0010100" when "01101100110001010", -- t[55690] = 20
      "0010100" when "01101100110001011", -- t[55691] = 20
      "0010100" when "01101100110001100", -- t[55692] = 20
      "0010100" when "01101100110001101", -- t[55693] = 20
      "0010100" when "01101100110001110", -- t[55694] = 20
      "0010100" when "01101100110001111", -- t[55695] = 20
      "0010100" when "01101100110010000", -- t[55696] = 20
      "0010100" when "01101100110010001", -- t[55697] = 20
      "0010100" when "01101100110010010", -- t[55698] = 20
      "0010100" when "01101100110010011", -- t[55699] = 20
      "0010100" when "01101100110010100", -- t[55700] = 20
      "0010100" when "01101100110010101", -- t[55701] = 20
      "0010100" when "01101100110010110", -- t[55702] = 20
      "0010100" when "01101100110010111", -- t[55703] = 20
      "0010100" when "01101100110011000", -- t[55704] = 20
      "0010100" when "01101100110011001", -- t[55705] = 20
      "0010100" when "01101100110011010", -- t[55706] = 20
      "0010100" when "01101100110011011", -- t[55707] = 20
      "0010100" when "01101100110011100", -- t[55708] = 20
      "0010100" when "01101100110011101", -- t[55709] = 20
      "0010100" when "01101100110011110", -- t[55710] = 20
      "0010100" when "01101100110011111", -- t[55711] = 20
      "0010100" when "01101100110100000", -- t[55712] = 20
      "0010100" when "01101100110100001", -- t[55713] = 20
      "0010100" when "01101100110100010", -- t[55714] = 20
      "0010100" when "01101100110100011", -- t[55715] = 20
      "0010100" when "01101100110100100", -- t[55716] = 20
      "0010100" when "01101100110100101", -- t[55717] = 20
      "0010100" when "01101100110100110", -- t[55718] = 20
      "0010100" when "01101100110100111", -- t[55719] = 20
      "0010100" when "01101100110101000", -- t[55720] = 20
      "0010100" when "01101100110101001", -- t[55721] = 20
      "0010100" when "01101100110101010", -- t[55722] = 20
      "0010100" when "01101100110101011", -- t[55723] = 20
      "0010100" when "01101100110101100", -- t[55724] = 20
      "0010100" when "01101100110101101", -- t[55725] = 20
      "0010100" when "01101100110101110", -- t[55726] = 20
      "0010100" when "01101100110101111", -- t[55727] = 20
      "0010100" when "01101100110110000", -- t[55728] = 20
      "0010100" when "01101100110110001", -- t[55729] = 20
      "0010100" when "01101100110110010", -- t[55730] = 20
      "0010100" when "01101100110110011", -- t[55731] = 20
      "0010100" when "01101100110110100", -- t[55732] = 20
      "0010100" when "01101100110110101", -- t[55733] = 20
      "0010100" when "01101100110110110", -- t[55734] = 20
      "0010100" when "01101100110110111", -- t[55735] = 20
      "0010100" when "01101100110111000", -- t[55736] = 20
      "0010100" when "01101100110111001", -- t[55737] = 20
      "0010100" when "01101100110111010", -- t[55738] = 20
      "0010100" when "01101100110111011", -- t[55739] = 20
      "0010100" when "01101100110111100", -- t[55740] = 20
      "0010100" when "01101100110111101", -- t[55741] = 20
      "0010100" when "01101100110111110", -- t[55742] = 20
      "0010100" when "01101100110111111", -- t[55743] = 20
      "0010100" when "01101100111000000", -- t[55744] = 20
      "0010100" when "01101100111000001", -- t[55745] = 20
      "0010100" when "01101100111000010", -- t[55746] = 20
      "0010100" when "01101100111000011", -- t[55747] = 20
      "0010100" when "01101100111000100", -- t[55748] = 20
      "0010100" when "01101100111000101", -- t[55749] = 20
      "0010100" when "01101100111000110", -- t[55750] = 20
      "0010100" when "01101100111000111", -- t[55751] = 20
      "0010100" when "01101100111001000", -- t[55752] = 20
      "0010100" when "01101100111001001", -- t[55753] = 20
      "0010100" when "01101100111001010", -- t[55754] = 20
      "0010100" when "01101100111001011", -- t[55755] = 20
      "0010100" when "01101100111001100", -- t[55756] = 20
      "0010100" when "01101100111001101", -- t[55757] = 20
      "0010100" when "01101100111001110", -- t[55758] = 20
      "0010100" when "01101100111001111", -- t[55759] = 20
      "0010100" when "01101100111010000", -- t[55760] = 20
      "0010100" when "01101100111010001", -- t[55761] = 20
      "0010100" when "01101100111010010", -- t[55762] = 20
      "0010100" when "01101100111010011", -- t[55763] = 20
      "0010100" when "01101100111010100", -- t[55764] = 20
      "0010100" when "01101100111010101", -- t[55765] = 20
      "0010100" when "01101100111010110", -- t[55766] = 20
      "0010100" when "01101100111010111", -- t[55767] = 20
      "0010100" when "01101100111011000", -- t[55768] = 20
      "0010100" when "01101100111011001", -- t[55769] = 20
      "0010100" when "01101100111011010", -- t[55770] = 20
      "0010100" when "01101100111011011", -- t[55771] = 20
      "0010100" when "01101100111011100", -- t[55772] = 20
      "0010100" when "01101100111011101", -- t[55773] = 20
      "0010100" when "01101100111011110", -- t[55774] = 20
      "0010100" when "01101100111011111", -- t[55775] = 20
      "0010100" when "01101100111100000", -- t[55776] = 20
      "0010100" when "01101100111100001", -- t[55777] = 20
      "0010100" when "01101100111100010", -- t[55778] = 20
      "0010100" when "01101100111100011", -- t[55779] = 20
      "0010100" when "01101100111100100", -- t[55780] = 20
      "0010100" when "01101100111100101", -- t[55781] = 20
      "0010100" when "01101100111100110", -- t[55782] = 20
      "0010100" when "01101100111100111", -- t[55783] = 20
      "0010100" when "01101100111101000", -- t[55784] = 20
      "0010100" when "01101100111101001", -- t[55785] = 20
      "0010100" when "01101100111101010", -- t[55786] = 20
      "0010100" when "01101100111101011", -- t[55787] = 20
      "0010100" when "01101100111101100", -- t[55788] = 20
      "0010100" when "01101100111101101", -- t[55789] = 20
      "0010100" when "01101100111101110", -- t[55790] = 20
      "0010100" when "01101100111101111", -- t[55791] = 20
      "0010100" when "01101100111110000", -- t[55792] = 20
      "0010100" when "01101100111110001", -- t[55793] = 20
      "0010100" when "01101100111110010", -- t[55794] = 20
      "0010100" when "01101100111110011", -- t[55795] = 20
      "0010100" when "01101100111110100", -- t[55796] = 20
      "0010100" when "01101100111110101", -- t[55797] = 20
      "0010100" when "01101100111110110", -- t[55798] = 20
      "0010100" when "01101100111110111", -- t[55799] = 20
      "0010100" when "01101100111111000", -- t[55800] = 20
      "0010100" when "01101100111111001", -- t[55801] = 20
      "0010100" when "01101100111111010", -- t[55802] = 20
      "0010100" when "01101100111111011", -- t[55803] = 20
      "0010100" when "01101100111111100", -- t[55804] = 20
      "0010100" when "01101100111111101", -- t[55805] = 20
      "0010100" when "01101100111111110", -- t[55806] = 20
      "0010100" when "01101100111111111", -- t[55807] = 20
      "0010100" when "01101101000000000", -- t[55808] = 20
      "0010100" when "01101101000000001", -- t[55809] = 20
      "0010100" when "01101101000000010", -- t[55810] = 20
      "0010100" when "01101101000000011", -- t[55811] = 20
      "0010100" when "01101101000000100", -- t[55812] = 20
      "0010100" when "01101101000000101", -- t[55813] = 20
      "0010100" when "01101101000000110", -- t[55814] = 20
      "0010100" when "01101101000000111", -- t[55815] = 20
      "0010100" when "01101101000001000", -- t[55816] = 20
      "0010100" when "01101101000001001", -- t[55817] = 20
      "0010100" when "01101101000001010", -- t[55818] = 20
      "0010100" when "01101101000001011", -- t[55819] = 20
      "0010100" when "01101101000001100", -- t[55820] = 20
      "0010100" when "01101101000001101", -- t[55821] = 20
      "0010100" when "01101101000001110", -- t[55822] = 20
      "0010100" when "01101101000001111", -- t[55823] = 20
      "0010100" when "01101101000010000", -- t[55824] = 20
      "0010100" when "01101101000010001", -- t[55825] = 20
      "0010100" when "01101101000010010", -- t[55826] = 20
      "0010100" when "01101101000010011", -- t[55827] = 20
      "0010100" when "01101101000010100", -- t[55828] = 20
      "0010100" when "01101101000010101", -- t[55829] = 20
      "0010100" when "01101101000010110", -- t[55830] = 20
      "0010100" when "01101101000010111", -- t[55831] = 20
      "0010100" when "01101101000011000", -- t[55832] = 20
      "0010100" when "01101101000011001", -- t[55833] = 20
      "0010100" when "01101101000011010", -- t[55834] = 20
      "0010100" when "01101101000011011", -- t[55835] = 20
      "0010100" when "01101101000011100", -- t[55836] = 20
      "0010100" when "01101101000011101", -- t[55837] = 20
      "0010100" when "01101101000011110", -- t[55838] = 20
      "0010100" when "01101101000011111", -- t[55839] = 20
      "0010100" when "01101101000100000", -- t[55840] = 20
      "0010100" when "01101101000100001", -- t[55841] = 20
      "0010100" when "01101101000100010", -- t[55842] = 20
      "0010100" when "01101101000100011", -- t[55843] = 20
      "0010100" when "01101101000100100", -- t[55844] = 20
      "0010100" when "01101101000100101", -- t[55845] = 20
      "0010100" when "01101101000100110", -- t[55846] = 20
      "0010100" when "01101101000100111", -- t[55847] = 20
      "0010100" when "01101101000101000", -- t[55848] = 20
      "0010100" when "01101101000101001", -- t[55849] = 20
      "0010100" when "01101101000101010", -- t[55850] = 20
      "0010100" when "01101101000101011", -- t[55851] = 20
      "0010100" when "01101101000101100", -- t[55852] = 20
      "0010100" when "01101101000101101", -- t[55853] = 20
      "0010100" when "01101101000101110", -- t[55854] = 20
      "0010100" when "01101101000101111", -- t[55855] = 20
      "0010100" when "01101101000110000", -- t[55856] = 20
      "0010100" when "01101101000110001", -- t[55857] = 20
      "0010100" when "01101101000110010", -- t[55858] = 20
      "0010100" when "01101101000110011", -- t[55859] = 20
      "0010100" when "01101101000110100", -- t[55860] = 20
      "0010100" when "01101101000110101", -- t[55861] = 20
      "0010100" when "01101101000110110", -- t[55862] = 20
      "0010100" when "01101101000110111", -- t[55863] = 20
      "0010100" when "01101101000111000", -- t[55864] = 20
      "0010100" when "01101101000111001", -- t[55865] = 20
      "0010100" when "01101101000111010", -- t[55866] = 20
      "0010100" when "01101101000111011", -- t[55867] = 20
      "0010100" when "01101101000111100", -- t[55868] = 20
      "0010100" when "01101101000111101", -- t[55869] = 20
      "0010100" when "01101101000111110", -- t[55870] = 20
      "0010100" when "01101101000111111", -- t[55871] = 20
      "0010100" when "01101101001000000", -- t[55872] = 20
      "0010100" when "01101101001000001", -- t[55873] = 20
      "0010100" when "01101101001000010", -- t[55874] = 20
      "0010100" when "01101101001000011", -- t[55875] = 20
      "0010100" when "01101101001000100", -- t[55876] = 20
      "0010100" when "01101101001000101", -- t[55877] = 20
      "0010100" when "01101101001000110", -- t[55878] = 20
      "0010100" when "01101101001000111", -- t[55879] = 20
      "0010100" when "01101101001001000", -- t[55880] = 20
      "0010100" when "01101101001001001", -- t[55881] = 20
      "0010100" when "01101101001001010", -- t[55882] = 20
      "0010100" when "01101101001001011", -- t[55883] = 20
      "0010100" when "01101101001001100", -- t[55884] = 20
      "0010100" when "01101101001001101", -- t[55885] = 20
      "0010100" when "01101101001001110", -- t[55886] = 20
      "0010100" when "01101101001001111", -- t[55887] = 20
      "0010100" when "01101101001010000", -- t[55888] = 20
      "0010100" when "01101101001010001", -- t[55889] = 20
      "0010100" when "01101101001010010", -- t[55890] = 20
      "0010100" when "01101101001010011", -- t[55891] = 20
      "0010100" when "01101101001010100", -- t[55892] = 20
      "0010100" when "01101101001010101", -- t[55893] = 20
      "0010100" when "01101101001010110", -- t[55894] = 20
      "0010100" when "01101101001010111", -- t[55895] = 20
      "0010100" when "01101101001011000", -- t[55896] = 20
      "0010100" when "01101101001011001", -- t[55897] = 20
      "0010100" when "01101101001011010", -- t[55898] = 20
      "0010100" when "01101101001011011", -- t[55899] = 20
      "0010100" when "01101101001011100", -- t[55900] = 20
      "0010100" when "01101101001011101", -- t[55901] = 20
      "0010100" when "01101101001011110", -- t[55902] = 20
      "0010100" when "01101101001011111", -- t[55903] = 20
      "0010100" when "01101101001100000", -- t[55904] = 20
      "0010100" when "01101101001100001", -- t[55905] = 20
      "0010100" when "01101101001100010", -- t[55906] = 20
      "0010100" when "01101101001100011", -- t[55907] = 20
      "0010100" when "01101101001100100", -- t[55908] = 20
      "0010100" when "01101101001100101", -- t[55909] = 20
      "0010100" when "01101101001100110", -- t[55910] = 20
      "0010100" when "01101101001100111", -- t[55911] = 20
      "0010100" when "01101101001101000", -- t[55912] = 20
      "0010100" when "01101101001101001", -- t[55913] = 20
      "0010100" when "01101101001101010", -- t[55914] = 20
      "0010100" when "01101101001101011", -- t[55915] = 20
      "0010100" when "01101101001101100", -- t[55916] = 20
      "0010100" when "01101101001101101", -- t[55917] = 20
      "0010100" when "01101101001101110", -- t[55918] = 20
      "0010100" when "01101101001101111", -- t[55919] = 20
      "0010100" when "01101101001110000", -- t[55920] = 20
      "0010100" when "01101101001110001", -- t[55921] = 20
      "0010100" when "01101101001110010", -- t[55922] = 20
      "0010100" when "01101101001110011", -- t[55923] = 20
      "0010100" when "01101101001110100", -- t[55924] = 20
      "0010100" when "01101101001110101", -- t[55925] = 20
      "0010100" when "01101101001110110", -- t[55926] = 20
      "0010100" when "01101101001110111", -- t[55927] = 20
      "0010100" when "01101101001111000", -- t[55928] = 20
      "0010100" when "01101101001111001", -- t[55929] = 20
      "0010100" when "01101101001111010", -- t[55930] = 20
      "0010100" when "01101101001111011", -- t[55931] = 20
      "0010101" when "01101101001111100", -- t[55932] = 21
      "0010101" when "01101101001111101", -- t[55933] = 21
      "0010101" when "01101101001111110", -- t[55934] = 21
      "0010101" when "01101101001111111", -- t[55935] = 21
      "0010101" when "01101101010000000", -- t[55936] = 21
      "0010101" when "01101101010000001", -- t[55937] = 21
      "0010101" when "01101101010000010", -- t[55938] = 21
      "0010101" when "01101101010000011", -- t[55939] = 21
      "0010101" when "01101101010000100", -- t[55940] = 21
      "0010101" when "01101101010000101", -- t[55941] = 21
      "0010101" when "01101101010000110", -- t[55942] = 21
      "0010101" when "01101101010000111", -- t[55943] = 21
      "0010101" when "01101101010001000", -- t[55944] = 21
      "0010101" when "01101101010001001", -- t[55945] = 21
      "0010101" when "01101101010001010", -- t[55946] = 21
      "0010101" when "01101101010001011", -- t[55947] = 21
      "0010101" when "01101101010001100", -- t[55948] = 21
      "0010101" when "01101101010001101", -- t[55949] = 21
      "0010101" when "01101101010001110", -- t[55950] = 21
      "0010101" when "01101101010001111", -- t[55951] = 21
      "0010101" when "01101101010010000", -- t[55952] = 21
      "0010101" when "01101101010010001", -- t[55953] = 21
      "0010101" when "01101101010010010", -- t[55954] = 21
      "0010101" when "01101101010010011", -- t[55955] = 21
      "0010101" when "01101101010010100", -- t[55956] = 21
      "0010101" when "01101101010010101", -- t[55957] = 21
      "0010101" when "01101101010010110", -- t[55958] = 21
      "0010101" when "01101101010010111", -- t[55959] = 21
      "0010101" when "01101101010011000", -- t[55960] = 21
      "0010101" when "01101101010011001", -- t[55961] = 21
      "0010101" when "01101101010011010", -- t[55962] = 21
      "0010101" when "01101101010011011", -- t[55963] = 21
      "0010101" when "01101101010011100", -- t[55964] = 21
      "0010101" when "01101101010011101", -- t[55965] = 21
      "0010101" when "01101101010011110", -- t[55966] = 21
      "0010101" when "01101101010011111", -- t[55967] = 21
      "0010101" when "01101101010100000", -- t[55968] = 21
      "0010101" when "01101101010100001", -- t[55969] = 21
      "0010101" when "01101101010100010", -- t[55970] = 21
      "0010101" when "01101101010100011", -- t[55971] = 21
      "0010101" when "01101101010100100", -- t[55972] = 21
      "0010101" when "01101101010100101", -- t[55973] = 21
      "0010101" when "01101101010100110", -- t[55974] = 21
      "0010101" when "01101101010100111", -- t[55975] = 21
      "0010101" when "01101101010101000", -- t[55976] = 21
      "0010101" when "01101101010101001", -- t[55977] = 21
      "0010101" when "01101101010101010", -- t[55978] = 21
      "0010101" when "01101101010101011", -- t[55979] = 21
      "0010101" when "01101101010101100", -- t[55980] = 21
      "0010101" when "01101101010101101", -- t[55981] = 21
      "0010101" when "01101101010101110", -- t[55982] = 21
      "0010101" when "01101101010101111", -- t[55983] = 21
      "0010101" when "01101101010110000", -- t[55984] = 21
      "0010101" when "01101101010110001", -- t[55985] = 21
      "0010101" when "01101101010110010", -- t[55986] = 21
      "0010101" when "01101101010110011", -- t[55987] = 21
      "0010101" when "01101101010110100", -- t[55988] = 21
      "0010101" when "01101101010110101", -- t[55989] = 21
      "0010101" when "01101101010110110", -- t[55990] = 21
      "0010101" when "01101101010110111", -- t[55991] = 21
      "0010101" when "01101101010111000", -- t[55992] = 21
      "0010101" when "01101101010111001", -- t[55993] = 21
      "0010101" when "01101101010111010", -- t[55994] = 21
      "0010101" when "01101101010111011", -- t[55995] = 21
      "0010101" when "01101101010111100", -- t[55996] = 21
      "0010101" when "01101101010111101", -- t[55997] = 21
      "0010101" when "01101101010111110", -- t[55998] = 21
      "0010101" when "01101101010111111", -- t[55999] = 21
      "0010101" when "01101101011000000", -- t[56000] = 21
      "0010101" when "01101101011000001", -- t[56001] = 21
      "0010101" when "01101101011000010", -- t[56002] = 21
      "0010101" when "01101101011000011", -- t[56003] = 21
      "0010101" when "01101101011000100", -- t[56004] = 21
      "0010101" when "01101101011000101", -- t[56005] = 21
      "0010101" when "01101101011000110", -- t[56006] = 21
      "0010101" when "01101101011000111", -- t[56007] = 21
      "0010101" when "01101101011001000", -- t[56008] = 21
      "0010101" when "01101101011001001", -- t[56009] = 21
      "0010101" when "01101101011001010", -- t[56010] = 21
      "0010101" when "01101101011001011", -- t[56011] = 21
      "0010101" when "01101101011001100", -- t[56012] = 21
      "0010101" when "01101101011001101", -- t[56013] = 21
      "0010101" when "01101101011001110", -- t[56014] = 21
      "0010101" when "01101101011001111", -- t[56015] = 21
      "0010101" when "01101101011010000", -- t[56016] = 21
      "0010101" when "01101101011010001", -- t[56017] = 21
      "0010101" when "01101101011010010", -- t[56018] = 21
      "0010101" when "01101101011010011", -- t[56019] = 21
      "0010101" when "01101101011010100", -- t[56020] = 21
      "0010101" when "01101101011010101", -- t[56021] = 21
      "0010101" when "01101101011010110", -- t[56022] = 21
      "0010101" when "01101101011010111", -- t[56023] = 21
      "0010101" when "01101101011011000", -- t[56024] = 21
      "0010101" when "01101101011011001", -- t[56025] = 21
      "0010101" when "01101101011011010", -- t[56026] = 21
      "0010101" when "01101101011011011", -- t[56027] = 21
      "0010101" when "01101101011011100", -- t[56028] = 21
      "0010101" when "01101101011011101", -- t[56029] = 21
      "0010101" when "01101101011011110", -- t[56030] = 21
      "0010101" when "01101101011011111", -- t[56031] = 21
      "0010101" when "01101101011100000", -- t[56032] = 21
      "0010101" when "01101101011100001", -- t[56033] = 21
      "0010101" when "01101101011100010", -- t[56034] = 21
      "0010101" when "01101101011100011", -- t[56035] = 21
      "0010101" when "01101101011100100", -- t[56036] = 21
      "0010101" when "01101101011100101", -- t[56037] = 21
      "0010101" when "01101101011100110", -- t[56038] = 21
      "0010101" when "01101101011100111", -- t[56039] = 21
      "0010101" when "01101101011101000", -- t[56040] = 21
      "0010101" when "01101101011101001", -- t[56041] = 21
      "0010101" when "01101101011101010", -- t[56042] = 21
      "0010101" when "01101101011101011", -- t[56043] = 21
      "0010101" when "01101101011101100", -- t[56044] = 21
      "0010101" when "01101101011101101", -- t[56045] = 21
      "0010101" when "01101101011101110", -- t[56046] = 21
      "0010101" when "01101101011101111", -- t[56047] = 21
      "0010101" when "01101101011110000", -- t[56048] = 21
      "0010101" when "01101101011110001", -- t[56049] = 21
      "0010101" when "01101101011110010", -- t[56050] = 21
      "0010101" when "01101101011110011", -- t[56051] = 21
      "0010101" when "01101101011110100", -- t[56052] = 21
      "0010101" when "01101101011110101", -- t[56053] = 21
      "0010101" when "01101101011110110", -- t[56054] = 21
      "0010101" when "01101101011110111", -- t[56055] = 21
      "0010101" when "01101101011111000", -- t[56056] = 21
      "0010101" when "01101101011111001", -- t[56057] = 21
      "0010101" when "01101101011111010", -- t[56058] = 21
      "0010101" when "01101101011111011", -- t[56059] = 21
      "0010101" when "01101101011111100", -- t[56060] = 21
      "0010101" when "01101101011111101", -- t[56061] = 21
      "0010101" when "01101101011111110", -- t[56062] = 21
      "0010101" when "01101101011111111", -- t[56063] = 21
      "0010101" when "01101101100000000", -- t[56064] = 21
      "0010101" when "01101101100000001", -- t[56065] = 21
      "0010101" when "01101101100000010", -- t[56066] = 21
      "0010101" when "01101101100000011", -- t[56067] = 21
      "0010101" when "01101101100000100", -- t[56068] = 21
      "0010101" when "01101101100000101", -- t[56069] = 21
      "0010101" when "01101101100000110", -- t[56070] = 21
      "0010101" when "01101101100000111", -- t[56071] = 21
      "0010101" when "01101101100001000", -- t[56072] = 21
      "0010101" when "01101101100001001", -- t[56073] = 21
      "0010101" when "01101101100001010", -- t[56074] = 21
      "0010101" when "01101101100001011", -- t[56075] = 21
      "0010101" when "01101101100001100", -- t[56076] = 21
      "0010101" when "01101101100001101", -- t[56077] = 21
      "0010101" when "01101101100001110", -- t[56078] = 21
      "0010101" when "01101101100001111", -- t[56079] = 21
      "0010101" when "01101101100010000", -- t[56080] = 21
      "0010101" when "01101101100010001", -- t[56081] = 21
      "0010101" when "01101101100010010", -- t[56082] = 21
      "0010101" when "01101101100010011", -- t[56083] = 21
      "0010101" when "01101101100010100", -- t[56084] = 21
      "0010101" when "01101101100010101", -- t[56085] = 21
      "0010101" when "01101101100010110", -- t[56086] = 21
      "0010101" when "01101101100010111", -- t[56087] = 21
      "0010101" when "01101101100011000", -- t[56088] = 21
      "0010101" when "01101101100011001", -- t[56089] = 21
      "0010101" when "01101101100011010", -- t[56090] = 21
      "0010101" when "01101101100011011", -- t[56091] = 21
      "0010101" when "01101101100011100", -- t[56092] = 21
      "0010101" when "01101101100011101", -- t[56093] = 21
      "0010101" when "01101101100011110", -- t[56094] = 21
      "0010101" when "01101101100011111", -- t[56095] = 21
      "0010101" when "01101101100100000", -- t[56096] = 21
      "0010101" when "01101101100100001", -- t[56097] = 21
      "0010101" when "01101101100100010", -- t[56098] = 21
      "0010101" when "01101101100100011", -- t[56099] = 21
      "0010101" when "01101101100100100", -- t[56100] = 21
      "0010101" when "01101101100100101", -- t[56101] = 21
      "0010101" when "01101101100100110", -- t[56102] = 21
      "0010101" when "01101101100100111", -- t[56103] = 21
      "0010101" when "01101101100101000", -- t[56104] = 21
      "0010101" when "01101101100101001", -- t[56105] = 21
      "0010101" when "01101101100101010", -- t[56106] = 21
      "0010101" when "01101101100101011", -- t[56107] = 21
      "0010101" when "01101101100101100", -- t[56108] = 21
      "0010101" when "01101101100101101", -- t[56109] = 21
      "0010101" when "01101101100101110", -- t[56110] = 21
      "0010101" when "01101101100101111", -- t[56111] = 21
      "0010101" when "01101101100110000", -- t[56112] = 21
      "0010101" when "01101101100110001", -- t[56113] = 21
      "0010101" when "01101101100110010", -- t[56114] = 21
      "0010101" when "01101101100110011", -- t[56115] = 21
      "0010101" when "01101101100110100", -- t[56116] = 21
      "0010101" when "01101101100110101", -- t[56117] = 21
      "0010101" when "01101101100110110", -- t[56118] = 21
      "0010101" when "01101101100110111", -- t[56119] = 21
      "0010101" when "01101101100111000", -- t[56120] = 21
      "0010101" when "01101101100111001", -- t[56121] = 21
      "0010101" when "01101101100111010", -- t[56122] = 21
      "0010101" when "01101101100111011", -- t[56123] = 21
      "0010101" when "01101101100111100", -- t[56124] = 21
      "0010101" when "01101101100111101", -- t[56125] = 21
      "0010101" when "01101101100111110", -- t[56126] = 21
      "0010101" when "01101101100111111", -- t[56127] = 21
      "0010101" when "01101101101000000", -- t[56128] = 21
      "0010101" when "01101101101000001", -- t[56129] = 21
      "0010101" when "01101101101000010", -- t[56130] = 21
      "0010101" when "01101101101000011", -- t[56131] = 21
      "0010101" when "01101101101000100", -- t[56132] = 21
      "0010101" when "01101101101000101", -- t[56133] = 21
      "0010101" when "01101101101000110", -- t[56134] = 21
      "0010101" when "01101101101000111", -- t[56135] = 21
      "0010101" when "01101101101001000", -- t[56136] = 21
      "0010101" when "01101101101001001", -- t[56137] = 21
      "0010101" when "01101101101001010", -- t[56138] = 21
      "0010101" when "01101101101001011", -- t[56139] = 21
      "0010101" when "01101101101001100", -- t[56140] = 21
      "0010101" when "01101101101001101", -- t[56141] = 21
      "0010101" when "01101101101001110", -- t[56142] = 21
      "0010101" when "01101101101001111", -- t[56143] = 21
      "0010101" when "01101101101010000", -- t[56144] = 21
      "0010101" when "01101101101010001", -- t[56145] = 21
      "0010101" when "01101101101010010", -- t[56146] = 21
      "0010101" when "01101101101010011", -- t[56147] = 21
      "0010101" when "01101101101010100", -- t[56148] = 21
      "0010101" when "01101101101010101", -- t[56149] = 21
      "0010101" when "01101101101010110", -- t[56150] = 21
      "0010101" when "01101101101010111", -- t[56151] = 21
      "0010101" when "01101101101011000", -- t[56152] = 21
      "0010101" when "01101101101011001", -- t[56153] = 21
      "0010101" when "01101101101011010", -- t[56154] = 21
      "0010101" when "01101101101011011", -- t[56155] = 21
      "0010101" when "01101101101011100", -- t[56156] = 21
      "0010101" when "01101101101011101", -- t[56157] = 21
      "0010101" when "01101101101011110", -- t[56158] = 21
      "0010101" when "01101101101011111", -- t[56159] = 21
      "0010101" when "01101101101100000", -- t[56160] = 21
      "0010101" when "01101101101100001", -- t[56161] = 21
      "0010101" when "01101101101100010", -- t[56162] = 21
      "0010101" when "01101101101100011", -- t[56163] = 21
      "0010101" when "01101101101100100", -- t[56164] = 21
      "0010101" when "01101101101100101", -- t[56165] = 21
      "0010101" when "01101101101100110", -- t[56166] = 21
      "0010101" when "01101101101100111", -- t[56167] = 21
      "0010101" when "01101101101101000", -- t[56168] = 21
      "0010101" when "01101101101101001", -- t[56169] = 21
      "0010101" when "01101101101101010", -- t[56170] = 21
      "0010101" when "01101101101101011", -- t[56171] = 21
      "0010101" when "01101101101101100", -- t[56172] = 21
      "0010101" when "01101101101101101", -- t[56173] = 21
      "0010101" when "01101101101101110", -- t[56174] = 21
      "0010101" when "01101101101101111", -- t[56175] = 21
      "0010101" when "01101101101110000", -- t[56176] = 21
      "0010101" when "01101101101110001", -- t[56177] = 21
      "0010101" when "01101101101110010", -- t[56178] = 21
      "0010101" when "01101101101110011", -- t[56179] = 21
      "0010101" when "01101101101110100", -- t[56180] = 21
      "0010101" when "01101101101110101", -- t[56181] = 21
      "0010101" when "01101101101110110", -- t[56182] = 21
      "0010101" when "01101101101110111", -- t[56183] = 21
      "0010101" when "01101101101111000", -- t[56184] = 21
      "0010101" when "01101101101111001", -- t[56185] = 21
      "0010101" when "01101101101111010", -- t[56186] = 21
      "0010101" when "01101101101111011", -- t[56187] = 21
      "0010101" when "01101101101111100", -- t[56188] = 21
      "0010101" when "01101101101111101", -- t[56189] = 21
      "0010101" when "01101101101111110", -- t[56190] = 21
      "0010101" when "01101101101111111", -- t[56191] = 21
      "0010101" when "01101101110000000", -- t[56192] = 21
      "0010101" when "01101101110000001", -- t[56193] = 21
      "0010101" when "01101101110000010", -- t[56194] = 21
      "0010101" when "01101101110000011", -- t[56195] = 21
      "0010101" when "01101101110000100", -- t[56196] = 21
      "0010101" when "01101101110000101", -- t[56197] = 21
      "0010101" when "01101101110000110", -- t[56198] = 21
      "0010101" when "01101101110000111", -- t[56199] = 21
      "0010101" when "01101101110001000", -- t[56200] = 21
      "0010101" when "01101101110001001", -- t[56201] = 21
      "0010101" when "01101101110001010", -- t[56202] = 21
      "0010101" when "01101101110001011", -- t[56203] = 21
      "0010101" when "01101101110001100", -- t[56204] = 21
      "0010101" when "01101101110001101", -- t[56205] = 21
      "0010101" when "01101101110001110", -- t[56206] = 21
      "0010101" when "01101101110001111", -- t[56207] = 21
      "0010101" when "01101101110010000", -- t[56208] = 21
      "0010101" when "01101101110010001", -- t[56209] = 21
      "0010101" when "01101101110010010", -- t[56210] = 21
      "0010101" when "01101101110010011", -- t[56211] = 21
      "0010101" when "01101101110010100", -- t[56212] = 21
      "0010101" when "01101101110010101", -- t[56213] = 21
      "0010101" when "01101101110010110", -- t[56214] = 21
      "0010101" when "01101101110010111", -- t[56215] = 21
      "0010101" when "01101101110011000", -- t[56216] = 21
      "0010101" when "01101101110011001", -- t[56217] = 21
      "0010101" when "01101101110011010", -- t[56218] = 21
      "0010101" when "01101101110011011", -- t[56219] = 21
      "0010101" when "01101101110011100", -- t[56220] = 21
      "0010101" when "01101101110011101", -- t[56221] = 21
      "0010101" when "01101101110011110", -- t[56222] = 21
      "0010101" when "01101101110011111", -- t[56223] = 21
      "0010101" when "01101101110100000", -- t[56224] = 21
      "0010101" when "01101101110100001", -- t[56225] = 21
      "0010101" when "01101101110100010", -- t[56226] = 21
      "0010101" when "01101101110100011", -- t[56227] = 21
      "0010101" when "01101101110100100", -- t[56228] = 21
      "0010101" when "01101101110100101", -- t[56229] = 21
      "0010101" when "01101101110100110", -- t[56230] = 21
      "0010101" when "01101101110100111", -- t[56231] = 21
      "0010101" when "01101101110101000", -- t[56232] = 21
      "0010101" when "01101101110101001", -- t[56233] = 21
      "0010101" when "01101101110101010", -- t[56234] = 21
      "0010101" when "01101101110101011", -- t[56235] = 21
      "0010101" when "01101101110101100", -- t[56236] = 21
      "0010101" when "01101101110101101", -- t[56237] = 21
      "0010101" when "01101101110101110", -- t[56238] = 21
      "0010101" when "01101101110101111", -- t[56239] = 21
      "0010101" when "01101101110110000", -- t[56240] = 21
      "0010101" when "01101101110110001", -- t[56241] = 21
      "0010101" when "01101101110110010", -- t[56242] = 21
      "0010101" when "01101101110110011", -- t[56243] = 21
      "0010101" when "01101101110110100", -- t[56244] = 21
      "0010101" when "01101101110110101", -- t[56245] = 21
      "0010101" when "01101101110110110", -- t[56246] = 21
      "0010101" when "01101101110110111", -- t[56247] = 21
      "0010101" when "01101101110111000", -- t[56248] = 21
      "0010101" when "01101101110111001", -- t[56249] = 21
      "0010101" when "01101101110111010", -- t[56250] = 21
      "0010101" when "01101101110111011", -- t[56251] = 21
      "0010101" when "01101101110111100", -- t[56252] = 21
      "0010101" when "01101101110111101", -- t[56253] = 21
      "0010101" when "01101101110111110", -- t[56254] = 21
      "0010101" when "01101101110111111", -- t[56255] = 21
      "0010101" when "01101101111000000", -- t[56256] = 21
      "0010101" when "01101101111000001", -- t[56257] = 21
      "0010101" when "01101101111000010", -- t[56258] = 21
      "0010101" when "01101101111000011", -- t[56259] = 21
      "0010101" when "01101101111000100", -- t[56260] = 21
      "0010101" when "01101101111000101", -- t[56261] = 21
      "0010101" when "01101101111000110", -- t[56262] = 21
      "0010101" when "01101101111000111", -- t[56263] = 21
      "0010101" when "01101101111001000", -- t[56264] = 21
      "0010101" when "01101101111001001", -- t[56265] = 21
      "0010101" when "01101101111001010", -- t[56266] = 21
      "0010101" when "01101101111001011", -- t[56267] = 21
      "0010101" when "01101101111001100", -- t[56268] = 21
      "0010101" when "01101101111001101", -- t[56269] = 21
      "0010101" when "01101101111001110", -- t[56270] = 21
      "0010101" when "01101101111001111", -- t[56271] = 21
      "0010101" when "01101101111010000", -- t[56272] = 21
      "0010101" when "01101101111010001", -- t[56273] = 21
      "0010101" when "01101101111010010", -- t[56274] = 21
      "0010101" when "01101101111010011", -- t[56275] = 21
      "0010101" when "01101101111010100", -- t[56276] = 21
      "0010101" when "01101101111010101", -- t[56277] = 21
      "0010101" when "01101101111010110", -- t[56278] = 21
      "0010101" when "01101101111010111", -- t[56279] = 21
      "0010101" when "01101101111011000", -- t[56280] = 21
      "0010101" when "01101101111011001", -- t[56281] = 21
      "0010101" when "01101101111011010", -- t[56282] = 21
      "0010101" when "01101101111011011", -- t[56283] = 21
      "0010101" when "01101101111011100", -- t[56284] = 21
      "0010101" when "01101101111011101", -- t[56285] = 21
      "0010101" when "01101101111011110", -- t[56286] = 21
      "0010101" when "01101101111011111", -- t[56287] = 21
      "0010101" when "01101101111100000", -- t[56288] = 21
      "0010101" when "01101101111100001", -- t[56289] = 21
      "0010101" when "01101101111100010", -- t[56290] = 21
      "0010101" when "01101101111100011", -- t[56291] = 21
      "0010101" when "01101101111100100", -- t[56292] = 21
      "0010101" when "01101101111100101", -- t[56293] = 21
      "0010101" when "01101101111100110", -- t[56294] = 21
      "0010101" when "01101101111100111", -- t[56295] = 21
      "0010101" when "01101101111101000", -- t[56296] = 21
      "0010101" when "01101101111101001", -- t[56297] = 21
      "0010101" when "01101101111101010", -- t[56298] = 21
      "0010101" when "01101101111101011", -- t[56299] = 21
      "0010101" when "01101101111101100", -- t[56300] = 21
      "0010101" when "01101101111101101", -- t[56301] = 21
      "0010101" when "01101101111101110", -- t[56302] = 21
      "0010101" when "01101101111101111", -- t[56303] = 21
      "0010101" when "01101101111110000", -- t[56304] = 21
      "0010101" when "01101101111110001", -- t[56305] = 21
      "0010101" when "01101101111110010", -- t[56306] = 21
      "0010101" when "01101101111110011", -- t[56307] = 21
      "0010101" when "01101101111110100", -- t[56308] = 21
      "0010101" when "01101101111110101", -- t[56309] = 21
      "0010101" when "01101101111110110", -- t[56310] = 21
      "0010101" when "01101101111110111", -- t[56311] = 21
      "0010101" when "01101101111111000", -- t[56312] = 21
      "0010101" when "01101101111111001", -- t[56313] = 21
      "0010101" when "01101101111111010", -- t[56314] = 21
      "0010101" when "01101101111111011", -- t[56315] = 21
      "0010101" when "01101101111111100", -- t[56316] = 21
      "0010101" when "01101101111111101", -- t[56317] = 21
      "0010101" when "01101101111111110", -- t[56318] = 21
      "0010101" when "01101101111111111", -- t[56319] = 21
      "0010101" when "01101110000000000", -- t[56320] = 21
      "0010101" when "01101110000000001", -- t[56321] = 21
      "0010101" when "01101110000000010", -- t[56322] = 21
      "0010101" when "01101110000000011", -- t[56323] = 21
      "0010101" when "01101110000000100", -- t[56324] = 21
      "0010101" when "01101110000000101", -- t[56325] = 21
      "0010101" when "01101110000000110", -- t[56326] = 21
      "0010101" when "01101110000000111", -- t[56327] = 21
      "0010101" when "01101110000001000", -- t[56328] = 21
      "0010101" when "01101110000001001", -- t[56329] = 21
      "0010101" when "01101110000001010", -- t[56330] = 21
      "0010101" when "01101110000001011", -- t[56331] = 21
      "0010101" when "01101110000001100", -- t[56332] = 21
      "0010101" when "01101110000001101", -- t[56333] = 21
      "0010101" when "01101110000001110", -- t[56334] = 21
      "0010101" when "01101110000001111", -- t[56335] = 21
      "0010101" when "01101110000010000", -- t[56336] = 21
      "0010101" when "01101110000010001", -- t[56337] = 21
      "0010101" when "01101110000010010", -- t[56338] = 21
      "0010101" when "01101110000010011", -- t[56339] = 21
      "0010101" when "01101110000010100", -- t[56340] = 21
      "0010101" when "01101110000010101", -- t[56341] = 21
      "0010101" when "01101110000010110", -- t[56342] = 21
      "0010101" when "01101110000010111", -- t[56343] = 21
      "0010101" when "01101110000011000", -- t[56344] = 21
      "0010101" when "01101110000011001", -- t[56345] = 21
      "0010101" when "01101110000011010", -- t[56346] = 21
      "0010101" when "01101110000011011", -- t[56347] = 21
      "0010101" when "01101110000011100", -- t[56348] = 21
      "0010101" when "01101110000011101", -- t[56349] = 21
      "0010101" when "01101110000011110", -- t[56350] = 21
      "0010101" when "01101110000011111", -- t[56351] = 21
      "0010101" when "01101110000100000", -- t[56352] = 21
      "0010101" when "01101110000100001", -- t[56353] = 21
      "0010101" when "01101110000100010", -- t[56354] = 21
      "0010101" when "01101110000100011", -- t[56355] = 21
      "0010101" when "01101110000100100", -- t[56356] = 21
      "0010101" when "01101110000100101", -- t[56357] = 21
      "0010101" when "01101110000100110", -- t[56358] = 21
      "0010101" when "01101110000100111", -- t[56359] = 21
      "0010101" when "01101110000101000", -- t[56360] = 21
      "0010101" when "01101110000101001", -- t[56361] = 21
      "0010101" when "01101110000101010", -- t[56362] = 21
      "0010101" when "01101110000101011", -- t[56363] = 21
      "0010101" when "01101110000101100", -- t[56364] = 21
      "0010101" when "01101110000101101", -- t[56365] = 21
      "0010101" when "01101110000101110", -- t[56366] = 21
      "0010101" when "01101110000101111", -- t[56367] = 21
      "0010101" when "01101110000110000", -- t[56368] = 21
      "0010101" when "01101110000110001", -- t[56369] = 21
      "0010101" when "01101110000110010", -- t[56370] = 21
      "0010101" when "01101110000110011", -- t[56371] = 21
      "0010101" when "01101110000110100", -- t[56372] = 21
      "0010101" when "01101110000110101", -- t[56373] = 21
      "0010101" when "01101110000110110", -- t[56374] = 21
      "0010101" when "01101110000110111", -- t[56375] = 21
      "0010101" when "01101110000111000", -- t[56376] = 21
      "0010101" when "01101110000111001", -- t[56377] = 21
      "0010101" when "01101110000111010", -- t[56378] = 21
      "0010101" when "01101110000111011", -- t[56379] = 21
      "0010101" when "01101110000111100", -- t[56380] = 21
      "0010101" when "01101110000111101", -- t[56381] = 21
      "0010101" when "01101110000111110", -- t[56382] = 21
      "0010101" when "01101110000111111", -- t[56383] = 21
      "0010101" when "01101110001000000", -- t[56384] = 21
      "0010101" when "01101110001000001", -- t[56385] = 21
      "0010101" when "01101110001000010", -- t[56386] = 21
      "0010101" when "01101110001000011", -- t[56387] = 21
      "0010101" when "01101110001000100", -- t[56388] = 21
      "0010101" when "01101110001000101", -- t[56389] = 21
      "0010101" when "01101110001000110", -- t[56390] = 21
      "0010101" when "01101110001000111", -- t[56391] = 21
      "0010101" when "01101110001001000", -- t[56392] = 21
      "0010101" when "01101110001001001", -- t[56393] = 21
      "0010101" when "01101110001001010", -- t[56394] = 21
      "0010101" when "01101110001001011", -- t[56395] = 21
      "0010101" when "01101110001001100", -- t[56396] = 21
      "0010101" when "01101110001001101", -- t[56397] = 21
      "0010101" when "01101110001001110", -- t[56398] = 21
      "0010101" when "01101110001001111", -- t[56399] = 21
      "0010101" when "01101110001010000", -- t[56400] = 21
      "0010101" when "01101110001010001", -- t[56401] = 21
      "0010101" when "01101110001010010", -- t[56402] = 21
      "0010101" when "01101110001010011", -- t[56403] = 21
      "0010101" when "01101110001010100", -- t[56404] = 21
      "0010101" when "01101110001010101", -- t[56405] = 21
      "0010101" when "01101110001010110", -- t[56406] = 21
      "0010101" when "01101110001010111", -- t[56407] = 21
      "0010101" when "01101110001011000", -- t[56408] = 21
      "0010101" when "01101110001011001", -- t[56409] = 21
      "0010101" when "01101110001011010", -- t[56410] = 21
      "0010101" when "01101110001011011", -- t[56411] = 21
      "0010101" when "01101110001011100", -- t[56412] = 21
      "0010101" when "01101110001011101", -- t[56413] = 21
      "0010101" when "01101110001011110", -- t[56414] = 21
      "0010101" when "01101110001011111", -- t[56415] = 21
      "0010101" when "01101110001100000", -- t[56416] = 21
      "0010101" when "01101110001100001", -- t[56417] = 21
      "0010101" when "01101110001100010", -- t[56418] = 21
      "0010101" when "01101110001100011", -- t[56419] = 21
      "0010101" when "01101110001100100", -- t[56420] = 21
      "0010101" when "01101110001100101", -- t[56421] = 21
      "0010101" when "01101110001100110", -- t[56422] = 21
      "0010101" when "01101110001100111", -- t[56423] = 21
      "0010101" when "01101110001101000", -- t[56424] = 21
      "0010101" when "01101110001101001", -- t[56425] = 21
      "0010101" when "01101110001101010", -- t[56426] = 21
      "0010101" when "01101110001101011", -- t[56427] = 21
      "0010101" when "01101110001101100", -- t[56428] = 21
      "0010101" when "01101110001101101", -- t[56429] = 21
      "0010101" when "01101110001101110", -- t[56430] = 21
      "0010101" when "01101110001101111", -- t[56431] = 21
      "0010101" when "01101110001110000", -- t[56432] = 21
      "0010101" when "01101110001110001", -- t[56433] = 21
      "0010101" when "01101110001110010", -- t[56434] = 21
      "0010101" when "01101110001110011", -- t[56435] = 21
      "0010101" when "01101110001110100", -- t[56436] = 21
      "0010101" when "01101110001110101", -- t[56437] = 21
      "0010101" when "01101110001110110", -- t[56438] = 21
      "0010101" when "01101110001110111", -- t[56439] = 21
      "0010101" when "01101110001111000", -- t[56440] = 21
      "0010101" when "01101110001111001", -- t[56441] = 21
      "0010101" when "01101110001111010", -- t[56442] = 21
      "0010101" when "01101110001111011", -- t[56443] = 21
      "0010101" when "01101110001111100", -- t[56444] = 21
      "0010101" when "01101110001111101", -- t[56445] = 21
      "0010101" when "01101110001111110", -- t[56446] = 21
      "0010101" when "01101110001111111", -- t[56447] = 21
      "0010101" when "01101110010000000", -- t[56448] = 21
      "0010101" when "01101110010000001", -- t[56449] = 21
      "0010101" when "01101110010000010", -- t[56450] = 21
      "0010101" when "01101110010000011", -- t[56451] = 21
      "0010101" when "01101110010000100", -- t[56452] = 21
      "0010101" when "01101110010000101", -- t[56453] = 21
      "0010101" when "01101110010000110", -- t[56454] = 21
      "0010101" when "01101110010000111", -- t[56455] = 21
      "0010101" when "01101110010001000", -- t[56456] = 21
      "0010101" when "01101110010001001", -- t[56457] = 21
      "0010101" when "01101110010001010", -- t[56458] = 21
      "0010101" when "01101110010001011", -- t[56459] = 21
      "0010101" when "01101110010001100", -- t[56460] = 21
      "0010101" when "01101110010001101", -- t[56461] = 21
      "0010101" when "01101110010001110", -- t[56462] = 21
      "0010101" when "01101110010001111", -- t[56463] = 21
      "0010101" when "01101110010010000", -- t[56464] = 21
      "0010101" when "01101110010010001", -- t[56465] = 21
      "0010101" when "01101110010010010", -- t[56466] = 21
      "0010101" when "01101110010010011", -- t[56467] = 21
      "0010101" when "01101110010010100", -- t[56468] = 21
      "0010101" when "01101110010010101", -- t[56469] = 21
      "0010101" when "01101110010010110", -- t[56470] = 21
      "0010101" when "01101110010010111", -- t[56471] = 21
      "0010101" when "01101110010011000", -- t[56472] = 21
      "0010101" when "01101110010011001", -- t[56473] = 21
      "0010101" when "01101110010011010", -- t[56474] = 21
      "0010101" when "01101110010011011", -- t[56475] = 21
      "0010101" when "01101110010011100", -- t[56476] = 21
      "0010101" when "01101110010011101", -- t[56477] = 21
      "0010101" when "01101110010011110", -- t[56478] = 21
      "0010101" when "01101110010011111", -- t[56479] = 21
      "0010101" when "01101110010100000", -- t[56480] = 21
      "0010101" when "01101110010100001", -- t[56481] = 21
      "0010101" when "01101110010100010", -- t[56482] = 21
      "0010101" when "01101110010100011", -- t[56483] = 21
      "0010101" when "01101110010100100", -- t[56484] = 21
      "0010101" when "01101110010100101", -- t[56485] = 21
      "0010101" when "01101110010100110", -- t[56486] = 21
      "0010101" when "01101110010100111", -- t[56487] = 21
      "0010101" when "01101110010101000", -- t[56488] = 21
      "0010101" when "01101110010101001", -- t[56489] = 21
      "0010101" when "01101110010101010", -- t[56490] = 21
      "0010101" when "01101110010101011", -- t[56491] = 21
      "0010101" when "01101110010101100", -- t[56492] = 21
      "0010101" when "01101110010101101", -- t[56493] = 21
      "0010110" when "01101110010101110", -- t[56494] = 22
      "0010110" when "01101110010101111", -- t[56495] = 22
      "0010110" when "01101110010110000", -- t[56496] = 22
      "0010110" when "01101110010110001", -- t[56497] = 22
      "0010110" when "01101110010110010", -- t[56498] = 22
      "0010110" when "01101110010110011", -- t[56499] = 22
      "0010110" when "01101110010110100", -- t[56500] = 22
      "0010110" when "01101110010110101", -- t[56501] = 22
      "0010110" when "01101110010110110", -- t[56502] = 22
      "0010110" when "01101110010110111", -- t[56503] = 22
      "0010110" when "01101110010111000", -- t[56504] = 22
      "0010110" when "01101110010111001", -- t[56505] = 22
      "0010110" when "01101110010111010", -- t[56506] = 22
      "0010110" when "01101110010111011", -- t[56507] = 22
      "0010110" when "01101110010111100", -- t[56508] = 22
      "0010110" when "01101110010111101", -- t[56509] = 22
      "0010110" when "01101110010111110", -- t[56510] = 22
      "0010110" when "01101110010111111", -- t[56511] = 22
      "0010110" when "01101110011000000", -- t[56512] = 22
      "0010110" when "01101110011000001", -- t[56513] = 22
      "0010110" when "01101110011000010", -- t[56514] = 22
      "0010110" when "01101110011000011", -- t[56515] = 22
      "0010110" when "01101110011000100", -- t[56516] = 22
      "0010110" when "01101110011000101", -- t[56517] = 22
      "0010110" when "01101110011000110", -- t[56518] = 22
      "0010110" when "01101110011000111", -- t[56519] = 22
      "0010110" when "01101110011001000", -- t[56520] = 22
      "0010110" when "01101110011001001", -- t[56521] = 22
      "0010110" when "01101110011001010", -- t[56522] = 22
      "0010110" when "01101110011001011", -- t[56523] = 22
      "0010110" when "01101110011001100", -- t[56524] = 22
      "0010110" when "01101110011001101", -- t[56525] = 22
      "0010110" when "01101110011001110", -- t[56526] = 22
      "0010110" when "01101110011001111", -- t[56527] = 22
      "0010110" when "01101110011010000", -- t[56528] = 22
      "0010110" when "01101110011010001", -- t[56529] = 22
      "0010110" when "01101110011010010", -- t[56530] = 22
      "0010110" when "01101110011010011", -- t[56531] = 22
      "0010110" when "01101110011010100", -- t[56532] = 22
      "0010110" when "01101110011010101", -- t[56533] = 22
      "0010110" when "01101110011010110", -- t[56534] = 22
      "0010110" when "01101110011010111", -- t[56535] = 22
      "0010110" when "01101110011011000", -- t[56536] = 22
      "0010110" when "01101110011011001", -- t[56537] = 22
      "0010110" when "01101110011011010", -- t[56538] = 22
      "0010110" when "01101110011011011", -- t[56539] = 22
      "0010110" when "01101110011011100", -- t[56540] = 22
      "0010110" when "01101110011011101", -- t[56541] = 22
      "0010110" when "01101110011011110", -- t[56542] = 22
      "0010110" when "01101110011011111", -- t[56543] = 22
      "0010110" when "01101110011100000", -- t[56544] = 22
      "0010110" when "01101110011100001", -- t[56545] = 22
      "0010110" when "01101110011100010", -- t[56546] = 22
      "0010110" when "01101110011100011", -- t[56547] = 22
      "0010110" when "01101110011100100", -- t[56548] = 22
      "0010110" when "01101110011100101", -- t[56549] = 22
      "0010110" when "01101110011100110", -- t[56550] = 22
      "0010110" when "01101110011100111", -- t[56551] = 22
      "0010110" when "01101110011101000", -- t[56552] = 22
      "0010110" when "01101110011101001", -- t[56553] = 22
      "0010110" when "01101110011101010", -- t[56554] = 22
      "0010110" when "01101110011101011", -- t[56555] = 22
      "0010110" when "01101110011101100", -- t[56556] = 22
      "0010110" when "01101110011101101", -- t[56557] = 22
      "0010110" when "01101110011101110", -- t[56558] = 22
      "0010110" when "01101110011101111", -- t[56559] = 22
      "0010110" when "01101110011110000", -- t[56560] = 22
      "0010110" when "01101110011110001", -- t[56561] = 22
      "0010110" when "01101110011110010", -- t[56562] = 22
      "0010110" when "01101110011110011", -- t[56563] = 22
      "0010110" when "01101110011110100", -- t[56564] = 22
      "0010110" when "01101110011110101", -- t[56565] = 22
      "0010110" when "01101110011110110", -- t[56566] = 22
      "0010110" when "01101110011110111", -- t[56567] = 22
      "0010110" when "01101110011111000", -- t[56568] = 22
      "0010110" when "01101110011111001", -- t[56569] = 22
      "0010110" when "01101110011111010", -- t[56570] = 22
      "0010110" when "01101110011111011", -- t[56571] = 22
      "0010110" when "01101110011111100", -- t[56572] = 22
      "0010110" when "01101110011111101", -- t[56573] = 22
      "0010110" when "01101110011111110", -- t[56574] = 22
      "0010110" when "01101110011111111", -- t[56575] = 22
      "0010110" when "01101110100000000", -- t[56576] = 22
      "0010110" when "01101110100000001", -- t[56577] = 22
      "0010110" when "01101110100000010", -- t[56578] = 22
      "0010110" when "01101110100000011", -- t[56579] = 22
      "0010110" when "01101110100000100", -- t[56580] = 22
      "0010110" when "01101110100000101", -- t[56581] = 22
      "0010110" when "01101110100000110", -- t[56582] = 22
      "0010110" when "01101110100000111", -- t[56583] = 22
      "0010110" when "01101110100001000", -- t[56584] = 22
      "0010110" when "01101110100001001", -- t[56585] = 22
      "0010110" when "01101110100001010", -- t[56586] = 22
      "0010110" when "01101110100001011", -- t[56587] = 22
      "0010110" when "01101110100001100", -- t[56588] = 22
      "0010110" when "01101110100001101", -- t[56589] = 22
      "0010110" when "01101110100001110", -- t[56590] = 22
      "0010110" when "01101110100001111", -- t[56591] = 22
      "0010110" when "01101110100010000", -- t[56592] = 22
      "0010110" when "01101110100010001", -- t[56593] = 22
      "0010110" when "01101110100010010", -- t[56594] = 22
      "0010110" when "01101110100010011", -- t[56595] = 22
      "0010110" when "01101110100010100", -- t[56596] = 22
      "0010110" when "01101110100010101", -- t[56597] = 22
      "0010110" when "01101110100010110", -- t[56598] = 22
      "0010110" when "01101110100010111", -- t[56599] = 22
      "0010110" when "01101110100011000", -- t[56600] = 22
      "0010110" when "01101110100011001", -- t[56601] = 22
      "0010110" when "01101110100011010", -- t[56602] = 22
      "0010110" when "01101110100011011", -- t[56603] = 22
      "0010110" when "01101110100011100", -- t[56604] = 22
      "0010110" when "01101110100011101", -- t[56605] = 22
      "0010110" when "01101110100011110", -- t[56606] = 22
      "0010110" when "01101110100011111", -- t[56607] = 22
      "0010110" when "01101110100100000", -- t[56608] = 22
      "0010110" when "01101110100100001", -- t[56609] = 22
      "0010110" when "01101110100100010", -- t[56610] = 22
      "0010110" when "01101110100100011", -- t[56611] = 22
      "0010110" when "01101110100100100", -- t[56612] = 22
      "0010110" when "01101110100100101", -- t[56613] = 22
      "0010110" when "01101110100100110", -- t[56614] = 22
      "0010110" when "01101110100100111", -- t[56615] = 22
      "0010110" when "01101110100101000", -- t[56616] = 22
      "0010110" when "01101110100101001", -- t[56617] = 22
      "0010110" when "01101110100101010", -- t[56618] = 22
      "0010110" when "01101110100101011", -- t[56619] = 22
      "0010110" when "01101110100101100", -- t[56620] = 22
      "0010110" when "01101110100101101", -- t[56621] = 22
      "0010110" when "01101110100101110", -- t[56622] = 22
      "0010110" when "01101110100101111", -- t[56623] = 22
      "0010110" when "01101110100110000", -- t[56624] = 22
      "0010110" when "01101110100110001", -- t[56625] = 22
      "0010110" when "01101110100110010", -- t[56626] = 22
      "0010110" when "01101110100110011", -- t[56627] = 22
      "0010110" when "01101110100110100", -- t[56628] = 22
      "0010110" when "01101110100110101", -- t[56629] = 22
      "0010110" when "01101110100110110", -- t[56630] = 22
      "0010110" when "01101110100110111", -- t[56631] = 22
      "0010110" when "01101110100111000", -- t[56632] = 22
      "0010110" when "01101110100111001", -- t[56633] = 22
      "0010110" when "01101110100111010", -- t[56634] = 22
      "0010110" when "01101110100111011", -- t[56635] = 22
      "0010110" when "01101110100111100", -- t[56636] = 22
      "0010110" when "01101110100111101", -- t[56637] = 22
      "0010110" when "01101110100111110", -- t[56638] = 22
      "0010110" when "01101110100111111", -- t[56639] = 22
      "0010110" when "01101110101000000", -- t[56640] = 22
      "0010110" when "01101110101000001", -- t[56641] = 22
      "0010110" when "01101110101000010", -- t[56642] = 22
      "0010110" when "01101110101000011", -- t[56643] = 22
      "0010110" when "01101110101000100", -- t[56644] = 22
      "0010110" when "01101110101000101", -- t[56645] = 22
      "0010110" when "01101110101000110", -- t[56646] = 22
      "0010110" when "01101110101000111", -- t[56647] = 22
      "0010110" when "01101110101001000", -- t[56648] = 22
      "0010110" when "01101110101001001", -- t[56649] = 22
      "0010110" when "01101110101001010", -- t[56650] = 22
      "0010110" when "01101110101001011", -- t[56651] = 22
      "0010110" when "01101110101001100", -- t[56652] = 22
      "0010110" when "01101110101001101", -- t[56653] = 22
      "0010110" when "01101110101001110", -- t[56654] = 22
      "0010110" when "01101110101001111", -- t[56655] = 22
      "0010110" when "01101110101010000", -- t[56656] = 22
      "0010110" when "01101110101010001", -- t[56657] = 22
      "0010110" when "01101110101010010", -- t[56658] = 22
      "0010110" when "01101110101010011", -- t[56659] = 22
      "0010110" when "01101110101010100", -- t[56660] = 22
      "0010110" when "01101110101010101", -- t[56661] = 22
      "0010110" when "01101110101010110", -- t[56662] = 22
      "0010110" when "01101110101010111", -- t[56663] = 22
      "0010110" when "01101110101011000", -- t[56664] = 22
      "0010110" when "01101110101011001", -- t[56665] = 22
      "0010110" when "01101110101011010", -- t[56666] = 22
      "0010110" when "01101110101011011", -- t[56667] = 22
      "0010110" when "01101110101011100", -- t[56668] = 22
      "0010110" when "01101110101011101", -- t[56669] = 22
      "0010110" when "01101110101011110", -- t[56670] = 22
      "0010110" when "01101110101011111", -- t[56671] = 22
      "0010110" when "01101110101100000", -- t[56672] = 22
      "0010110" when "01101110101100001", -- t[56673] = 22
      "0010110" when "01101110101100010", -- t[56674] = 22
      "0010110" when "01101110101100011", -- t[56675] = 22
      "0010110" when "01101110101100100", -- t[56676] = 22
      "0010110" when "01101110101100101", -- t[56677] = 22
      "0010110" when "01101110101100110", -- t[56678] = 22
      "0010110" when "01101110101100111", -- t[56679] = 22
      "0010110" when "01101110101101000", -- t[56680] = 22
      "0010110" when "01101110101101001", -- t[56681] = 22
      "0010110" when "01101110101101010", -- t[56682] = 22
      "0010110" when "01101110101101011", -- t[56683] = 22
      "0010110" when "01101110101101100", -- t[56684] = 22
      "0010110" when "01101110101101101", -- t[56685] = 22
      "0010110" when "01101110101101110", -- t[56686] = 22
      "0010110" when "01101110101101111", -- t[56687] = 22
      "0010110" when "01101110101110000", -- t[56688] = 22
      "0010110" when "01101110101110001", -- t[56689] = 22
      "0010110" when "01101110101110010", -- t[56690] = 22
      "0010110" when "01101110101110011", -- t[56691] = 22
      "0010110" when "01101110101110100", -- t[56692] = 22
      "0010110" when "01101110101110101", -- t[56693] = 22
      "0010110" when "01101110101110110", -- t[56694] = 22
      "0010110" when "01101110101110111", -- t[56695] = 22
      "0010110" when "01101110101111000", -- t[56696] = 22
      "0010110" when "01101110101111001", -- t[56697] = 22
      "0010110" when "01101110101111010", -- t[56698] = 22
      "0010110" when "01101110101111011", -- t[56699] = 22
      "0010110" when "01101110101111100", -- t[56700] = 22
      "0010110" when "01101110101111101", -- t[56701] = 22
      "0010110" when "01101110101111110", -- t[56702] = 22
      "0010110" when "01101110101111111", -- t[56703] = 22
      "0010110" when "01101110110000000", -- t[56704] = 22
      "0010110" when "01101110110000001", -- t[56705] = 22
      "0010110" when "01101110110000010", -- t[56706] = 22
      "0010110" when "01101110110000011", -- t[56707] = 22
      "0010110" when "01101110110000100", -- t[56708] = 22
      "0010110" when "01101110110000101", -- t[56709] = 22
      "0010110" when "01101110110000110", -- t[56710] = 22
      "0010110" when "01101110110000111", -- t[56711] = 22
      "0010110" when "01101110110001000", -- t[56712] = 22
      "0010110" when "01101110110001001", -- t[56713] = 22
      "0010110" when "01101110110001010", -- t[56714] = 22
      "0010110" when "01101110110001011", -- t[56715] = 22
      "0010110" when "01101110110001100", -- t[56716] = 22
      "0010110" when "01101110110001101", -- t[56717] = 22
      "0010110" when "01101110110001110", -- t[56718] = 22
      "0010110" when "01101110110001111", -- t[56719] = 22
      "0010110" when "01101110110010000", -- t[56720] = 22
      "0010110" when "01101110110010001", -- t[56721] = 22
      "0010110" when "01101110110010010", -- t[56722] = 22
      "0010110" when "01101110110010011", -- t[56723] = 22
      "0010110" when "01101110110010100", -- t[56724] = 22
      "0010110" when "01101110110010101", -- t[56725] = 22
      "0010110" when "01101110110010110", -- t[56726] = 22
      "0010110" when "01101110110010111", -- t[56727] = 22
      "0010110" when "01101110110011000", -- t[56728] = 22
      "0010110" when "01101110110011001", -- t[56729] = 22
      "0010110" when "01101110110011010", -- t[56730] = 22
      "0010110" when "01101110110011011", -- t[56731] = 22
      "0010110" when "01101110110011100", -- t[56732] = 22
      "0010110" when "01101110110011101", -- t[56733] = 22
      "0010110" when "01101110110011110", -- t[56734] = 22
      "0010110" when "01101110110011111", -- t[56735] = 22
      "0010110" when "01101110110100000", -- t[56736] = 22
      "0010110" when "01101110110100001", -- t[56737] = 22
      "0010110" when "01101110110100010", -- t[56738] = 22
      "0010110" when "01101110110100011", -- t[56739] = 22
      "0010110" when "01101110110100100", -- t[56740] = 22
      "0010110" when "01101110110100101", -- t[56741] = 22
      "0010110" when "01101110110100110", -- t[56742] = 22
      "0010110" when "01101110110100111", -- t[56743] = 22
      "0010110" when "01101110110101000", -- t[56744] = 22
      "0010110" when "01101110110101001", -- t[56745] = 22
      "0010110" when "01101110110101010", -- t[56746] = 22
      "0010110" when "01101110110101011", -- t[56747] = 22
      "0010110" when "01101110110101100", -- t[56748] = 22
      "0010110" when "01101110110101101", -- t[56749] = 22
      "0010110" when "01101110110101110", -- t[56750] = 22
      "0010110" when "01101110110101111", -- t[56751] = 22
      "0010110" when "01101110110110000", -- t[56752] = 22
      "0010110" when "01101110110110001", -- t[56753] = 22
      "0010110" when "01101110110110010", -- t[56754] = 22
      "0010110" when "01101110110110011", -- t[56755] = 22
      "0010110" when "01101110110110100", -- t[56756] = 22
      "0010110" when "01101110110110101", -- t[56757] = 22
      "0010110" when "01101110110110110", -- t[56758] = 22
      "0010110" when "01101110110110111", -- t[56759] = 22
      "0010110" when "01101110110111000", -- t[56760] = 22
      "0010110" when "01101110110111001", -- t[56761] = 22
      "0010110" when "01101110110111010", -- t[56762] = 22
      "0010110" when "01101110110111011", -- t[56763] = 22
      "0010110" when "01101110110111100", -- t[56764] = 22
      "0010110" when "01101110110111101", -- t[56765] = 22
      "0010110" when "01101110110111110", -- t[56766] = 22
      "0010110" when "01101110110111111", -- t[56767] = 22
      "0010110" when "01101110111000000", -- t[56768] = 22
      "0010110" when "01101110111000001", -- t[56769] = 22
      "0010110" when "01101110111000010", -- t[56770] = 22
      "0010110" when "01101110111000011", -- t[56771] = 22
      "0010110" when "01101110111000100", -- t[56772] = 22
      "0010110" when "01101110111000101", -- t[56773] = 22
      "0010110" when "01101110111000110", -- t[56774] = 22
      "0010110" when "01101110111000111", -- t[56775] = 22
      "0010110" when "01101110111001000", -- t[56776] = 22
      "0010110" when "01101110111001001", -- t[56777] = 22
      "0010110" when "01101110111001010", -- t[56778] = 22
      "0010110" when "01101110111001011", -- t[56779] = 22
      "0010110" when "01101110111001100", -- t[56780] = 22
      "0010110" when "01101110111001101", -- t[56781] = 22
      "0010110" when "01101110111001110", -- t[56782] = 22
      "0010110" when "01101110111001111", -- t[56783] = 22
      "0010110" when "01101110111010000", -- t[56784] = 22
      "0010110" when "01101110111010001", -- t[56785] = 22
      "0010110" when "01101110111010010", -- t[56786] = 22
      "0010110" when "01101110111010011", -- t[56787] = 22
      "0010110" when "01101110111010100", -- t[56788] = 22
      "0010110" when "01101110111010101", -- t[56789] = 22
      "0010110" when "01101110111010110", -- t[56790] = 22
      "0010110" when "01101110111010111", -- t[56791] = 22
      "0010110" when "01101110111011000", -- t[56792] = 22
      "0010110" when "01101110111011001", -- t[56793] = 22
      "0010110" when "01101110111011010", -- t[56794] = 22
      "0010110" when "01101110111011011", -- t[56795] = 22
      "0010110" when "01101110111011100", -- t[56796] = 22
      "0010110" when "01101110111011101", -- t[56797] = 22
      "0010110" when "01101110111011110", -- t[56798] = 22
      "0010110" when "01101110111011111", -- t[56799] = 22
      "0010110" when "01101110111100000", -- t[56800] = 22
      "0010110" when "01101110111100001", -- t[56801] = 22
      "0010110" when "01101110111100010", -- t[56802] = 22
      "0010110" when "01101110111100011", -- t[56803] = 22
      "0010110" when "01101110111100100", -- t[56804] = 22
      "0010110" when "01101110111100101", -- t[56805] = 22
      "0010110" when "01101110111100110", -- t[56806] = 22
      "0010110" when "01101110111100111", -- t[56807] = 22
      "0010110" when "01101110111101000", -- t[56808] = 22
      "0010110" when "01101110111101001", -- t[56809] = 22
      "0010110" when "01101110111101010", -- t[56810] = 22
      "0010110" when "01101110111101011", -- t[56811] = 22
      "0010110" when "01101110111101100", -- t[56812] = 22
      "0010110" when "01101110111101101", -- t[56813] = 22
      "0010110" when "01101110111101110", -- t[56814] = 22
      "0010110" when "01101110111101111", -- t[56815] = 22
      "0010110" when "01101110111110000", -- t[56816] = 22
      "0010110" when "01101110111110001", -- t[56817] = 22
      "0010110" when "01101110111110010", -- t[56818] = 22
      "0010110" when "01101110111110011", -- t[56819] = 22
      "0010110" when "01101110111110100", -- t[56820] = 22
      "0010110" when "01101110111110101", -- t[56821] = 22
      "0010110" when "01101110111110110", -- t[56822] = 22
      "0010110" when "01101110111110111", -- t[56823] = 22
      "0010110" when "01101110111111000", -- t[56824] = 22
      "0010110" when "01101110111111001", -- t[56825] = 22
      "0010110" when "01101110111111010", -- t[56826] = 22
      "0010110" when "01101110111111011", -- t[56827] = 22
      "0010110" when "01101110111111100", -- t[56828] = 22
      "0010110" when "01101110111111101", -- t[56829] = 22
      "0010110" when "01101110111111110", -- t[56830] = 22
      "0010110" when "01101110111111111", -- t[56831] = 22
      "0010110" when "01101111000000000", -- t[56832] = 22
      "0010110" when "01101111000000001", -- t[56833] = 22
      "0010110" when "01101111000000010", -- t[56834] = 22
      "0010110" when "01101111000000011", -- t[56835] = 22
      "0010110" when "01101111000000100", -- t[56836] = 22
      "0010110" when "01101111000000101", -- t[56837] = 22
      "0010110" when "01101111000000110", -- t[56838] = 22
      "0010110" when "01101111000000111", -- t[56839] = 22
      "0010110" when "01101111000001000", -- t[56840] = 22
      "0010110" when "01101111000001001", -- t[56841] = 22
      "0010110" when "01101111000001010", -- t[56842] = 22
      "0010110" when "01101111000001011", -- t[56843] = 22
      "0010110" when "01101111000001100", -- t[56844] = 22
      "0010110" when "01101111000001101", -- t[56845] = 22
      "0010110" when "01101111000001110", -- t[56846] = 22
      "0010110" when "01101111000001111", -- t[56847] = 22
      "0010110" when "01101111000010000", -- t[56848] = 22
      "0010110" when "01101111000010001", -- t[56849] = 22
      "0010110" when "01101111000010010", -- t[56850] = 22
      "0010110" when "01101111000010011", -- t[56851] = 22
      "0010110" when "01101111000010100", -- t[56852] = 22
      "0010110" when "01101111000010101", -- t[56853] = 22
      "0010110" when "01101111000010110", -- t[56854] = 22
      "0010110" when "01101111000010111", -- t[56855] = 22
      "0010110" when "01101111000011000", -- t[56856] = 22
      "0010110" when "01101111000011001", -- t[56857] = 22
      "0010110" when "01101111000011010", -- t[56858] = 22
      "0010110" when "01101111000011011", -- t[56859] = 22
      "0010110" when "01101111000011100", -- t[56860] = 22
      "0010110" when "01101111000011101", -- t[56861] = 22
      "0010110" when "01101111000011110", -- t[56862] = 22
      "0010110" when "01101111000011111", -- t[56863] = 22
      "0010110" when "01101111000100000", -- t[56864] = 22
      "0010110" when "01101111000100001", -- t[56865] = 22
      "0010110" when "01101111000100010", -- t[56866] = 22
      "0010110" when "01101111000100011", -- t[56867] = 22
      "0010110" when "01101111000100100", -- t[56868] = 22
      "0010110" when "01101111000100101", -- t[56869] = 22
      "0010110" when "01101111000100110", -- t[56870] = 22
      "0010110" when "01101111000100111", -- t[56871] = 22
      "0010110" when "01101111000101000", -- t[56872] = 22
      "0010110" when "01101111000101001", -- t[56873] = 22
      "0010110" when "01101111000101010", -- t[56874] = 22
      "0010110" when "01101111000101011", -- t[56875] = 22
      "0010110" when "01101111000101100", -- t[56876] = 22
      "0010110" when "01101111000101101", -- t[56877] = 22
      "0010110" when "01101111000101110", -- t[56878] = 22
      "0010110" when "01101111000101111", -- t[56879] = 22
      "0010110" when "01101111000110000", -- t[56880] = 22
      "0010110" when "01101111000110001", -- t[56881] = 22
      "0010110" when "01101111000110010", -- t[56882] = 22
      "0010110" when "01101111000110011", -- t[56883] = 22
      "0010110" when "01101111000110100", -- t[56884] = 22
      "0010110" when "01101111000110101", -- t[56885] = 22
      "0010110" when "01101111000110110", -- t[56886] = 22
      "0010110" when "01101111000110111", -- t[56887] = 22
      "0010110" when "01101111000111000", -- t[56888] = 22
      "0010110" when "01101111000111001", -- t[56889] = 22
      "0010110" when "01101111000111010", -- t[56890] = 22
      "0010110" when "01101111000111011", -- t[56891] = 22
      "0010110" when "01101111000111100", -- t[56892] = 22
      "0010110" when "01101111000111101", -- t[56893] = 22
      "0010110" when "01101111000111110", -- t[56894] = 22
      "0010110" when "01101111000111111", -- t[56895] = 22
      "0010110" when "01101111001000000", -- t[56896] = 22
      "0010110" when "01101111001000001", -- t[56897] = 22
      "0010110" when "01101111001000010", -- t[56898] = 22
      "0010110" when "01101111001000011", -- t[56899] = 22
      "0010110" when "01101111001000100", -- t[56900] = 22
      "0010110" when "01101111001000101", -- t[56901] = 22
      "0010110" when "01101111001000110", -- t[56902] = 22
      "0010110" when "01101111001000111", -- t[56903] = 22
      "0010110" when "01101111001001000", -- t[56904] = 22
      "0010110" when "01101111001001001", -- t[56905] = 22
      "0010110" when "01101111001001010", -- t[56906] = 22
      "0010110" when "01101111001001011", -- t[56907] = 22
      "0010110" when "01101111001001100", -- t[56908] = 22
      "0010110" when "01101111001001101", -- t[56909] = 22
      "0010110" when "01101111001001110", -- t[56910] = 22
      "0010110" when "01101111001001111", -- t[56911] = 22
      "0010110" when "01101111001010000", -- t[56912] = 22
      "0010110" when "01101111001010001", -- t[56913] = 22
      "0010110" when "01101111001010010", -- t[56914] = 22
      "0010110" when "01101111001010011", -- t[56915] = 22
      "0010110" when "01101111001010100", -- t[56916] = 22
      "0010110" when "01101111001010101", -- t[56917] = 22
      "0010110" when "01101111001010110", -- t[56918] = 22
      "0010110" when "01101111001010111", -- t[56919] = 22
      "0010110" when "01101111001011000", -- t[56920] = 22
      "0010110" when "01101111001011001", -- t[56921] = 22
      "0010110" when "01101111001011010", -- t[56922] = 22
      "0010110" when "01101111001011011", -- t[56923] = 22
      "0010110" when "01101111001011100", -- t[56924] = 22
      "0010110" when "01101111001011101", -- t[56925] = 22
      "0010110" when "01101111001011110", -- t[56926] = 22
      "0010110" when "01101111001011111", -- t[56927] = 22
      "0010110" when "01101111001100000", -- t[56928] = 22
      "0010110" when "01101111001100001", -- t[56929] = 22
      "0010110" when "01101111001100010", -- t[56930] = 22
      "0010110" when "01101111001100011", -- t[56931] = 22
      "0010110" when "01101111001100100", -- t[56932] = 22
      "0010110" when "01101111001100101", -- t[56933] = 22
      "0010110" when "01101111001100110", -- t[56934] = 22
      "0010110" when "01101111001100111", -- t[56935] = 22
      "0010110" when "01101111001101000", -- t[56936] = 22
      "0010110" when "01101111001101001", -- t[56937] = 22
      "0010110" when "01101111001101010", -- t[56938] = 22
      "0010110" when "01101111001101011", -- t[56939] = 22
      "0010110" when "01101111001101100", -- t[56940] = 22
      "0010110" when "01101111001101101", -- t[56941] = 22
      "0010110" when "01101111001101110", -- t[56942] = 22
      "0010110" when "01101111001101111", -- t[56943] = 22
      "0010110" when "01101111001110000", -- t[56944] = 22
      "0010110" when "01101111001110001", -- t[56945] = 22
      "0010110" when "01101111001110010", -- t[56946] = 22
      "0010110" when "01101111001110011", -- t[56947] = 22
      "0010110" when "01101111001110100", -- t[56948] = 22
      "0010110" when "01101111001110101", -- t[56949] = 22
      "0010110" when "01101111001110110", -- t[56950] = 22
      "0010110" when "01101111001110111", -- t[56951] = 22
      "0010110" when "01101111001111000", -- t[56952] = 22
      "0010110" when "01101111001111001", -- t[56953] = 22
      "0010110" when "01101111001111010", -- t[56954] = 22
      "0010110" when "01101111001111011", -- t[56955] = 22
      "0010110" when "01101111001111100", -- t[56956] = 22
      "0010110" when "01101111001111101", -- t[56957] = 22
      "0010110" when "01101111001111110", -- t[56958] = 22
      "0010110" when "01101111001111111", -- t[56959] = 22
      "0010110" when "01101111010000000", -- t[56960] = 22
      "0010110" when "01101111010000001", -- t[56961] = 22
      "0010110" when "01101111010000010", -- t[56962] = 22
      "0010110" when "01101111010000011", -- t[56963] = 22
      "0010110" when "01101111010000100", -- t[56964] = 22
      "0010110" when "01101111010000101", -- t[56965] = 22
      "0010110" when "01101111010000110", -- t[56966] = 22
      "0010110" when "01101111010000111", -- t[56967] = 22
      "0010110" when "01101111010001000", -- t[56968] = 22
      "0010110" when "01101111010001001", -- t[56969] = 22
      "0010110" when "01101111010001010", -- t[56970] = 22
      "0010110" when "01101111010001011", -- t[56971] = 22
      "0010110" when "01101111010001100", -- t[56972] = 22
      "0010110" when "01101111010001101", -- t[56973] = 22
      "0010110" when "01101111010001110", -- t[56974] = 22
      "0010110" when "01101111010001111", -- t[56975] = 22
      "0010110" when "01101111010010000", -- t[56976] = 22
      "0010110" when "01101111010010001", -- t[56977] = 22
      "0010110" when "01101111010010010", -- t[56978] = 22
      "0010110" when "01101111010010011", -- t[56979] = 22
      "0010110" when "01101111010010100", -- t[56980] = 22
      "0010110" when "01101111010010101", -- t[56981] = 22
      "0010110" when "01101111010010110", -- t[56982] = 22
      "0010110" when "01101111010010111", -- t[56983] = 22
      "0010110" when "01101111010011000", -- t[56984] = 22
      "0010110" when "01101111010011001", -- t[56985] = 22
      "0010110" when "01101111010011010", -- t[56986] = 22
      "0010110" when "01101111010011011", -- t[56987] = 22
      "0010110" when "01101111010011100", -- t[56988] = 22
      "0010110" when "01101111010011101", -- t[56989] = 22
      "0010110" when "01101111010011110", -- t[56990] = 22
      "0010110" when "01101111010011111", -- t[56991] = 22
      "0010110" when "01101111010100000", -- t[56992] = 22
      "0010110" when "01101111010100001", -- t[56993] = 22
      "0010110" when "01101111010100010", -- t[56994] = 22
      "0010110" when "01101111010100011", -- t[56995] = 22
      "0010110" when "01101111010100100", -- t[56996] = 22
      "0010110" when "01101111010100101", -- t[56997] = 22
      "0010110" when "01101111010100110", -- t[56998] = 22
      "0010110" when "01101111010100111", -- t[56999] = 22
      "0010110" when "01101111010101000", -- t[57000] = 22
      "0010110" when "01101111010101001", -- t[57001] = 22
      "0010110" when "01101111010101010", -- t[57002] = 22
      "0010110" when "01101111010101011", -- t[57003] = 22
      "0010110" when "01101111010101100", -- t[57004] = 22
      "0010110" when "01101111010101101", -- t[57005] = 22
      "0010110" when "01101111010101110", -- t[57006] = 22
      "0010110" when "01101111010101111", -- t[57007] = 22
      "0010110" when "01101111010110000", -- t[57008] = 22
      "0010110" when "01101111010110001", -- t[57009] = 22
      "0010110" when "01101111010110010", -- t[57010] = 22
      "0010110" when "01101111010110011", -- t[57011] = 22
      "0010110" when "01101111010110100", -- t[57012] = 22
      "0010110" when "01101111010110101", -- t[57013] = 22
      "0010110" when "01101111010110110", -- t[57014] = 22
      "0010110" when "01101111010110111", -- t[57015] = 22
      "0010110" when "01101111010111000", -- t[57016] = 22
      "0010110" when "01101111010111001", -- t[57017] = 22
      "0010110" when "01101111010111010", -- t[57018] = 22
      "0010110" when "01101111010111011", -- t[57019] = 22
      "0010110" when "01101111010111100", -- t[57020] = 22
      "0010110" when "01101111010111101", -- t[57021] = 22
      "0010110" when "01101111010111110", -- t[57022] = 22
      "0010110" when "01101111010111111", -- t[57023] = 22
      "0010110" when "01101111011000000", -- t[57024] = 22
      "0010110" when "01101111011000001", -- t[57025] = 22
      "0010110" when "01101111011000010", -- t[57026] = 22
      "0010110" when "01101111011000011", -- t[57027] = 22
      "0010110" when "01101111011000100", -- t[57028] = 22
      "0010110" when "01101111011000101", -- t[57029] = 22
      "0010110" when "01101111011000110", -- t[57030] = 22
      "0010111" when "01101111011000111", -- t[57031] = 23
      "0010111" when "01101111011001000", -- t[57032] = 23
      "0010111" when "01101111011001001", -- t[57033] = 23
      "0010111" when "01101111011001010", -- t[57034] = 23
      "0010111" when "01101111011001011", -- t[57035] = 23
      "0010111" when "01101111011001100", -- t[57036] = 23
      "0010111" when "01101111011001101", -- t[57037] = 23
      "0010111" when "01101111011001110", -- t[57038] = 23
      "0010111" when "01101111011001111", -- t[57039] = 23
      "0010111" when "01101111011010000", -- t[57040] = 23
      "0010111" when "01101111011010001", -- t[57041] = 23
      "0010111" when "01101111011010010", -- t[57042] = 23
      "0010111" when "01101111011010011", -- t[57043] = 23
      "0010111" when "01101111011010100", -- t[57044] = 23
      "0010111" when "01101111011010101", -- t[57045] = 23
      "0010111" when "01101111011010110", -- t[57046] = 23
      "0010111" when "01101111011010111", -- t[57047] = 23
      "0010111" when "01101111011011000", -- t[57048] = 23
      "0010111" when "01101111011011001", -- t[57049] = 23
      "0010111" when "01101111011011010", -- t[57050] = 23
      "0010111" when "01101111011011011", -- t[57051] = 23
      "0010111" when "01101111011011100", -- t[57052] = 23
      "0010111" when "01101111011011101", -- t[57053] = 23
      "0010111" when "01101111011011110", -- t[57054] = 23
      "0010111" when "01101111011011111", -- t[57055] = 23
      "0010111" when "01101111011100000", -- t[57056] = 23
      "0010111" when "01101111011100001", -- t[57057] = 23
      "0010111" when "01101111011100010", -- t[57058] = 23
      "0010111" when "01101111011100011", -- t[57059] = 23
      "0010111" when "01101111011100100", -- t[57060] = 23
      "0010111" when "01101111011100101", -- t[57061] = 23
      "0010111" when "01101111011100110", -- t[57062] = 23
      "0010111" when "01101111011100111", -- t[57063] = 23
      "0010111" when "01101111011101000", -- t[57064] = 23
      "0010111" when "01101111011101001", -- t[57065] = 23
      "0010111" when "01101111011101010", -- t[57066] = 23
      "0010111" when "01101111011101011", -- t[57067] = 23
      "0010111" when "01101111011101100", -- t[57068] = 23
      "0010111" when "01101111011101101", -- t[57069] = 23
      "0010111" when "01101111011101110", -- t[57070] = 23
      "0010111" when "01101111011101111", -- t[57071] = 23
      "0010111" when "01101111011110000", -- t[57072] = 23
      "0010111" when "01101111011110001", -- t[57073] = 23
      "0010111" when "01101111011110010", -- t[57074] = 23
      "0010111" when "01101111011110011", -- t[57075] = 23
      "0010111" when "01101111011110100", -- t[57076] = 23
      "0010111" when "01101111011110101", -- t[57077] = 23
      "0010111" when "01101111011110110", -- t[57078] = 23
      "0010111" when "01101111011110111", -- t[57079] = 23
      "0010111" when "01101111011111000", -- t[57080] = 23
      "0010111" when "01101111011111001", -- t[57081] = 23
      "0010111" when "01101111011111010", -- t[57082] = 23
      "0010111" when "01101111011111011", -- t[57083] = 23
      "0010111" when "01101111011111100", -- t[57084] = 23
      "0010111" when "01101111011111101", -- t[57085] = 23
      "0010111" when "01101111011111110", -- t[57086] = 23
      "0010111" when "01101111011111111", -- t[57087] = 23
      "0010111" when "01101111100000000", -- t[57088] = 23
      "0010111" when "01101111100000001", -- t[57089] = 23
      "0010111" when "01101111100000010", -- t[57090] = 23
      "0010111" when "01101111100000011", -- t[57091] = 23
      "0010111" when "01101111100000100", -- t[57092] = 23
      "0010111" when "01101111100000101", -- t[57093] = 23
      "0010111" when "01101111100000110", -- t[57094] = 23
      "0010111" when "01101111100000111", -- t[57095] = 23
      "0010111" when "01101111100001000", -- t[57096] = 23
      "0010111" when "01101111100001001", -- t[57097] = 23
      "0010111" when "01101111100001010", -- t[57098] = 23
      "0010111" when "01101111100001011", -- t[57099] = 23
      "0010111" when "01101111100001100", -- t[57100] = 23
      "0010111" when "01101111100001101", -- t[57101] = 23
      "0010111" when "01101111100001110", -- t[57102] = 23
      "0010111" when "01101111100001111", -- t[57103] = 23
      "0010111" when "01101111100010000", -- t[57104] = 23
      "0010111" when "01101111100010001", -- t[57105] = 23
      "0010111" when "01101111100010010", -- t[57106] = 23
      "0010111" when "01101111100010011", -- t[57107] = 23
      "0010111" when "01101111100010100", -- t[57108] = 23
      "0010111" when "01101111100010101", -- t[57109] = 23
      "0010111" when "01101111100010110", -- t[57110] = 23
      "0010111" when "01101111100010111", -- t[57111] = 23
      "0010111" when "01101111100011000", -- t[57112] = 23
      "0010111" when "01101111100011001", -- t[57113] = 23
      "0010111" when "01101111100011010", -- t[57114] = 23
      "0010111" when "01101111100011011", -- t[57115] = 23
      "0010111" when "01101111100011100", -- t[57116] = 23
      "0010111" when "01101111100011101", -- t[57117] = 23
      "0010111" when "01101111100011110", -- t[57118] = 23
      "0010111" when "01101111100011111", -- t[57119] = 23
      "0010111" when "01101111100100000", -- t[57120] = 23
      "0010111" when "01101111100100001", -- t[57121] = 23
      "0010111" when "01101111100100010", -- t[57122] = 23
      "0010111" when "01101111100100011", -- t[57123] = 23
      "0010111" when "01101111100100100", -- t[57124] = 23
      "0010111" when "01101111100100101", -- t[57125] = 23
      "0010111" when "01101111100100110", -- t[57126] = 23
      "0010111" when "01101111100100111", -- t[57127] = 23
      "0010111" when "01101111100101000", -- t[57128] = 23
      "0010111" when "01101111100101001", -- t[57129] = 23
      "0010111" when "01101111100101010", -- t[57130] = 23
      "0010111" when "01101111100101011", -- t[57131] = 23
      "0010111" when "01101111100101100", -- t[57132] = 23
      "0010111" when "01101111100101101", -- t[57133] = 23
      "0010111" when "01101111100101110", -- t[57134] = 23
      "0010111" when "01101111100101111", -- t[57135] = 23
      "0010111" when "01101111100110000", -- t[57136] = 23
      "0010111" when "01101111100110001", -- t[57137] = 23
      "0010111" when "01101111100110010", -- t[57138] = 23
      "0010111" when "01101111100110011", -- t[57139] = 23
      "0010111" when "01101111100110100", -- t[57140] = 23
      "0010111" when "01101111100110101", -- t[57141] = 23
      "0010111" when "01101111100110110", -- t[57142] = 23
      "0010111" when "01101111100110111", -- t[57143] = 23
      "0010111" when "01101111100111000", -- t[57144] = 23
      "0010111" when "01101111100111001", -- t[57145] = 23
      "0010111" when "01101111100111010", -- t[57146] = 23
      "0010111" when "01101111100111011", -- t[57147] = 23
      "0010111" when "01101111100111100", -- t[57148] = 23
      "0010111" when "01101111100111101", -- t[57149] = 23
      "0010111" when "01101111100111110", -- t[57150] = 23
      "0010111" when "01101111100111111", -- t[57151] = 23
      "0010111" when "01101111101000000", -- t[57152] = 23
      "0010111" when "01101111101000001", -- t[57153] = 23
      "0010111" when "01101111101000010", -- t[57154] = 23
      "0010111" when "01101111101000011", -- t[57155] = 23
      "0010111" when "01101111101000100", -- t[57156] = 23
      "0010111" when "01101111101000101", -- t[57157] = 23
      "0010111" when "01101111101000110", -- t[57158] = 23
      "0010111" when "01101111101000111", -- t[57159] = 23
      "0010111" when "01101111101001000", -- t[57160] = 23
      "0010111" when "01101111101001001", -- t[57161] = 23
      "0010111" when "01101111101001010", -- t[57162] = 23
      "0010111" when "01101111101001011", -- t[57163] = 23
      "0010111" when "01101111101001100", -- t[57164] = 23
      "0010111" when "01101111101001101", -- t[57165] = 23
      "0010111" when "01101111101001110", -- t[57166] = 23
      "0010111" when "01101111101001111", -- t[57167] = 23
      "0010111" when "01101111101010000", -- t[57168] = 23
      "0010111" when "01101111101010001", -- t[57169] = 23
      "0010111" when "01101111101010010", -- t[57170] = 23
      "0010111" when "01101111101010011", -- t[57171] = 23
      "0010111" when "01101111101010100", -- t[57172] = 23
      "0010111" when "01101111101010101", -- t[57173] = 23
      "0010111" when "01101111101010110", -- t[57174] = 23
      "0010111" when "01101111101010111", -- t[57175] = 23
      "0010111" when "01101111101011000", -- t[57176] = 23
      "0010111" when "01101111101011001", -- t[57177] = 23
      "0010111" when "01101111101011010", -- t[57178] = 23
      "0010111" when "01101111101011011", -- t[57179] = 23
      "0010111" when "01101111101011100", -- t[57180] = 23
      "0010111" when "01101111101011101", -- t[57181] = 23
      "0010111" when "01101111101011110", -- t[57182] = 23
      "0010111" when "01101111101011111", -- t[57183] = 23
      "0010111" when "01101111101100000", -- t[57184] = 23
      "0010111" when "01101111101100001", -- t[57185] = 23
      "0010111" when "01101111101100010", -- t[57186] = 23
      "0010111" when "01101111101100011", -- t[57187] = 23
      "0010111" when "01101111101100100", -- t[57188] = 23
      "0010111" when "01101111101100101", -- t[57189] = 23
      "0010111" when "01101111101100110", -- t[57190] = 23
      "0010111" when "01101111101100111", -- t[57191] = 23
      "0010111" when "01101111101101000", -- t[57192] = 23
      "0010111" when "01101111101101001", -- t[57193] = 23
      "0010111" when "01101111101101010", -- t[57194] = 23
      "0010111" when "01101111101101011", -- t[57195] = 23
      "0010111" when "01101111101101100", -- t[57196] = 23
      "0010111" when "01101111101101101", -- t[57197] = 23
      "0010111" when "01101111101101110", -- t[57198] = 23
      "0010111" when "01101111101101111", -- t[57199] = 23
      "0010111" when "01101111101110000", -- t[57200] = 23
      "0010111" when "01101111101110001", -- t[57201] = 23
      "0010111" when "01101111101110010", -- t[57202] = 23
      "0010111" when "01101111101110011", -- t[57203] = 23
      "0010111" when "01101111101110100", -- t[57204] = 23
      "0010111" when "01101111101110101", -- t[57205] = 23
      "0010111" when "01101111101110110", -- t[57206] = 23
      "0010111" when "01101111101110111", -- t[57207] = 23
      "0010111" when "01101111101111000", -- t[57208] = 23
      "0010111" when "01101111101111001", -- t[57209] = 23
      "0010111" when "01101111101111010", -- t[57210] = 23
      "0010111" when "01101111101111011", -- t[57211] = 23
      "0010111" when "01101111101111100", -- t[57212] = 23
      "0010111" when "01101111101111101", -- t[57213] = 23
      "0010111" when "01101111101111110", -- t[57214] = 23
      "0010111" when "01101111101111111", -- t[57215] = 23
      "0010111" when "01101111110000000", -- t[57216] = 23
      "0010111" when "01101111110000001", -- t[57217] = 23
      "0010111" when "01101111110000010", -- t[57218] = 23
      "0010111" when "01101111110000011", -- t[57219] = 23
      "0010111" when "01101111110000100", -- t[57220] = 23
      "0010111" when "01101111110000101", -- t[57221] = 23
      "0010111" when "01101111110000110", -- t[57222] = 23
      "0010111" when "01101111110000111", -- t[57223] = 23
      "0010111" when "01101111110001000", -- t[57224] = 23
      "0010111" when "01101111110001001", -- t[57225] = 23
      "0010111" when "01101111110001010", -- t[57226] = 23
      "0010111" when "01101111110001011", -- t[57227] = 23
      "0010111" when "01101111110001100", -- t[57228] = 23
      "0010111" when "01101111110001101", -- t[57229] = 23
      "0010111" when "01101111110001110", -- t[57230] = 23
      "0010111" when "01101111110001111", -- t[57231] = 23
      "0010111" when "01101111110010000", -- t[57232] = 23
      "0010111" when "01101111110010001", -- t[57233] = 23
      "0010111" when "01101111110010010", -- t[57234] = 23
      "0010111" when "01101111110010011", -- t[57235] = 23
      "0010111" when "01101111110010100", -- t[57236] = 23
      "0010111" when "01101111110010101", -- t[57237] = 23
      "0010111" when "01101111110010110", -- t[57238] = 23
      "0010111" when "01101111110010111", -- t[57239] = 23
      "0010111" when "01101111110011000", -- t[57240] = 23
      "0010111" when "01101111110011001", -- t[57241] = 23
      "0010111" when "01101111110011010", -- t[57242] = 23
      "0010111" when "01101111110011011", -- t[57243] = 23
      "0010111" when "01101111110011100", -- t[57244] = 23
      "0010111" when "01101111110011101", -- t[57245] = 23
      "0010111" when "01101111110011110", -- t[57246] = 23
      "0010111" when "01101111110011111", -- t[57247] = 23
      "0010111" when "01101111110100000", -- t[57248] = 23
      "0010111" when "01101111110100001", -- t[57249] = 23
      "0010111" when "01101111110100010", -- t[57250] = 23
      "0010111" when "01101111110100011", -- t[57251] = 23
      "0010111" when "01101111110100100", -- t[57252] = 23
      "0010111" when "01101111110100101", -- t[57253] = 23
      "0010111" when "01101111110100110", -- t[57254] = 23
      "0010111" when "01101111110100111", -- t[57255] = 23
      "0010111" when "01101111110101000", -- t[57256] = 23
      "0010111" when "01101111110101001", -- t[57257] = 23
      "0010111" when "01101111110101010", -- t[57258] = 23
      "0010111" when "01101111110101011", -- t[57259] = 23
      "0010111" when "01101111110101100", -- t[57260] = 23
      "0010111" when "01101111110101101", -- t[57261] = 23
      "0010111" when "01101111110101110", -- t[57262] = 23
      "0010111" when "01101111110101111", -- t[57263] = 23
      "0010111" when "01101111110110000", -- t[57264] = 23
      "0010111" when "01101111110110001", -- t[57265] = 23
      "0010111" when "01101111110110010", -- t[57266] = 23
      "0010111" when "01101111110110011", -- t[57267] = 23
      "0010111" when "01101111110110100", -- t[57268] = 23
      "0010111" when "01101111110110101", -- t[57269] = 23
      "0010111" when "01101111110110110", -- t[57270] = 23
      "0010111" when "01101111110110111", -- t[57271] = 23
      "0010111" when "01101111110111000", -- t[57272] = 23
      "0010111" when "01101111110111001", -- t[57273] = 23
      "0010111" when "01101111110111010", -- t[57274] = 23
      "0010111" when "01101111110111011", -- t[57275] = 23
      "0010111" when "01101111110111100", -- t[57276] = 23
      "0010111" when "01101111110111101", -- t[57277] = 23
      "0010111" when "01101111110111110", -- t[57278] = 23
      "0010111" when "01101111110111111", -- t[57279] = 23
      "0010111" when "01101111111000000", -- t[57280] = 23
      "0010111" when "01101111111000001", -- t[57281] = 23
      "0010111" when "01101111111000010", -- t[57282] = 23
      "0010111" when "01101111111000011", -- t[57283] = 23
      "0010111" when "01101111111000100", -- t[57284] = 23
      "0010111" when "01101111111000101", -- t[57285] = 23
      "0010111" when "01101111111000110", -- t[57286] = 23
      "0010111" when "01101111111000111", -- t[57287] = 23
      "0010111" when "01101111111001000", -- t[57288] = 23
      "0010111" when "01101111111001001", -- t[57289] = 23
      "0010111" when "01101111111001010", -- t[57290] = 23
      "0010111" when "01101111111001011", -- t[57291] = 23
      "0010111" when "01101111111001100", -- t[57292] = 23
      "0010111" when "01101111111001101", -- t[57293] = 23
      "0010111" when "01101111111001110", -- t[57294] = 23
      "0010111" when "01101111111001111", -- t[57295] = 23
      "0010111" when "01101111111010000", -- t[57296] = 23
      "0010111" when "01101111111010001", -- t[57297] = 23
      "0010111" when "01101111111010010", -- t[57298] = 23
      "0010111" when "01101111111010011", -- t[57299] = 23
      "0010111" when "01101111111010100", -- t[57300] = 23
      "0010111" when "01101111111010101", -- t[57301] = 23
      "0010111" when "01101111111010110", -- t[57302] = 23
      "0010111" when "01101111111010111", -- t[57303] = 23
      "0010111" when "01101111111011000", -- t[57304] = 23
      "0010111" when "01101111111011001", -- t[57305] = 23
      "0010111" when "01101111111011010", -- t[57306] = 23
      "0010111" when "01101111111011011", -- t[57307] = 23
      "0010111" when "01101111111011100", -- t[57308] = 23
      "0010111" when "01101111111011101", -- t[57309] = 23
      "0010111" when "01101111111011110", -- t[57310] = 23
      "0010111" when "01101111111011111", -- t[57311] = 23
      "0010111" when "01101111111100000", -- t[57312] = 23
      "0010111" when "01101111111100001", -- t[57313] = 23
      "0010111" when "01101111111100010", -- t[57314] = 23
      "0010111" when "01101111111100011", -- t[57315] = 23
      "0010111" when "01101111111100100", -- t[57316] = 23
      "0010111" when "01101111111100101", -- t[57317] = 23
      "0010111" when "01101111111100110", -- t[57318] = 23
      "0010111" when "01101111111100111", -- t[57319] = 23
      "0010111" when "01101111111101000", -- t[57320] = 23
      "0010111" when "01101111111101001", -- t[57321] = 23
      "0010111" when "01101111111101010", -- t[57322] = 23
      "0010111" when "01101111111101011", -- t[57323] = 23
      "0010111" when "01101111111101100", -- t[57324] = 23
      "0010111" when "01101111111101101", -- t[57325] = 23
      "0010111" when "01101111111101110", -- t[57326] = 23
      "0010111" when "01101111111101111", -- t[57327] = 23
      "0010111" when "01101111111110000", -- t[57328] = 23
      "0010111" when "01101111111110001", -- t[57329] = 23
      "0010111" when "01101111111110010", -- t[57330] = 23
      "0010111" when "01101111111110011", -- t[57331] = 23
      "0010111" when "01101111111110100", -- t[57332] = 23
      "0010111" when "01101111111110101", -- t[57333] = 23
      "0010111" when "01101111111110110", -- t[57334] = 23
      "0010111" when "01101111111110111", -- t[57335] = 23
      "0010111" when "01101111111111000", -- t[57336] = 23
      "0010111" when "01101111111111001", -- t[57337] = 23
      "0010111" when "01101111111111010", -- t[57338] = 23
      "0010111" when "01101111111111011", -- t[57339] = 23
      "0010111" when "01101111111111100", -- t[57340] = 23
      "0010111" when "01101111111111101", -- t[57341] = 23
      "0010111" when "01101111111111110", -- t[57342] = 23
      "0010111" when "01101111111111111", -- t[57343] = 23
      "0010111" when "01110000000000000", -- t[57344] = 23
      "0010111" when "01110000000000001", -- t[57345] = 23
      "0010111" when "01110000000000010", -- t[57346] = 23
      "0010111" when "01110000000000011", -- t[57347] = 23
      "0010111" when "01110000000000100", -- t[57348] = 23
      "0010111" when "01110000000000101", -- t[57349] = 23
      "0010111" when "01110000000000110", -- t[57350] = 23
      "0010111" when "01110000000000111", -- t[57351] = 23
      "0010111" when "01110000000001000", -- t[57352] = 23
      "0010111" when "01110000000001001", -- t[57353] = 23
      "0010111" when "01110000000001010", -- t[57354] = 23
      "0010111" when "01110000000001011", -- t[57355] = 23
      "0010111" when "01110000000001100", -- t[57356] = 23
      "0010111" when "01110000000001101", -- t[57357] = 23
      "0010111" when "01110000000001110", -- t[57358] = 23
      "0010111" when "01110000000001111", -- t[57359] = 23
      "0010111" when "01110000000010000", -- t[57360] = 23
      "0010111" when "01110000000010001", -- t[57361] = 23
      "0010111" when "01110000000010010", -- t[57362] = 23
      "0010111" when "01110000000010011", -- t[57363] = 23
      "0010111" when "01110000000010100", -- t[57364] = 23
      "0010111" when "01110000000010101", -- t[57365] = 23
      "0010111" when "01110000000010110", -- t[57366] = 23
      "0010111" when "01110000000010111", -- t[57367] = 23
      "0010111" when "01110000000011000", -- t[57368] = 23
      "0010111" when "01110000000011001", -- t[57369] = 23
      "0010111" when "01110000000011010", -- t[57370] = 23
      "0010111" when "01110000000011011", -- t[57371] = 23
      "0010111" when "01110000000011100", -- t[57372] = 23
      "0010111" when "01110000000011101", -- t[57373] = 23
      "0010111" when "01110000000011110", -- t[57374] = 23
      "0010111" when "01110000000011111", -- t[57375] = 23
      "0010111" when "01110000000100000", -- t[57376] = 23
      "0010111" when "01110000000100001", -- t[57377] = 23
      "0010111" when "01110000000100010", -- t[57378] = 23
      "0010111" when "01110000000100011", -- t[57379] = 23
      "0010111" when "01110000000100100", -- t[57380] = 23
      "0010111" when "01110000000100101", -- t[57381] = 23
      "0010111" when "01110000000100110", -- t[57382] = 23
      "0010111" when "01110000000100111", -- t[57383] = 23
      "0010111" when "01110000000101000", -- t[57384] = 23
      "0010111" when "01110000000101001", -- t[57385] = 23
      "0010111" when "01110000000101010", -- t[57386] = 23
      "0010111" when "01110000000101011", -- t[57387] = 23
      "0010111" when "01110000000101100", -- t[57388] = 23
      "0010111" when "01110000000101101", -- t[57389] = 23
      "0010111" when "01110000000101110", -- t[57390] = 23
      "0010111" when "01110000000101111", -- t[57391] = 23
      "0010111" when "01110000000110000", -- t[57392] = 23
      "0010111" when "01110000000110001", -- t[57393] = 23
      "0010111" when "01110000000110010", -- t[57394] = 23
      "0010111" when "01110000000110011", -- t[57395] = 23
      "0010111" when "01110000000110100", -- t[57396] = 23
      "0010111" when "01110000000110101", -- t[57397] = 23
      "0010111" when "01110000000110110", -- t[57398] = 23
      "0010111" when "01110000000110111", -- t[57399] = 23
      "0010111" when "01110000000111000", -- t[57400] = 23
      "0010111" when "01110000000111001", -- t[57401] = 23
      "0010111" when "01110000000111010", -- t[57402] = 23
      "0010111" when "01110000000111011", -- t[57403] = 23
      "0010111" when "01110000000111100", -- t[57404] = 23
      "0010111" when "01110000000111101", -- t[57405] = 23
      "0010111" when "01110000000111110", -- t[57406] = 23
      "0010111" when "01110000000111111", -- t[57407] = 23
      "0010111" when "01110000001000000", -- t[57408] = 23
      "0010111" when "01110000001000001", -- t[57409] = 23
      "0010111" when "01110000001000010", -- t[57410] = 23
      "0010111" when "01110000001000011", -- t[57411] = 23
      "0010111" when "01110000001000100", -- t[57412] = 23
      "0010111" when "01110000001000101", -- t[57413] = 23
      "0010111" when "01110000001000110", -- t[57414] = 23
      "0010111" when "01110000001000111", -- t[57415] = 23
      "0010111" when "01110000001001000", -- t[57416] = 23
      "0010111" when "01110000001001001", -- t[57417] = 23
      "0010111" when "01110000001001010", -- t[57418] = 23
      "0010111" when "01110000001001011", -- t[57419] = 23
      "0010111" when "01110000001001100", -- t[57420] = 23
      "0010111" when "01110000001001101", -- t[57421] = 23
      "0010111" when "01110000001001110", -- t[57422] = 23
      "0010111" when "01110000001001111", -- t[57423] = 23
      "0010111" when "01110000001010000", -- t[57424] = 23
      "0010111" when "01110000001010001", -- t[57425] = 23
      "0010111" when "01110000001010010", -- t[57426] = 23
      "0010111" when "01110000001010011", -- t[57427] = 23
      "0010111" when "01110000001010100", -- t[57428] = 23
      "0010111" when "01110000001010101", -- t[57429] = 23
      "0010111" when "01110000001010110", -- t[57430] = 23
      "0010111" when "01110000001010111", -- t[57431] = 23
      "0010111" when "01110000001011000", -- t[57432] = 23
      "0010111" when "01110000001011001", -- t[57433] = 23
      "0010111" when "01110000001011010", -- t[57434] = 23
      "0010111" when "01110000001011011", -- t[57435] = 23
      "0010111" when "01110000001011100", -- t[57436] = 23
      "0010111" when "01110000001011101", -- t[57437] = 23
      "0010111" when "01110000001011110", -- t[57438] = 23
      "0010111" when "01110000001011111", -- t[57439] = 23
      "0010111" when "01110000001100000", -- t[57440] = 23
      "0010111" when "01110000001100001", -- t[57441] = 23
      "0010111" when "01110000001100010", -- t[57442] = 23
      "0010111" when "01110000001100011", -- t[57443] = 23
      "0010111" when "01110000001100100", -- t[57444] = 23
      "0010111" when "01110000001100101", -- t[57445] = 23
      "0010111" when "01110000001100110", -- t[57446] = 23
      "0010111" when "01110000001100111", -- t[57447] = 23
      "0010111" when "01110000001101000", -- t[57448] = 23
      "0010111" when "01110000001101001", -- t[57449] = 23
      "0010111" when "01110000001101010", -- t[57450] = 23
      "0010111" when "01110000001101011", -- t[57451] = 23
      "0010111" when "01110000001101100", -- t[57452] = 23
      "0010111" when "01110000001101101", -- t[57453] = 23
      "0010111" when "01110000001101110", -- t[57454] = 23
      "0010111" when "01110000001101111", -- t[57455] = 23
      "0010111" when "01110000001110000", -- t[57456] = 23
      "0010111" when "01110000001110001", -- t[57457] = 23
      "0010111" when "01110000001110010", -- t[57458] = 23
      "0010111" when "01110000001110011", -- t[57459] = 23
      "0010111" when "01110000001110100", -- t[57460] = 23
      "0010111" when "01110000001110101", -- t[57461] = 23
      "0010111" when "01110000001110110", -- t[57462] = 23
      "0010111" when "01110000001110111", -- t[57463] = 23
      "0010111" when "01110000001111000", -- t[57464] = 23
      "0010111" when "01110000001111001", -- t[57465] = 23
      "0010111" when "01110000001111010", -- t[57466] = 23
      "0010111" when "01110000001111011", -- t[57467] = 23
      "0010111" when "01110000001111100", -- t[57468] = 23
      "0010111" when "01110000001111101", -- t[57469] = 23
      "0010111" when "01110000001111110", -- t[57470] = 23
      "0010111" when "01110000001111111", -- t[57471] = 23
      "0010111" when "01110000010000000", -- t[57472] = 23
      "0010111" when "01110000010000001", -- t[57473] = 23
      "0010111" when "01110000010000010", -- t[57474] = 23
      "0010111" when "01110000010000011", -- t[57475] = 23
      "0010111" when "01110000010000100", -- t[57476] = 23
      "0010111" when "01110000010000101", -- t[57477] = 23
      "0010111" when "01110000010000110", -- t[57478] = 23
      "0010111" when "01110000010000111", -- t[57479] = 23
      "0010111" when "01110000010001000", -- t[57480] = 23
      "0010111" when "01110000010001001", -- t[57481] = 23
      "0010111" when "01110000010001010", -- t[57482] = 23
      "0010111" when "01110000010001011", -- t[57483] = 23
      "0010111" when "01110000010001100", -- t[57484] = 23
      "0010111" when "01110000010001101", -- t[57485] = 23
      "0010111" when "01110000010001110", -- t[57486] = 23
      "0010111" when "01110000010001111", -- t[57487] = 23
      "0010111" when "01110000010010000", -- t[57488] = 23
      "0010111" when "01110000010010001", -- t[57489] = 23
      "0010111" when "01110000010010010", -- t[57490] = 23
      "0010111" when "01110000010010011", -- t[57491] = 23
      "0010111" when "01110000010010100", -- t[57492] = 23
      "0010111" when "01110000010010101", -- t[57493] = 23
      "0010111" when "01110000010010110", -- t[57494] = 23
      "0010111" when "01110000010010111", -- t[57495] = 23
      "0010111" when "01110000010011000", -- t[57496] = 23
      "0010111" when "01110000010011001", -- t[57497] = 23
      "0010111" when "01110000010011010", -- t[57498] = 23
      "0010111" when "01110000010011011", -- t[57499] = 23
      "0010111" when "01110000010011100", -- t[57500] = 23
      "0010111" when "01110000010011101", -- t[57501] = 23
      "0010111" when "01110000010011110", -- t[57502] = 23
      "0010111" when "01110000010011111", -- t[57503] = 23
      "0010111" when "01110000010100000", -- t[57504] = 23
      "0010111" when "01110000010100001", -- t[57505] = 23
      "0010111" when "01110000010100010", -- t[57506] = 23
      "0010111" when "01110000010100011", -- t[57507] = 23
      "0010111" when "01110000010100100", -- t[57508] = 23
      "0010111" when "01110000010100101", -- t[57509] = 23
      "0010111" when "01110000010100110", -- t[57510] = 23
      "0010111" when "01110000010100111", -- t[57511] = 23
      "0010111" when "01110000010101000", -- t[57512] = 23
      "0010111" when "01110000010101001", -- t[57513] = 23
      "0010111" when "01110000010101010", -- t[57514] = 23
      "0010111" when "01110000010101011", -- t[57515] = 23
      "0010111" when "01110000010101100", -- t[57516] = 23
      "0010111" when "01110000010101101", -- t[57517] = 23
      "0010111" when "01110000010101110", -- t[57518] = 23
      "0010111" when "01110000010101111", -- t[57519] = 23
      "0010111" when "01110000010110000", -- t[57520] = 23
      "0010111" when "01110000010110001", -- t[57521] = 23
      "0010111" when "01110000010110010", -- t[57522] = 23
      "0010111" when "01110000010110011", -- t[57523] = 23
      "0010111" when "01110000010110100", -- t[57524] = 23
      "0010111" when "01110000010110101", -- t[57525] = 23
      "0010111" when "01110000010110110", -- t[57526] = 23
      "0010111" when "01110000010110111", -- t[57527] = 23
      "0010111" when "01110000010111000", -- t[57528] = 23
      "0010111" when "01110000010111001", -- t[57529] = 23
      "0010111" when "01110000010111010", -- t[57530] = 23
      "0010111" when "01110000010111011", -- t[57531] = 23
      "0010111" when "01110000010111100", -- t[57532] = 23
      "0010111" when "01110000010111101", -- t[57533] = 23
      "0010111" when "01110000010111110", -- t[57534] = 23
      "0010111" when "01110000010111111", -- t[57535] = 23
      "0010111" when "01110000011000000", -- t[57536] = 23
      "0010111" when "01110000011000001", -- t[57537] = 23
      "0010111" when "01110000011000010", -- t[57538] = 23
      "0010111" when "01110000011000011", -- t[57539] = 23
      "0010111" when "01110000011000100", -- t[57540] = 23
      "0010111" when "01110000011000101", -- t[57541] = 23
      "0010111" when "01110000011000110", -- t[57542] = 23
      "0010111" when "01110000011000111", -- t[57543] = 23
      "0011000" when "01110000011001000", -- t[57544] = 24
      "0011000" when "01110000011001001", -- t[57545] = 24
      "0011000" when "01110000011001010", -- t[57546] = 24
      "0011000" when "01110000011001011", -- t[57547] = 24
      "0011000" when "01110000011001100", -- t[57548] = 24
      "0011000" when "01110000011001101", -- t[57549] = 24
      "0011000" when "01110000011001110", -- t[57550] = 24
      "0011000" when "01110000011001111", -- t[57551] = 24
      "0011000" when "01110000011010000", -- t[57552] = 24
      "0011000" when "01110000011010001", -- t[57553] = 24
      "0011000" when "01110000011010010", -- t[57554] = 24
      "0011000" when "01110000011010011", -- t[57555] = 24
      "0011000" when "01110000011010100", -- t[57556] = 24
      "0011000" when "01110000011010101", -- t[57557] = 24
      "0011000" when "01110000011010110", -- t[57558] = 24
      "0011000" when "01110000011010111", -- t[57559] = 24
      "0011000" when "01110000011011000", -- t[57560] = 24
      "0011000" when "01110000011011001", -- t[57561] = 24
      "0011000" when "01110000011011010", -- t[57562] = 24
      "0011000" when "01110000011011011", -- t[57563] = 24
      "0011000" when "01110000011011100", -- t[57564] = 24
      "0011000" when "01110000011011101", -- t[57565] = 24
      "0011000" when "01110000011011110", -- t[57566] = 24
      "0011000" when "01110000011011111", -- t[57567] = 24
      "0011000" when "01110000011100000", -- t[57568] = 24
      "0011000" when "01110000011100001", -- t[57569] = 24
      "0011000" when "01110000011100010", -- t[57570] = 24
      "0011000" when "01110000011100011", -- t[57571] = 24
      "0011000" when "01110000011100100", -- t[57572] = 24
      "0011000" when "01110000011100101", -- t[57573] = 24
      "0011000" when "01110000011100110", -- t[57574] = 24
      "0011000" when "01110000011100111", -- t[57575] = 24
      "0011000" when "01110000011101000", -- t[57576] = 24
      "0011000" when "01110000011101001", -- t[57577] = 24
      "0011000" when "01110000011101010", -- t[57578] = 24
      "0011000" when "01110000011101011", -- t[57579] = 24
      "0011000" when "01110000011101100", -- t[57580] = 24
      "0011000" when "01110000011101101", -- t[57581] = 24
      "0011000" when "01110000011101110", -- t[57582] = 24
      "0011000" when "01110000011101111", -- t[57583] = 24
      "0011000" when "01110000011110000", -- t[57584] = 24
      "0011000" when "01110000011110001", -- t[57585] = 24
      "0011000" when "01110000011110010", -- t[57586] = 24
      "0011000" when "01110000011110011", -- t[57587] = 24
      "0011000" when "01110000011110100", -- t[57588] = 24
      "0011000" when "01110000011110101", -- t[57589] = 24
      "0011000" when "01110000011110110", -- t[57590] = 24
      "0011000" when "01110000011110111", -- t[57591] = 24
      "0011000" when "01110000011111000", -- t[57592] = 24
      "0011000" when "01110000011111001", -- t[57593] = 24
      "0011000" when "01110000011111010", -- t[57594] = 24
      "0011000" when "01110000011111011", -- t[57595] = 24
      "0011000" when "01110000011111100", -- t[57596] = 24
      "0011000" when "01110000011111101", -- t[57597] = 24
      "0011000" when "01110000011111110", -- t[57598] = 24
      "0011000" when "01110000011111111", -- t[57599] = 24
      "0011000" when "01110000100000000", -- t[57600] = 24
      "0011000" when "01110000100000001", -- t[57601] = 24
      "0011000" when "01110000100000010", -- t[57602] = 24
      "0011000" when "01110000100000011", -- t[57603] = 24
      "0011000" when "01110000100000100", -- t[57604] = 24
      "0011000" when "01110000100000101", -- t[57605] = 24
      "0011000" when "01110000100000110", -- t[57606] = 24
      "0011000" when "01110000100000111", -- t[57607] = 24
      "0011000" when "01110000100001000", -- t[57608] = 24
      "0011000" when "01110000100001001", -- t[57609] = 24
      "0011000" when "01110000100001010", -- t[57610] = 24
      "0011000" when "01110000100001011", -- t[57611] = 24
      "0011000" when "01110000100001100", -- t[57612] = 24
      "0011000" when "01110000100001101", -- t[57613] = 24
      "0011000" when "01110000100001110", -- t[57614] = 24
      "0011000" when "01110000100001111", -- t[57615] = 24
      "0011000" when "01110000100010000", -- t[57616] = 24
      "0011000" when "01110000100010001", -- t[57617] = 24
      "0011000" when "01110000100010010", -- t[57618] = 24
      "0011000" when "01110000100010011", -- t[57619] = 24
      "0011000" when "01110000100010100", -- t[57620] = 24
      "0011000" when "01110000100010101", -- t[57621] = 24
      "0011000" when "01110000100010110", -- t[57622] = 24
      "0011000" when "01110000100010111", -- t[57623] = 24
      "0011000" when "01110000100011000", -- t[57624] = 24
      "0011000" when "01110000100011001", -- t[57625] = 24
      "0011000" when "01110000100011010", -- t[57626] = 24
      "0011000" when "01110000100011011", -- t[57627] = 24
      "0011000" when "01110000100011100", -- t[57628] = 24
      "0011000" when "01110000100011101", -- t[57629] = 24
      "0011000" when "01110000100011110", -- t[57630] = 24
      "0011000" when "01110000100011111", -- t[57631] = 24
      "0011000" when "01110000100100000", -- t[57632] = 24
      "0011000" when "01110000100100001", -- t[57633] = 24
      "0011000" when "01110000100100010", -- t[57634] = 24
      "0011000" when "01110000100100011", -- t[57635] = 24
      "0011000" when "01110000100100100", -- t[57636] = 24
      "0011000" when "01110000100100101", -- t[57637] = 24
      "0011000" when "01110000100100110", -- t[57638] = 24
      "0011000" when "01110000100100111", -- t[57639] = 24
      "0011000" when "01110000100101000", -- t[57640] = 24
      "0011000" when "01110000100101001", -- t[57641] = 24
      "0011000" when "01110000100101010", -- t[57642] = 24
      "0011000" when "01110000100101011", -- t[57643] = 24
      "0011000" when "01110000100101100", -- t[57644] = 24
      "0011000" when "01110000100101101", -- t[57645] = 24
      "0011000" when "01110000100101110", -- t[57646] = 24
      "0011000" when "01110000100101111", -- t[57647] = 24
      "0011000" when "01110000100110000", -- t[57648] = 24
      "0011000" when "01110000100110001", -- t[57649] = 24
      "0011000" when "01110000100110010", -- t[57650] = 24
      "0011000" when "01110000100110011", -- t[57651] = 24
      "0011000" when "01110000100110100", -- t[57652] = 24
      "0011000" when "01110000100110101", -- t[57653] = 24
      "0011000" when "01110000100110110", -- t[57654] = 24
      "0011000" when "01110000100110111", -- t[57655] = 24
      "0011000" when "01110000100111000", -- t[57656] = 24
      "0011000" when "01110000100111001", -- t[57657] = 24
      "0011000" when "01110000100111010", -- t[57658] = 24
      "0011000" when "01110000100111011", -- t[57659] = 24
      "0011000" when "01110000100111100", -- t[57660] = 24
      "0011000" when "01110000100111101", -- t[57661] = 24
      "0011000" when "01110000100111110", -- t[57662] = 24
      "0011000" when "01110000100111111", -- t[57663] = 24
      "0011000" when "01110000101000000", -- t[57664] = 24
      "0011000" when "01110000101000001", -- t[57665] = 24
      "0011000" when "01110000101000010", -- t[57666] = 24
      "0011000" when "01110000101000011", -- t[57667] = 24
      "0011000" when "01110000101000100", -- t[57668] = 24
      "0011000" when "01110000101000101", -- t[57669] = 24
      "0011000" when "01110000101000110", -- t[57670] = 24
      "0011000" when "01110000101000111", -- t[57671] = 24
      "0011000" when "01110000101001000", -- t[57672] = 24
      "0011000" when "01110000101001001", -- t[57673] = 24
      "0011000" when "01110000101001010", -- t[57674] = 24
      "0011000" when "01110000101001011", -- t[57675] = 24
      "0011000" when "01110000101001100", -- t[57676] = 24
      "0011000" when "01110000101001101", -- t[57677] = 24
      "0011000" when "01110000101001110", -- t[57678] = 24
      "0011000" when "01110000101001111", -- t[57679] = 24
      "0011000" when "01110000101010000", -- t[57680] = 24
      "0011000" when "01110000101010001", -- t[57681] = 24
      "0011000" when "01110000101010010", -- t[57682] = 24
      "0011000" when "01110000101010011", -- t[57683] = 24
      "0011000" when "01110000101010100", -- t[57684] = 24
      "0011000" when "01110000101010101", -- t[57685] = 24
      "0011000" when "01110000101010110", -- t[57686] = 24
      "0011000" when "01110000101010111", -- t[57687] = 24
      "0011000" when "01110000101011000", -- t[57688] = 24
      "0011000" when "01110000101011001", -- t[57689] = 24
      "0011000" when "01110000101011010", -- t[57690] = 24
      "0011000" when "01110000101011011", -- t[57691] = 24
      "0011000" when "01110000101011100", -- t[57692] = 24
      "0011000" when "01110000101011101", -- t[57693] = 24
      "0011000" when "01110000101011110", -- t[57694] = 24
      "0011000" when "01110000101011111", -- t[57695] = 24
      "0011000" when "01110000101100000", -- t[57696] = 24
      "0011000" when "01110000101100001", -- t[57697] = 24
      "0011000" when "01110000101100010", -- t[57698] = 24
      "0011000" when "01110000101100011", -- t[57699] = 24
      "0011000" when "01110000101100100", -- t[57700] = 24
      "0011000" when "01110000101100101", -- t[57701] = 24
      "0011000" when "01110000101100110", -- t[57702] = 24
      "0011000" when "01110000101100111", -- t[57703] = 24
      "0011000" when "01110000101101000", -- t[57704] = 24
      "0011000" when "01110000101101001", -- t[57705] = 24
      "0011000" when "01110000101101010", -- t[57706] = 24
      "0011000" when "01110000101101011", -- t[57707] = 24
      "0011000" when "01110000101101100", -- t[57708] = 24
      "0011000" when "01110000101101101", -- t[57709] = 24
      "0011000" when "01110000101101110", -- t[57710] = 24
      "0011000" when "01110000101101111", -- t[57711] = 24
      "0011000" when "01110000101110000", -- t[57712] = 24
      "0011000" when "01110000101110001", -- t[57713] = 24
      "0011000" when "01110000101110010", -- t[57714] = 24
      "0011000" when "01110000101110011", -- t[57715] = 24
      "0011000" when "01110000101110100", -- t[57716] = 24
      "0011000" when "01110000101110101", -- t[57717] = 24
      "0011000" when "01110000101110110", -- t[57718] = 24
      "0011000" when "01110000101110111", -- t[57719] = 24
      "0011000" when "01110000101111000", -- t[57720] = 24
      "0011000" when "01110000101111001", -- t[57721] = 24
      "0011000" when "01110000101111010", -- t[57722] = 24
      "0011000" when "01110000101111011", -- t[57723] = 24
      "0011000" when "01110000101111100", -- t[57724] = 24
      "0011000" when "01110000101111101", -- t[57725] = 24
      "0011000" when "01110000101111110", -- t[57726] = 24
      "0011000" when "01110000101111111", -- t[57727] = 24
      "0011000" when "01110000110000000", -- t[57728] = 24
      "0011000" when "01110000110000001", -- t[57729] = 24
      "0011000" when "01110000110000010", -- t[57730] = 24
      "0011000" when "01110000110000011", -- t[57731] = 24
      "0011000" when "01110000110000100", -- t[57732] = 24
      "0011000" when "01110000110000101", -- t[57733] = 24
      "0011000" when "01110000110000110", -- t[57734] = 24
      "0011000" when "01110000110000111", -- t[57735] = 24
      "0011000" when "01110000110001000", -- t[57736] = 24
      "0011000" when "01110000110001001", -- t[57737] = 24
      "0011000" when "01110000110001010", -- t[57738] = 24
      "0011000" when "01110000110001011", -- t[57739] = 24
      "0011000" when "01110000110001100", -- t[57740] = 24
      "0011000" when "01110000110001101", -- t[57741] = 24
      "0011000" when "01110000110001110", -- t[57742] = 24
      "0011000" when "01110000110001111", -- t[57743] = 24
      "0011000" when "01110000110010000", -- t[57744] = 24
      "0011000" when "01110000110010001", -- t[57745] = 24
      "0011000" when "01110000110010010", -- t[57746] = 24
      "0011000" when "01110000110010011", -- t[57747] = 24
      "0011000" when "01110000110010100", -- t[57748] = 24
      "0011000" when "01110000110010101", -- t[57749] = 24
      "0011000" when "01110000110010110", -- t[57750] = 24
      "0011000" when "01110000110010111", -- t[57751] = 24
      "0011000" when "01110000110011000", -- t[57752] = 24
      "0011000" when "01110000110011001", -- t[57753] = 24
      "0011000" when "01110000110011010", -- t[57754] = 24
      "0011000" when "01110000110011011", -- t[57755] = 24
      "0011000" when "01110000110011100", -- t[57756] = 24
      "0011000" when "01110000110011101", -- t[57757] = 24
      "0011000" when "01110000110011110", -- t[57758] = 24
      "0011000" when "01110000110011111", -- t[57759] = 24
      "0011000" when "01110000110100000", -- t[57760] = 24
      "0011000" when "01110000110100001", -- t[57761] = 24
      "0011000" when "01110000110100010", -- t[57762] = 24
      "0011000" when "01110000110100011", -- t[57763] = 24
      "0011000" when "01110000110100100", -- t[57764] = 24
      "0011000" when "01110000110100101", -- t[57765] = 24
      "0011000" when "01110000110100110", -- t[57766] = 24
      "0011000" when "01110000110100111", -- t[57767] = 24
      "0011000" when "01110000110101000", -- t[57768] = 24
      "0011000" when "01110000110101001", -- t[57769] = 24
      "0011000" when "01110000110101010", -- t[57770] = 24
      "0011000" when "01110000110101011", -- t[57771] = 24
      "0011000" when "01110000110101100", -- t[57772] = 24
      "0011000" when "01110000110101101", -- t[57773] = 24
      "0011000" when "01110000110101110", -- t[57774] = 24
      "0011000" when "01110000110101111", -- t[57775] = 24
      "0011000" when "01110000110110000", -- t[57776] = 24
      "0011000" when "01110000110110001", -- t[57777] = 24
      "0011000" when "01110000110110010", -- t[57778] = 24
      "0011000" when "01110000110110011", -- t[57779] = 24
      "0011000" when "01110000110110100", -- t[57780] = 24
      "0011000" when "01110000110110101", -- t[57781] = 24
      "0011000" when "01110000110110110", -- t[57782] = 24
      "0011000" when "01110000110110111", -- t[57783] = 24
      "0011000" when "01110000110111000", -- t[57784] = 24
      "0011000" when "01110000110111001", -- t[57785] = 24
      "0011000" when "01110000110111010", -- t[57786] = 24
      "0011000" when "01110000110111011", -- t[57787] = 24
      "0011000" when "01110000110111100", -- t[57788] = 24
      "0011000" when "01110000110111101", -- t[57789] = 24
      "0011000" when "01110000110111110", -- t[57790] = 24
      "0011000" when "01110000110111111", -- t[57791] = 24
      "0011000" when "01110000111000000", -- t[57792] = 24
      "0011000" when "01110000111000001", -- t[57793] = 24
      "0011000" when "01110000111000010", -- t[57794] = 24
      "0011000" when "01110000111000011", -- t[57795] = 24
      "0011000" when "01110000111000100", -- t[57796] = 24
      "0011000" when "01110000111000101", -- t[57797] = 24
      "0011000" when "01110000111000110", -- t[57798] = 24
      "0011000" when "01110000111000111", -- t[57799] = 24
      "0011000" when "01110000111001000", -- t[57800] = 24
      "0011000" when "01110000111001001", -- t[57801] = 24
      "0011000" when "01110000111001010", -- t[57802] = 24
      "0011000" when "01110000111001011", -- t[57803] = 24
      "0011000" when "01110000111001100", -- t[57804] = 24
      "0011000" when "01110000111001101", -- t[57805] = 24
      "0011000" when "01110000111001110", -- t[57806] = 24
      "0011000" when "01110000111001111", -- t[57807] = 24
      "0011000" when "01110000111010000", -- t[57808] = 24
      "0011000" when "01110000111010001", -- t[57809] = 24
      "0011000" when "01110000111010010", -- t[57810] = 24
      "0011000" when "01110000111010011", -- t[57811] = 24
      "0011000" when "01110000111010100", -- t[57812] = 24
      "0011000" when "01110000111010101", -- t[57813] = 24
      "0011000" when "01110000111010110", -- t[57814] = 24
      "0011000" when "01110000111010111", -- t[57815] = 24
      "0011000" when "01110000111011000", -- t[57816] = 24
      "0011000" when "01110000111011001", -- t[57817] = 24
      "0011000" when "01110000111011010", -- t[57818] = 24
      "0011000" when "01110000111011011", -- t[57819] = 24
      "0011000" when "01110000111011100", -- t[57820] = 24
      "0011000" when "01110000111011101", -- t[57821] = 24
      "0011000" when "01110000111011110", -- t[57822] = 24
      "0011000" when "01110000111011111", -- t[57823] = 24
      "0011000" when "01110000111100000", -- t[57824] = 24
      "0011000" when "01110000111100001", -- t[57825] = 24
      "0011000" when "01110000111100010", -- t[57826] = 24
      "0011000" when "01110000111100011", -- t[57827] = 24
      "0011000" when "01110000111100100", -- t[57828] = 24
      "0011000" when "01110000111100101", -- t[57829] = 24
      "0011000" when "01110000111100110", -- t[57830] = 24
      "0011000" when "01110000111100111", -- t[57831] = 24
      "0011000" when "01110000111101000", -- t[57832] = 24
      "0011000" when "01110000111101001", -- t[57833] = 24
      "0011000" when "01110000111101010", -- t[57834] = 24
      "0011000" when "01110000111101011", -- t[57835] = 24
      "0011000" when "01110000111101100", -- t[57836] = 24
      "0011000" when "01110000111101101", -- t[57837] = 24
      "0011000" when "01110000111101110", -- t[57838] = 24
      "0011000" when "01110000111101111", -- t[57839] = 24
      "0011000" when "01110000111110000", -- t[57840] = 24
      "0011000" when "01110000111110001", -- t[57841] = 24
      "0011000" when "01110000111110010", -- t[57842] = 24
      "0011000" when "01110000111110011", -- t[57843] = 24
      "0011000" when "01110000111110100", -- t[57844] = 24
      "0011000" when "01110000111110101", -- t[57845] = 24
      "0011000" when "01110000111110110", -- t[57846] = 24
      "0011000" when "01110000111110111", -- t[57847] = 24
      "0011000" when "01110000111111000", -- t[57848] = 24
      "0011000" when "01110000111111001", -- t[57849] = 24
      "0011000" when "01110000111111010", -- t[57850] = 24
      "0011000" when "01110000111111011", -- t[57851] = 24
      "0011000" when "01110000111111100", -- t[57852] = 24
      "0011000" when "01110000111111101", -- t[57853] = 24
      "0011000" when "01110000111111110", -- t[57854] = 24
      "0011000" when "01110000111111111", -- t[57855] = 24
      "0011000" when "01110001000000000", -- t[57856] = 24
      "0011000" when "01110001000000001", -- t[57857] = 24
      "0011000" when "01110001000000010", -- t[57858] = 24
      "0011000" when "01110001000000011", -- t[57859] = 24
      "0011000" when "01110001000000100", -- t[57860] = 24
      "0011000" when "01110001000000101", -- t[57861] = 24
      "0011000" when "01110001000000110", -- t[57862] = 24
      "0011000" when "01110001000000111", -- t[57863] = 24
      "0011000" when "01110001000001000", -- t[57864] = 24
      "0011000" when "01110001000001001", -- t[57865] = 24
      "0011000" when "01110001000001010", -- t[57866] = 24
      "0011000" when "01110001000001011", -- t[57867] = 24
      "0011000" when "01110001000001100", -- t[57868] = 24
      "0011000" when "01110001000001101", -- t[57869] = 24
      "0011000" when "01110001000001110", -- t[57870] = 24
      "0011000" when "01110001000001111", -- t[57871] = 24
      "0011000" when "01110001000010000", -- t[57872] = 24
      "0011000" when "01110001000010001", -- t[57873] = 24
      "0011000" when "01110001000010010", -- t[57874] = 24
      "0011000" when "01110001000010011", -- t[57875] = 24
      "0011000" when "01110001000010100", -- t[57876] = 24
      "0011000" when "01110001000010101", -- t[57877] = 24
      "0011000" when "01110001000010110", -- t[57878] = 24
      "0011000" when "01110001000010111", -- t[57879] = 24
      "0011000" when "01110001000011000", -- t[57880] = 24
      "0011000" when "01110001000011001", -- t[57881] = 24
      "0011000" when "01110001000011010", -- t[57882] = 24
      "0011000" when "01110001000011011", -- t[57883] = 24
      "0011000" when "01110001000011100", -- t[57884] = 24
      "0011000" when "01110001000011101", -- t[57885] = 24
      "0011000" when "01110001000011110", -- t[57886] = 24
      "0011000" when "01110001000011111", -- t[57887] = 24
      "0011000" when "01110001000100000", -- t[57888] = 24
      "0011000" when "01110001000100001", -- t[57889] = 24
      "0011000" when "01110001000100010", -- t[57890] = 24
      "0011000" when "01110001000100011", -- t[57891] = 24
      "0011000" when "01110001000100100", -- t[57892] = 24
      "0011000" when "01110001000100101", -- t[57893] = 24
      "0011000" when "01110001000100110", -- t[57894] = 24
      "0011000" when "01110001000100111", -- t[57895] = 24
      "0011000" when "01110001000101000", -- t[57896] = 24
      "0011000" when "01110001000101001", -- t[57897] = 24
      "0011000" when "01110001000101010", -- t[57898] = 24
      "0011000" when "01110001000101011", -- t[57899] = 24
      "0011000" when "01110001000101100", -- t[57900] = 24
      "0011000" when "01110001000101101", -- t[57901] = 24
      "0011000" when "01110001000101110", -- t[57902] = 24
      "0011000" when "01110001000101111", -- t[57903] = 24
      "0011000" when "01110001000110000", -- t[57904] = 24
      "0011000" when "01110001000110001", -- t[57905] = 24
      "0011000" when "01110001000110010", -- t[57906] = 24
      "0011000" when "01110001000110011", -- t[57907] = 24
      "0011000" when "01110001000110100", -- t[57908] = 24
      "0011000" when "01110001000110101", -- t[57909] = 24
      "0011000" when "01110001000110110", -- t[57910] = 24
      "0011000" when "01110001000110111", -- t[57911] = 24
      "0011000" when "01110001000111000", -- t[57912] = 24
      "0011000" when "01110001000111001", -- t[57913] = 24
      "0011000" when "01110001000111010", -- t[57914] = 24
      "0011000" when "01110001000111011", -- t[57915] = 24
      "0011000" when "01110001000111100", -- t[57916] = 24
      "0011000" when "01110001000111101", -- t[57917] = 24
      "0011000" when "01110001000111110", -- t[57918] = 24
      "0011000" when "01110001000111111", -- t[57919] = 24
      "0011000" when "01110001001000000", -- t[57920] = 24
      "0011000" when "01110001001000001", -- t[57921] = 24
      "0011000" when "01110001001000010", -- t[57922] = 24
      "0011000" when "01110001001000011", -- t[57923] = 24
      "0011000" when "01110001001000100", -- t[57924] = 24
      "0011000" when "01110001001000101", -- t[57925] = 24
      "0011000" when "01110001001000110", -- t[57926] = 24
      "0011000" when "01110001001000111", -- t[57927] = 24
      "0011000" when "01110001001001000", -- t[57928] = 24
      "0011000" when "01110001001001001", -- t[57929] = 24
      "0011000" when "01110001001001010", -- t[57930] = 24
      "0011000" when "01110001001001011", -- t[57931] = 24
      "0011000" when "01110001001001100", -- t[57932] = 24
      "0011000" when "01110001001001101", -- t[57933] = 24
      "0011000" when "01110001001001110", -- t[57934] = 24
      "0011000" when "01110001001001111", -- t[57935] = 24
      "0011000" when "01110001001010000", -- t[57936] = 24
      "0011000" when "01110001001010001", -- t[57937] = 24
      "0011000" when "01110001001010010", -- t[57938] = 24
      "0011000" when "01110001001010011", -- t[57939] = 24
      "0011000" when "01110001001010100", -- t[57940] = 24
      "0011000" when "01110001001010101", -- t[57941] = 24
      "0011000" when "01110001001010110", -- t[57942] = 24
      "0011000" when "01110001001010111", -- t[57943] = 24
      "0011000" when "01110001001011000", -- t[57944] = 24
      "0011000" when "01110001001011001", -- t[57945] = 24
      "0011000" when "01110001001011010", -- t[57946] = 24
      "0011000" when "01110001001011011", -- t[57947] = 24
      "0011000" when "01110001001011100", -- t[57948] = 24
      "0011000" when "01110001001011101", -- t[57949] = 24
      "0011000" when "01110001001011110", -- t[57950] = 24
      "0011000" when "01110001001011111", -- t[57951] = 24
      "0011000" when "01110001001100000", -- t[57952] = 24
      "0011000" when "01110001001100001", -- t[57953] = 24
      "0011000" when "01110001001100010", -- t[57954] = 24
      "0011000" when "01110001001100011", -- t[57955] = 24
      "0011000" when "01110001001100100", -- t[57956] = 24
      "0011000" when "01110001001100101", -- t[57957] = 24
      "0011000" when "01110001001100110", -- t[57958] = 24
      "0011000" when "01110001001100111", -- t[57959] = 24
      "0011000" when "01110001001101000", -- t[57960] = 24
      "0011000" when "01110001001101001", -- t[57961] = 24
      "0011000" when "01110001001101010", -- t[57962] = 24
      "0011000" when "01110001001101011", -- t[57963] = 24
      "0011000" when "01110001001101100", -- t[57964] = 24
      "0011000" when "01110001001101101", -- t[57965] = 24
      "0011000" when "01110001001101110", -- t[57966] = 24
      "0011000" when "01110001001101111", -- t[57967] = 24
      "0011000" when "01110001001110000", -- t[57968] = 24
      "0011000" when "01110001001110001", -- t[57969] = 24
      "0011000" when "01110001001110010", -- t[57970] = 24
      "0011000" when "01110001001110011", -- t[57971] = 24
      "0011000" when "01110001001110100", -- t[57972] = 24
      "0011000" when "01110001001110101", -- t[57973] = 24
      "0011000" when "01110001001110110", -- t[57974] = 24
      "0011000" when "01110001001110111", -- t[57975] = 24
      "0011000" when "01110001001111000", -- t[57976] = 24
      "0011000" when "01110001001111001", -- t[57977] = 24
      "0011000" when "01110001001111010", -- t[57978] = 24
      "0011000" when "01110001001111011", -- t[57979] = 24
      "0011000" when "01110001001111100", -- t[57980] = 24
      "0011000" when "01110001001111101", -- t[57981] = 24
      "0011000" when "01110001001111110", -- t[57982] = 24
      "0011000" when "01110001001111111", -- t[57983] = 24
      "0011000" when "01110001010000000", -- t[57984] = 24
      "0011000" when "01110001010000001", -- t[57985] = 24
      "0011000" when "01110001010000010", -- t[57986] = 24
      "0011000" when "01110001010000011", -- t[57987] = 24
      "0011000" when "01110001010000100", -- t[57988] = 24
      "0011000" when "01110001010000101", -- t[57989] = 24
      "0011000" when "01110001010000110", -- t[57990] = 24
      "0011000" when "01110001010000111", -- t[57991] = 24
      "0011000" when "01110001010001000", -- t[57992] = 24
      "0011000" when "01110001010001001", -- t[57993] = 24
      "0011000" when "01110001010001010", -- t[57994] = 24
      "0011000" when "01110001010001011", -- t[57995] = 24
      "0011000" when "01110001010001100", -- t[57996] = 24
      "0011000" when "01110001010001101", -- t[57997] = 24
      "0011000" when "01110001010001110", -- t[57998] = 24
      "0011000" when "01110001010001111", -- t[57999] = 24
      "0011000" when "01110001010010000", -- t[58000] = 24
      "0011000" when "01110001010010001", -- t[58001] = 24
      "0011000" when "01110001010010010", -- t[58002] = 24
      "0011000" when "01110001010010011", -- t[58003] = 24
      "0011000" when "01110001010010100", -- t[58004] = 24
      "0011000" when "01110001010010101", -- t[58005] = 24
      "0011000" when "01110001010010110", -- t[58006] = 24
      "0011000" when "01110001010010111", -- t[58007] = 24
      "0011000" when "01110001010011000", -- t[58008] = 24
      "0011000" when "01110001010011001", -- t[58009] = 24
      "0011000" when "01110001010011010", -- t[58010] = 24
      "0011000" when "01110001010011011", -- t[58011] = 24
      "0011000" when "01110001010011100", -- t[58012] = 24
      "0011000" when "01110001010011101", -- t[58013] = 24
      "0011000" when "01110001010011110", -- t[58014] = 24
      "0011000" when "01110001010011111", -- t[58015] = 24
      "0011000" when "01110001010100000", -- t[58016] = 24
      "0011000" when "01110001010100001", -- t[58017] = 24
      "0011000" when "01110001010100010", -- t[58018] = 24
      "0011000" when "01110001010100011", -- t[58019] = 24
      "0011000" when "01110001010100100", -- t[58020] = 24
      "0011000" when "01110001010100101", -- t[58021] = 24
      "0011000" when "01110001010100110", -- t[58022] = 24
      "0011000" when "01110001010100111", -- t[58023] = 24
      "0011000" when "01110001010101000", -- t[58024] = 24
      "0011000" when "01110001010101001", -- t[58025] = 24
      "0011000" when "01110001010101010", -- t[58026] = 24
      "0011000" when "01110001010101011", -- t[58027] = 24
      "0011000" when "01110001010101100", -- t[58028] = 24
      "0011000" when "01110001010101101", -- t[58029] = 24
      "0011000" when "01110001010101110", -- t[58030] = 24
      "0011000" when "01110001010101111", -- t[58031] = 24
      "0011000" when "01110001010110000", -- t[58032] = 24
      "0011000" when "01110001010110001", -- t[58033] = 24
      "0011000" when "01110001010110010", -- t[58034] = 24
      "0011000" when "01110001010110011", -- t[58035] = 24
      "0011001" when "01110001010110100", -- t[58036] = 25
      "0011001" when "01110001010110101", -- t[58037] = 25
      "0011001" when "01110001010110110", -- t[58038] = 25
      "0011001" when "01110001010110111", -- t[58039] = 25
      "0011001" when "01110001010111000", -- t[58040] = 25
      "0011001" when "01110001010111001", -- t[58041] = 25
      "0011001" when "01110001010111010", -- t[58042] = 25
      "0011001" when "01110001010111011", -- t[58043] = 25
      "0011001" when "01110001010111100", -- t[58044] = 25
      "0011001" when "01110001010111101", -- t[58045] = 25
      "0011001" when "01110001010111110", -- t[58046] = 25
      "0011001" when "01110001010111111", -- t[58047] = 25
      "0011001" when "01110001011000000", -- t[58048] = 25
      "0011001" when "01110001011000001", -- t[58049] = 25
      "0011001" when "01110001011000010", -- t[58050] = 25
      "0011001" when "01110001011000011", -- t[58051] = 25
      "0011001" when "01110001011000100", -- t[58052] = 25
      "0011001" when "01110001011000101", -- t[58053] = 25
      "0011001" when "01110001011000110", -- t[58054] = 25
      "0011001" when "01110001011000111", -- t[58055] = 25
      "0011001" when "01110001011001000", -- t[58056] = 25
      "0011001" when "01110001011001001", -- t[58057] = 25
      "0011001" when "01110001011001010", -- t[58058] = 25
      "0011001" when "01110001011001011", -- t[58059] = 25
      "0011001" when "01110001011001100", -- t[58060] = 25
      "0011001" when "01110001011001101", -- t[58061] = 25
      "0011001" when "01110001011001110", -- t[58062] = 25
      "0011001" when "01110001011001111", -- t[58063] = 25
      "0011001" when "01110001011010000", -- t[58064] = 25
      "0011001" when "01110001011010001", -- t[58065] = 25
      "0011001" when "01110001011010010", -- t[58066] = 25
      "0011001" when "01110001011010011", -- t[58067] = 25
      "0011001" when "01110001011010100", -- t[58068] = 25
      "0011001" when "01110001011010101", -- t[58069] = 25
      "0011001" when "01110001011010110", -- t[58070] = 25
      "0011001" when "01110001011010111", -- t[58071] = 25
      "0011001" when "01110001011011000", -- t[58072] = 25
      "0011001" when "01110001011011001", -- t[58073] = 25
      "0011001" when "01110001011011010", -- t[58074] = 25
      "0011001" when "01110001011011011", -- t[58075] = 25
      "0011001" when "01110001011011100", -- t[58076] = 25
      "0011001" when "01110001011011101", -- t[58077] = 25
      "0011001" when "01110001011011110", -- t[58078] = 25
      "0011001" when "01110001011011111", -- t[58079] = 25
      "0011001" when "01110001011100000", -- t[58080] = 25
      "0011001" when "01110001011100001", -- t[58081] = 25
      "0011001" when "01110001011100010", -- t[58082] = 25
      "0011001" when "01110001011100011", -- t[58083] = 25
      "0011001" when "01110001011100100", -- t[58084] = 25
      "0011001" when "01110001011100101", -- t[58085] = 25
      "0011001" when "01110001011100110", -- t[58086] = 25
      "0011001" when "01110001011100111", -- t[58087] = 25
      "0011001" when "01110001011101000", -- t[58088] = 25
      "0011001" when "01110001011101001", -- t[58089] = 25
      "0011001" when "01110001011101010", -- t[58090] = 25
      "0011001" when "01110001011101011", -- t[58091] = 25
      "0011001" when "01110001011101100", -- t[58092] = 25
      "0011001" when "01110001011101101", -- t[58093] = 25
      "0011001" when "01110001011101110", -- t[58094] = 25
      "0011001" when "01110001011101111", -- t[58095] = 25
      "0011001" when "01110001011110000", -- t[58096] = 25
      "0011001" when "01110001011110001", -- t[58097] = 25
      "0011001" when "01110001011110010", -- t[58098] = 25
      "0011001" when "01110001011110011", -- t[58099] = 25
      "0011001" when "01110001011110100", -- t[58100] = 25
      "0011001" when "01110001011110101", -- t[58101] = 25
      "0011001" when "01110001011110110", -- t[58102] = 25
      "0011001" when "01110001011110111", -- t[58103] = 25
      "0011001" when "01110001011111000", -- t[58104] = 25
      "0011001" when "01110001011111001", -- t[58105] = 25
      "0011001" when "01110001011111010", -- t[58106] = 25
      "0011001" when "01110001011111011", -- t[58107] = 25
      "0011001" when "01110001011111100", -- t[58108] = 25
      "0011001" when "01110001011111101", -- t[58109] = 25
      "0011001" when "01110001011111110", -- t[58110] = 25
      "0011001" when "01110001011111111", -- t[58111] = 25
      "0011001" when "01110001100000000", -- t[58112] = 25
      "0011001" when "01110001100000001", -- t[58113] = 25
      "0011001" when "01110001100000010", -- t[58114] = 25
      "0011001" when "01110001100000011", -- t[58115] = 25
      "0011001" when "01110001100000100", -- t[58116] = 25
      "0011001" when "01110001100000101", -- t[58117] = 25
      "0011001" when "01110001100000110", -- t[58118] = 25
      "0011001" when "01110001100000111", -- t[58119] = 25
      "0011001" when "01110001100001000", -- t[58120] = 25
      "0011001" when "01110001100001001", -- t[58121] = 25
      "0011001" when "01110001100001010", -- t[58122] = 25
      "0011001" when "01110001100001011", -- t[58123] = 25
      "0011001" when "01110001100001100", -- t[58124] = 25
      "0011001" when "01110001100001101", -- t[58125] = 25
      "0011001" when "01110001100001110", -- t[58126] = 25
      "0011001" when "01110001100001111", -- t[58127] = 25
      "0011001" when "01110001100010000", -- t[58128] = 25
      "0011001" when "01110001100010001", -- t[58129] = 25
      "0011001" when "01110001100010010", -- t[58130] = 25
      "0011001" when "01110001100010011", -- t[58131] = 25
      "0011001" when "01110001100010100", -- t[58132] = 25
      "0011001" when "01110001100010101", -- t[58133] = 25
      "0011001" when "01110001100010110", -- t[58134] = 25
      "0011001" when "01110001100010111", -- t[58135] = 25
      "0011001" when "01110001100011000", -- t[58136] = 25
      "0011001" when "01110001100011001", -- t[58137] = 25
      "0011001" when "01110001100011010", -- t[58138] = 25
      "0011001" when "01110001100011011", -- t[58139] = 25
      "0011001" when "01110001100011100", -- t[58140] = 25
      "0011001" when "01110001100011101", -- t[58141] = 25
      "0011001" when "01110001100011110", -- t[58142] = 25
      "0011001" when "01110001100011111", -- t[58143] = 25
      "0011001" when "01110001100100000", -- t[58144] = 25
      "0011001" when "01110001100100001", -- t[58145] = 25
      "0011001" when "01110001100100010", -- t[58146] = 25
      "0011001" when "01110001100100011", -- t[58147] = 25
      "0011001" when "01110001100100100", -- t[58148] = 25
      "0011001" when "01110001100100101", -- t[58149] = 25
      "0011001" when "01110001100100110", -- t[58150] = 25
      "0011001" when "01110001100100111", -- t[58151] = 25
      "0011001" when "01110001100101000", -- t[58152] = 25
      "0011001" when "01110001100101001", -- t[58153] = 25
      "0011001" when "01110001100101010", -- t[58154] = 25
      "0011001" when "01110001100101011", -- t[58155] = 25
      "0011001" when "01110001100101100", -- t[58156] = 25
      "0011001" when "01110001100101101", -- t[58157] = 25
      "0011001" when "01110001100101110", -- t[58158] = 25
      "0011001" when "01110001100101111", -- t[58159] = 25
      "0011001" when "01110001100110000", -- t[58160] = 25
      "0011001" when "01110001100110001", -- t[58161] = 25
      "0011001" when "01110001100110010", -- t[58162] = 25
      "0011001" when "01110001100110011", -- t[58163] = 25
      "0011001" when "01110001100110100", -- t[58164] = 25
      "0011001" when "01110001100110101", -- t[58165] = 25
      "0011001" when "01110001100110110", -- t[58166] = 25
      "0011001" when "01110001100110111", -- t[58167] = 25
      "0011001" when "01110001100111000", -- t[58168] = 25
      "0011001" when "01110001100111001", -- t[58169] = 25
      "0011001" when "01110001100111010", -- t[58170] = 25
      "0011001" when "01110001100111011", -- t[58171] = 25
      "0011001" when "01110001100111100", -- t[58172] = 25
      "0011001" when "01110001100111101", -- t[58173] = 25
      "0011001" when "01110001100111110", -- t[58174] = 25
      "0011001" when "01110001100111111", -- t[58175] = 25
      "0011001" when "01110001101000000", -- t[58176] = 25
      "0011001" when "01110001101000001", -- t[58177] = 25
      "0011001" when "01110001101000010", -- t[58178] = 25
      "0011001" when "01110001101000011", -- t[58179] = 25
      "0011001" when "01110001101000100", -- t[58180] = 25
      "0011001" when "01110001101000101", -- t[58181] = 25
      "0011001" when "01110001101000110", -- t[58182] = 25
      "0011001" when "01110001101000111", -- t[58183] = 25
      "0011001" when "01110001101001000", -- t[58184] = 25
      "0011001" when "01110001101001001", -- t[58185] = 25
      "0011001" when "01110001101001010", -- t[58186] = 25
      "0011001" when "01110001101001011", -- t[58187] = 25
      "0011001" when "01110001101001100", -- t[58188] = 25
      "0011001" when "01110001101001101", -- t[58189] = 25
      "0011001" when "01110001101001110", -- t[58190] = 25
      "0011001" when "01110001101001111", -- t[58191] = 25
      "0011001" when "01110001101010000", -- t[58192] = 25
      "0011001" when "01110001101010001", -- t[58193] = 25
      "0011001" when "01110001101010010", -- t[58194] = 25
      "0011001" when "01110001101010011", -- t[58195] = 25
      "0011001" when "01110001101010100", -- t[58196] = 25
      "0011001" when "01110001101010101", -- t[58197] = 25
      "0011001" when "01110001101010110", -- t[58198] = 25
      "0011001" when "01110001101010111", -- t[58199] = 25
      "0011001" when "01110001101011000", -- t[58200] = 25
      "0011001" when "01110001101011001", -- t[58201] = 25
      "0011001" when "01110001101011010", -- t[58202] = 25
      "0011001" when "01110001101011011", -- t[58203] = 25
      "0011001" when "01110001101011100", -- t[58204] = 25
      "0011001" when "01110001101011101", -- t[58205] = 25
      "0011001" when "01110001101011110", -- t[58206] = 25
      "0011001" when "01110001101011111", -- t[58207] = 25
      "0011001" when "01110001101100000", -- t[58208] = 25
      "0011001" when "01110001101100001", -- t[58209] = 25
      "0011001" when "01110001101100010", -- t[58210] = 25
      "0011001" when "01110001101100011", -- t[58211] = 25
      "0011001" when "01110001101100100", -- t[58212] = 25
      "0011001" when "01110001101100101", -- t[58213] = 25
      "0011001" when "01110001101100110", -- t[58214] = 25
      "0011001" when "01110001101100111", -- t[58215] = 25
      "0011001" when "01110001101101000", -- t[58216] = 25
      "0011001" when "01110001101101001", -- t[58217] = 25
      "0011001" when "01110001101101010", -- t[58218] = 25
      "0011001" when "01110001101101011", -- t[58219] = 25
      "0011001" when "01110001101101100", -- t[58220] = 25
      "0011001" when "01110001101101101", -- t[58221] = 25
      "0011001" when "01110001101101110", -- t[58222] = 25
      "0011001" when "01110001101101111", -- t[58223] = 25
      "0011001" when "01110001101110000", -- t[58224] = 25
      "0011001" when "01110001101110001", -- t[58225] = 25
      "0011001" when "01110001101110010", -- t[58226] = 25
      "0011001" when "01110001101110011", -- t[58227] = 25
      "0011001" when "01110001101110100", -- t[58228] = 25
      "0011001" when "01110001101110101", -- t[58229] = 25
      "0011001" when "01110001101110110", -- t[58230] = 25
      "0011001" when "01110001101110111", -- t[58231] = 25
      "0011001" when "01110001101111000", -- t[58232] = 25
      "0011001" when "01110001101111001", -- t[58233] = 25
      "0011001" when "01110001101111010", -- t[58234] = 25
      "0011001" when "01110001101111011", -- t[58235] = 25
      "0011001" when "01110001101111100", -- t[58236] = 25
      "0011001" when "01110001101111101", -- t[58237] = 25
      "0011001" when "01110001101111110", -- t[58238] = 25
      "0011001" when "01110001101111111", -- t[58239] = 25
      "0011001" when "01110001110000000", -- t[58240] = 25
      "0011001" when "01110001110000001", -- t[58241] = 25
      "0011001" when "01110001110000010", -- t[58242] = 25
      "0011001" when "01110001110000011", -- t[58243] = 25
      "0011001" when "01110001110000100", -- t[58244] = 25
      "0011001" when "01110001110000101", -- t[58245] = 25
      "0011001" when "01110001110000110", -- t[58246] = 25
      "0011001" when "01110001110000111", -- t[58247] = 25
      "0011001" when "01110001110001000", -- t[58248] = 25
      "0011001" when "01110001110001001", -- t[58249] = 25
      "0011001" when "01110001110001010", -- t[58250] = 25
      "0011001" when "01110001110001011", -- t[58251] = 25
      "0011001" when "01110001110001100", -- t[58252] = 25
      "0011001" when "01110001110001101", -- t[58253] = 25
      "0011001" when "01110001110001110", -- t[58254] = 25
      "0011001" when "01110001110001111", -- t[58255] = 25
      "0011001" when "01110001110010000", -- t[58256] = 25
      "0011001" when "01110001110010001", -- t[58257] = 25
      "0011001" when "01110001110010010", -- t[58258] = 25
      "0011001" when "01110001110010011", -- t[58259] = 25
      "0011001" when "01110001110010100", -- t[58260] = 25
      "0011001" when "01110001110010101", -- t[58261] = 25
      "0011001" when "01110001110010110", -- t[58262] = 25
      "0011001" when "01110001110010111", -- t[58263] = 25
      "0011001" when "01110001110011000", -- t[58264] = 25
      "0011001" when "01110001110011001", -- t[58265] = 25
      "0011001" when "01110001110011010", -- t[58266] = 25
      "0011001" when "01110001110011011", -- t[58267] = 25
      "0011001" when "01110001110011100", -- t[58268] = 25
      "0011001" when "01110001110011101", -- t[58269] = 25
      "0011001" when "01110001110011110", -- t[58270] = 25
      "0011001" when "01110001110011111", -- t[58271] = 25
      "0011001" when "01110001110100000", -- t[58272] = 25
      "0011001" when "01110001110100001", -- t[58273] = 25
      "0011001" when "01110001110100010", -- t[58274] = 25
      "0011001" when "01110001110100011", -- t[58275] = 25
      "0011001" when "01110001110100100", -- t[58276] = 25
      "0011001" when "01110001110100101", -- t[58277] = 25
      "0011001" when "01110001110100110", -- t[58278] = 25
      "0011001" when "01110001110100111", -- t[58279] = 25
      "0011001" when "01110001110101000", -- t[58280] = 25
      "0011001" when "01110001110101001", -- t[58281] = 25
      "0011001" when "01110001110101010", -- t[58282] = 25
      "0011001" when "01110001110101011", -- t[58283] = 25
      "0011001" when "01110001110101100", -- t[58284] = 25
      "0011001" when "01110001110101101", -- t[58285] = 25
      "0011001" when "01110001110101110", -- t[58286] = 25
      "0011001" when "01110001110101111", -- t[58287] = 25
      "0011001" when "01110001110110000", -- t[58288] = 25
      "0011001" when "01110001110110001", -- t[58289] = 25
      "0011001" when "01110001110110010", -- t[58290] = 25
      "0011001" when "01110001110110011", -- t[58291] = 25
      "0011001" when "01110001110110100", -- t[58292] = 25
      "0011001" when "01110001110110101", -- t[58293] = 25
      "0011001" when "01110001110110110", -- t[58294] = 25
      "0011001" when "01110001110110111", -- t[58295] = 25
      "0011001" when "01110001110111000", -- t[58296] = 25
      "0011001" when "01110001110111001", -- t[58297] = 25
      "0011001" when "01110001110111010", -- t[58298] = 25
      "0011001" when "01110001110111011", -- t[58299] = 25
      "0011001" when "01110001110111100", -- t[58300] = 25
      "0011001" when "01110001110111101", -- t[58301] = 25
      "0011001" when "01110001110111110", -- t[58302] = 25
      "0011001" when "01110001110111111", -- t[58303] = 25
      "0011001" when "01110001111000000", -- t[58304] = 25
      "0011001" when "01110001111000001", -- t[58305] = 25
      "0011001" when "01110001111000010", -- t[58306] = 25
      "0011001" when "01110001111000011", -- t[58307] = 25
      "0011001" when "01110001111000100", -- t[58308] = 25
      "0011001" when "01110001111000101", -- t[58309] = 25
      "0011001" when "01110001111000110", -- t[58310] = 25
      "0011001" when "01110001111000111", -- t[58311] = 25
      "0011001" when "01110001111001000", -- t[58312] = 25
      "0011001" when "01110001111001001", -- t[58313] = 25
      "0011001" when "01110001111001010", -- t[58314] = 25
      "0011001" when "01110001111001011", -- t[58315] = 25
      "0011001" when "01110001111001100", -- t[58316] = 25
      "0011001" when "01110001111001101", -- t[58317] = 25
      "0011001" when "01110001111001110", -- t[58318] = 25
      "0011001" when "01110001111001111", -- t[58319] = 25
      "0011001" when "01110001111010000", -- t[58320] = 25
      "0011001" when "01110001111010001", -- t[58321] = 25
      "0011001" when "01110001111010010", -- t[58322] = 25
      "0011001" when "01110001111010011", -- t[58323] = 25
      "0011001" when "01110001111010100", -- t[58324] = 25
      "0011001" when "01110001111010101", -- t[58325] = 25
      "0011001" when "01110001111010110", -- t[58326] = 25
      "0011001" when "01110001111010111", -- t[58327] = 25
      "0011001" when "01110001111011000", -- t[58328] = 25
      "0011001" when "01110001111011001", -- t[58329] = 25
      "0011001" when "01110001111011010", -- t[58330] = 25
      "0011001" when "01110001111011011", -- t[58331] = 25
      "0011001" when "01110001111011100", -- t[58332] = 25
      "0011001" when "01110001111011101", -- t[58333] = 25
      "0011001" when "01110001111011110", -- t[58334] = 25
      "0011001" when "01110001111011111", -- t[58335] = 25
      "0011001" when "01110001111100000", -- t[58336] = 25
      "0011001" when "01110001111100001", -- t[58337] = 25
      "0011001" when "01110001111100010", -- t[58338] = 25
      "0011001" when "01110001111100011", -- t[58339] = 25
      "0011001" when "01110001111100100", -- t[58340] = 25
      "0011001" when "01110001111100101", -- t[58341] = 25
      "0011001" when "01110001111100110", -- t[58342] = 25
      "0011001" when "01110001111100111", -- t[58343] = 25
      "0011001" when "01110001111101000", -- t[58344] = 25
      "0011001" when "01110001111101001", -- t[58345] = 25
      "0011001" when "01110001111101010", -- t[58346] = 25
      "0011001" when "01110001111101011", -- t[58347] = 25
      "0011001" when "01110001111101100", -- t[58348] = 25
      "0011001" when "01110001111101101", -- t[58349] = 25
      "0011001" when "01110001111101110", -- t[58350] = 25
      "0011001" when "01110001111101111", -- t[58351] = 25
      "0011001" when "01110001111110000", -- t[58352] = 25
      "0011001" when "01110001111110001", -- t[58353] = 25
      "0011001" when "01110001111110010", -- t[58354] = 25
      "0011001" when "01110001111110011", -- t[58355] = 25
      "0011001" when "01110001111110100", -- t[58356] = 25
      "0011001" when "01110001111110101", -- t[58357] = 25
      "0011001" when "01110001111110110", -- t[58358] = 25
      "0011001" when "01110001111110111", -- t[58359] = 25
      "0011001" when "01110001111111000", -- t[58360] = 25
      "0011001" when "01110001111111001", -- t[58361] = 25
      "0011001" when "01110001111111010", -- t[58362] = 25
      "0011001" when "01110001111111011", -- t[58363] = 25
      "0011001" when "01110001111111100", -- t[58364] = 25
      "0011001" when "01110001111111101", -- t[58365] = 25
      "0011001" when "01110001111111110", -- t[58366] = 25
      "0011001" when "01110001111111111", -- t[58367] = 25
      "0011001" when "01110010000000000", -- t[58368] = 25
      "0011001" when "01110010000000001", -- t[58369] = 25
      "0011001" when "01110010000000010", -- t[58370] = 25
      "0011001" when "01110010000000011", -- t[58371] = 25
      "0011001" when "01110010000000100", -- t[58372] = 25
      "0011001" when "01110010000000101", -- t[58373] = 25
      "0011001" when "01110010000000110", -- t[58374] = 25
      "0011001" when "01110010000000111", -- t[58375] = 25
      "0011001" when "01110010000001000", -- t[58376] = 25
      "0011001" when "01110010000001001", -- t[58377] = 25
      "0011001" when "01110010000001010", -- t[58378] = 25
      "0011001" when "01110010000001011", -- t[58379] = 25
      "0011001" when "01110010000001100", -- t[58380] = 25
      "0011001" when "01110010000001101", -- t[58381] = 25
      "0011001" when "01110010000001110", -- t[58382] = 25
      "0011001" when "01110010000001111", -- t[58383] = 25
      "0011001" when "01110010000010000", -- t[58384] = 25
      "0011001" when "01110010000010001", -- t[58385] = 25
      "0011001" when "01110010000010010", -- t[58386] = 25
      "0011001" when "01110010000010011", -- t[58387] = 25
      "0011001" when "01110010000010100", -- t[58388] = 25
      "0011001" when "01110010000010101", -- t[58389] = 25
      "0011001" when "01110010000010110", -- t[58390] = 25
      "0011001" when "01110010000010111", -- t[58391] = 25
      "0011001" when "01110010000011000", -- t[58392] = 25
      "0011001" when "01110010000011001", -- t[58393] = 25
      "0011001" when "01110010000011010", -- t[58394] = 25
      "0011001" when "01110010000011011", -- t[58395] = 25
      "0011001" when "01110010000011100", -- t[58396] = 25
      "0011001" when "01110010000011101", -- t[58397] = 25
      "0011001" when "01110010000011110", -- t[58398] = 25
      "0011001" when "01110010000011111", -- t[58399] = 25
      "0011001" when "01110010000100000", -- t[58400] = 25
      "0011001" when "01110010000100001", -- t[58401] = 25
      "0011001" when "01110010000100010", -- t[58402] = 25
      "0011001" when "01110010000100011", -- t[58403] = 25
      "0011001" when "01110010000100100", -- t[58404] = 25
      "0011001" when "01110010000100101", -- t[58405] = 25
      "0011001" when "01110010000100110", -- t[58406] = 25
      "0011001" when "01110010000100111", -- t[58407] = 25
      "0011001" when "01110010000101000", -- t[58408] = 25
      "0011001" when "01110010000101001", -- t[58409] = 25
      "0011001" when "01110010000101010", -- t[58410] = 25
      "0011001" when "01110010000101011", -- t[58411] = 25
      "0011001" when "01110010000101100", -- t[58412] = 25
      "0011001" when "01110010000101101", -- t[58413] = 25
      "0011001" when "01110010000101110", -- t[58414] = 25
      "0011001" when "01110010000101111", -- t[58415] = 25
      "0011001" when "01110010000110000", -- t[58416] = 25
      "0011001" when "01110010000110001", -- t[58417] = 25
      "0011001" when "01110010000110010", -- t[58418] = 25
      "0011001" when "01110010000110011", -- t[58419] = 25
      "0011001" when "01110010000110100", -- t[58420] = 25
      "0011001" when "01110010000110101", -- t[58421] = 25
      "0011001" when "01110010000110110", -- t[58422] = 25
      "0011001" when "01110010000110111", -- t[58423] = 25
      "0011001" when "01110010000111000", -- t[58424] = 25
      "0011001" when "01110010000111001", -- t[58425] = 25
      "0011001" when "01110010000111010", -- t[58426] = 25
      "0011001" when "01110010000111011", -- t[58427] = 25
      "0011001" when "01110010000111100", -- t[58428] = 25
      "0011001" when "01110010000111101", -- t[58429] = 25
      "0011001" when "01110010000111110", -- t[58430] = 25
      "0011001" when "01110010000111111", -- t[58431] = 25
      "0011001" when "01110010001000000", -- t[58432] = 25
      "0011001" when "01110010001000001", -- t[58433] = 25
      "0011001" when "01110010001000010", -- t[58434] = 25
      "0011001" when "01110010001000011", -- t[58435] = 25
      "0011001" when "01110010001000100", -- t[58436] = 25
      "0011001" when "01110010001000101", -- t[58437] = 25
      "0011001" when "01110010001000110", -- t[58438] = 25
      "0011001" when "01110010001000111", -- t[58439] = 25
      "0011001" when "01110010001001000", -- t[58440] = 25
      "0011001" when "01110010001001001", -- t[58441] = 25
      "0011001" when "01110010001001010", -- t[58442] = 25
      "0011001" when "01110010001001011", -- t[58443] = 25
      "0011001" when "01110010001001100", -- t[58444] = 25
      "0011001" when "01110010001001101", -- t[58445] = 25
      "0011001" when "01110010001001110", -- t[58446] = 25
      "0011001" when "01110010001001111", -- t[58447] = 25
      "0011001" when "01110010001010000", -- t[58448] = 25
      "0011001" when "01110010001010001", -- t[58449] = 25
      "0011001" when "01110010001010010", -- t[58450] = 25
      "0011001" when "01110010001010011", -- t[58451] = 25
      "0011001" when "01110010001010100", -- t[58452] = 25
      "0011001" when "01110010001010101", -- t[58453] = 25
      "0011001" when "01110010001010110", -- t[58454] = 25
      "0011001" when "01110010001010111", -- t[58455] = 25
      "0011001" when "01110010001011000", -- t[58456] = 25
      "0011001" when "01110010001011001", -- t[58457] = 25
      "0011001" when "01110010001011010", -- t[58458] = 25
      "0011001" when "01110010001011011", -- t[58459] = 25
      "0011001" when "01110010001011100", -- t[58460] = 25
      "0011001" when "01110010001011101", -- t[58461] = 25
      "0011001" when "01110010001011110", -- t[58462] = 25
      "0011001" when "01110010001011111", -- t[58463] = 25
      "0011001" when "01110010001100000", -- t[58464] = 25
      "0011001" when "01110010001100001", -- t[58465] = 25
      "0011001" when "01110010001100010", -- t[58466] = 25
      "0011001" when "01110010001100011", -- t[58467] = 25
      "0011001" when "01110010001100100", -- t[58468] = 25
      "0011001" when "01110010001100101", -- t[58469] = 25
      "0011001" when "01110010001100110", -- t[58470] = 25
      "0011001" when "01110010001100111", -- t[58471] = 25
      "0011001" when "01110010001101000", -- t[58472] = 25
      "0011001" when "01110010001101001", -- t[58473] = 25
      "0011001" when "01110010001101010", -- t[58474] = 25
      "0011001" when "01110010001101011", -- t[58475] = 25
      "0011001" when "01110010001101100", -- t[58476] = 25
      "0011001" when "01110010001101101", -- t[58477] = 25
      "0011001" when "01110010001101110", -- t[58478] = 25
      "0011001" when "01110010001101111", -- t[58479] = 25
      "0011001" when "01110010001110000", -- t[58480] = 25
      "0011001" when "01110010001110001", -- t[58481] = 25
      "0011001" when "01110010001110010", -- t[58482] = 25
      "0011001" when "01110010001110011", -- t[58483] = 25
      "0011001" when "01110010001110100", -- t[58484] = 25
      "0011001" when "01110010001110101", -- t[58485] = 25
      "0011001" when "01110010001110110", -- t[58486] = 25
      "0011001" when "01110010001110111", -- t[58487] = 25
      "0011001" when "01110010001111000", -- t[58488] = 25
      "0011001" when "01110010001111001", -- t[58489] = 25
      "0011001" when "01110010001111010", -- t[58490] = 25
      "0011001" when "01110010001111011", -- t[58491] = 25
      "0011001" when "01110010001111100", -- t[58492] = 25
      "0011001" when "01110010001111101", -- t[58493] = 25
      "0011001" when "01110010001111110", -- t[58494] = 25
      "0011001" when "01110010001111111", -- t[58495] = 25
      "0011001" when "01110010010000000", -- t[58496] = 25
      "0011001" when "01110010010000001", -- t[58497] = 25
      "0011001" when "01110010010000010", -- t[58498] = 25
      "0011001" when "01110010010000011", -- t[58499] = 25
      "0011001" when "01110010010000100", -- t[58500] = 25
      "0011001" when "01110010010000101", -- t[58501] = 25
      "0011001" when "01110010010000110", -- t[58502] = 25
      "0011001" when "01110010010000111", -- t[58503] = 25
      "0011001" when "01110010010001000", -- t[58504] = 25
      "0011001" when "01110010010001001", -- t[58505] = 25
      "0011001" when "01110010010001010", -- t[58506] = 25
      "0011001" when "01110010010001011", -- t[58507] = 25
      "0011001" when "01110010010001100", -- t[58508] = 25
      "0011010" when "01110010010001101", -- t[58509] = 26
      "0011010" when "01110010010001110", -- t[58510] = 26
      "0011010" when "01110010010001111", -- t[58511] = 26
      "0011010" when "01110010010010000", -- t[58512] = 26
      "0011010" when "01110010010010001", -- t[58513] = 26
      "0011010" when "01110010010010010", -- t[58514] = 26
      "0011010" when "01110010010010011", -- t[58515] = 26
      "0011010" when "01110010010010100", -- t[58516] = 26
      "0011010" when "01110010010010101", -- t[58517] = 26
      "0011010" when "01110010010010110", -- t[58518] = 26
      "0011010" when "01110010010010111", -- t[58519] = 26
      "0011010" when "01110010010011000", -- t[58520] = 26
      "0011010" when "01110010010011001", -- t[58521] = 26
      "0011010" when "01110010010011010", -- t[58522] = 26
      "0011010" when "01110010010011011", -- t[58523] = 26
      "0011010" when "01110010010011100", -- t[58524] = 26
      "0011010" when "01110010010011101", -- t[58525] = 26
      "0011010" when "01110010010011110", -- t[58526] = 26
      "0011010" when "01110010010011111", -- t[58527] = 26
      "0011010" when "01110010010100000", -- t[58528] = 26
      "0011010" when "01110010010100001", -- t[58529] = 26
      "0011010" when "01110010010100010", -- t[58530] = 26
      "0011010" when "01110010010100011", -- t[58531] = 26
      "0011010" when "01110010010100100", -- t[58532] = 26
      "0011010" when "01110010010100101", -- t[58533] = 26
      "0011010" when "01110010010100110", -- t[58534] = 26
      "0011010" when "01110010010100111", -- t[58535] = 26
      "0011010" when "01110010010101000", -- t[58536] = 26
      "0011010" when "01110010010101001", -- t[58537] = 26
      "0011010" when "01110010010101010", -- t[58538] = 26
      "0011010" when "01110010010101011", -- t[58539] = 26
      "0011010" when "01110010010101100", -- t[58540] = 26
      "0011010" when "01110010010101101", -- t[58541] = 26
      "0011010" when "01110010010101110", -- t[58542] = 26
      "0011010" when "01110010010101111", -- t[58543] = 26
      "0011010" when "01110010010110000", -- t[58544] = 26
      "0011010" when "01110010010110001", -- t[58545] = 26
      "0011010" when "01110010010110010", -- t[58546] = 26
      "0011010" when "01110010010110011", -- t[58547] = 26
      "0011010" when "01110010010110100", -- t[58548] = 26
      "0011010" when "01110010010110101", -- t[58549] = 26
      "0011010" when "01110010010110110", -- t[58550] = 26
      "0011010" when "01110010010110111", -- t[58551] = 26
      "0011010" when "01110010010111000", -- t[58552] = 26
      "0011010" when "01110010010111001", -- t[58553] = 26
      "0011010" when "01110010010111010", -- t[58554] = 26
      "0011010" when "01110010010111011", -- t[58555] = 26
      "0011010" when "01110010010111100", -- t[58556] = 26
      "0011010" when "01110010010111101", -- t[58557] = 26
      "0011010" when "01110010010111110", -- t[58558] = 26
      "0011010" when "01110010010111111", -- t[58559] = 26
      "0011010" when "01110010011000000", -- t[58560] = 26
      "0011010" when "01110010011000001", -- t[58561] = 26
      "0011010" when "01110010011000010", -- t[58562] = 26
      "0011010" when "01110010011000011", -- t[58563] = 26
      "0011010" when "01110010011000100", -- t[58564] = 26
      "0011010" when "01110010011000101", -- t[58565] = 26
      "0011010" when "01110010011000110", -- t[58566] = 26
      "0011010" when "01110010011000111", -- t[58567] = 26
      "0011010" when "01110010011001000", -- t[58568] = 26
      "0011010" when "01110010011001001", -- t[58569] = 26
      "0011010" when "01110010011001010", -- t[58570] = 26
      "0011010" when "01110010011001011", -- t[58571] = 26
      "0011010" when "01110010011001100", -- t[58572] = 26
      "0011010" when "01110010011001101", -- t[58573] = 26
      "0011010" when "01110010011001110", -- t[58574] = 26
      "0011010" when "01110010011001111", -- t[58575] = 26
      "0011010" when "01110010011010000", -- t[58576] = 26
      "0011010" when "01110010011010001", -- t[58577] = 26
      "0011010" when "01110010011010010", -- t[58578] = 26
      "0011010" when "01110010011010011", -- t[58579] = 26
      "0011010" when "01110010011010100", -- t[58580] = 26
      "0011010" when "01110010011010101", -- t[58581] = 26
      "0011010" when "01110010011010110", -- t[58582] = 26
      "0011010" when "01110010011010111", -- t[58583] = 26
      "0011010" when "01110010011011000", -- t[58584] = 26
      "0011010" when "01110010011011001", -- t[58585] = 26
      "0011010" when "01110010011011010", -- t[58586] = 26
      "0011010" when "01110010011011011", -- t[58587] = 26
      "0011010" when "01110010011011100", -- t[58588] = 26
      "0011010" when "01110010011011101", -- t[58589] = 26
      "0011010" when "01110010011011110", -- t[58590] = 26
      "0011010" when "01110010011011111", -- t[58591] = 26
      "0011010" when "01110010011100000", -- t[58592] = 26
      "0011010" when "01110010011100001", -- t[58593] = 26
      "0011010" when "01110010011100010", -- t[58594] = 26
      "0011010" when "01110010011100011", -- t[58595] = 26
      "0011010" when "01110010011100100", -- t[58596] = 26
      "0011010" when "01110010011100101", -- t[58597] = 26
      "0011010" when "01110010011100110", -- t[58598] = 26
      "0011010" when "01110010011100111", -- t[58599] = 26
      "0011010" when "01110010011101000", -- t[58600] = 26
      "0011010" when "01110010011101001", -- t[58601] = 26
      "0011010" when "01110010011101010", -- t[58602] = 26
      "0011010" when "01110010011101011", -- t[58603] = 26
      "0011010" when "01110010011101100", -- t[58604] = 26
      "0011010" when "01110010011101101", -- t[58605] = 26
      "0011010" when "01110010011101110", -- t[58606] = 26
      "0011010" when "01110010011101111", -- t[58607] = 26
      "0011010" when "01110010011110000", -- t[58608] = 26
      "0011010" when "01110010011110001", -- t[58609] = 26
      "0011010" when "01110010011110010", -- t[58610] = 26
      "0011010" when "01110010011110011", -- t[58611] = 26
      "0011010" when "01110010011110100", -- t[58612] = 26
      "0011010" when "01110010011110101", -- t[58613] = 26
      "0011010" when "01110010011110110", -- t[58614] = 26
      "0011010" when "01110010011110111", -- t[58615] = 26
      "0011010" when "01110010011111000", -- t[58616] = 26
      "0011010" when "01110010011111001", -- t[58617] = 26
      "0011010" when "01110010011111010", -- t[58618] = 26
      "0011010" when "01110010011111011", -- t[58619] = 26
      "0011010" when "01110010011111100", -- t[58620] = 26
      "0011010" when "01110010011111101", -- t[58621] = 26
      "0011010" when "01110010011111110", -- t[58622] = 26
      "0011010" when "01110010011111111", -- t[58623] = 26
      "0011010" when "01110010100000000", -- t[58624] = 26
      "0011010" when "01110010100000001", -- t[58625] = 26
      "0011010" when "01110010100000010", -- t[58626] = 26
      "0011010" when "01110010100000011", -- t[58627] = 26
      "0011010" when "01110010100000100", -- t[58628] = 26
      "0011010" when "01110010100000101", -- t[58629] = 26
      "0011010" when "01110010100000110", -- t[58630] = 26
      "0011010" when "01110010100000111", -- t[58631] = 26
      "0011010" when "01110010100001000", -- t[58632] = 26
      "0011010" when "01110010100001001", -- t[58633] = 26
      "0011010" when "01110010100001010", -- t[58634] = 26
      "0011010" when "01110010100001011", -- t[58635] = 26
      "0011010" when "01110010100001100", -- t[58636] = 26
      "0011010" when "01110010100001101", -- t[58637] = 26
      "0011010" when "01110010100001110", -- t[58638] = 26
      "0011010" when "01110010100001111", -- t[58639] = 26
      "0011010" when "01110010100010000", -- t[58640] = 26
      "0011010" when "01110010100010001", -- t[58641] = 26
      "0011010" when "01110010100010010", -- t[58642] = 26
      "0011010" when "01110010100010011", -- t[58643] = 26
      "0011010" when "01110010100010100", -- t[58644] = 26
      "0011010" when "01110010100010101", -- t[58645] = 26
      "0011010" when "01110010100010110", -- t[58646] = 26
      "0011010" when "01110010100010111", -- t[58647] = 26
      "0011010" when "01110010100011000", -- t[58648] = 26
      "0011010" when "01110010100011001", -- t[58649] = 26
      "0011010" when "01110010100011010", -- t[58650] = 26
      "0011010" when "01110010100011011", -- t[58651] = 26
      "0011010" when "01110010100011100", -- t[58652] = 26
      "0011010" when "01110010100011101", -- t[58653] = 26
      "0011010" when "01110010100011110", -- t[58654] = 26
      "0011010" when "01110010100011111", -- t[58655] = 26
      "0011010" when "01110010100100000", -- t[58656] = 26
      "0011010" when "01110010100100001", -- t[58657] = 26
      "0011010" when "01110010100100010", -- t[58658] = 26
      "0011010" when "01110010100100011", -- t[58659] = 26
      "0011010" when "01110010100100100", -- t[58660] = 26
      "0011010" when "01110010100100101", -- t[58661] = 26
      "0011010" when "01110010100100110", -- t[58662] = 26
      "0011010" when "01110010100100111", -- t[58663] = 26
      "0011010" when "01110010100101000", -- t[58664] = 26
      "0011010" when "01110010100101001", -- t[58665] = 26
      "0011010" when "01110010100101010", -- t[58666] = 26
      "0011010" when "01110010100101011", -- t[58667] = 26
      "0011010" when "01110010100101100", -- t[58668] = 26
      "0011010" when "01110010100101101", -- t[58669] = 26
      "0011010" when "01110010100101110", -- t[58670] = 26
      "0011010" when "01110010100101111", -- t[58671] = 26
      "0011010" when "01110010100110000", -- t[58672] = 26
      "0011010" when "01110010100110001", -- t[58673] = 26
      "0011010" when "01110010100110010", -- t[58674] = 26
      "0011010" when "01110010100110011", -- t[58675] = 26
      "0011010" when "01110010100110100", -- t[58676] = 26
      "0011010" when "01110010100110101", -- t[58677] = 26
      "0011010" when "01110010100110110", -- t[58678] = 26
      "0011010" when "01110010100110111", -- t[58679] = 26
      "0011010" when "01110010100111000", -- t[58680] = 26
      "0011010" when "01110010100111001", -- t[58681] = 26
      "0011010" when "01110010100111010", -- t[58682] = 26
      "0011010" when "01110010100111011", -- t[58683] = 26
      "0011010" when "01110010100111100", -- t[58684] = 26
      "0011010" when "01110010100111101", -- t[58685] = 26
      "0011010" when "01110010100111110", -- t[58686] = 26
      "0011010" when "01110010100111111", -- t[58687] = 26
      "0011010" when "01110010101000000", -- t[58688] = 26
      "0011010" when "01110010101000001", -- t[58689] = 26
      "0011010" when "01110010101000010", -- t[58690] = 26
      "0011010" when "01110010101000011", -- t[58691] = 26
      "0011010" when "01110010101000100", -- t[58692] = 26
      "0011010" when "01110010101000101", -- t[58693] = 26
      "0011010" when "01110010101000110", -- t[58694] = 26
      "0011010" when "01110010101000111", -- t[58695] = 26
      "0011010" when "01110010101001000", -- t[58696] = 26
      "0011010" when "01110010101001001", -- t[58697] = 26
      "0011010" when "01110010101001010", -- t[58698] = 26
      "0011010" when "01110010101001011", -- t[58699] = 26
      "0011010" when "01110010101001100", -- t[58700] = 26
      "0011010" when "01110010101001101", -- t[58701] = 26
      "0011010" when "01110010101001110", -- t[58702] = 26
      "0011010" when "01110010101001111", -- t[58703] = 26
      "0011010" when "01110010101010000", -- t[58704] = 26
      "0011010" when "01110010101010001", -- t[58705] = 26
      "0011010" when "01110010101010010", -- t[58706] = 26
      "0011010" when "01110010101010011", -- t[58707] = 26
      "0011010" when "01110010101010100", -- t[58708] = 26
      "0011010" when "01110010101010101", -- t[58709] = 26
      "0011010" when "01110010101010110", -- t[58710] = 26
      "0011010" when "01110010101010111", -- t[58711] = 26
      "0011010" when "01110010101011000", -- t[58712] = 26
      "0011010" when "01110010101011001", -- t[58713] = 26
      "0011010" when "01110010101011010", -- t[58714] = 26
      "0011010" when "01110010101011011", -- t[58715] = 26
      "0011010" when "01110010101011100", -- t[58716] = 26
      "0011010" when "01110010101011101", -- t[58717] = 26
      "0011010" when "01110010101011110", -- t[58718] = 26
      "0011010" when "01110010101011111", -- t[58719] = 26
      "0011010" when "01110010101100000", -- t[58720] = 26
      "0011010" when "01110010101100001", -- t[58721] = 26
      "0011010" when "01110010101100010", -- t[58722] = 26
      "0011010" when "01110010101100011", -- t[58723] = 26
      "0011010" when "01110010101100100", -- t[58724] = 26
      "0011010" when "01110010101100101", -- t[58725] = 26
      "0011010" when "01110010101100110", -- t[58726] = 26
      "0011010" when "01110010101100111", -- t[58727] = 26
      "0011010" when "01110010101101000", -- t[58728] = 26
      "0011010" when "01110010101101001", -- t[58729] = 26
      "0011010" when "01110010101101010", -- t[58730] = 26
      "0011010" when "01110010101101011", -- t[58731] = 26
      "0011010" when "01110010101101100", -- t[58732] = 26
      "0011010" when "01110010101101101", -- t[58733] = 26
      "0011010" when "01110010101101110", -- t[58734] = 26
      "0011010" when "01110010101101111", -- t[58735] = 26
      "0011010" when "01110010101110000", -- t[58736] = 26
      "0011010" when "01110010101110001", -- t[58737] = 26
      "0011010" when "01110010101110010", -- t[58738] = 26
      "0011010" when "01110010101110011", -- t[58739] = 26
      "0011010" when "01110010101110100", -- t[58740] = 26
      "0011010" when "01110010101110101", -- t[58741] = 26
      "0011010" when "01110010101110110", -- t[58742] = 26
      "0011010" when "01110010101110111", -- t[58743] = 26
      "0011010" when "01110010101111000", -- t[58744] = 26
      "0011010" when "01110010101111001", -- t[58745] = 26
      "0011010" when "01110010101111010", -- t[58746] = 26
      "0011010" when "01110010101111011", -- t[58747] = 26
      "0011010" when "01110010101111100", -- t[58748] = 26
      "0011010" when "01110010101111101", -- t[58749] = 26
      "0011010" when "01110010101111110", -- t[58750] = 26
      "0011010" when "01110010101111111", -- t[58751] = 26
      "0011010" when "01110010110000000", -- t[58752] = 26
      "0011010" when "01110010110000001", -- t[58753] = 26
      "0011010" when "01110010110000010", -- t[58754] = 26
      "0011010" when "01110010110000011", -- t[58755] = 26
      "0011010" when "01110010110000100", -- t[58756] = 26
      "0011010" when "01110010110000101", -- t[58757] = 26
      "0011010" when "01110010110000110", -- t[58758] = 26
      "0011010" when "01110010110000111", -- t[58759] = 26
      "0011010" when "01110010110001000", -- t[58760] = 26
      "0011010" when "01110010110001001", -- t[58761] = 26
      "0011010" when "01110010110001010", -- t[58762] = 26
      "0011010" when "01110010110001011", -- t[58763] = 26
      "0011010" when "01110010110001100", -- t[58764] = 26
      "0011010" when "01110010110001101", -- t[58765] = 26
      "0011010" when "01110010110001110", -- t[58766] = 26
      "0011010" when "01110010110001111", -- t[58767] = 26
      "0011010" when "01110010110010000", -- t[58768] = 26
      "0011010" when "01110010110010001", -- t[58769] = 26
      "0011010" when "01110010110010010", -- t[58770] = 26
      "0011010" when "01110010110010011", -- t[58771] = 26
      "0011010" when "01110010110010100", -- t[58772] = 26
      "0011010" when "01110010110010101", -- t[58773] = 26
      "0011010" when "01110010110010110", -- t[58774] = 26
      "0011010" when "01110010110010111", -- t[58775] = 26
      "0011010" when "01110010110011000", -- t[58776] = 26
      "0011010" when "01110010110011001", -- t[58777] = 26
      "0011010" when "01110010110011010", -- t[58778] = 26
      "0011010" when "01110010110011011", -- t[58779] = 26
      "0011010" when "01110010110011100", -- t[58780] = 26
      "0011010" when "01110010110011101", -- t[58781] = 26
      "0011010" when "01110010110011110", -- t[58782] = 26
      "0011010" when "01110010110011111", -- t[58783] = 26
      "0011010" when "01110010110100000", -- t[58784] = 26
      "0011010" when "01110010110100001", -- t[58785] = 26
      "0011010" when "01110010110100010", -- t[58786] = 26
      "0011010" when "01110010110100011", -- t[58787] = 26
      "0011010" when "01110010110100100", -- t[58788] = 26
      "0011010" when "01110010110100101", -- t[58789] = 26
      "0011010" when "01110010110100110", -- t[58790] = 26
      "0011010" when "01110010110100111", -- t[58791] = 26
      "0011010" when "01110010110101000", -- t[58792] = 26
      "0011010" when "01110010110101001", -- t[58793] = 26
      "0011010" when "01110010110101010", -- t[58794] = 26
      "0011010" when "01110010110101011", -- t[58795] = 26
      "0011010" when "01110010110101100", -- t[58796] = 26
      "0011010" when "01110010110101101", -- t[58797] = 26
      "0011010" when "01110010110101110", -- t[58798] = 26
      "0011010" when "01110010110101111", -- t[58799] = 26
      "0011010" when "01110010110110000", -- t[58800] = 26
      "0011010" when "01110010110110001", -- t[58801] = 26
      "0011010" when "01110010110110010", -- t[58802] = 26
      "0011010" when "01110010110110011", -- t[58803] = 26
      "0011010" when "01110010110110100", -- t[58804] = 26
      "0011010" when "01110010110110101", -- t[58805] = 26
      "0011010" when "01110010110110110", -- t[58806] = 26
      "0011010" when "01110010110110111", -- t[58807] = 26
      "0011010" when "01110010110111000", -- t[58808] = 26
      "0011010" when "01110010110111001", -- t[58809] = 26
      "0011010" when "01110010110111010", -- t[58810] = 26
      "0011010" when "01110010110111011", -- t[58811] = 26
      "0011010" when "01110010110111100", -- t[58812] = 26
      "0011010" when "01110010110111101", -- t[58813] = 26
      "0011010" when "01110010110111110", -- t[58814] = 26
      "0011010" when "01110010110111111", -- t[58815] = 26
      "0011010" when "01110010111000000", -- t[58816] = 26
      "0011010" when "01110010111000001", -- t[58817] = 26
      "0011010" when "01110010111000010", -- t[58818] = 26
      "0011010" when "01110010111000011", -- t[58819] = 26
      "0011010" when "01110010111000100", -- t[58820] = 26
      "0011010" when "01110010111000101", -- t[58821] = 26
      "0011010" when "01110010111000110", -- t[58822] = 26
      "0011010" when "01110010111000111", -- t[58823] = 26
      "0011010" when "01110010111001000", -- t[58824] = 26
      "0011010" when "01110010111001001", -- t[58825] = 26
      "0011010" when "01110010111001010", -- t[58826] = 26
      "0011010" when "01110010111001011", -- t[58827] = 26
      "0011010" when "01110010111001100", -- t[58828] = 26
      "0011010" when "01110010111001101", -- t[58829] = 26
      "0011010" when "01110010111001110", -- t[58830] = 26
      "0011010" when "01110010111001111", -- t[58831] = 26
      "0011010" when "01110010111010000", -- t[58832] = 26
      "0011010" when "01110010111010001", -- t[58833] = 26
      "0011010" when "01110010111010010", -- t[58834] = 26
      "0011010" when "01110010111010011", -- t[58835] = 26
      "0011010" when "01110010111010100", -- t[58836] = 26
      "0011010" when "01110010111010101", -- t[58837] = 26
      "0011010" when "01110010111010110", -- t[58838] = 26
      "0011010" when "01110010111010111", -- t[58839] = 26
      "0011010" when "01110010111011000", -- t[58840] = 26
      "0011010" when "01110010111011001", -- t[58841] = 26
      "0011010" when "01110010111011010", -- t[58842] = 26
      "0011010" when "01110010111011011", -- t[58843] = 26
      "0011010" when "01110010111011100", -- t[58844] = 26
      "0011010" when "01110010111011101", -- t[58845] = 26
      "0011010" when "01110010111011110", -- t[58846] = 26
      "0011010" when "01110010111011111", -- t[58847] = 26
      "0011010" when "01110010111100000", -- t[58848] = 26
      "0011010" when "01110010111100001", -- t[58849] = 26
      "0011010" when "01110010111100010", -- t[58850] = 26
      "0011010" when "01110010111100011", -- t[58851] = 26
      "0011010" when "01110010111100100", -- t[58852] = 26
      "0011010" when "01110010111100101", -- t[58853] = 26
      "0011010" when "01110010111100110", -- t[58854] = 26
      "0011010" when "01110010111100111", -- t[58855] = 26
      "0011010" when "01110010111101000", -- t[58856] = 26
      "0011010" when "01110010111101001", -- t[58857] = 26
      "0011010" when "01110010111101010", -- t[58858] = 26
      "0011010" when "01110010111101011", -- t[58859] = 26
      "0011010" when "01110010111101100", -- t[58860] = 26
      "0011010" when "01110010111101101", -- t[58861] = 26
      "0011010" when "01110010111101110", -- t[58862] = 26
      "0011010" when "01110010111101111", -- t[58863] = 26
      "0011010" when "01110010111110000", -- t[58864] = 26
      "0011010" when "01110010111110001", -- t[58865] = 26
      "0011010" when "01110010111110010", -- t[58866] = 26
      "0011010" when "01110010111110011", -- t[58867] = 26
      "0011010" when "01110010111110100", -- t[58868] = 26
      "0011010" when "01110010111110101", -- t[58869] = 26
      "0011010" when "01110010111110110", -- t[58870] = 26
      "0011010" when "01110010111110111", -- t[58871] = 26
      "0011010" when "01110010111111000", -- t[58872] = 26
      "0011010" when "01110010111111001", -- t[58873] = 26
      "0011010" when "01110010111111010", -- t[58874] = 26
      "0011010" when "01110010111111011", -- t[58875] = 26
      "0011010" when "01110010111111100", -- t[58876] = 26
      "0011010" when "01110010111111101", -- t[58877] = 26
      "0011010" when "01110010111111110", -- t[58878] = 26
      "0011010" when "01110010111111111", -- t[58879] = 26
      "0011010" when "01110011000000000", -- t[58880] = 26
      "0011010" when "01110011000000001", -- t[58881] = 26
      "0011010" when "01110011000000010", -- t[58882] = 26
      "0011010" when "01110011000000011", -- t[58883] = 26
      "0011010" when "01110011000000100", -- t[58884] = 26
      "0011010" when "01110011000000101", -- t[58885] = 26
      "0011010" when "01110011000000110", -- t[58886] = 26
      "0011010" when "01110011000000111", -- t[58887] = 26
      "0011010" when "01110011000001000", -- t[58888] = 26
      "0011010" when "01110011000001001", -- t[58889] = 26
      "0011010" when "01110011000001010", -- t[58890] = 26
      "0011010" when "01110011000001011", -- t[58891] = 26
      "0011010" when "01110011000001100", -- t[58892] = 26
      "0011010" when "01110011000001101", -- t[58893] = 26
      "0011010" when "01110011000001110", -- t[58894] = 26
      "0011010" when "01110011000001111", -- t[58895] = 26
      "0011010" when "01110011000010000", -- t[58896] = 26
      "0011010" when "01110011000010001", -- t[58897] = 26
      "0011010" when "01110011000010010", -- t[58898] = 26
      "0011010" when "01110011000010011", -- t[58899] = 26
      "0011010" when "01110011000010100", -- t[58900] = 26
      "0011010" when "01110011000010101", -- t[58901] = 26
      "0011010" when "01110011000010110", -- t[58902] = 26
      "0011010" when "01110011000010111", -- t[58903] = 26
      "0011010" when "01110011000011000", -- t[58904] = 26
      "0011010" when "01110011000011001", -- t[58905] = 26
      "0011010" when "01110011000011010", -- t[58906] = 26
      "0011010" when "01110011000011011", -- t[58907] = 26
      "0011010" when "01110011000011100", -- t[58908] = 26
      "0011010" when "01110011000011101", -- t[58909] = 26
      "0011010" when "01110011000011110", -- t[58910] = 26
      "0011010" when "01110011000011111", -- t[58911] = 26
      "0011010" when "01110011000100000", -- t[58912] = 26
      "0011010" when "01110011000100001", -- t[58913] = 26
      "0011010" when "01110011000100010", -- t[58914] = 26
      "0011010" when "01110011000100011", -- t[58915] = 26
      "0011010" when "01110011000100100", -- t[58916] = 26
      "0011010" when "01110011000100101", -- t[58917] = 26
      "0011010" when "01110011000100110", -- t[58918] = 26
      "0011010" when "01110011000100111", -- t[58919] = 26
      "0011010" when "01110011000101000", -- t[58920] = 26
      "0011010" when "01110011000101001", -- t[58921] = 26
      "0011010" when "01110011000101010", -- t[58922] = 26
      "0011010" when "01110011000101011", -- t[58923] = 26
      "0011010" when "01110011000101100", -- t[58924] = 26
      "0011010" when "01110011000101101", -- t[58925] = 26
      "0011010" when "01110011000101110", -- t[58926] = 26
      "0011010" when "01110011000101111", -- t[58927] = 26
      "0011010" when "01110011000110000", -- t[58928] = 26
      "0011010" when "01110011000110001", -- t[58929] = 26
      "0011010" when "01110011000110010", -- t[58930] = 26
      "0011010" when "01110011000110011", -- t[58931] = 26
      "0011010" when "01110011000110100", -- t[58932] = 26
      "0011010" when "01110011000110101", -- t[58933] = 26
      "0011010" when "01110011000110110", -- t[58934] = 26
      "0011010" when "01110011000110111", -- t[58935] = 26
      "0011010" when "01110011000111000", -- t[58936] = 26
      "0011010" when "01110011000111001", -- t[58937] = 26
      "0011010" when "01110011000111010", -- t[58938] = 26
      "0011010" when "01110011000111011", -- t[58939] = 26
      "0011010" when "01110011000111100", -- t[58940] = 26
      "0011010" when "01110011000111101", -- t[58941] = 26
      "0011010" when "01110011000111110", -- t[58942] = 26
      "0011010" when "01110011000111111", -- t[58943] = 26
      "0011010" when "01110011001000000", -- t[58944] = 26
      "0011010" when "01110011001000001", -- t[58945] = 26
      "0011010" when "01110011001000010", -- t[58946] = 26
      "0011010" when "01110011001000011", -- t[58947] = 26
      "0011010" when "01110011001000100", -- t[58948] = 26
      "0011010" when "01110011001000101", -- t[58949] = 26
      "0011010" when "01110011001000110", -- t[58950] = 26
      "0011010" when "01110011001000111", -- t[58951] = 26
      "0011010" when "01110011001001000", -- t[58952] = 26
      "0011010" when "01110011001001001", -- t[58953] = 26
      "0011010" when "01110011001001010", -- t[58954] = 26
      "0011010" when "01110011001001011", -- t[58955] = 26
      "0011010" when "01110011001001100", -- t[58956] = 26
      "0011010" when "01110011001001101", -- t[58957] = 26
      "0011010" when "01110011001001110", -- t[58958] = 26
      "0011010" when "01110011001001111", -- t[58959] = 26
      "0011010" when "01110011001010000", -- t[58960] = 26
      "0011010" when "01110011001010001", -- t[58961] = 26
      "0011010" when "01110011001010010", -- t[58962] = 26
      "0011011" when "01110011001010011", -- t[58963] = 27
      "0011011" when "01110011001010100", -- t[58964] = 27
      "0011011" when "01110011001010101", -- t[58965] = 27
      "0011011" when "01110011001010110", -- t[58966] = 27
      "0011011" when "01110011001010111", -- t[58967] = 27
      "0011011" when "01110011001011000", -- t[58968] = 27
      "0011011" when "01110011001011001", -- t[58969] = 27
      "0011011" when "01110011001011010", -- t[58970] = 27
      "0011011" when "01110011001011011", -- t[58971] = 27
      "0011011" when "01110011001011100", -- t[58972] = 27
      "0011011" when "01110011001011101", -- t[58973] = 27
      "0011011" when "01110011001011110", -- t[58974] = 27
      "0011011" when "01110011001011111", -- t[58975] = 27
      "0011011" when "01110011001100000", -- t[58976] = 27
      "0011011" when "01110011001100001", -- t[58977] = 27
      "0011011" when "01110011001100010", -- t[58978] = 27
      "0011011" when "01110011001100011", -- t[58979] = 27
      "0011011" when "01110011001100100", -- t[58980] = 27
      "0011011" when "01110011001100101", -- t[58981] = 27
      "0011011" when "01110011001100110", -- t[58982] = 27
      "0011011" when "01110011001100111", -- t[58983] = 27
      "0011011" when "01110011001101000", -- t[58984] = 27
      "0011011" when "01110011001101001", -- t[58985] = 27
      "0011011" when "01110011001101010", -- t[58986] = 27
      "0011011" when "01110011001101011", -- t[58987] = 27
      "0011011" when "01110011001101100", -- t[58988] = 27
      "0011011" when "01110011001101101", -- t[58989] = 27
      "0011011" when "01110011001101110", -- t[58990] = 27
      "0011011" when "01110011001101111", -- t[58991] = 27
      "0011011" when "01110011001110000", -- t[58992] = 27
      "0011011" when "01110011001110001", -- t[58993] = 27
      "0011011" when "01110011001110010", -- t[58994] = 27
      "0011011" when "01110011001110011", -- t[58995] = 27
      "0011011" when "01110011001110100", -- t[58996] = 27
      "0011011" when "01110011001110101", -- t[58997] = 27
      "0011011" when "01110011001110110", -- t[58998] = 27
      "0011011" when "01110011001110111", -- t[58999] = 27
      "0011011" when "01110011001111000", -- t[59000] = 27
      "0011011" when "01110011001111001", -- t[59001] = 27
      "0011011" when "01110011001111010", -- t[59002] = 27
      "0011011" when "01110011001111011", -- t[59003] = 27
      "0011011" when "01110011001111100", -- t[59004] = 27
      "0011011" when "01110011001111101", -- t[59005] = 27
      "0011011" when "01110011001111110", -- t[59006] = 27
      "0011011" when "01110011001111111", -- t[59007] = 27
      "0011011" when "01110011010000000", -- t[59008] = 27
      "0011011" when "01110011010000001", -- t[59009] = 27
      "0011011" when "01110011010000010", -- t[59010] = 27
      "0011011" when "01110011010000011", -- t[59011] = 27
      "0011011" when "01110011010000100", -- t[59012] = 27
      "0011011" when "01110011010000101", -- t[59013] = 27
      "0011011" when "01110011010000110", -- t[59014] = 27
      "0011011" when "01110011010000111", -- t[59015] = 27
      "0011011" when "01110011010001000", -- t[59016] = 27
      "0011011" when "01110011010001001", -- t[59017] = 27
      "0011011" when "01110011010001010", -- t[59018] = 27
      "0011011" when "01110011010001011", -- t[59019] = 27
      "0011011" when "01110011010001100", -- t[59020] = 27
      "0011011" when "01110011010001101", -- t[59021] = 27
      "0011011" when "01110011010001110", -- t[59022] = 27
      "0011011" when "01110011010001111", -- t[59023] = 27
      "0011011" when "01110011010010000", -- t[59024] = 27
      "0011011" when "01110011010010001", -- t[59025] = 27
      "0011011" when "01110011010010010", -- t[59026] = 27
      "0011011" when "01110011010010011", -- t[59027] = 27
      "0011011" when "01110011010010100", -- t[59028] = 27
      "0011011" when "01110011010010101", -- t[59029] = 27
      "0011011" when "01110011010010110", -- t[59030] = 27
      "0011011" when "01110011010010111", -- t[59031] = 27
      "0011011" when "01110011010011000", -- t[59032] = 27
      "0011011" when "01110011010011001", -- t[59033] = 27
      "0011011" when "01110011010011010", -- t[59034] = 27
      "0011011" when "01110011010011011", -- t[59035] = 27
      "0011011" when "01110011010011100", -- t[59036] = 27
      "0011011" when "01110011010011101", -- t[59037] = 27
      "0011011" when "01110011010011110", -- t[59038] = 27
      "0011011" when "01110011010011111", -- t[59039] = 27
      "0011011" when "01110011010100000", -- t[59040] = 27
      "0011011" when "01110011010100001", -- t[59041] = 27
      "0011011" when "01110011010100010", -- t[59042] = 27
      "0011011" when "01110011010100011", -- t[59043] = 27
      "0011011" when "01110011010100100", -- t[59044] = 27
      "0011011" when "01110011010100101", -- t[59045] = 27
      "0011011" when "01110011010100110", -- t[59046] = 27
      "0011011" when "01110011010100111", -- t[59047] = 27
      "0011011" when "01110011010101000", -- t[59048] = 27
      "0011011" when "01110011010101001", -- t[59049] = 27
      "0011011" when "01110011010101010", -- t[59050] = 27
      "0011011" when "01110011010101011", -- t[59051] = 27
      "0011011" when "01110011010101100", -- t[59052] = 27
      "0011011" when "01110011010101101", -- t[59053] = 27
      "0011011" when "01110011010101110", -- t[59054] = 27
      "0011011" when "01110011010101111", -- t[59055] = 27
      "0011011" when "01110011010110000", -- t[59056] = 27
      "0011011" when "01110011010110001", -- t[59057] = 27
      "0011011" when "01110011010110010", -- t[59058] = 27
      "0011011" when "01110011010110011", -- t[59059] = 27
      "0011011" when "01110011010110100", -- t[59060] = 27
      "0011011" when "01110011010110101", -- t[59061] = 27
      "0011011" when "01110011010110110", -- t[59062] = 27
      "0011011" when "01110011010110111", -- t[59063] = 27
      "0011011" when "01110011010111000", -- t[59064] = 27
      "0011011" when "01110011010111001", -- t[59065] = 27
      "0011011" when "01110011010111010", -- t[59066] = 27
      "0011011" when "01110011010111011", -- t[59067] = 27
      "0011011" when "01110011010111100", -- t[59068] = 27
      "0011011" when "01110011010111101", -- t[59069] = 27
      "0011011" when "01110011010111110", -- t[59070] = 27
      "0011011" when "01110011010111111", -- t[59071] = 27
      "0011011" when "01110011011000000", -- t[59072] = 27
      "0011011" when "01110011011000001", -- t[59073] = 27
      "0011011" when "01110011011000010", -- t[59074] = 27
      "0011011" when "01110011011000011", -- t[59075] = 27
      "0011011" when "01110011011000100", -- t[59076] = 27
      "0011011" when "01110011011000101", -- t[59077] = 27
      "0011011" when "01110011011000110", -- t[59078] = 27
      "0011011" when "01110011011000111", -- t[59079] = 27
      "0011011" when "01110011011001000", -- t[59080] = 27
      "0011011" when "01110011011001001", -- t[59081] = 27
      "0011011" when "01110011011001010", -- t[59082] = 27
      "0011011" when "01110011011001011", -- t[59083] = 27
      "0011011" when "01110011011001100", -- t[59084] = 27
      "0011011" when "01110011011001101", -- t[59085] = 27
      "0011011" when "01110011011001110", -- t[59086] = 27
      "0011011" when "01110011011001111", -- t[59087] = 27
      "0011011" when "01110011011010000", -- t[59088] = 27
      "0011011" when "01110011011010001", -- t[59089] = 27
      "0011011" when "01110011011010010", -- t[59090] = 27
      "0011011" when "01110011011010011", -- t[59091] = 27
      "0011011" when "01110011011010100", -- t[59092] = 27
      "0011011" when "01110011011010101", -- t[59093] = 27
      "0011011" when "01110011011010110", -- t[59094] = 27
      "0011011" when "01110011011010111", -- t[59095] = 27
      "0011011" when "01110011011011000", -- t[59096] = 27
      "0011011" when "01110011011011001", -- t[59097] = 27
      "0011011" when "01110011011011010", -- t[59098] = 27
      "0011011" when "01110011011011011", -- t[59099] = 27
      "0011011" when "01110011011011100", -- t[59100] = 27
      "0011011" when "01110011011011101", -- t[59101] = 27
      "0011011" when "01110011011011110", -- t[59102] = 27
      "0011011" when "01110011011011111", -- t[59103] = 27
      "0011011" when "01110011011100000", -- t[59104] = 27
      "0011011" when "01110011011100001", -- t[59105] = 27
      "0011011" when "01110011011100010", -- t[59106] = 27
      "0011011" when "01110011011100011", -- t[59107] = 27
      "0011011" when "01110011011100100", -- t[59108] = 27
      "0011011" when "01110011011100101", -- t[59109] = 27
      "0011011" when "01110011011100110", -- t[59110] = 27
      "0011011" when "01110011011100111", -- t[59111] = 27
      "0011011" when "01110011011101000", -- t[59112] = 27
      "0011011" when "01110011011101001", -- t[59113] = 27
      "0011011" when "01110011011101010", -- t[59114] = 27
      "0011011" when "01110011011101011", -- t[59115] = 27
      "0011011" when "01110011011101100", -- t[59116] = 27
      "0011011" when "01110011011101101", -- t[59117] = 27
      "0011011" when "01110011011101110", -- t[59118] = 27
      "0011011" when "01110011011101111", -- t[59119] = 27
      "0011011" when "01110011011110000", -- t[59120] = 27
      "0011011" when "01110011011110001", -- t[59121] = 27
      "0011011" when "01110011011110010", -- t[59122] = 27
      "0011011" when "01110011011110011", -- t[59123] = 27
      "0011011" when "01110011011110100", -- t[59124] = 27
      "0011011" when "01110011011110101", -- t[59125] = 27
      "0011011" when "01110011011110110", -- t[59126] = 27
      "0011011" when "01110011011110111", -- t[59127] = 27
      "0011011" when "01110011011111000", -- t[59128] = 27
      "0011011" when "01110011011111001", -- t[59129] = 27
      "0011011" when "01110011011111010", -- t[59130] = 27
      "0011011" when "01110011011111011", -- t[59131] = 27
      "0011011" when "01110011011111100", -- t[59132] = 27
      "0011011" when "01110011011111101", -- t[59133] = 27
      "0011011" when "01110011011111110", -- t[59134] = 27
      "0011011" when "01110011011111111", -- t[59135] = 27
      "0011011" when "01110011100000000", -- t[59136] = 27
      "0011011" when "01110011100000001", -- t[59137] = 27
      "0011011" when "01110011100000010", -- t[59138] = 27
      "0011011" when "01110011100000011", -- t[59139] = 27
      "0011011" when "01110011100000100", -- t[59140] = 27
      "0011011" when "01110011100000101", -- t[59141] = 27
      "0011011" when "01110011100000110", -- t[59142] = 27
      "0011011" when "01110011100000111", -- t[59143] = 27
      "0011011" when "01110011100001000", -- t[59144] = 27
      "0011011" when "01110011100001001", -- t[59145] = 27
      "0011011" when "01110011100001010", -- t[59146] = 27
      "0011011" when "01110011100001011", -- t[59147] = 27
      "0011011" when "01110011100001100", -- t[59148] = 27
      "0011011" when "01110011100001101", -- t[59149] = 27
      "0011011" when "01110011100001110", -- t[59150] = 27
      "0011011" when "01110011100001111", -- t[59151] = 27
      "0011011" when "01110011100010000", -- t[59152] = 27
      "0011011" when "01110011100010001", -- t[59153] = 27
      "0011011" when "01110011100010010", -- t[59154] = 27
      "0011011" when "01110011100010011", -- t[59155] = 27
      "0011011" when "01110011100010100", -- t[59156] = 27
      "0011011" when "01110011100010101", -- t[59157] = 27
      "0011011" when "01110011100010110", -- t[59158] = 27
      "0011011" when "01110011100010111", -- t[59159] = 27
      "0011011" when "01110011100011000", -- t[59160] = 27
      "0011011" when "01110011100011001", -- t[59161] = 27
      "0011011" when "01110011100011010", -- t[59162] = 27
      "0011011" when "01110011100011011", -- t[59163] = 27
      "0011011" when "01110011100011100", -- t[59164] = 27
      "0011011" when "01110011100011101", -- t[59165] = 27
      "0011011" when "01110011100011110", -- t[59166] = 27
      "0011011" when "01110011100011111", -- t[59167] = 27
      "0011011" when "01110011100100000", -- t[59168] = 27
      "0011011" when "01110011100100001", -- t[59169] = 27
      "0011011" when "01110011100100010", -- t[59170] = 27
      "0011011" when "01110011100100011", -- t[59171] = 27
      "0011011" when "01110011100100100", -- t[59172] = 27
      "0011011" when "01110011100100101", -- t[59173] = 27
      "0011011" when "01110011100100110", -- t[59174] = 27
      "0011011" when "01110011100100111", -- t[59175] = 27
      "0011011" when "01110011100101000", -- t[59176] = 27
      "0011011" when "01110011100101001", -- t[59177] = 27
      "0011011" when "01110011100101010", -- t[59178] = 27
      "0011011" when "01110011100101011", -- t[59179] = 27
      "0011011" when "01110011100101100", -- t[59180] = 27
      "0011011" when "01110011100101101", -- t[59181] = 27
      "0011011" when "01110011100101110", -- t[59182] = 27
      "0011011" when "01110011100101111", -- t[59183] = 27
      "0011011" when "01110011100110000", -- t[59184] = 27
      "0011011" when "01110011100110001", -- t[59185] = 27
      "0011011" when "01110011100110010", -- t[59186] = 27
      "0011011" when "01110011100110011", -- t[59187] = 27
      "0011011" when "01110011100110100", -- t[59188] = 27
      "0011011" when "01110011100110101", -- t[59189] = 27
      "0011011" when "01110011100110110", -- t[59190] = 27
      "0011011" when "01110011100110111", -- t[59191] = 27
      "0011011" when "01110011100111000", -- t[59192] = 27
      "0011011" when "01110011100111001", -- t[59193] = 27
      "0011011" when "01110011100111010", -- t[59194] = 27
      "0011011" when "01110011100111011", -- t[59195] = 27
      "0011011" when "01110011100111100", -- t[59196] = 27
      "0011011" when "01110011100111101", -- t[59197] = 27
      "0011011" when "01110011100111110", -- t[59198] = 27
      "0011011" when "01110011100111111", -- t[59199] = 27
      "0011011" when "01110011101000000", -- t[59200] = 27
      "0011011" when "01110011101000001", -- t[59201] = 27
      "0011011" when "01110011101000010", -- t[59202] = 27
      "0011011" when "01110011101000011", -- t[59203] = 27
      "0011011" when "01110011101000100", -- t[59204] = 27
      "0011011" when "01110011101000101", -- t[59205] = 27
      "0011011" when "01110011101000110", -- t[59206] = 27
      "0011011" when "01110011101000111", -- t[59207] = 27
      "0011011" when "01110011101001000", -- t[59208] = 27
      "0011011" when "01110011101001001", -- t[59209] = 27
      "0011011" when "01110011101001010", -- t[59210] = 27
      "0011011" when "01110011101001011", -- t[59211] = 27
      "0011011" when "01110011101001100", -- t[59212] = 27
      "0011011" when "01110011101001101", -- t[59213] = 27
      "0011011" when "01110011101001110", -- t[59214] = 27
      "0011011" when "01110011101001111", -- t[59215] = 27
      "0011011" when "01110011101010000", -- t[59216] = 27
      "0011011" when "01110011101010001", -- t[59217] = 27
      "0011011" when "01110011101010010", -- t[59218] = 27
      "0011011" when "01110011101010011", -- t[59219] = 27
      "0011011" when "01110011101010100", -- t[59220] = 27
      "0011011" when "01110011101010101", -- t[59221] = 27
      "0011011" when "01110011101010110", -- t[59222] = 27
      "0011011" when "01110011101010111", -- t[59223] = 27
      "0011011" when "01110011101011000", -- t[59224] = 27
      "0011011" when "01110011101011001", -- t[59225] = 27
      "0011011" when "01110011101011010", -- t[59226] = 27
      "0011011" when "01110011101011011", -- t[59227] = 27
      "0011011" when "01110011101011100", -- t[59228] = 27
      "0011011" when "01110011101011101", -- t[59229] = 27
      "0011011" when "01110011101011110", -- t[59230] = 27
      "0011011" when "01110011101011111", -- t[59231] = 27
      "0011011" when "01110011101100000", -- t[59232] = 27
      "0011011" when "01110011101100001", -- t[59233] = 27
      "0011011" when "01110011101100010", -- t[59234] = 27
      "0011011" when "01110011101100011", -- t[59235] = 27
      "0011011" when "01110011101100100", -- t[59236] = 27
      "0011011" when "01110011101100101", -- t[59237] = 27
      "0011011" when "01110011101100110", -- t[59238] = 27
      "0011011" when "01110011101100111", -- t[59239] = 27
      "0011011" when "01110011101101000", -- t[59240] = 27
      "0011011" when "01110011101101001", -- t[59241] = 27
      "0011011" when "01110011101101010", -- t[59242] = 27
      "0011011" when "01110011101101011", -- t[59243] = 27
      "0011011" when "01110011101101100", -- t[59244] = 27
      "0011011" when "01110011101101101", -- t[59245] = 27
      "0011011" when "01110011101101110", -- t[59246] = 27
      "0011011" when "01110011101101111", -- t[59247] = 27
      "0011011" when "01110011101110000", -- t[59248] = 27
      "0011011" when "01110011101110001", -- t[59249] = 27
      "0011011" when "01110011101110010", -- t[59250] = 27
      "0011011" when "01110011101110011", -- t[59251] = 27
      "0011011" when "01110011101110100", -- t[59252] = 27
      "0011011" when "01110011101110101", -- t[59253] = 27
      "0011011" when "01110011101110110", -- t[59254] = 27
      "0011011" when "01110011101110111", -- t[59255] = 27
      "0011011" when "01110011101111000", -- t[59256] = 27
      "0011011" when "01110011101111001", -- t[59257] = 27
      "0011011" when "01110011101111010", -- t[59258] = 27
      "0011011" when "01110011101111011", -- t[59259] = 27
      "0011011" when "01110011101111100", -- t[59260] = 27
      "0011011" when "01110011101111101", -- t[59261] = 27
      "0011011" when "01110011101111110", -- t[59262] = 27
      "0011011" when "01110011101111111", -- t[59263] = 27
      "0011011" when "01110011110000000", -- t[59264] = 27
      "0011011" when "01110011110000001", -- t[59265] = 27
      "0011011" when "01110011110000010", -- t[59266] = 27
      "0011011" when "01110011110000011", -- t[59267] = 27
      "0011011" when "01110011110000100", -- t[59268] = 27
      "0011011" when "01110011110000101", -- t[59269] = 27
      "0011011" when "01110011110000110", -- t[59270] = 27
      "0011011" when "01110011110000111", -- t[59271] = 27
      "0011011" when "01110011110001000", -- t[59272] = 27
      "0011011" when "01110011110001001", -- t[59273] = 27
      "0011011" when "01110011110001010", -- t[59274] = 27
      "0011011" when "01110011110001011", -- t[59275] = 27
      "0011011" when "01110011110001100", -- t[59276] = 27
      "0011011" when "01110011110001101", -- t[59277] = 27
      "0011011" when "01110011110001110", -- t[59278] = 27
      "0011011" when "01110011110001111", -- t[59279] = 27
      "0011011" when "01110011110010000", -- t[59280] = 27
      "0011011" when "01110011110010001", -- t[59281] = 27
      "0011011" when "01110011110010010", -- t[59282] = 27
      "0011011" when "01110011110010011", -- t[59283] = 27
      "0011011" when "01110011110010100", -- t[59284] = 27
      "0011011" when "01110011110010101", -- t[59285] = 27
      "0011011" when "01110011110010110", -- t[59286] = 27
      "0011011" when "01110011110010111", -- t[59287] = 27
      "0011011" when "01110011110011000", -- t[59288] = 27
      "0011011" when "01110011110011001", -- t[59289] = 27
      "0011011" when "01110011110011010", -- t[59290] = 27
      "0011011" when "01110011110011011", -- t[59291] = 27
      "0011011" when "01110011110011100", -- t[59292] = 27
      "0011011" when "01110011110011101", -- t[59293] = 27
      "0011011" when "01110011110011110", -- t[59294] = 27
      "0011011" when "01110011110011111", -- t[59295] = 27
      "0011011" when "01110011110100000", -- t[59296] = 27
      "0011011" when "01110011110100001", -- t[59297] = 27
      "0011011" when "01110011110100010", -- t[59298] = 27
      "0011011" when "01110011110100011", -- t[59299] = 27
      "0011011" when "01110011110100100", -- t[59300] = 27
      "0011011" when "01110011110100101", -- t[59301] = 27
      "0011011" when "01110011110100110", -- t[59302] = 27
      "0011011" when "01110011110100111", -- t[59303] = 27
      "0011011" when "01110011110101000", -- t[59304] = 27
      "0011011" when "01110011110101001", -- t[59305] = 27
      "0011011" when "01110011110101010", -- t[59306] = 27
      "0011011" when "01110011110101011", -- t[59307] = 27
      "0011011" when "01110011110101100", -- t[59308] = 27
      "0011011" when "01110011110101101", -- t[59309] = 27
      "0011011" when "01110011110101110", -- t[59310] = 27
      "0011011" when "01110011110101111", -- t[59311] = 27
      "0011011" when "01110011110110000", -- t[59312] = 27
      "0011011" when "01110011110110001", -- t[59313] = 27
      "0011011" when "01110011110110010", -- t[59314] = 27
      "0011011" when "01110011110110011", -- t[59315] = 27
      "0011011" when "01110011110110100", -- t[59316] = 27
      "0011011" when "01110011110110101", -- t[59317] = 27
      "0011011" when "01110011110110110", -- t[59318] = 27
      "0011011" when "01110011110110111", -- t[59319] = 27
      "0011011" when "01110011110111000", -- t[59320] = 27
      "0011011" when "01110011110111001", -- t[59321] = 27
      "0011011" when "01110011110111010", -- t[59322] = 27
      "0011011" when "01110011110111011", -- t[59323] = 27
      "0011011" when "01110011110111100", -- t[59324] = 27
      "0011011" when "01110011110111101", -- t[59325] = 27
      "0011011" when "01110011110111110", -- t[59326] = 27
      "0011011" when "01110011110111111", -- t[59327] = 27
      "0011011" when "01110011111000000", -- t[59328] = 27
      "0011011" when "01110011111000001", -- t[59329] = 27
      "0011011" when "01110011111000010", -- t[59330] = 27
      "0011011" when "01110011111000011", -- t[59331] = 27
      "0011011" when "01110011111000100", -- t[59332] = 27
      "0011011" when "01110011111000101", -- t[59333] = 27
      "0011011" when "01110011111000110", -- t[59334] = 27
      "0011011" when "01110011111000111", -- t[59335] = 27
      "0011011" when "01110011111001000", -- t[59336] = 27
      "0011011" when "01110011111001001", -- t[59337] = 27
      "0011011" when "01110011111001010", -- t[59338] = 27
      "0011011" when "01110011111001011", -- t[59339] = 27
      "0011011" when "01110011111001100", -- t[59340] = 27
      "0011011" when "01110011111001101", -- t[59341] = 27
      "0011011" when "01110011111001110", -- t[59342] = 27
      "0011011" when "01110011111001111", -- t[59343] = 27
      "0011011" when "01110011111010000", -- t[59344] = 27
      "0011011" when "01110011111010001", -- t[59345] = 27
      "0011011" when "01110011111010010", -- t[59346] = 27
      "0011011" when "01110011111010011", -- t[59347] = 27
      "0011011" when "01110011111010100", -- t[59348] = 27
      "0011011" when "01110011111010101", -- t[59349] = 27
      "0011011" when "01110011111010110", -- t[59350] = 27
      "0011011" when "01110011111010111", -- t[59351] = 27
      "0011011" when "01110011111011000", -- t[59352] = 27
      "0011011" when "01110011111011001", -- t[59353] = 27
      "0011011" when "01110011111011010", -- t[59354] = 27
      "0011011" when "01110011111011011", -- t[59355] = 27
      "0011011" when "01110011111011100", -- t[59356] = 27
      "0011011" when "01110011111011101", -- t[59357] = 27
      "0011011" when "01110011111011110", -- t[59358] = 27
      "0011011" when "01110011111011111", -- t[59359] = 27
      "0011011" when "01110011111100000", -- t[59360] = 27
      "0011011" when "01110011111100001", -- t[59361] = 27
      "0011011" when "01110011111100010", -- t[59362] = 27
      "0011011" when "01110011111100011", -- t[59363] = 27
      "0011011" when "01110011111100100", -- t[59364] = 27
      "0011011" when "01110011111100101", -- t[59365] = 27
      "0011011" when "01110011111100110", -- t[59366] = 27
      "0011011" when "01110011111100111", -- t[59367] = 27
      "0011011" when "01110011111101000", -- t[59368] = 27
      "0011011" when "01110011111101001", -- t[59369] = 27
      "0011011" when "01110011111101010", -- t[59370] = 27
      "0011011" when "01110011111101011", -- t[59371] = 27
      "0011011" when "01110011111101100", -- t[59372] = 27
      "0011011" when "01110011111101101", -- t[59373] = 27
      "0011011" when "01110011111101110", -- t[59374] = 27
      "0011011" when "01110011111101111", -- t[59375] = 27
      "0011011" when "01110011111110000", -- t[59376] = 27
      "0011011" when "01110011111110001", -- t[59377] = 27
      "0011011" when "01110011111110010", -- t[59378] = 27
      "0011011" when "01110011111110011", -- t[59379] = 27
      "0011011" when "01110011111110100", -- t[59380] = 27
      "0011011" when "01110011111110101", -- t[59381] = 27
      "0011011" when "01110011111110110", -- t[59382] = 27
      "0011011" when "01110011111110111", -- t[59383] = 27
      "0011011" when "01110011111111000", -- t[59384] = 27
      "0011011" when "01110011111111001", -- t[59385] = 27
      "0011011" when "01110011111111010", -- t[59386] = 27
      "0011011" when "01110011111111011", -- t[59387] = 27
      "0011011" when "01110011111111100", -- t[59388] = 27
      "0011011" when "01110011111111101", -- t[59389] = 27
      "0011011" when "01110011111111110", -- t[59390] = 27
      "0011011" when "01110011111111111", -- t[59391] = 27
      "0011011" when "01110100000000000", -- t[59392] = 27
      "0011011" when "01110100000000001", -- t[59393] = 27
      "0011011" when "01110100000000010", -- t[59394] = 27
      "0011011" when "01110100000000011", -- t[59395] = 27
      "0011011" when "01110100000000100", -- t[59396] = 27
      "0011011" when "01110100000000101", -- t[59397] = 27
      "0011011" when "01110100000000110", -- t[59398] = 27
      "0011011" when "01110100000000111", -- t[59399] = 27
      "0011100" when "01110100000001000", -- t[59400] = 28
      "0011100" when "01110100000001001", -- t[59401] = 28
      "0011100" when "01110100000001010", -- t[59402] = 28
      "0011100" when "01110100000001011", -- t[59403] = 28
      "0011100" when "01110100000001100", -- t[59404] = 28
      "0011100" when "01110100000001101", -- t[59405] = 28
      "0011100" when "01110100000001110", -- t[59406] = 28
      "0011100" when "01110100000001111", -- t[59407] = 28
      "0011100" when "01110100000010000", -- t[59408] = 28
      "0011100" when "01110100000010001", -- t[59409] = 28
      "0011100" when "01110100000010010", -- t[59410] = 28
      "0011100" when "01110100000010011", -- t[59411] = 28
      "0011100" when "01110100000010100", -- t[59412] = 28
      "0011100" when "01110100000010101", -- t[59413] = 28
      "0011100" when "01110100000010110", -- t[59414] = 28
      "0011100" when "01110100000010111", -- t[59415] = 28
      "0011100" when "01110100000011000", -- t[59416] = 28
      "0011100" when "01110100000011001", -- t[59417] = 28
      "0011100" when "01110100000011010", -- t[59418] = 28
      "0011100" when "01110100000011011", -- t[59419] = 28
      "0011100" when "01110100000011100", -- t[59420] = 28
      "0011100" when "01110100000011101", -- t[59421] = 28
      "0011100" when "01110100000011110", -- t[59422] = 28
      "0011100" when "01110100000011111", -- t[59423] = 28
      "0011100" when "01110100000100000", -- t[59424] = 28
      "0011100" when "01110100000100001", -- t[59425] = 28
      "0011100" when "01110100000100010", -- t[59426] = 28
      "0011100" when "01110100000100011", -- t[59427] = 28
      "0011100" when "01110100000100100", -- t[59428] = 28
      "0011100" when "01110100000100101", -- t[59429] = 28
      "0011100" when "01110100000100110", -- t[59430] = 28
      "0011100" when "01110100000100111", -- t[59431] = 28
      "0011100" when "01110100000101000", -- t[59432] = 28
      "0011100" when "01110100000101001", -- t[59433] = 28
      "0011100" when "01110100000101010", -- t[59434] = 28
      "0011100" when "01110100000101011", -- t[59435] = 28
      "0011100" when "01110100000101100", -- t[59436] = 28
      "0011100" when "01110100000101101", -- t[59437] = 28
      "0011100" when "01110100000101110", -- t[59438] = 28
      "0011100" when "01110100000101111", -- t[59439] = 28
      "0011100" when "01110100000110000", -- t[59440] = 28
      "0011100" when "01110100000110001", -- t[59441] = 28
      "0011100" when "01110100000110010", -- t[59442] = 28
      "0011100" when "01110100000110011", -- t[59443] = 28
      "0011100" when "01110100000110100", -- t[59444] = 28
      "0011100" when "01110100000110101", -- t[59445] = 28
      "0011100" when "01110100000110110", -- t[59446] = 28
      "0011100" when "01110100000110111", -- t[59447] = 28
      "0011100" when "01110100000111000", -- t[59448] = 28
      "0011100" when "01110100000111001", -- t[59449] = 28
      "0011100" when "01110100000111010", -- t[59450] = 28
      "0011100" when "01110100000111011", -- t[59451] = 28
      "0011100" when "01110100000111100", -- t[59452] = 28
      "0011100" when "01110100000111101", -- t[59453] = 28
      "0011100" when "01110100000111110", -- t[59454] = 28
      "0011100" when "01110100000111111", -- t[59455] = 28
      "0011100" when "01110100001000000", -- t[59456] = 28
      "0011100" when "01110100001000001", -- t[59457] = 28
      "0011100" when "01110100001000010", -- t[59458] = 28
      "0011100" when "01110100001000011", -- t[59459] = 28
      "0011100" when "01110100001000100", -- t[59460] = 28
      "0011100" when "01110100001000101", -- t[59461] = 28
      "0011100" when "01110100001000110", -- t[59462] = 28
      "0011100" when "01110100001000111", -- t[59463] = 28
      "0011100" when "01110100001001000", -- t[59464] = 28
      "0011100" when "01110100001001001", -- t[59465] = 28
      "0011100" when "01110100001001010", -- t[59466] = 28
      "0011100" when "01110100001001011", -- t[59467] = 28
      "0011100" when "01110100001001100", -- t[59468] = 28
      "0011100" when "01110100001001101", -- t[59469] = 28
      "0011100" when "01110100001001110", -- t[59470] = 28
      "0011100" when "01110100001001111", -- t[59471] = 28
      "0011100" when "01110100001010000", -- t[59472] = 28
      "0011100" when "01110100001010001", -- t[59473] = 28
      "0011100" when "01110100001010010", -- t[59474] = 28
      "0011100" when "01110100001010011", -- t[59475] = 28
      "0011100" when "01110100001010100", -- t[59476] = 28
      "0011100" when "01110100001010101", -- t[59477] = 28
      "0011100" when "01110100001010110", -- t[59478] = 28
      "0011100" when "01110100001010111", -- t[59479] = 28
      "0011100" when "01110100001011000", -- t[59480] = 28
      "0011100" when "01110100001011001", -- t[59481] = 28
      "0011100" when "01110100001011010", -- t[59482] = 28
      "0011100" when "01110100001011011", -- t[59483] = 28
      "0011100" when "01110100001011100", -- t[59484] = 28
      "0011100" when "01110100001011101", -- t[59485] = 28
      "0011100" when "01110100001011110", -- t[59486] = 28
      "0011100" when "01110100001011111", -- t[59487] = 28
      "0011100" when "01110100001100000", -- t[59488] = 28
      "0011100" when "01110100001100001", -- t[59489] = 28
      "0011100" when "01110100001100010", -- t[59490] = 28
      "0011100" when "01110100001100011", -- t[59491] = 28
      "0011100" when "01110100001100100", -- t[59492] = 28
      "0011100" when "01110100001100101", -- t[59493] = 28
      "0011100" when "01110100001100110", -- t[59494] = 28
      "0011100" when "01110100001100111", -- t[59495] = 28
      "0011100" when "01110100001101000", -- t[59496] = 28
      "0011100" when "01110100001101001", -- t[59497] = 28
      "0011100" when "01110100001101010", -- t[59498] = 28
      "0011100" when "01110100001101011", -- t[59499] = 28
      "0011100" when "01110100001101100", -- t[59500] = 28
      "0011100" when "01110100001101101", -- t[59501] = 28
      "0011100" when "01110100001101110", -- t[59502] = 28
      "0011100" when "01110100001101111", -- t[59503] = 28
      "0011100" when "01110100001110000", -- t[59504] = 28
      "0011100" when "01110100001110001", -- t[59505] = 28
      "0011100" when "01110100001110010", -- t[59506] = 28
      "0011100" when "01110100001110011", -- t[59507] = 28
      "0011100" when "01110100001110100", -- t[59508] = 28
      "0011100" when "01110100001110101", -- t[59509] = 28
      "0011100" when "01110100001110110", -- t[59510] = 28
      "0011100" when "01110100001110111", -- t[59511] = 28
      "0011100" when "01110100001111000", -- t[59512] = 28
      "0011100" when "01110100001111001", -- t[59513] = 28
      "0011100" when "01110100001111010", -- t[59514] = 28
      "0011100" when "01110100001111011", -- t[59515] = 28
      "0011100" when "01110100001111100", -- t[59516] = 28
      "0011100" when "01110100001111101", -- t[59517] = 28
      "0011100" when "01110100001111110", -- t[59518] = 28
      "0011100" when "01110100001111111", -- t[59519] = 28
      "0011100" when "01110100010000000", -- t[59520] = 28
      "0011100" when "01110100010000001", -- t[59521] = 28
      "0011100" when "01110100010000010", -- t[59522] = 28
      "0011100" when "01110100010000011", -- t[59523] = 28
      "0011100" when "01110100010000100", -- t[59524] = 28
      "0011100" when "01110100010000101", -- t[59525] = 28
      "0011100" when "01110100010000110", -- t[59526] = 28
      "0011100" when "01110100010000111", -- t[59527] = 28
      "0011100" when "01110100010001000", -- t[59528] = 28
      "0011100" when "01110100010001001", -- t[59529] = 28
      "0011100" when "01110100010001010", -- t[59530] = 28
      "0011100" when "01110100010001011", -- t[59531] = 28
      "0011100" when "01110100010001100", -- t[59532] = 28
      "0011100" when "01110100010001101", -- t[59533] = 28
      "0011100" when "01110100010001110", -- t[59534] = 28
      "0011100" when "01110100010001111", -- t[59535] = 28
      "0011100" when "01110100010010000", -- t[59536] = 28
      "0011100" when "01110100010010001", -- t[59537] = 28
      "0011100" when "01110100010010010", -- t[59538] = 28
      "0011100" when "01110100010010011", -- t[59539] = 28
      "0011100" when "01110100010010100", -- t[59540] = 28
      "0011100" when "01110100010010101", -- t[59541] = 28
      "0011100" when "01110100010010110", -- t[59542] = 28
      "0011100" when "01110100010010111", -- t[59543] = 28
      "0011100" when "01110100010011000", -- t[59544] = 28
      "0011100" when "01110100010011001", -- t[59545] = 28
      "0011100" when "01110100010011010", -- t[59546] = 28
      "0011100" when "01110100010011011", -- t[59547] = 28
      "0011100" when "01110100010011100", -- t[59548] = 28
      "0011100" when "01110100010011101", -- t[59549] = 28
      "0011100" when "01110100010011110", -- t[59550] = 28
      "0011100" when "01110100010011111", -- t[59551] = 28
      "0011100" when "01110100010100000", -- t[59552] = 28
      "0011100" when "01110100010100001", -- t[59553] = 28
      "0011100" when "01110100010100010", -- t[59554] = 28
      "0011100" when "01110100010100011", -- t[59555] = 28
      "0011100" when "01110100010100100", -- t[59556] = 28
      "0011100" when "01110100010100101", -- t[59557] = 28
      "0011100" when "01110100010100110", -- t[59558] = 28
      "0011100" when "01110100010100111", -- t[59559] = 28
      "0011100" when "01110100010101000", -- t[59560] = 28
      "0011100" when "01110100010101001", -- t[59561] = 28
      "0011100" when "01110100010101010", -- t[59562] = 28
      "0011100" when "01110100010101011", -- t[59563] = 28
      "0011100" when "01110100010101100", -- t[59564] = 28
      "0011100" when "01110100010101101", -- t[59565] = 28
      "0011100" when "01110100010101110", -- t[59566] = 28
      "0011100" when "01110100010101111", -- t[59567] = 28
      "0011100" when "01110100010110000", -- t[59568] = 28
      "0011100" when "01110100010110001", -- t[59569] = 28
      "0011100" when "01110100010110010", -- t[59570] = 28
      "0011100" when "01110100010110011", -- t[59571] = 28
      "0011100" when "01110100010110100", -- t[59572] = 28
      "0011100" when "01110100010110101", -- t[59573] = 28
      "0011100" when "01110100010110110", -- t[59574] = 28
      "0011100" when "01110100010110111", -- t[59575] = 28
      "0011100" when "01110100010111000", -- t[59576] = 28
      "0011100" when "01110100010111001", -- t[59577] = 28
      "0011100" when "01110100010111010", -- t[59578] = 28
      "0011100" when "01110100010111011", -- t[59579] = 28
      "0011100" when "01110100010111100", -- t[59580] = 28
      "0011100" when "01110100010111101", -- t[59581] = 28
      "0011100" when "01110100010111110", -- t[59582] = 28
      "0011100" when "01110100010111111", -- t[59583] = 28
      "0011100" when "01110100011000000", -- t[59584] = 28
      "0011100" when "01110100011000001", -- t[59585] = 28
      "0011100" when "01110100011000010", -- t[59586] = 28
      "0011100" when "01110100011000011", -- t[59587] = 28
      "0011100" when "01110100011000100", -- t[59588] = 28
      "0011100" when "01110100011000101", -- t[59589] = 28
      "0011100" when "01110100011000110", -- t[59590] = 28
      "0011100" when "01110100011000111", -- t[59591] = 28
      "0011100" when "01110100011001000", -- t[59592] = 28
      "0011100" when "01110100011001001", -- t[59593] = 28
      "0011100" when "01110100011001010", -- t[59594] = 28
      "0011100" when "01110100011001011", -- t[59595] = 28
      "0011100" when "01110100011001100", -- t[59596] = 28
      "0011100" when "01110100011001101", -- t[59597] = 28
      "0011100" when "01110100011001110", -- t[59598] = 28
      "0011100" when "01110100011001111", -- t[59599] = 28
      "0011100" when "01110100011010000", -- t[59600] = 28
      "0011100" when "01110100011010001", -- t[59601] = 28
      "0011100" when "01110100011010010", -- t[59602] = 28
      "0011100" when "01110100011010011", -- t[59603] = 28
      "0011100" when "01110100011010100", -- t[59604] = 28
      "0011100" when "01110100011010101", -- t[59605] = 28
      "0011100" when "01110100011010110", -- t[59606] = 28
      "0011100" when "01110100011010111", -- t[59607] = 28
      "0011100" when "01110100011011000", -- t[59608] = 28
      "0011100" when "01110100011011001", -- t[59609] = 28
      "0011100" when "01110100011011010", -- t[59610] = 28
      "0011100" when "01110100011011011", -- t[59611] = 28
      "0011100" when "01110100011011100", -- t[59612] = 28
      "0011100" when "01110100011011101", -- t[59613] = 28
      "0011100" when "01110100011011110", -- t[59614] = 28
      "0011100" when "01110100011011111", -- t[59615] = 28
      "0011100" when "01110100011100000", -- t[59616] = 28
      "0011100" when "01110100011100001", -- t[59617] = 28
      "0011100" when "01110100011100010", -- t[59618] = 28
      "0011100" when "01110100011100011", -- t[59619] = 28
      "0011100" when "01110100011100100", -- t[59620] = 28
      "0011100" when "01110100011100101", -- t[59621] = 28
      "0011100" when "01110100011100110", -- t[59622] = 28
      "0011100" when "01110100011100111", -- t[59623] = 28
      "0011100" when "01110100011101000", -- t[59624] = 28
      "0011100" when "01110100011101001", -- t[59625] = 28
      "0011100" when "01110100011101010", -- t[59626] = 28
      "0011100" when "01110100011101011", -- t[59627] = 28
      "0011100" when "01110100011101100", -- t[59628] = 28
      "0011100" when "01110100011101101", -- t[59629] = 28
      "0011100" when "01110100011101110", -- t[59630] = 28
      "0011100" when "01110100011101111", -- t[59631] = 28
      "0011100" when "01110100011110000", -- t[59632] = 28
      "0011100" when "01110100011110001", -- t[59633] = 28
      "0011100" when "01110100011110010", -- t[59634] = 28
      "0011100" when "01110100011110011", -- t[59635] = 28
      "0011100" when "01110100011110100", -- t[59636] = 28
      "0011100" when "01110100011110101", -- t[59637] = 28
      "0011100" when "01110100011110110", -- t[59638] = 28
      "0011100" when "01110100011110111", -- t[59639] = 28
      "0011100" when "01110100011111000", -- t[59640] = 28
      "0011100" when "01110100011111001", -- t[59641] = 28
      "0011100" when "01110100011111010", -- t[59642] = 28
      "0011100" when "01110100011111011", -- t[59643] = 28
      "0011100" when "01110100011111100", -- t[59644] = 28
      "0011100" when "01110100011111101", -- t[59645] = 28
      "0011100" when "01110100011111110", -- t[59646] = 28
      "0011100" when "01110100011111111", -- t[59647] = 28
      "0011100" when "01110100100000000", -- t[59648] = 28
      "0011100" when "01110100100000001", -- t[59649] = 28
      "0011100" when "01110100100000010", -- t[59650] = 28
      "0011100" when "01110100100000011", -- t[59651] = 28
      "0011100" when "01110100100000100", -- t[59652] = 28
      "0011100" when "01110100100000101", -- t[59653] = 28
      "0011100" when "01110100100000110", -- t[59654] = 28
      "0011100" when "01110100100000111", -- t[59655] = 28
      "0011100" when "01110100100001000", -- t[59656] = 28
      "0011100" when "01110100100001001", -- t[59657] = 28
      "0011100" when "01110100100001010", -- t[59658] = 28
      "0011100" when "01110100100001011", -- t[59659] = 28
      "0011100" when "01110100100001100", -- t[59660] = 28
      "0011100" when "01110100100001101", -- t[59661] = 28
      "0011100" when "01110100100001110", -- t[59662] = 28
      "0011100" when "01110100100001111", -- t[59663] = 28
      "0011100" when "01110100100010000", -- t[59664] = 28
      "0011100" when "01110100100010001", -- t[59665] = 28
      "0011100" when "01110100100010010", -- t[59666] = 28
      "0011100" when "01110100100010011", -- t[59667] = 28
      "0011100" when "01110100100010100", -- t[59668] = 28
      "0011100" when "01110100100010101", -- t[59669] = 28
      "0011100" when "01110100100010110", -- t[59670] = 28
      "0011100" when "01110100100010111", -- t[59671] = 28
      "0011100" when "01110100100011000", -- t[59672] = 28
      "0011100" when "01110100100011001", -- t[59673] = 28
      "0011100" when "01110100100011010", -- t[59674] = 28
      "0011100" when "01110100100011011", -- t[59675] = 28
      "0011100" when "01110100100011100", -- t[59676] = 28
      "0011100" when "01110100100011101", -- t[59677] = 28
      "0011100" when "01110100100011110", -- t[59678] = 28
      "0011100" when "01110100100011111", -- t[59679] = 28
      "0011100" when "01110100100100000", -- t[59680] = 28
      "0011100" when "01110100100100001", -- t[59681] = 28
      "0011100" when "01110100100100010", -- t[59682] = 28
      "0011100" when "01110100100100011", -- t[59683] = 28
      "0011100" when "01110100100100100", -- t[59684] = 28
      "0011100" when "01110100100100101", -- t[59685] = 28
      "0011100" when "01110100100100110", -- t[59686] = 28
      "0011100" when "01110100100100111", -- t[59687] = 28
      "0011100" when "01110100100101000", -- t[59688] = 28
      "0011100" when "01110100100101001", -- t[59689] = 28
      "0011100" when "01110100100101010", -- t[59690] = 28
      "0011100" when "01110100100101011", -- t[59691] = 28
      "0011100" when "01110100100101100", -- t[59692] = 28
      "0011100" when "01110100100101101", -- t[59693] = 28
      "0011100" when "01110100100101110", -- t[59694] = 28
      "0011100" when "01110100100101111", -- t[59695] = 28
      "0011100" when "01110100100110000", -- t[59696] = 28
      "0011100" when "01110100100110001", -- t[59697] = 28
      "0011100" when "01110100100110010", -- t[59698] = 28
      "0011100" when "01110100100110011", -- t[59699] = 28
      "0011100" when "01110100100110100", -- t[59700] = 28
      "0011100" when "01110100100110101", -- t[59701] = 28
      "0011100" when "01110100100110110", -- t[59702] = 28
      "0011100" when "01110100100110111", -- t[59703] = 28
      "0011100" when "01110100100111000", -- t[59704] = 28
      "0011100" when "01110100100111001", -- t[59705] = 28
      "0011100" when "01110100100111010", -- t[59706] = 28
      "0011100" when "01110100100111011", -- t[59707] = 28
      "0011100" when "01110100100111100", -- t[59708] = 28
      "0011100" when "01110100100111101", -- t[59709] = 28
      "0011100" when "01110100100111110", -- t[59710] = 28
      "0011100" when "01110100100111111", -- t[59711] = 28
      "0011100" when "01110100101000000", -- t[59712] = 28
      "0011100" when "01110100101000001", -- t[59713] = 28
      "0011100" when "01110100101000010", -- t[59714] = 28
      "0011100" when "01110100101000011", -- t[59715] = 28
      "0011100" when "01110100101000100", -- t[59716] = 28
      "0011100" when "01110100101000101", -- t[59717] = 28
      "0011100" when "01110100101000110", -- t[59718] = 28
      "0011100" when "01110100101000111", -- t[59719] = 28
      "0011100" when "01110100101001000", -- t[59720] = 28
      "0011100" when "01110100101001001", -- t[59721] = 28
      "0011100" when "01110100101001010", -- t[59722] = 28
      "0011100" when "01110100101001011", -- t[59723] = 28
      "0011100" when "01110100101001100", -- t[59724] = 28
      "0011100" when "01110100101001101", -- t[59725] = 28
      "0011100" when "01110100101001110", -- t[59726] = 28
      "0011100" when "01110100101001111", -- t[59727] = 28
      "0011100" when "01110100101010000", -- t[59728] = 28
      "0011100" when "01110100101010001", -- t[59729] = 28
      "0011100" when "01110100101010010", -- t[59730] = 28
      "0011100" when "01110100101010011", -- t[59731] = 28
      "0011100" when "01110100101010100", -- t[59732] = 28
      "0011100" when "01110100101010101", -- t[59733] = 28
      "0011100" when "01110100101010110", -- t[59734] = 28
      "0011100" when "01110100101010111", -- t[59735] = 28
      "0011100" when "01110100101011000", -- t[59736] = 28
      "0011100" when "01110100101011001", -- t[59737] = 28
      "0011100" when "01110100101011010", -- t[59738] = 28
      "0011100" when "01110100101011011", -- t[59739] = 28
      "0011100" when "01110100101011100", -- t[59740] = 28
      "0011100" when "01110100101011101", -- t[59741] = 28
      "0011100" when "01110100101011110", -- t[59742] = 28
      "0011100" when "01110100101011111", -- t[59743] = 28
      "0011100" when "01110100101100000", -- t[59744] = 28
      "0011100" when "01110100101100001", -- t[59745] = 28
      "0011100" when "01110100101100010", -- t[59746] = 28
      "0011100" when "01110100101100011", -- t[59747] = 28
      "0011100" when "01110100101100100", -- t[59748] = 28
      "0011100" when "01110100101100101", -- t[59749] = 28
      "0011100" when "01110100101100110", -- t[59750] = 28
      "0011100" when "01110100101100111", -- t[59751] = 28
      "0011100" when "01110100101101000", -- t[59752] = 28
      "0011100" when "01110100101101001", -- t[59753] = 28
      "0011100" when "01110100101101010", -- t[59754] = 28
      "0011100" when "01110100101101011", -- t[59755] = 28
      "0011100" when "01110100101101100", -- t[59756] = 28
      "0011100" when "01110100101101101", -- t[59757] = 28
      "0011100" when "01110100101101110", -- t[59758] = 28
      "0011100" when "01110100101101111", -- t[59759] = 28
      "0011100" when "01110100101110000", -- t[59760] = 28
      "0011100" when "01110100101110001", -- t[59761] = 28
      "0011100" when "01110100101110010", -- t[59762] = 28
      "0011100" when "01110100101110011", -- t[59763] = 28
      "0011100" when "01110100101110100", -- t[59764] = 28
      "0011100" when "01110100101110101", -- t[59765] = 28
      "0011100" when "01110100101110110", -- t[59766] = 28
      "0011100" when "01110100101110111", -- t[59767] = 28
      "0011100" when "01110100101111000", -- t[59768] = 28
      "0011100" when "01110100101111001", -- t[59769] = 28
      "0011100" when "01110100101111010", -- t[59770] = 28
      "0011100" when "01110100101111011", -- t[59771] = 28
      "0011100" when "01110100101111100", -- t[59772] = 28
      "0011100" when "01110100101111101", -- t[59773] = 28
      "0011100" when "01110100101111110", -- t[59774] = 28
      "0011100" when "01110100101111111", -- t[59775] = 28
      "0011100" when "01110100110000000", -- t[59776] = 28
      "0011100" when "01110100110000001", -- t[59777] = 28
      "0011100" when "01110100110000010", -- t[59778] = 28
      "0011100" when "01110100110000011", -- t[59779] = 28
      "0011100" when "01110100110000100", -- t[59780] = 28
      "0011100" when "01110100110000101", -- t[59781] = 28
      "0011100" when "01110100110000110", -- t[59782] = 28
      "0011100" when "01110100110000111", -- t[59783] = 28
      "0011100" when "01110100110001000", -- t[59784] = 28
      "0011100" when "01110100110001001", -- t[59785] = 28
      "0011100" when "01110100110001010", -- t[59786] = 28
      "0011100" when "01110100110001011", -- t[59787] = 28
      "0011100" when "01110100110001100", -- t[59788] = 28
      "0011100" when "01110100110001101", -- t[59789] = 28
      "0011100" when "01110100110001110", -- t[59790] = 28
      "0011100" when "01110100110001111", -- t[59791] = 28
      "0011100" when "01110100110010000", -- t[59792] = 28
      "0011100" when "01110100110010001", -- t[59793] = 28
      "0011100" when "01110100110010010", -- t[59794] = 28
      "0011100" when "01110100110010011", -- t[59795] = 28
      "0011100" when "01110100110010100", -- t[59796] = 28
      "0011100" when "01110100110010101", -- t[59797] = 28
      "0011100" when "01110100110010110", -- t[59798] = 28
      "0011100" when "01110100110010111", -- t[59799] = 28
      "0011100" when "01110100110011000", -- t[59800] = 28
      "0011100" when "01110100110011001", -- t[59801] = 28
      "0011100" when "01110100110011010", -- t[59802] = 28
      "0011100" when "01110100110011011", -- t[59803] = 28
      "0011100" when "01110100110011100", -- t[59804] = 28
      "0011100" when "01110100110011101", -- t[59805] = 28
      "0011100" when "01110100110011110", -- t[59806] = 28
      "0011100" when "01110100110011111", -- t[59807] = 28
      "0011100" when "01110100110100000", -- t[59808] = 28
      "0011100" when "01110100110100001", -- t[59809] = 28
      "0011100" when "01110100110100010", -- t[59810] = 28
      "0011100" when "01110100110100011", -- t[59811] = 28
      "0011100" when "01110100110100100", -- t[59812] = 28
      "0011100" when "01110100110100101", -- t[59813] = 28
      "0011100" when "01110100110100110", -- t[59814] = 28
      "0011100" when "01110100110100111", -- t[59815] = 28
      "0011100" when "01110100110101000", -- t[59816] = 28
      "0011100" when "01110100110101001", -- t[59817] = 28
      "0011100" when "01110100110101010", -- t[59818] = 28
      "0011100" when "01110100110101011", -- t[59819] = 28
      "0011100" when "01110100110101100", -- t[59820] = 28
      "0011100" when "01110100110101101", -- t[59821] = 28
      "0011101" when "01110100110101110", -- t[59822] = 29
      "0011101" when "01110100110101111", -- t[59823] = 29
      "0011101" when "01110100110110000", -- t[59824] = 29
      "0011101" when "01110100110110001", -- t[59825] = 29
      "0011101" when "01110100110110010", -- t[59826] = 29
      "0011101" when "01110100110110011", -- t[59827] = 29
      "0011101" when "01110100110110100", -- t[59828] = 29
      "0011101" when "01110100110110101", -- t[59829] = 29
      "0011101" when "01110100110110110", -- t[59830] = 29
      "0011101" when "01110100110110111", -- t[59831] = 29
      "0011101" when "01110100110111000", -- t[59832] = 29
      "0011101" when "01110100110111001", -- t[59833] = 29
      "0011101" when "01110100110111010", -- t[59834] = 29
      "0011101" when "01110100110111011", -- t[59835] = 29
      "0011101" when "01110100110111100", -- t[59836] = 29
      "0011101" when "01110100110111101", -- t[59837] = 29
      "0011101" when "01110100110111110", -- t[59838] = 29
      "0011101" when "01110100110111111", -- t[59839] = 29
      "0011101" when "01110100111000000", -- t[59840] = 29
      "0011101" when "01110100111000001", -- t[59841] = 29
      "0011101" when "01110100111000010", -- t[59842] = 29
      "0011101" when "01110100111000011", -- t[59843] = 29
      "0011101" when "01110100111000100", -- t[59844] = 29
      "0011101" when "01110100111000101", -- t[59845] = 29
      "0011101" when "01110100111000110", -- t[59846] = 29
      "0011101" when "01110100111000111", -- t[59847] = 29
      "0011101" when "01110100111001000", -- t[59848] = 29
      "0011101" when "01110100111001001", -- t[59849] = 29
      "0011101" when "01110100111001010", -- t[59850] = 29
      "0011101" when "01110100111001011", -- t[59851] = 29
      "0011101" when "01110100111001100", -- t[59852] = 29
      "0011101" when "01110100111001101", -- t[59853] = 29
      "0011101" when "01110100111001110", -- t[59854] = 29
      "0011101" when "01110100111001111", -- t[59855] = 29
      "0011101" when "01110100111010000", -- t[59856] = 29
      "0011101" when "01110100111010001", -- t[59857] = 29
      "0011101" when "01110100111010010", -- t[59858] = 29
      "0011101" when "01110100111010011", -- t[59859] = 29
      "0011101" when "01110100111010100", -- t[59860] = 29
      "0011101" when "01110100111010101", -- t[59861] = 29
      "0011101" when "01110100111010110", -- t[59862] = 29
      "0011101" when "01110100111010111", -- t[59863] = 29
      "0011101" when "01110100111011000", -- t[59864] = 29
      "0011101" when "01110100111011001", -- t[59865] = 29
      "0011101" when "01110100111011010", -- t[59866] = 29
      "0011101" when "01110100111011011", -- t[59867] = 29
      "0011101" when "01110100111011100", -- t[59868] = 29
      "0011101" when "01110100111011101", -- t[59869] = 29
      "0011101" when "01110100111011110", -- t[59870] = 29
      "0011101" when "01110100111011111", -- t[59871] = 29
      "0011101" when "01110100111100000", -- t[59872] = 29
      "0011101" when "01110100111100001", -- t[59873] = 29
      "0011101" when "01110100111100010", -- t[59874] = 29
      "0011101" when "01110100111100011", -- t[59875] = 29
      "0011101" when "01110100111100100", -- t[59876] = 29
      "0011101" when "01110100111100101", -- t[59877] = 29
      "0011101" when "01110100111100110", -- t[59878] = 29
      "0011101" when "01110100111100111", -- t[59879] = 29
      "0011101" when "01110100111101000", -- t[59880] = 29
      "0011101" when "01110100111101001", -- t[59881] = 29
      "0011101" when "01110100111101010", -- t[59882] = 29
      "0011101" when "01110100111101011", -- t[59883] = 29
      "0011101" when "01110100111101100", -- t[59884] = 29
      "0011101" when "01110100111101101", -- t[59885] = 29
      "0011101" when "01110100111101110", -- t[59886] = 29
      "0011101" when "01110100111101111", -- t[59887] = 29
      "0011101" when "01110100111110000", -- t[59888] = 29
      "0011101" when "01110100111110001", -- t[59889] = 29
      "0011101" when "01110100111110010", -- t[59890] = 29
      "0011101" when "01110100111110011", -- t[59891] = 29
      "0011101" when "01110100111110100", -- t[59892] = 29
      "0011101" when "01110100111110101", -- t[59893] = 29
      "0011101" when "01110100111110110", -- t[59894] = 29
      "0011101" when "01110100111110111", -- t[59895] = 29
      "0011101" when "01110100111111000", -- t[59896] = 29
      "0011101" when "01110100111111001", -- t[59897] = 29
      "0011101" when "01110100111111010", -- t[59898] = 29
      "0011101" when "01110100111111011", -- t[59899] = 29
      "0011101" when "01110100111111100", -- t[59900] = 29
      "0011101" when "01110100111111101", -- t[59901] = 29
      "0011101" when "01110100111111110", -- t[59902] = 29
      "0011101" when "01110100111111111", -- t[59903] = 29
      "0011101" when "01110101000000000", -- t[59904] = 29
      "0011101" when "01110101000000001", -- t[59905] = 29
      "0011101" when "01110101000000010", -- t[59906] = 29
      "0011101" when "01110101000000011", -- t[59907] = 29
      "0011101" when "01110101000000100", -- t[59908] = 29
      "0011101" when "01110101000000101", -- t[59909] = 29
      "0011101" when "01110101000000110", -- t[59910] = 29
      "0011101" when "01110101000000111", -- t[59911] = 29
      "0011101" when "01110101000001000", -- t[59912] = 29
      "0011101" when "01110101000001001", -- t[59913] = 29
      "0011101" when "01110101000001010", -- t[59914] = 29
      "0011101" when "01110101000001011", -- t[59915] = 29
      "0011101" when "01110101000001100", -- t[59916] = 29
      "0011101" when "01110101000001101", -- t[59917] = 29
      "0011101" when "01110101000001110", -- t[59918] = 29
      "0011101" when "01110101000001111", -- t[59919] = 29
      "0011101" when "01110101000010000", -- t[59920] = 29
      "0011101" when "01110101000010001", -- t[59921] = 29
      "0011101" when "01110101000010010", -- t[59922] = 29
      "0011101" when "01110101000010011", -- t[59923] = 29
      "0011101" when "01110101000010100", -- t[59924] = 29
      "0011101" when "01110101000010101", -- t[59925] = 29
      "0011101" when "01110101000010110", -- t[59926] = 29
      "0011101" when "01110101000010111", -- t[59927] = 29
      "0011101" when "01110101000011000", -- t[59928] = 29
      "0011101" when "01110101000011001", -- t[59929] = 29
      "0011101" when "01110101000011010", -- t[59930] = 29
      "0011101" when "01110101000011011", -- t[59931] = 29
      "0011101" when "01110101000011100", -- t[59932] = 29
      "0011101" when "01110101000011101", -- t[59933] = 29
      "0011101" when "01110101000011110", -- t[59934] = 29
      "0011101" when "01110101000011111", -- t[59935] = 29
      "0011101" when "01110101000100000", -- t[59936] = 29
      "0011101" when "01110101000100001", -- t[59937] = 29
      "0011101" when "01110101000100010", -- t[59938] = 29
      "0011101" when "01110101000100011", -- t[59939] = 29
      "0011101" when "01110101000100100", -- t[59940] = 29
      "0011101" when "01110101000100101", -- t[59941] = 29
      "0011101" when "01110101000100110", -- t[59942] = 29
      "0011101" when "01110101000100111", -- t[59943] = 29
      "0011101" when "01110101000101000", -- t[59944] = 29
      "0011101" when "01110101000101001", -- t[59945] = 29
      "0011101" when "01110101000101010", -- t[59946] = 29
      "0011101" when "01110101000101011", -- t[59947] = 29
      "0011101" when "01110101000101100", -- t[59948] = 29
      "0011101" when "01110101000101101", -- t[59949] = 29
      "0011101" when "01110101000101110", -- t[59950] = 29
      "0011101" when "01110101000101111", -- t[59951] = 29
      "0011101" when "01110101000110000", -- t[59952] = 29
      "0011101" when "01110101000110001", -- t[59953] = 29
      "0011101" when "01110101000110010", -- t[59954] = 29
      "0011101" when "01110101000110011", -- t[59955] = 29
      "0011101" when "01110101000110100", -- t[59956] = 29
      "0011101" when "01110101000110101", -- t[59957] = 29
      "0011101" when "01110101000110110", -- t[59958] = 29
      "0011101" when "01110101000110111", -- t[59959] = 29
      "0011101" when "01110101000111000", -- t[59960] = 29
      "0011101" when "01110101000111001", -- t[59961] = 29
      "0011101" when "01110101000111010", -- t[59962] = 29
      "0011101" when "01110101000111011", -- t[59963] = 29
      "0011101" when "01110101000111100", -- t[59964] = 29
      "0011101" when "01110101000111101", -- t[59965] = 29
      "0011101" when "01110101000111110", -- t[59966] = 29
      "0011101" when "01110101000111111", -- t[59967] = 29
      "0011101" when "01110101001000000", -- t[59968] = 29
      "0011101" when "01110101001000001", -- t[59969] = 29
      "0011101" when "01110101001000010", -- t[59970] = 29
      "0011101" when "01110101001000011", -- t[59971] = 29
      "0011101" when "01110101001000100", -- t[59972] = 29
      "0011101" when "01110101001000101", -- t[59973] = 29
      "0011101" when "01110101001000110", -- t[59974] = 29
      "0011101" when "01110101001000111", -- t[59975] = 29
      "0011101" when "01110101001001000", -- t[59976] = 29
      "0011101" when "01110101001001001", -- t[59977] = 29
      "0011101" when "01110101001001010", -- t[59978] = 29
      "0011101" when "01110101001001011", -- t[59979] = 29
      "0011101" when "01110101001001100", -- t[59980] = 29
      "0011101" when "01110101001001101", -- t[59981] = 29
      "0011101" when "01110101001001110", -- t[59982] = 29
      "0011101" when "01110101001001111", -- t[59983] = 29
      "0011101" when "01110101001010000", -- t[59984] = 29
      "0011101" when "01110101001010001", -- t[59985] = 29
      "0011101" when "01110101001010010", -- t[59986] = 29
      "0011101" when "01110101001010011", -- t[59987] = 29
      "0011101" when "01110101001010100", -- t[59988] = 29
      "0011101" when "01110101001010101", -- t[59989] = 29
      "0011101" when "01110101001010110", -- t[59990] = 29
      "0011101" when "01110101001010111", -- t[59991] = 29
      "0011101" when "01110101001011000", -- t[59992] = 29
      "0011101" when "01110101001011001", -- t[59993] = 29
      "0011101" when "01110101001011010", -- t[59994] = 29
      "0011101" when "01110101001011011", -- t[59995] = 29
      "0011101" when "01110101001011100", -- t[59996] = 29
      "0011101" when "01110101001011101", -- t[59997] = 29
      "0011101" when "01110101001011110", -- t[59998] = 29
      "0011101" when "01110101001011111", -- t[59999] = 29
      "0011101" when "01110101001100000", -- t[60000] = 29
      "0011101" when "01110101001100001", -- t[60001] = 29
      "0011101" when "01110101001100010", -- t[60002] = 29
      "0011101" when "01110101001100011", -- t[60003] = 29
      "0011101" when "01110101001100100", -- t[60004] = 29
      "0011101" when "01110101001100101", -- t[60005] = 29
      "0011101" when "01110101001100110", -- t[60006] = 29
      "0011101" when "01110101001100111", -- t[60007] = 29
      "0011101" when "01110101001101000", -- t[60008] = 29
      "0011101" when "01110101001101001", -- t[60009] = 29
      "0011101" when "01110101001101010", -- t[60010] = 29
      "0011101" when "01110101001101011", -- t[60011] = 29
      "0011101" when "01110101001101100", -- t[60012] = 29
      "0011101" when "01110101001101101", -- t[60013] = 29
      "0011101" when "01110101001101110", -- t[60014] = 29
      "0011101" when "01110101001101111", -- t[60015] = 29
      "0011101" when "01110101001110000", -- t[60016] = 29
      "0011101" when "01110101001110001", -- t[60017] = 29
      "0011101" when "01110101001110010", -- t[60018] = 29
      "0011101" when "01110101001110011", -- t[60019] = 29
      "0011101" when "01110101001110100", -- t[60020] = 29
      "0011101" when "01110101001110101", -- t[60021] = 29
      "0011101" when "01110101001110110", -- t[60022] = 29
      "0011101" when "01110101001110111", -- t[60023] = 29
      "0011101" when "01110101001111000", -- t[60024] = 29
      "0011101" when "01110101001111001", -- t[60025] = 29
      "0011101" when "01110101001111010", -- t[60026] = 29
      "0011101" when "01110101001111011", -- t[60027] = 29
      "0011101" when "01110101001111100", -- t[60028] = 29
      "0011101" when "01110101001111101", -- t[60029] = 29
      "0011101" when "01110101001111110", -- t[60030] = 29
      "0011101" when "01110101001111111", -- t[60031] = 29
      "0011101" when "01110101010000000", -- t[60032] = 29
      "0011101" when "01110101010000001", -- t[60033] = 29
      "0011101" when "01110101010000010", -- t[60034] = 29
      "0011101" when "01110101010000011", -- t[60035] = 29
      "0011101" when "01110101010000100", -- t[60036] = 29
      "0011101" when "01110101010000101", -- t[60037] = 29
      "0011101" when "01110101010000110", -- t[60038] = 29
      "0011101" when "01110101010000111", -- t[60039] = 29
      "0011101" when "01110101010001000", -- t[60040] = 29
      "0011101" when "01110101010001001", -- t[60041] = 29
      "0011101" when "01110101010001010", -- t[60042] = 29
      "0011101" when "01110101010001011", -- t[60043] = 29
      "0011101" when "01110101010001100", -- t[60044] = 29
      "0011101" when "01110101010001101", -- t[60045] = 29
      "0011101" when "01110101010001110", -- t[60046] = 29
      "0011101" when "01110101010001111", -- t[60047] = 29
      "0011101" when "01110101010010000", -- t[60048] = 29
      "0011101" when "01110101010010001", -- t[60049] = 29
      "0011101" when "01110101010010010", -- t[60050] = 29
      "0011101" when "01110101010010011", -- t[60051] = 29
      "0011101" when "01110101010010100", -- t[60052] = 29
      "0011101" when "01110101010010101", -- t[60053] = 29
      "0011101" when "01110101010010110", -- t[60054] = 29
      "0011101" when "01110101010010111", -- t[60055] = 29
      "0011101" when "01110101010011000", -- t[60056] = 29
      "0011101" when "01110101010011001", -- t[60057] = 29
      "0011101" when "01110101010011010", -- t[60058] = 29
      "0011101" when "01110101010011011", -- t[60059] = 29
      "0011101" when "01110101010011100", -- t[60060] = 29
      "0011101" when "01110101010011101", -- t[60061] = 29
      "0011101" when "01110101010011110", -- t[60062] = 29
      "0011101" when "01110101010011111", -- t[60063] = 29
      "0011101" when "01110101010100000", -- t[60064] = 29
      "0011101" when "01110101010100001", -- t[60065] = 29
      "0011101" when "01110101010100010", -- t[60066] = 29
      "0011101" when "01110101010100011", -- t[60067] = 29
      "0011101" when "01110101010100100", -- t[60068] = 29
      "0011101" when "01110101010100101", -- t[60069] = 29
      "0011101" when "01110101010100110", -- t[60070] = 29
      "0011101" when "01110101010100111", -- t[60071] = 29
      "0011101" when "01110101010101000", -- t[60072] = 29
      "0011101" when "01110101010101001", -- t[60073] = 29
      "0011101" when "01110101010101010", -- t[60074] = 29
      "0011101" when "01110101010101011", -- t[60075] = 29
      "0011101" when "01110101010101100", -- t[60076] = 29
      "0011101" when "01110101010101101", -- t[60077] = 29
      "0011101" when "01110101010101110", -- t[60078] = 29
      "0011101" when "01110101010101111", -- t[60079] = 29
      "0011101" when "01110101010110000", -- t[60080] = 29
      "0011101" when "01110101010110001", -- t[60081] = 29
      "0011101" when "01110101010110010", -- t[60082] = 29
      "0011101" when "01110101010110011", -- t[60083] = 29
      "0011101" when "01110101010110100", -- t[60084] = 29
      "0011101" when "01110101010110101", -- t[60085] = 29
      "0011101" when "01110101010110110", -- t[60086] = 29
      "0011101" when "01110101010110111", -- t[60087] = 29
      "0011101" when "01110101010111000", -- t[60088] = 29
      "0011101" when "01110101010111001", -- t[60089] = 29
      "0011101" when "01110101010111010", -- t[60090] = 29
      "0011101" when "01110101010111011", -- t[60091] = 29
      "0011101" when "01110101010111100", -- t[60092] = 29
      "0011101" when "01110101010111101", -- t[60093] = 29
      "0011101" when "01110101010111110", -- t[60094] = 29
      "0011101" when "01110101010111111", -- t[60095] = 29
      "0011101" when "01110101011000000", -- t[60096] = 29
      "0011101" when "01110101011000001", -- t[60097] = 29
      "0011101" when "01110101011000010", -- t[60098] = 29
      "0011101" when "01110101011000011", -- t[60099] = 29
      "0011101" when "01110101011000100", -- t[60100] = 29
      "0011101" when "01110101011000101", -- t[60101] = 29
      "0011101" when "01110101011000110", -- t[60102] = 29
      "0011101" when "01110101011000111", -- t[60103] = 29
      "0011101" when "01110101011001000", -- t[60104] = 29
      "0011101" when "01110101011001001", -- t[60105] = 29
      "0011101" when "01110101011001010", -- t[60106] = 29
      "0011101" when "01110101011001011", -- t[60107] = 29
      "0011101" when "01110101011001100", -- t[60108] = 29
      "0011101" when "01110101011001101", -- t[60109] = 29
      "0011101" when "01110101011001110", -- t[60110] = 29
      "0011101" when "01110101011001111", -- t[60111] = 29
      "0011101" when "01110101011010000", -- t[60112] = 29
      "0011101" when "01110101011010001", -- t[60113] = 29
      "0011101" when "01110101011010010", -- t[60114] = 29
      "0011101" when "01110101011010011", -- t[60115] = 29
      "0011101" when "01110101011010100", -- t[60116] = 29
      "0011101" when "01110101011010101", -- t[60117] = 29
      "0011101" when "01110101011010110", -- t[60118] = 29
      "0011101" when "01110101011010111", -- t[60119] = 29
      "0011101" when "01110101011011000", -- t[60120] = 29
      "0011101" when "01110101011011001", -- t[60121] = 29
      "0011101" when "01110101011011010", -- t[60122] = 29
      "0011101" when "01110101011011011", -- t[60123] = 29
      "0011101" when "01110101011011100", -- t[60124] = 29
      "0011101" when "01110101011011101", -- t[60125] = 29
      "0011101" when "01110101011011110", -- t[60126] = 29
      "0011101" when "01110101011011111", -- t[60127] = 29
      "0011101" when "01110101011100000", -- t[60128] = 29
      "0011101" when "01110101011100001", -- t[60129] = 29
      "0011101" when "01110101011100010", -- t[60130] = 29
      "0011101" when "01110101011100011", -- t[60131] = 29
      "0011101" when "01110101011100100", -- t[60132] = 29
      "0011101" when "01110101011100101", -- t[60133] = 29
      "0011101" when "01110101011100110", -- t[60134] = 29
      "0011101" when "01110101011100111", -- t[60135] = 29
      "0011101" when "01110101011101000", -- t[60136] = 29
      "0011101" when "01110101011101001", -- t[60137] = 29
      "0011101" when "01110101011101010", -- t[60138] = 29
      "0011101" when "01110101011101011", -- t[60139] = 29
      "0011101" when "01110101011101100", -- t[60140] = 29
      "0011101" when "01110101011101101", -- t[60141] = 29
      "0011101" when "01110101011101110", -- t[60142] = 29
      "0011101" when "01110101011101111", -- t[60143] = 29
      "0011101" when "01110101011110000", -- t[60144] = 29
      "0011101" when "01110101011110001", -- t[60145] = 29
      "0011101" when "01110101011110010", -- t[60146] = 29
      "0011101" when "01110101011110011", -- t[60147] = 29
      "0011101" when "01110101011110100", -- t[60148] = 29
      "0011101" when "01110101011110101", -- t[60149] = 29
      "0011101" when "01110101011110110", -- t[60150] = 29
      "0011101" when "01110101011110111", -- t[60151] = 29
      "0011101" when "01110101011111000", -- t[60152] = 29
      "0011101" when "01110101011111001", -- t[60153] = 29
      "0011101" when "01110101011111010", -- t[60154] = 29
      "0011101" when "01110101011111011", -- t[60155] = 29
      "0011101" when "01110101011111100", -- t[60156] = 29
      "0011101" when "01110101011111101", -- t[60157] = 29
      "0011101" when "01110101011111110", -- t[60158] = 29
      "0011101" when "01110101011111111", -- t[60159] = 29
      "0011101" when "01110101100000000", -- t[60160] = 29
      "0011101" when "01110101100000001", -- t[60161] = 29
      "0011101" when "01110101100000010", -- t[60162] = 29
      "0011101" when "01110101100000011", -- t[60163] = 29
      "0011101" when "01110101100000100", -- t[60164] = 29
      "0011101" when "01110101100000101", -- t[60165] = 29
      "0011101" when "01110101100000110", -- t[60166] = 29
      "0011101" when "01110101100000111", -- t[60167] = 29
      "0011101" when "01110101100001000", -- t[60168] = 29
      "0011101" when "01110101100001001", -- t[60169] = 29
      "0011101" when "01110101100001010", -- t[60170] = 29
      "0011101" when "01110101100001011", -- t[60171] = 29
      "0011101" when "01110101100001100", -- t[60172] = 29
      "0011101" when "01110101100001101", -- t[60173] = 29
      "0011101" when "01110101100001110", -- t[60174] = 29
      "0011101" when "01110101100001111", -- t[60175] = 29
      "0011101" when "01110101100010000", -- t[60176] = 29
      "0011101" when "01110101100010001", -- t[60177] = 29
      "0011101" when "01110101100010010", -- t[60178] = 29
      "0011101" when "01110101100010011", -- t[60179] = 29
      "0011101" when "01110101100010100", -- t[60180] = 29
      "0011101" when "01110101100010101", -- t[60181] = 29
      "0011101" when "01110101100010110", -- t[60182] = 29
      "0011101" when "01110101100010111", -- t[60183] = 29
      "0011101" when "01110101100011000", -- t[60184] = 29
      "0011101" when "01110101100011001", -- t[60185] = 29
      "0011101" when "01110101100011010", -- t[60186] = 29
      "0011101" when "01110101100011011", -- t[60187] = 29
      "0011101" when "01110101100011100", -- t[60188] = 29
      "0011101" when "01110101100011101", -- t[60189] = 29
      "0011101" when "01110101100011110", -- t[60190] = 29
      "0011101" when "01110101100011111", -- t[60191] = 29
      "0011101" when "01110101100100000", -- t[60192] = 29
      "0011101" when "01110101100100001", -- t[60193] = 29
      "0011101" when "01110101100100010", -- t[60194] = 29
      "0011101" when "01110101100100011", -- t[60195] = 29
      "0011101" when "01110101100100100", -- t[60196] = 29
      "0011101" when "01110101100100101", -- t[60197] = 29
      "0011101" when "01110101100100110", -- t[60198] = 29
      "0011101" when "01110101100100111", -- t[60199] = 29
      "0011101" when "01110101100101000", -- t[60200] = 29
      "0011101" when "01110101100101001", -- t[60201] = 29
      "0011101" when "01110101100101010", -- t[60202] = 29
      "0011101" when "01110101100101011", -- t[60203] = 29
      "0011101" when "01110101100101100", -- t[60204] = 29
      "0011101" when "01110101100101101", -- t[60205] = 29
      "0011101" when "01110101100101110", -- t[60206] = 29
      "0011101" when "01110101100101111", -- t[60207] = 29
      "0011101" when "01110101100110000", -- t[60208] = 29
      "0011101" when "01110101100110001", -- t[60209] = 29
      "0011101" when "01110101100110010", -- t[60210] = 29
      "0011101" when "01110101100110011", -- t[60211] = 29
      "0011101" when "01110101100110100", -- t[60212] = 29
      "0011101" when "01110101100110101", -- t[60213] = 29
      "0011101" when "01110101100110110", -- t[60214] = 29
      "0011101" when "01110101100110111", -- t[60215] = 29
      "0011101" when "01110101100111000", -- t[60216] = 29
      "0011101" when "01110101100111001", -- t[60217] = 29
      "0011101" when "01110101100111010", -- t[60218] = 29
      "0011101" when "01110101100111011", -- t[60219] = 29
      "0011101" when "01110101100111100", -- t[60220] = 29
      "0011101" when "01110101100111101", -- t[60221] = 29
      "0011101" when "01110101100111110", -- t[60222] = 29
      "0011101" when "01110101100111111", -- t[60223] = 29
      "0011101" when "01110101101000000", -- t[60224] = 29
      "0011101" when "01110101101000001", -- t[60225] = 29
      "0011101" when "01110101101000010", -- t[60226] = 29
      "0011101" when "01110101101000011", -- t[60227] = 29
      "0011101" when "01110101101000100", -- t[60228] = 29
      "0011110" when "01110101101000101", -- t[60229] = 30
      "0011110" when "01110101101000110", -- t[60230] = 30
      "0011110" when "01110101101000111", -- t[60231] = 30
      "0011110" when "01110101101001000", -- t[60232] = 30
      "0011110" when "01110101101001001", -- t[60233] = 30
      "0011110" when "01110101101001010", -- t[60234] = 30
      "0011110" when "01110101101001011", -- t[60235] = 30
      "0011110" when "01110101101001100", -- t[60236] = 30
      "0011110" when "01110101101001101", -- t[60237] = 30
      "0011110" when "01110101101001110", -- t[60238] = 30
      "0011110" when "01110101101001111", -- t[60239] = 30
      "0011110" when "01110101101010000", -- t[60240] = 30
      "0011110" when "01110101101010001", -- t[60241] = 30
      "0011110" when "01110101101010010", -- t[60242] = 30
      "0011110" when "01110101101010011", -- t[60243] = 30
      "0011110" when "01110101101010100", -- t[60244] = 30
      "0011110" when "01110101101010101", -- t[60245] = 30
      "0011110" when "01110101101010110", -- t[60246] = 30
      "0011110" when "01110101101010111", -- t[60247] = 30
      "0011110" when "01110101101011000", -- t[60248] = 30
      "0011110" when "01110101101011001", -- t[60249] = 30
      "0011110" when "01110101101011010", -- t[60250] = 30
      "0011110" when "01110101101011011", -- t[60251] = 30
      "0011110" when "01110101101011100", -- t[60252] = 30
      "0011110" when "01110101101011101", -- t[60253] = 30
      "0011110" when "01110101101011110", -- t[60254] = 30
      "0011110" when "01110101101011111", -- t[60255] = 30
      "0011110" when "01110101101100000", -- t[60256] = 30
      "0011110" when "01110101101100001", -- t[60257] = 30
      "0011110" when "01110101101100010", -- t[60258] = 30
      "0011110" when "01110101101100011", -- t[60259] = 30
      "0011110" when "01110101101100100", -- t[60260] = 30
      "0011110" when "01110101101100101", -- t[60261] = 30
      "0011110" when "01110101101100110", -- t[60262] = 30
      "0011110" when "01110101101100111", -- t[60263] = 30
      "0011110" when "01110101101101000", -- t[60264] = 30
      "0011110" when "01110101101101001", -- t[60265] = 30
      "0011110" when "01110101101101010", -- t[60266] = 30
      "0011110" when "01110101101101011", -- t[60267] = 30
      "0011110" when "01110101101101100", -- t[60268] = 30
      "0011110" when "01110101101101101", -- t[60269] = 30
      "0011110" when "01110101101101110", -- t[60270] = 30
      "0011110" when "01110101101101111", -- t[60271] = 30
      "0011110" when "01110101101110000", -- t[60272] = 30
      "0011110" when "01110101101110001", -- t[60273] = 30
      "0011110" when "01110101101110010", -- t[60274] = 30
      "0011110" when "01110101101110011", -- t[60275] = 30
      "0011110" when "01110101101110100", -- t[60276] = 30
      "0011110" when "01110101101110101", -- t[60277] = 30
      "0011110" when "01110101101110110", -- t[60278] = 30
      "0011110" when "01110101101110111", -- t[60279] = 30
      "0011110" when "01110101101111000", -- t[60280] = 30
      "0011110" when "01110101101111001", -- t[60281] = 30
      "0011110" when "01110101101111010", -- t[60282] = 30
      "0011110" when "01110101101111011", -- t[60283] = 30
      "0011110" when "01110101101111100", -- t[60284] = 30
      "0011110" when "01110101101111101", -- t[60285] = 30
      "0011110" when "01110101101111110", -- t[60286] = 30
      "0011110" when "01110101101111111", -- t[60287] = 30
      "0011110" when "01110101110000000", -- t[60288] = 30
      "0011110" when "01110101110000001", -- t[60289] = 30
      "0011110" when "01110101110000010", -- t[60290] = 30
      "0011110" when "01110101110000011", -- t[60291] = 30
      "0011110" when "01110101110000100", -- t[60292] = 30
      "0011110" when "01110101110000101", -- t[60293] = 30
      "0011110" when "01110101110000110", -- t[60294] = 30
      "0011110" when "01110101110000111", -- t[60295] = 30
      "0011110" when "01110101110001000", -- t[60296] = 30
      "0011110" when "01110101110001001", -- t[60297] = 30
      "0011110" when "01110101110001010", -- t[60298] = 30
      "0011110" when "01110101110001011", -- t[60299] = 30
      "0011110" when "01110101110001100", -- t[60300] = 30
      "0011110" when "01110101110001101", -- t[60301] = 30
      "0011110" when "01110101110001110", -- t[60302] = 30
      "0011110" when "01110101110001111", -- t[60303] = 30
      "0011110" when "01110101110010000", -- t[60304] = 30
      "0011110" when "01110101110010001", -- t[60305] = 30
      "0011110" when "01110101110010010", -- t[60306] = 30
      "0011110" when "01110101110010011", -- t[60307] = 30
      "0011110" when "01110101110010100", -- t[60308] = 30
      "0011110" when "01110101110010101", -- t[60309] = 30
      "0011110" when "01110101110010110", -- t[60310] = 30
      "0011110" when "01110101110010111", -- t[60311] = 30
      "0011110" when "01110101110011000", -- t[60312] = 30
      "0011110" when "01110101110011001", -- t[60313] = 30
      "0011110" when "01110101110011010", -- t[60314] = 30
      "0011110" when "01110101110011011", -- t[60315] = 30
      "0011110" when "01110101110011100", -- t[60316] = 30
      "0011110" when "01110101110011101", -- t[60317] = 30
      "0011110" when "01110101110011110", -- t[60318] = 30
      "0011110" when "01110101110011111", -- t[60319] = 30
      "0011110" when "01110101110100000", -- t[60320] = 30
      "0011110" when "01110101110100001", -- t[60321] = 30
      "0011110" when "01110101110100010", -- t[60322] = 30
      "0011110" when "01110101110100011", -- t[60323] = 30
      "0011110" when "01110101110100100", -- t[60324] = 30
      "0011110" when "01110101110100101", -- t[60325] = 30
      "0011110" when "01110101110100110", -- t[60326] = 30
      "0011110" when "01110101110100111", -- t[60327] = 30
      "0011110" when "01110101110101000", -- t[60328] = 30
      "0011110" when "01110101110101001", -- t[60329] = 30
      "0011110" when "01110101110101010", -- t[60330] = 30
      "0011110" when "01110101110101011", -- t[60331] = 30
      "0011110" when "01110101110101100", -- t[60332] = 30
      "0011110" when "01110101110101101", -- t[60333] = 30
      "0011110" when "01110101110101110", -- t[60334] = 30
      "0011110" when "01110101110101111", -- t[60335] = 30
      "0011110" when "01110101110110000", -- t[60336] = 30
      "0011110" when "01110101110110001", -- t[60337] = 30
      "0011110" when "01110101110110010", -- t[60338] = 30
      "0011110" when "01110101110110011", -- t[60339] = 30
      "0011110" when "01110101110110100", -- t[60340] = 30
      "0011110" when "01110101110110101", -- t[60341] = 30
      "0011110" when "01110101110110110", -- t[60342] = 30
      "0011110" when "01110101110110111", -- t[60343] = 30
      "0011110" when "01110101110111000", -- t[60344] = 30
      "0011110" when "01110101110111001", -- t[60345] = 30
      "0011110" when "01110101110111010", -- t[60346] = 30
      "0011110" when "01110101110111011", -- t[60347] = 30
      "0011110" when "01110101110111100", -- t[60348] = 30
      "0011110" when "01110101110111101", -- t[60349] = 30
      "0011110" when "01110101110111110", -- t[60350] = 30
      "0011110" when "01110101110111111", -- t[60351] = 30
      "0011110" when "01110101111000000", -- t[60352] = 30
      "0011110" when "01110101111000001", -- t[60353] = 30
      "0011110" when "01110101111000010", -- t[60354] = 30
      "0011110" when "01110101111000011", -- t[60355] = 30
      "0011110" when "01110101111000100", -- t[60356] = 30
      "0011110" when "01110101111000101", -- t[60357] = 30
      "0011110" when "01110101111000110", -- t[60358] = 30
      "0011110" when "01110101111000111", -- t[60359] = 30
      "0011110" when "01110101111001000", -- t[60360] = 30
      "0011110" when "01110101111001001", -- t[60361] = 30
      "0011110" when "01110101111001010", -- t[60362] = 30
      "0011110" when "01110101111001011", -- t[60363] = 30
      "0011110" when "01110101111001100", -- t[60364] = 30
      "0011110" when "01110101111001101", -- t[60365] = 30
      "0011110" when "01110101111001110", -- t[60366] = 30
      "0011110" when "01110101111001111", -- t[60367] = 30
      "0011110" when "01110101111010000", -- t[60368] = 30
      "0011110" when "01110101111010001", -- t[60369] = 30
      "0011110" when "01110101111010010", -- t[60370] = 30
      "0011110" when "01110101111010011", -- t[60371] = 30
      "0011110" when "01110101111010100", -- t[60372] = 30
      "0011110" when "01110101111010101", -- t[60373] = 30
      "0011110" when "01110101111010110", -- t[60374] = 30
      "0011110" when "01110101111010111", -- t[60375] = 30
      "0011110" when "01110101111011000", -- t[60376] = 30
      "0011110" when "01110101111011001", -- t[60377] = 30
      "0011110" when "01110101111011010", -- t[60378] = 30
      "0011110" when "01110101111011011", -- t[60379] = 30
      "0011110" when "01110101111011100", -- t[60380] = 30
      "0011110" when "01110101111011101", -- t[60381] = 30
      "0011110" when "01110101111011110", -- t[60382] = 30
      "0011110" when "01110101111011111", -- t[60383] = 30
      "0011110" when "01110101111100000", -- t[60384] = 30
      "0011110" when "01110101111100001", -- t[60385] = 30
      "0011110" when "01110101111100010", -- t[60386] = 30
      "0011110" when "01110101111100011", -- t[60387] = 30
      "0011110" when "01110101111100100", -- t[60388] = 30
      "0011110" when "01110101111100101", -- t[60389] = 30
      "0011110" when "01110101111100110", -- t[60390] = 30
      "0011110" when "01110101111100111", -- t[60391] = 30
      "0011110" when "01110101111101000", -- t[60392] = 30
      "0011110" when "01110101111101001", -- t[60393] = 30
      "0011110" when "01110101111101010", -- t[60394] = 30
      "0011110" when "01110101111101011", -- t[60395] = 30
      "0011110" when "01110101111101100", -- t[60396] = 30
      "0011110" when "01110101111101101", -- t[60397] = 30
      "0011110" when "01110101111101110", -- t[60398] = 30
      "0011110" when "01110101111101111", -- t[60399] = 30
      "0011110" when "01110101111110000", -- t[60400] = 30
      "0011110" when "01110101111110001", -- t[60401] = 30
      "0011110" when "01110101111110010", -- t[60402] = 30
      "0011110" when "01110101111110011", -- t[60403] = 30
      "0011110" when "01110101111110100", -- t[60404] = 30
      "0011110" when "01110101111110101", -- t[60405] = 30
      "0011110" when "01110101111110110", -- t[60406] = 30
      "0011110" when "01110101111110111", -- t[60407] = 30
      "0011110" when "01110101111111000", -- t[60408] = 30
      "0011110" when "01110101111111001", -- t[60409] = 30
      "0011110" when "01110101111111010", -- t[60410] = 30
      "0011110" when "01110101111111011", -- t[60411] = 30
      "0011110" when "01110101111111100", -- t[60412] = 30
      "0011110" when "01110101111111101", -- t[60413] = 30
      "0011110" when "01110101111111110", -- t[60414] = 30
      "0011110" when "01110101111111111", -- t[60415] = 30
      "0011110" when "01110110000000000", -- t[60416] = 30
      "0011110" when "01110110000000001", -- t[60417] = 30
      "0011110" when "01110110000000010", -- t[60418] = 30
      "0011110" when "01110110000000011", -- t[60419] = 30
      "0011110" when "01110110000000100", -- t[60420] = 30
      "0011110" when "01110110000000101", -- t[60421] = 30
      "0011110" when "01110110000000110", -- t[60422] = 30
      "0011110" when "01110110000000111", -- t[60423] = 30
      "0011110" when "01110110000001000", -- t[60424] = 30
      "0011110" when "01110110000001001", -- t[60425] = 30
      "0011110" when "01110110000001010", -- t[60426] = 30
      "0011110" when "01110110000001011", -- t[60427] = 30
      "0011110" when "01110110000001100", -- t[60428] = 30
      "0011110" when "01110110000001101", -- t[60429] = 30
      "0011110" when "01110110000001110", -- t[60430] = 30
      "0011110" when "01110110000001111", -- t[60431] = 30
      "0011110" when "01110110000010000", -- t[60432] = 30
      "0011110" when "01110110000010001", -- t[60433] = 30
      "0011110" when "01110110000010010", -- t[60434] = 30
      "0011110" when "01110110000010011", -- t[60435] = 30
      "0011110" when "01110110000010100", -- t[60436] = 30
      "0011110" when "01110110000010101", -- t[60437] = 30
      "0011110" when "01110110000010110", -- t[60438] = 30
      "0011110" when "01110110000010111", -- t[60439] = 30
      "0011110" when "01110110000011000", -- t[60440] = 30
      "0011110" when "01110110000011001", -- t[60441] = 30
      "0011110" when "01110110000011010", -- t[60442] = 30
      "0011110" when "01110110000011011", -- t[60443] = 30
      "0011110" when "01110110000011100", -- t[60444] = 30
      "0011110" when "01110110000011101", -- t[60445] = 30
      "0011110" when "01110110000011110", -- t[60446] = 30
      "0011110" when "01110110000011111", -- t[60447] = 30
      "0011110" when "01110110000100000", -- t[60448] = 30
      "0011110" when "01110110000100001", -- t[60449] = 30
      "0011110" when "01110110000100010", -- t[60450] = 30
      "0011110" when "01110110000100011", -- t[60451] = 30
      "0011110" when "01110110000100100", -- t[60452] = 30
      "0011110" when "01110110000100101", -- t[60453] = 30
      "0011110" when "01110110000100110", -- t[60454] = 30
      "0011110" when "01110110000100111", -- t[60455] = 30
      "0011110" when "01110110000101000", -- t[60456] = 30
      "0011110" when "01110110000101001", -- t[60457] = 30
      "0011110" when "01110110000101010", -- t[60458] = 30
      "0011110" when "01110110000101011", -- t[60459] = 30
      "0011110" when "01110110000101100", -- t[60460] = 30
      "0011110" when "01110110000101101", -- t[60461] = 30
      "0011110" when "01110110000101110", -- t[60462] = 30
      "0011110" when "01110110000101111", -- t[60463] = 30
      "0011110" when "01110110000110000", -- t[60464] = 30
      "0011110" when "01110110000110001", -- t[60465] = 30
      "0011110" when "01110110000110010", -- t[60466] = 30
      "0011110" when "01110110000110011", -- t[60467] = 30
      "0011110" when "01110110000110100", -- t[60468] = 30
      "0011110" when "01110110000110101", -- t[60469] = 30
      "0011110" when "01110110000110110", -- t[60470] = 30
      "0011110" when "01110110000110111", -- t[60471] = 30
      "0011110" when "01110110000111000", -- t[60472] = 30
      "0011110" when "01110110000111001", -- t[60473] = 30
      "0011110" when "01110110000111010", -- t[60474] = 30
      "0011110" when "01110110000111011", -- t[60475] = 30
      "0011110" when "01110110000111100", -- t[60476] = 30
      "0011110" when "01110110000111101", -- t[60477] = 30
      "0011110" when "01110110000111110", -- t[60478] = 30
      "0011110" when "01110110000111111", -- t[60479] = 30
      "0011110" when "01110110001000000", -- t[60480] = 30
      "0011110" when "01110110001000001", -- t[60481] = 30
      "0011110" when "01110110001000010", -- t[60482] = 30
      "0011110" when "01110110001000011", -- t[60483] = 30
      "0011110" when "01110110001000100", -- t[60484] = 30
      "0011110" when "01110110001000101", -- t[60485] = 30
      "0011110" when "01110110001000110", -- t[60486] = 30
      "0011110" when "01110110001000111", -- t[60487] = 30
      "0011110" when "01110110001001000", -- t[60488] = 30
      "0011110" when "01110110001001001", -- t[60489] = 30
      "0011110" when "01110110001001010", -- t[60490] = 30
      "0011110" when "01110110001001011", -- t[60491] = 30
      "0011110" when "01110110001001100", -- t[60492] = 30
      "0011110" when "01110110001001101", -- t[60493] = 30
      "0011110" when "01110110001001110", -- t[60494] = 30
      "0011110" when "01110110001001111", -- t[60495] = 30
      "0011110" when "01110110001010000", -- t[60496] = 30
      "0011110" when "01110110001010001", -- t[60497] = 30
      "0011110" when "01110110001010010", -- t[60498] = 30
      "0011110" when "01110110001010011", -- t[60499] = 30
      "0011110" when "01110110001010100", -- t[60500] = 30
      "0011110" when "01110110001010101", -- t[60501] = 30
      "0011110" when "01110110001010110", -- t[60502] = 30
      "0011110" when "01110110001010111", -- t[60503] = 30
      "0011110" when "01110110001011000", -- t[60504] = 30
      "0011110" when "01110110001011001", -- t[60505] = 30
      "0011110" when "01110110001011010", -- t[60506] = 30
      "0011110" when "01110110001011011", -- t[60507] = 30
      "0011110" when "01110110001011100", -- t[60508] = 30
      "0011110" when "01110110001011101", -- t[60509] = 30
      "0011110" when "01110110001011110", -- t[60510] = 30
      "0011110" when "01110110001011111", -- t[60511] = 30
      "0011110" when "01110110001100000", -- t[60512] = 30
      "0011110" when "01110110001100001", -- t[60513] = 30
      "0011110" when "01110110001100010", -- t[60514] = 30
      "0011110" when "01110110001100011", -- t[60515] = 30
      "0011110" when "01110110001100100", -- t[60516] = 30
      "0011110" when "01110110001100101", -- t[60517] = 30
      "0011110" when "01110110001100110", -- t[60518] = 30
      "0011110" when "01110110001100111", -- t[60519] = 30
      "0011110" when "01110110001101000", -- t[60520] = 30
      "0011110" when "01110110001101001", -- t[60521] = 30
      "0011110" when "01110110001101010", -- t[60522] = 30
      "0011110" when "01110110001101011", -- t[60523] = 30
      "0011110" when "01110110001101100", -- t[60524] = 30
      "0011110" when "01110110001101101", -- t[60525] = 30
      "0011110" when "01110110001101110", -- t[60526] = 30
      "0011110" when "01110110001101111", -- t[60527] = 30
      "0011110" when "01110110001110000", -- t[60528] = 30
      "0011110" when "01110110001110001", -- t[60529] = 30
      "0011110" when "01110110001110010", -- t[60530] = 30
      "0011110" when "01110110001110011", -- t[60531] = 30
      "0011110" when "01110110001110100", -- t[60532] = 30
      "0011110" when "01110110001110101", -- t[60533] = 30
      "0011110" when "01110110001110110", -- t[60534] = 30
      "0011110" when "01110110001110111", -- t[60535] = 30
      "0011110" when "01110110001111000", -- t[60536] = 30
      "0011110" when "01110110001111001", -- t[60537] = 30
      "0011110" when "01110110001111010", -- t[60538] = 30
      "0011110" when "01110110001111011", -- t[60539] = 30
      "0011110" when "01110110001111100", -- t[60540] = 30
      "0011110" when "01110110001111101", -- t[60541] = 30
      "0011110" when "01110110001111110", -- t[60542] = 30
      "0011110" when "01110110001111111", -- t[60543] = 30
      "0011110" when "01110110010000000", -- t[60544] = 30
      "0011110" when "01110110010000001", -- t[60545] = 30
      "0011110" when "01110110010000010", -- t[60546] = 30
      "0011110" when "01110110010000011", -- t[60547] = 30
      "0011110" when "01110110010000100", -- t[60548] = 30
      "0011110" when "01110110010000101", -- t[60549] = 30
      "0011110" when "01110110010000110", -- t[60550] = 30
      "0011110" when "01110110010000111", -- t[60551] = 30
      "0011110" when "01110110010001000", -- t[60552] = 30
      "0011110" when "01110110010001001", -- t[60553] = 30
      "0011110" when "01110110010001010", -- t[60554] = 30
      "0011110" when "01110110010001011", -- t[60555] = 30
      "0011110" when "01110110010001100", -- t[60556] = 30
      "0011110" when "01110110010001101", -- t[60557] = 30
      "0011110" when "01110110010001110", -- t[60558] = 30
      "0011110" when "01110110010001111", -- t[60559] = 30
      "0011110" when "01110110010010000", -- t[60560] = 30
      "0011110" when "01110110010010001", -- t[60561] = 30
      "0011110" when "01110110010010010", -- t[60562] = 30
      "0011110" when "01110110010010011", -- t[60563] = 30
      "0011110" when "01110110010010100", -- t[60564] = 30
      "0011110" when "01110110010010101", -- t[60565] = 30
      "0011110" when "01110110010010110", -- t[60566] = 30
      "0011110" when "01110110010010111", -- t[60567] = 30
      "0011110" when "01110110010011000", -- t[60568] = 30
      "0011110" when "01110110010011001", -- t[60569] = 30
      "0011110" when "01110110010011010", -- t[60570] = 30
      "0011110" when "01110110010011011", -- t[60571] = 30
      "0011110" when "01110110010011100", -- t[60572] = 30
      "0011110" when "01110110010011101", -- t[60573] = 30
      "0011110" when "01110110010011110", -- t[60574] = 30
      "0011110" when "01110110010011111", -- t[60575] = 30
      "0011110" when "01110110010100000", -- t[60576] = 30
      "0011110" when "01110110010100001", -- t[60577] = 30
      "0011110" when "01110110010100010", -- t[60578] = 30
      "0011110" when "01110110010100011", -- t[60579] = 30
      "0011110" when "01110110010100100", -- t[60580] = 30
      "0011110" when "01110110010100101", -- t[60581] = 30
      "0011110" when "01110110010100110", -- t[60582] = 30
      "0011110" when "01110110010100111", -- t[60583] = 30
      "0011110" when "01110110010101000", -- t[60584] = 30
      "0011110" when "01110110010101001", -- t[60585] = 30
      "0011110" when "01110110010101010", -- t[60586] = 30
      "0011110" when "01110110010101011", -- t[60587] = 30
      "0011110" when "01110110010101100", -- t[60588] = 30
      "0011110" when "01110110010101101", -- t[60589] = 30
      "0011110" when "01110110010101110", -- t[60590] = 30
      "0011110" when "01110110010101111", -- t[60591] = 30
      "0011110" when "01110110010110000", -- t[60592] = 30
      "0011110" when "01110110010110001", -- t[60593] = 30
      "0011110" when "01110110010110010", -- t[60594] = 30
      "0011110" when "01110110010110011", -- t[60595] = 30
      "0011110" when "01110110010110100", -- t[60596] = 30
      "0011110" when "01110110010110101", -- t[60597] = 30
      "0011110" when "01110110010110110", -- t[60598] = 30
      "0011110" when "01110110010110111", -- t[60599] = 30
      "0011110" when "01110110010111000", -- t[60600] = 30
      "0011110" when "01110110010111001", -- t[60601] = 30
      "0011110" when "01110110010111010", -- t[60602] = 30
      "0011110" when "01110110010111011", -- t[60603] = 30
      "0011110" when "01110110010111100", -- t[60604] = 30
      "0011110" when "01110110010111101", -- t[60605] = 30
      "0011110" when "01110110010111110", -- t[60606] = 30
      "0011110" when "01110110010111111", -- t[60607] = 30
      "0011110" when "01110110011000000", -- t[60608] = 30
      "0011110" when "01110110011000001", -- t[60609] = 30
      "0011110" when "01110110011000010", -- t[60610] = 30
      "0011110" when "01110110011000011", -- t[60611] = 30
      "0011110" when "01110110011000100", -- t[60612] = 30
      "0011110" when "01110110011000101", -- t[60613] = 30
      "0011110" when "01110110011000110", -- t[60614] = 30
      "0011110" when "01110110011000111", -- t[60615] = 30
      "0011110" when "01110110011001000", -- t[60616] = 30
      "0011110" when "01110110011001001", -- t[60617] = 30
      "0011110" when "01110110011001010", -- t[60618] = 30
      "0011110" when "01110110011001011", -- t[60619] = 30
      "0011110" when "01110110011001100", -- t[60620] = 30
      "0011110" when "01110110011001101", -- t[60621] = 30
      "0011111" when "01110110011001110", -- t[60622] = 31
      "0011111" when "01110110011001111", -- t[60623] = 31
      "0011111" when "01110110011010000", -- t[60624] = 31
      "0011111" when "01110110011010001", -- t[60625] = 31
      "0011111" when "01110110011010010", -- t[60626] = 31
      "0011111" when "01110110011010011", -- t[60627] = 31
      "0011111" when "01110110011010100", -- t[60628] = 31
      "0011111" when "01110110011010101", -- t[60629] = 31
      "0011111" when "01110110011010110", -- t[60630] = 31
      "0011111" when "01110110011010111", -- t[60631] = 31
      "0011111" when "01110110011011000", -- t[60632] = 31
      "0011111" when "01110110011011001", -- t[60633] = 31
      "0011111" when "01110110011011010", -- t[60634] = 31
      "0011111" when "01110110011011011", -- t[60635] = 31
      "0011111" when "01110110011011100", -- t[60636] = 31
      "0011111" when "01110110011011101", -- t[60637] = 31
      "0011111" when "01110110011011110", -- t[60638] = 31
      "0011111" when "01110110011011111", -- t[60639] = 31
      "0011111" when "01110110011100000", -- t[60640] = 31
      "0011111" when "01110110011100001", -- t[60641] = 31
      "0011111" when "01110110011100010", -- t[60642] = 31
      "0011111" when "01110110011100011", -- t[60643] = 31
      "0011111" when "01110110011100100", -- t[60644] = 31
      "0011111" when "01110110011100101", -- t[60645] = 31
      "0011111" when "01110110011100110", -- t[60646] = 31
      "0011111" when "01110110011100111", -- t[60647] = 31
      "0011111" when "01110110011101000", -- t[60648] = 31
      "0011111" when "01110110011101001", -- t[60649] = 31
      "0011111" when "01110110011101010", -- t[60650] = 31
      "0011111" when "01110110011101011", -- t[60651] = 31
      "0011111" when "01110110011101100", -- t[60652] = 31
      "0011111" when "01110110011101101", -- t[60653] = 31
      "0011111" when "01110110011101110", -- t[60654] = 31
      "0011111" when "01110110011101111", -- t[60655] = 31
      "0011111" when "01110110011110000", -- t[60656] = 31
      "0011111" when "01110110011110001", -- t[60657] = 31
      "0011111" when "01110110011110010", -- t[60658] = 31
      "0011111" when "01110110011110011", -- t[60659] = 31
      "0011111" when "01110110011110100", -- t[60660] = 31
      "0011111" when "01110110011110101", -- t[60661] = 31
      "0011111" when "01110110011110110", -- t[60662] = 31
      "0011111" when "01110110011110111", -- t[60663] = 31
      "0011111" when "01110110011111000", -- t[60664] = 31
      "0011111" when "01110110011111001", -- t[60665] = 31
      "0011111" when "01110110011111010", -- t[60666] = 31
      "0011111" when "01110110011111011", -- t[60667] = 31
      "0011111" when "01110110011111100", -- t[60668] = 31
      "0011111" when "01110110011111101", -- t[60669] = 31
      "0011111" when "01110110011111110", -- t[60670] = 31
      "0011111" when "01110110011111111", -- t[60671] = 31
      "0011111" when "01110110100000000", -- t[60672] = 31
      "0011111" when "01110110100000001", -- t[60673] = 31
      "0011111" when "01110110100000010", -- t[60674] = 31
      "0011111" when "01110110100000011", -- t[60675] = 31
      "0011111" when "01110110100000100", -- t[60676] = 31
      "0011111" when "01110110100000101", -- t[60677] = 31
      "0011111" when "01110110100000110", -- t[60678] = 31
      "0011111" when "01110110100000111", -- t[60679] = 31
      "0011111" when "01110110100001000", -- t[60680] = 31
      "0011111" when "01110110100001001", -- t[60681] = 31
      "0011111" when "01110110100001010", -- t[60682] = 31
      "0011111" when "01110110100001011", -- t[60683] = 31
      "0011111" when "01110110100001100", -- t[60684] = 31
      "0011111" when "01110110100001101", -- t[60685] = 31
      "0011111" when "01110110100001110", -- t[60686] = 31
      "0011111" when "01110110100001111", -- t[60687] = 31
      "0011111" when "01110110100010000", -- t[60688] = 31
      "0011111" when "01110110100010001", -- t[60689] = 31
      "0011111" when "01110110100010010", -- t[60690] = 31
      "0011111" when "01110110100010011", -- t[60691] = 31
      "0011111" when "01110110100010100", -- t[60692] = 31
      "0011111" when "01110110100010101", -- t[60693] = 31
      "0011111" when "01110110100010110", -- t[60694] = 31
      "0011111" when "01110110100010111", -- t[60695] = 31
      "0011111" when "01110110100011000", -- t[60696] = 31
      "0011111" when "01110110100011001", -- t[60697] = 31
      "0011111" when "01110110100011010", -- t[60698] = 31
      "0011111" when "01110110100011011", -- t[60699] = 31
      "0011111" when "01110110100011100", -- t[60700] = 31
      "0011111" when "01110110100011101", -- t[60701] = 31
      "0011111" when "01110110100011110", -- t[60702] = 31
      "0011111" when "01110110100011111", -- t[60703] = 31
      "0011111" when "01110110100100000", -- t[60704] = 31
      "0011111" when "01110110100100001", -- t[60705] = 31
      "0011111" when "01110110100100010", -- t[60706] = 31
      "0011111" when "01110110100100011", -- t[60707] = 31
      "0011111" when "01110110100100100", -- t[60708] = 31
      "0011111" when "01110110100100101", -- t[60709] = 31
      "0011111" when "01110110100100110", -- t[60710] = 31
      "0011111" when "01110110100100111", -- t[60711] = 31
      "0011111" when "01110110100101000", -- t[60712] = 31
      "0011111" when "01110110100101001", -- t[60713] = 31
      "0011111" when "01110110100101010", -- t[60714] = 31
      "0011111" when "01110110100101011", -- t[60715] = 31
      "0011111" when "01110110100101100", -- t[60716] = 31
      "0011111" when "01110110100101101", -- t[60717] = 31
      "0011111" when "01110110100101110", -- t[60718] = 31
      "0011111" when "01110110100101111", -- t[60719] = 31
      "0011111" when "01110110100110000", -- t[60720] = 31
      "0011111" when "01110110100110001", -- t[60721] = 31
      "0011111" when "01110110100110010", -- t[60722] = 31
      "0011111" when "01110110100110011", -- t[60723] = 31
      "0011111" when "01110110100110100", -- t[60724] = 31
      "0011111" when "01110110100110101", -- t[60725] = 31
      "0011111" when "01110110100110110", -- t[60726] = 31
      "0011111" when "01110110100110111", -- t[60727] = 31
      "0011111" when "01110110100111000", -- t[60728] = 31
      "0011111" when "01110110100111001", -- t[60729] = 31
      "0011111" when "01110110100111010", -- t[60730] = 31
      "0011111" when "01110110100111011", -- t[60731] = 31
      "0011111" when "01110110100111100", -- t[60732] = 31
      "0011111" when "01110110100111101", -- t[60733] = 31
      "0011111" when "01110110100111110", -- t[60734] = 31
      "0011111" when "01110110100111111", -- t[60735] = 31
      "0011111" when "01110110101000000", -- t[60736] = 31
      "0011111" when "01110110101000001", -- t[60737] = 31
      "0011111" when "01110110101000010", -- t[60738] = 31
      "0011111" when "01110110101000011", -- t[60739] = 31
      "0011111" when "01110110101000100", -- t[60740] = 31
      "0011111" when "01110110101000101", -- t[60741] = 31
      "0011111" when "01110110101000110", -- t[60742] = 31
      "0011111" when "01110110101000111", -- t[60743] = 31
      "0011111" when "01110110101001000", -- t[60744] = 31
      "0011111" when "01110110101001001", -- t[60745] = 31
      "0011111" when "01110110101001010", -- t[60746] = 31
      "0011111" when "01110110101001011", -- t[60747] = 31
      "0011111" when "01110110101001100", -- t[60748] = 31
      "0011111" when "01110110101001101", -- t[60749] = 31
      "0011111" when "01110110101001110", -- t[60750] = 31
      "0011111" when "01110110101001111", -- t[60751] = 31
      "0011111" when "01110110101010000", -- t[60752] = 31
      "0011111" when "01110110101010001", -- t[60753] = 31
      "0011111" when "01110110101010010", -- t[60754] = 31
      "0011111" when "01110110101010011", -- t[60755] = 31
      "0011111" when "01110110101010100", -- t[60756] = 31
      "0011111" when "01110110101010101", -- t[60757] = 31
      "0011111" when "01110110101010110", -- t[60758] = 31
      "0011111" when "01110110101010111", -- t[60759] = 31
      "0011111" when "01110110101011000", -- t[60760] = 31
      "0011111" when "01110110101011001", -- t[60761] = 31
      "0011111" when "01110110101011010", -- t[60762] = 31
      "0011111" when "01110110101011011", -- t[60763] = 31
      "0011111" when "01110110101011100", -- t[60764] = 31
      "0011111" when "01110110101011101", -- t[60765] = 31
      "0011111" when "01110110101011110", -- t[60766] = 31
      "0011111" when "01110110101011111", -- t[60767] = 31
      "0011111" when "01110110101100000", -- t[60768] = 31
      "0011111" when "01110110101100001", -- t[60769] = 31
      "0011111" when "01110110101100010", -- t[60770] = 31
      "0011111" when "01110110101100011", -- t[60771] = 31
      "0011111" when "01110110101100100", -- t[60772] = 31
      "0011111" when "01110110101100101", -- t[60773] = 31
      "0011111" when "01110110101100110", -- t[60774] = 31
      "0011111" when "01110110101100111", -- t[60775] = 31
      "0011111" when "01110110101101000", -- t[60776] = 31
      "0011111" when "01110110101101001", -- t[60777] = 31
      "0011111" when "01110110101101010", -- t[60778] = 31
      "0011111" when "01110110101101011", -- t[60779] = 31
      "0011111" when "01110110101101100", -- t[60780] = 31
      "0011111" when "01110110101101101", -- t[60781] = 31
      "0011111" when "01110110101101110", -- t[60782] = 31
      "0011111" when "01110110101101111", -- t[60783] = 31
      "0011111" when "01110110101110000", -- t[60784] = 31
      "0011111" when "01110110101110001", -- t[60785] = 31
      "0011111" when "01110110101110010", -- t[60786] = 31
      "0011111" when "01110110101110011", -- t[60787] = 31
      "0011111" when "01110110101110100", -- t[60788] = 31
      "0011111" when "01110110101110101", -- t[60789] = 31
      "0011111" when "01110110101110110", -- t[60790] = 31
      "0011111" when "01110110101110111", -- t[60791] = 31
      "0011111" when "01110110101111000", -- t[60792] = 31
      "0011111" when "01110110101111001", -- t[60793] = 31
      "0011111" when "01110110101111010", -- t[60794] = 31
      "0011111" when "01110110101111011", -- t[60795] = 31
      "0011111" when "01110110101111100", -- t[60796] = 31
      "0011111" when "01110110101111101", -- t[60797] = 31
      "0011111" when "01110110101111110", -- t[60798] = 31
      "0011111" when "01110110101111111", -- t[60799] = 31
      "0011111" when "01110110110000000", -- t[60800] = 31
      "0011111" when "01110110110000001", -- t[60801] = 31
      "0011111" when "01110110110000010", -- t[60802] = 31
      "0011111" when "01110110110000011", -- t[60803] = 31
      "0011111" when "01110110110000100", -- t[60804] = 31
      "0011111" when "01110110110000101", -- t[60805] = 31
      "0011111" when "01110110110000110", -- t[60806] = 31
      "0011111" when "01110110110000111", -- t[60807] = 31
      "0011111" when "01110110110001000", -- t[60808] = 31
      "0011111" when "01110110110001001", -- t[60809] = 31
      "0011111" when "01110110110001010", -- t[60810] = 31
      "0011111" when "01110110110001011", -- t[60811] = 31
      "0011111" when "01110110110001100", -- t[60812] = 31
      "0011111" when "01110110110001101", -- t[60813] = 31
      "0011111" when "01110110110001110", -- t[60814] = 31
      "0011111" when "01110110110001111", -- t[60815] = 31
      "0011111" when "01110110110010000", -- t[60816] = 31
      "0011111" when "01110110110010001", -- t[60817] = 31
      "0011111" when "01110110110010010", -- t[60818] = 31
      "0011111" when "01110110110010011", -- t[60819] = 31
      "0011111" when "01110110110010100", -- t[60820] = 31
      "0011111" when "01110110110010101", -- t[60821] = 31
      "0011111" when "01110110110010110", -- t[60822] = 31
      "0011111" when "01110110110010111", -- t[60823] = 31
      "0011111" when "01110110110011000", -- t[60824] = 31
      "0011111" when "01110110110011001", -- t[60825] = 31
      "0011111" when "01110110110011010", -- t[60826] = 31
      "0011111" when "01110110110011011", -- t[60827] = 31
      "0011111" when "01110110110011100", -- t[60828] = 31
      "0011111" when "01110110110011101", -- t[60829] = 31
      "0011111" when "01110110110011110", -- t[60830] = 31
      "0011111" when "01110110110011111", -- t[60831] = 31
      "0011111" when "01110110110100000", -- t[60832] = 31
      "0011111" when "01110110110100001", -- t[60833] = 31
      "0011111" when "01110110110100010", -- t[60834] = 31
      "0011111" when "01110110110100011", -- t[60835] = 31
      "0011111" when "01110110110100100", -- t[60836] = 31
      "0011111" when "01110110110100101", -- t[60837] = 31
      "0011111" when "01110110110100110", -- t[60838] = 31
      "0011111" when "01110110110100111", -- t[60839] = 31
      "0011111" when "01110110110101000", -- t[60840] = 31
      "0011111" when "01110110110101001", -- t[60841] = 31
      "0011111" when "01110110110101010", -- t[60842] = 31
      "0011111" when "01110110110101011", -- t[60843] = 31
      "0011111" when "01110110110101100", -- t[60844] = 31
      "0011111" when "01110110110101101", -- t[60845] = 31
      "0011111" when "01110110110101110", -- t[60846] = 31
      "0011111" when "01110110110101111", -- t[60847] = 31
      "0011111" when "01110110110110000", -- t[60848] = 31
      "0011111" when "01110110110110001", -- t[60849] = 31
      "0011111" when "01110110110110010", -- t[60850] = 31
      "0011111" when "01110110110110011", -- t[60851] = 31
      "0011111" when "01110110110110100", -- t[60852] = 31
      "0011111" when "01110110110110101", -- t[60853] = 31
      "0011111" when "01110110110110110", -- t[60854] = 31
      "0011111" when "01110110110110111", -- t[60855] = 31
      "0011111" when "01110110110111000", -- t[60856] = 31
      "0011111" when "01110110110111001", -- t[60857] = 31
      "0011111" when "01110110110111010", -- t[60858] = 31
      "0011111" when "01110110110111011", -- t[60859] = 31
      "0011111" when "01110110110111100", -- t[60860] = 31
      "0011111" when "01110110110111101", -- t[60861] = 31
      "0011111" when "01110110110111110", -- t[60862] = 31
      "0011111" when "01110110110111111", -- t[60863] = 31
      "0011111" when "01110110111000000", -- t[60864] = 31
      "0011111" when "01110110111000001", -- t[60865] = 31
      "0011111" when "01110110111000010", -- t[60866] = 31
      "0011111" when "01110110111000011", -- t[60867] = 31
      "0011111" when "01110110111000100", -- t[60868] = 31
      "0011111" when "01110110111000101", -- t[60869] = 31
      "0011111" when "01110110111000110", -- t[60870] = 31
      "0011111" when "01110110111000111", -- t[60871] = 31
      "0011111" when "01110110111001000", -- t[60872] = 31
      "0011111" when "01110110111001001", -- t[60873] = 31
      "0011111" when "01110110111001010", -- t[60874] = 31
      "0011111" when "01110110111001011", -- t[60875] = 31
      "0011111" when "01110110111001100", -- t[60876] = 31
      "0011111" when "01110110111001101", -- t[60877] = 31
      "0011111" when "01110110111001110", -- t[60878] = 31
      "0011111" when "01110110111001111", -- t[60879] = 31
      "0011111" when "01110110111010000", -- t[60880] = 31
      "0011111" when "01110110111010001", -- t[60881] = 31
      "0011111" when "01110110111010010", -- t[60882] = 31
      "0011111" when "01110110111010011", -- t[60883] = 31
      "0011111" when "01110110111010100", -- t[60884] = 31
      "0011111" when "01110110111010101", -- t[60885] = 31
      "0011111" when "01110110111010110", -- t[60886] = 31
      "0011111" when "01110110111010111", -- t[60887] = 31
      "0011111" when "01110110111011000", -- t[60888] = 31
      "0011111" when "01110110111011001", -- t[60889] = 31
      "0011111" when "01110110111011010", -- t[60890] = 31
      "0011111" when "01110110111011011", -- t[60891] = 31
      "0011111" when "01110110111011100", -- t[60892] = 31
      "0011111" when "01110110111011101", -- t[60893] = 31
      "0011111" when "01110110111011110", -- t[60894] = 31
      "0011111" when "01110110111011111", -- t[60895] = 31
      "0011111" when "01110110111100000", -- t[60896] = 31
      "0011111" when "01110110111100001", -- t[60897] = 31
      "0011111" when "01110110111100010", -- t[60898] = 31
      "0011111" when "01110110111100011", -- t[60899] = 31
      "0011111" when "01110110111100100", -- t[60900] = 31
      "0011111" when "01110110111100101", -- t[60901] = 31
      "0011111" when "01110110111100110", -- t[60902] = 31
      "0011111" when "01110110111100111", -- t[60903] = 31
      "0011111" when "01110110111101000", -- t[60904] = 31
      "0011111" when "01110110111101001", -- t[60905] = 31
      "0011111" when "01110110111101010", -- t[60906] = 31
      "0011111" when "01110110111101011", -- t[60907] = 31
      "0011111" when "01110110111101100", -- t[60908] = 31
      "0011111" when "01110110111101101", -- t[60909] = 31
      "0011111" when "01110110111101110", -- t[60910] = 31
      "0011111" when "01110110111101111", -- t[60911] = 31
      "0011111" when "01110110111110000", -- t[60912] = 31
      "0011111" when "01110110111110001", -- t[60913] = 31
      "0011111" when "01110110111110010", -- t[60914] = 31
      "0011111" when "01110110111110011", -- t[60915] = 31
      "0011111" when "01110110111110100", -- t[60916] = 31
      "0011111" when "01110110111110101", -- t[60917] = 31
      "0011111" when "01110110111110110", -- t[60918] = 31
      "0011111" when "01110110111110111", -- t[60919] = 31
      "0011111" when "01110110111111000", -- t[60920] = 31
      "0011111" when "01110110111111001", -- t[60921] = 31
      "0011111" when "01110110111111010", -- t[60922] = 31
      "0011111" when "01110110111111011", -- t[60923] = 31
      "0011111" when "01110110111111100", -- t[60924] = 31
      "0011111" when "01110110111111101", -- t[60925] = 31
      "0011111" when "01110110111111110", -- t[60926] = 31
      "0011111" when "01110110111111111", -- t[60927] = 31
      "0011111" when "01110111000000000", -- t[60928] = 31
      "0011111" when "01110111000000001", -- t[60929] = 31
      "0011111" when "01110111000000010", -- t[60930] = 31
      "0011111" when "01110111000000011", -- t[60931] = 31
      "0011111" when "01110111000000100", -- t[60932] = 31
      "0011111" when "01110111000000101", -- t[60933] = 31
      "0011111" when "01110111000000110", -- t[60934] = 31
      "0011111" when "01110111000000111", -- t[60935] = 31
      "0011111" when "01110111000001000", -- t[60936] = 31
      "0011111" when "01110111000001001", -- t[60937] = 31
      "0011111" when "01110111000001010", -- t[60938] = 31
      "0011111" when "01110111000001011", -- t[60939] = 31
      "0011111" when "01110111000001100", -- t[60940] = 31
      "0011111" when "01110111000001101", -- t[60941] = 31
      "0011111" when "01110111000001110", -- t[60942] = 31
      "0011111" when "01110111000001111", -- t[60943] = 31
      "0011111" when "01110111000010000", -- t[60944] = 31
      "0011111" when "01110111000010001", -- t[60945] = 31
      "0011111" when "01110111000010010", -- t[60946] = 31
      "0011111" when "01110111000010011", -- t[60947] = 31
      "0011111" when "01110111000010100", -- t[60948] = 31
      "0011111" when "01110111000010101", -- t[60949] = 31
      "0011111" when "01110111000010110", -- t[60950] = 31
      "0011111" when "01110111000010111", -- t[60951] = 31
      "0011111" when "01110111000011000", -- t[60952] = 31
      "0011111" when "01110111000011001", -- t[60953] = 31
      "0011111" when "01110111000011010", -- t[60954] = 31
      "0011111" when "01110111000011011", -- t[60955] = 31
      "0011111" when "01110111000011100", -- t[60956] = 31
      "0011111" when "01110111000011101", -- t[60957] = 31
      "0011111" when "01110111000011110", -- t[60958] = 31
      "0011111" when "01110111000011111", -- t[60959] = 31
      "0011111" when "01110111000100000", -- t[60960] = 31
      "0011111" when "01110111000100001", -- t[60961] = 31
      "0011111" when "01110111000100010", -- t[60962] = 31
      "0011111" when "01110111000100011", -- t[60963] = 31
      "0011111" when "01110111000100100", -- t[60964] = 31
      "0011111" when "01110111000100101", -- t[60965] = 31
      "0011111" when "01110111000100110", -- t[60966] = 31
      "0011111" when "01110111000100111", -- t[60967] = 31
      "0011111" when "01110111000101000", -- t[60968] = 31
      "0011111" when "01110111000101001", -- t[60969] = 31
      "0011111" when "01110111000101010", -- t[60970] = 31
      "0011111" when "01110111000101011", -- t[60971] = 31
      "0011111" when "01110111000101100", -- t[60972] = 31
      "0011111" when "01110111000101101", -- t[60973] = 31
      "0011111" when "01110111000101110", -- t[60974] = 31
      "0011111" when "01110111000101111", -- t[60975] = 31
      "0011111" when "01110111000110000", -- t[60976] = 31
      "0011111" when "01110111000110001", -- t[60977] = 31
      "0011111" when "01110111000110010", -- t[60978] = 31
      "0011111" when "01110111000110011", -- t[60979] = 31
      "0011111" when "01110111000110100", -- t[60980] = 31
      "0011111" when "01110111000110101", -- t[60981] = 31
      "0011111" when "01110111000110110", -- t[60982] = 31
      "0011111" when "01110111000110111", -- t[60983] = 31
      "0011111" when "01110111000111000", -- t[60984] = 31
      "0011111" when "01110111000111001", -- t[60985] = 31
      "0011111" when "01110111000111010", -- t[60986] = 31
      "0011111" when "01110111000111011", -- t[60987] = 31
      "0011111" when "01110111000111100", -- t[60988] = 31
      "0011111" when "01110111000111101", -- t[60989] = 31
      "0011111" when "01110111000111110", -- t[60990] = 31
      "0011111" when "01110111000111111", -- t[60991] = 31
      "0011111" when "01110111001000000", -- t[60992] = 31
      "0011111" when "01110111001000001", -- t[60993] = 31
      "0011111" when "01110111001000010", -- t[60994] = 31
      "0011111" when "01110111001000011", -- t[60995] = 31
      "0011111" when "01110111001000100", -- t[60996] = 31
      "0011111" when "01110111001000101", -- t[60997] = 31
      "0011111" when "01110111001000110", -- t[60998] = 31
      "0011111" when "01110111001000111", -- t[60999] = 31
      "0011111" when "01110111001001000", -- t[61000] = 31
      "0011111" when "01110111001001001", -- t[61001] = 31
      "0011111" when "01110111001001010", -- t[61002] = 31
      "0100000" when "01110111001001011", -- t[61003] = 32
      "0100000" when "01110111001001100", -- t[61004] = 32
      "0100000" when "01110111001001101", -- t[61005] = 32
      "0100000" when "01110111001001110", -- t[61006] = 32
      "0100000" when "01110111001001111", -- t[61007] = 32
      "0100000" when "01110111001010000", -- t[61008] = 32
      "0100000" when "01110111001010001", -- t[61009] = 32
      "0100000" when "01110111001010010", -- t[61010] = 32
      "0100000" when "01110111001010011", -- t[61011] = 32
      "0100000" when "01110111001010100", -- t[61012] = 32
      "0100000" when "01110111001010101", -- t[61013] = 32
      "0100000" when "01110111001010110", -- t[61014] = 32
      "0100000" when "01110111001010111", -- t[61015] = 32
      "0100000" when "01110111001011000", -- t[61016] = 32
      "0100000" when "01110111001011001", -- t[61017] = 32
      "0100000" when "01110111001011010", -- t[61018] = 32
      "0100000" when "01110111001011011", -- t[61019] = 32
      "0100000" when "01110111001011100", -- t[61020] = 32
      "0100000" when "01110111001011101", -- t[61021] = 32
      "0100000" when "01110111001011110", -- t[61022] = 32
      "0100000" when "01110111001011111", -- t[61023] = 32
      "0100000" when "01110111001100000", -- t[61024] = 32
      "0100000" when "01110111001100001", -- t[61025] = 32
      "0100000" when "01110111001100010", -- t[61026] = 32
      "0100000" when "01110111001100011", -- t[61027] = 32
      "0100000" when "01110111001100100", -- t[61028] = 32
      "0100000" when "01110111001100101", -- t[61029] = 32
      "0100000" when "01110111001100110", -- t[61030] = 32
      "0100000" when "01110111001100111", -- t[61031] = 32
      "0100000" when "01110111001101000", -- t[61032] = 32
      "0100000" when "01110111001101001", -- t[61033] = 32
      "0100000" when "01110111001101010", -- t[61034] = 32
      "0100000" when "01110111001101011", -- t[61035] = 32
      "0100000" when "01110111001101100", -- t[61036] = 32
      "0100000" when "01110111001101101", -- t[61037] = 32
      "0100000" when "01110111001101110", -- t[61038] = 32
      "0100000" when "01110111001101111", -- t[61039] = 32
      "0100000" when "01110111001110000", -- t[61040] = 32
      "0100000" when "01110111001110001", -- t[61041] = 32
      "0100000" when "01110111001110010", -- t[61042] = 32
      "0100000" when "01110111001110011", -- t[61043] = 32
      "0100000" when "01110111001110100", -- t[61044] = 32
      "0100000" when "01110111001110101", -- t[61045] = 32
      "0100000" when "01110111001110110", -- t[61046] = 32
      "0100000" when "01110111001110111", -- t[61047] = 32
      "0100000" when "01110111001111000", -- t[61048] = 32
      "0100000" when "01110111001111001", -- t[61049] = 32
      "0100000" when "01110111001111010", -- t[61050] = 32
      "0100000" when "01110111001111011", -- t[61051] = 32
      "0100000" when "01110111001111100", -- t[61052] = 32
      "0100000" when "01110111001111101", -- t[61053] = 32
      "0100000" when "01110111001111110", -- t[61054] = 32
      "0100000" when "01110111001111111", -- t[61055] = 32
      "0100000" when "01110111010000000", -- t[61056] = 32
      "0100000" when "01110111010000001", -- t[61057] = 32
      "0100000" when "01110111010000010", -- t[61058] = 32
      "0100000" when "01110111010000011", -- t[61059] = 32
      "0100000" when "01110111010000100", -- t[61060] = 32
      "0100000" when "01110111010000101", -- t[61061] = 32
      "0100000" when "01110111010000110", -- t[61062] = 32
      "0100000" when "01110111010000111", -- t[61063] = 32
      "0100000" when "01110111010001000", -- t[61064] = 32
      "0100000" when "01110111010001001", -- t[61065] = 32
      "0100000" when "01110111010001010", -- t[61066] = 32
      "0100000" when "01110111010001011", -- t[61067] = 32
      "0100000" when "01110111010001100", -- t[61068] = 32
      "0100000" when "01110111010001101", -- t[61069] = 32
      "0100000" when "01110111010001110", -- t[61070] = 32
      "0100000" when "01110111010001111", -- t[61071] = 32
      "0100000" when "01110111010010000", -- t[61072] = 32
      "0100000" when "01110111010010001", -- t[61073] = 32
      "0100000" when "01110111010010010", -- t[61074] = 32
      "0100000" when "01110111010010011", -- t[61075] = 32
      "0100000" when "01110111010010100", -- t[61076] = 32
      "0100000" when "01110111010010101", -- t[61077] = 32
      "0100000" when "01110111010010110", -- t[61078] = 32
      "0100000" when "01110111010010111", -- t[61079] = 32
      "0100000" when "01110111010011000", -- t[61080] = 32
      "0100000" when "01110111010011001", -- t[61081] = 32
      "0100000" when "01110111010011010", -- t[61082] = 32
      "0100000" when "01110111010011011", -- t[61083] = 32
      "0100000" when "01110111010011100", -- t[61084] = 32
      "0100000" when "01110111010011101", -- t[61085] = 32
      "0100000" when "01110111010011110", -- t[61086] = 32
      "0100000" when "01110111010011111", -- t[61087] = 32
      "0100000" when "01110111010100000", -- t[61088] = 32
      "0100000" when "01110111010100001", -- t[61089] = 32
      "0100000" when "01110111010100010", -- t[61090] = 32
      "0100000" when "01110111010100011", -- t[61091] = 32
      "0100000" when "01110111010100100", -- t[61092] = 32
      "0100000" when "01110111010100101", -- t[61093] = 32
      "0100000" when "01110111010100110", -- t[61094] = 32
      "0100000" when "01110111010100111", -- t[61095] = 32
      "0100000" when "01110111010101000", -- t[61096] = 32
      "0100000" when "01110111010101001", -- t[61097] = 32
      "0100000" when "01110111010101010", -- t[61098] = 32
      "0100000" when "01110111010101011", -- t[61099] = 32
      "0100000" when "01110111010101100", -- t[61100] = 32
      "0100000" when "01110111010101101", -- t[61101] = 32
      "0100000" when "01110111010101110", -- t[61102] = 32
      "0100000" when "01110111010101111", -- t[61103] = 32
      "0100000" when "01110111010110000", -- t[61104] = 32
      "0100000" when "01110111010110001", -- t[61105] = 32
      "0100000" when "01110111010110010", -- t[61106] = 32
      "0100000" when "01110111010110011", -- t[61107] = 32
      "0100000" when "01110111010110100", -- t[61108] = 32
      "0100000" when "01110111010110101", -- t[61109] = 32
      "0100000" when "01110111010110110", -- t[61110] = 32
      "0100000" when "01110111010110111", -- t[61111] = 32
      "0100000" when "01110111010111000", -- t[61112] = 32
      "0100000" when "01110111010111001", -- t[61113] = 32
      "0100000" when "01110111010111010", -- t[61114] = 32
      "0100000" when "01110111010111011", -- t[61115] = 32
      "0100000" when "01110111010111100", -- t[61116] = 32
      "0100000" when "01110111010111101", -- t[61117] = 32
      "0100000" when "01110111010111110", -- t[61118] = 32
      "0100000" when "01110111010111111", -- t[61119] = 32
      "0100000" when "01110111011000000", -- t[61120] = 32
      "0100000" when "01110111011000001", -- t[61121] = 32
      "0100000" when "01110111011000010", -- t[61122] = 32
      "0100000" when "01110111011000011", -- t[61123] = 32
      "0100000" when "01110111011000100", -- t[61124] = 32
      "0100000" when "01110111011000101", -- t[61125] = 32
      "0100000" when "01110111011000110", -- t[61126] = 32
      "0100000" when "01110111011000111", -- t[61127] = 32
      "0100000" when "01110111011001000", -- t[61128] = 32
      "0100000" when "01110111011001001", -- t[61129] = 32
      "0100000" when "01110111011001010", -- t[61130] = 32
      "0100000" when "01110111011001011", -- t[61131] = 32
      "0100000" when "01110111011001100", -- t[61132] = 32
      "0100000" when "01110111011001101", -- t[61133] = 32
      "0100000" when "01110111011001110", -- t[61134] = 32
      "0100000" when "01110111011001111", -- t[61135] = 32
      "0100000" when "01110111011010000", -- t[61136] = 32
      "0100000" when "01110111011010001", -- t[61137] = 32
      "0100000" when "01110111011010010", -- t[61138] = 32
      "0100000" when "01110111011010011", -- t[61139] = 32
      "0100000" when "01110111011010100", -- t[61140] = 32
      "0100000" when "01110111011010101", -- t[61141] = 32
      "0100000" when "01110111011010110", -- t[61142] = 32
      "0100000" when "01110111011010111", -- t[61143] = 32
      "0100000" when "01110111011011000", -- t[61144] = 32
      "0100000" when "01110111011011001", -- t[61145] = 32
      "0100000" when "01110111011011010", -- t[61146] = 32
      "0100000" when "01110111011011011", -- t[61147] = 32
      "0100000" when "01110111011011100", -- t[61148] = 32
      "0100000" when "01110111011011101", -- t[61149] = 32
      "0100000" when "01110111011011110", -- t[61150] = 32
      "0100000" when "01110111011011111", -- t[61151] = 32
      "0100000" when "01110111011100000", -- t[61152] = 32
      "0100000" when "01110111011100001", -- t[61153] = 32
      "0100000" when "01110111011100010", -- t[61154] = 32
      "0100000" when "01110111011100011", -- t[61155] = 32
      "0100000" when "01110111011100100", -- t[61156] = 32
      "0100000" when "01110111011100101", -- t[61157] = 32
      "0100000" when "01110111011100110", -- t[61158] = 32
      "0100000" when "01110111011100111", -- t[61159] = 32
      "0100000" when "01110111011101000", -- t[61160] = 32
      "0100000" when "01110111011101001", -- t[61161] = 32
      "0100000" when "01110111011101010", -- t[61162] = 32
      "0100000" when "01110111011101011", -- t[61163] = 32
      "0100000" when "01110111011101100", -- t[61164] = 32
      "0100000" when "01110111011101101", -- t[61165] = 32
      "0100000" when "01110111011101110", -- t[61166] = 32
      "0100000" when "01110111011101111", -- t[61167] = 32
      "0100000" when "01110111011110000", -- t[61168] = 32
      "0100000" when "01110111011110001", -- t[61169] = 32
      "0100000" when "01110111011110010", -- t[61170] = 32
      "0100000" when "01110111011110011", -- t[61171] = 32
      "0100000" when "01110111011110100", -- t[61172] = 32
      "0100000" when "01110111011110101", -- t[61173] = 32
      "0100000" when "01110111011110110", -- t[61174] = 32
      "0100000" when "01110111011110111", -- t[61175] = 32
      "0100000" when "01110111011111000", -- t[61176] = 32
      "0100000" when "01110111011111001", -- t[61177] = 32
      "0100000" when "01110111011111010", -- t[61178] = 32
      "0100000" when "01110111011111011", -- t[61179] = 32
      "0100000" when "01110111011111100", -- t[61180] = 32
      "0100000" when "01110111011111101", -- t[61181] = 32
      "0100000" when "01110111011111110", -- t[61182] = 32
      "0100000" when "01110111011111111", -- t[61183] = 32
      "0100000" when "01110111100000000", -- t[61184] = 32
      "0100000" when "01110111100000001", -- t[61185] = 32
      "0100000" when "01110111100000010", -- t[61186] = 32
      "0100000" when "01110111100000011", -- t[61187] = 32
      "0100000" when "01110111100000100", -- t[61188] = 32
      "0100000" when "01110111100000101", -- t[61189] = 32
      "0100000" when "01110111100000110", -- t[61190] = 32
      "0100000" when "01110111100000111", -- t[61191] = 32
      "0100000" when "01110111100001000", -- t[61192] = 32
      "0100000" when "01110111100001001", -- t[61193] = 32
      "0100000" when "01110111100001010", -- t[61194] = 32
      "0100000" when "01110111100001011", -- t[61195] = 32
      "0100000" when "01110111100001100", -- t[61196] = 32
      "0100000" when "01110111100001101", -- t[61197] = 32
      "0100000" when "01110111100001110", -- t[61198] = 32
      "0100000" when "01110111100001111", -- t[61199] = 32
      "0100000" when "01110111100010000", -- t[61200] = 32
      "0100000" when "01110111100010001", -- t[61201] = 32
      "0100000" when "01110111100010010", -- t[61202] = 32
      "0100000" when "01110111100010011", -- t[61203] = 32
      "0100000" when "01110111100010100", -- t[61204] = 32
      "0100000" when "01110111100010101", -- t[61205] = 32
      "0100000" when "01110111100010110", -- t[61206] = 32
      "0100000" when "01110111100010111", -- t[61207] = 32
      "0100000" when "01110111100011000", -- t[61208] = 32
      "0100000" when "01110111100011001", -- t[61209] = 32
      "0100000" when "01110111100011010", -- t[61210] = 32
      "0100000" when "01110111100011011", -- t[61211] = 32
      "0100000" when "01110111100011100", -- t[61212] = 32
      "0100000" when "01110111100011101", -- t[61213] = 32
      "0100000" when "01110111100011110", -- t[61214] = 32
      "0100000" when "01110111100011111", -- t[61215] = 32
      "0100000" when "01110111100100000", -- t[61216] = 32
      "0100000" when "01110111100100001", -- t[61217] = 32
      "0100000" when "01110111100100010", -- t[61218] = 32
      "0100000" when "01110111100100011", -- t[61219] = 32
      "0100000" when "01110111100100100", -- t[61220] = 32
      "0100000" when "01110111100100101", -- t[61221] = 32
      "0100000" when "01110111100100110", -- t[61222] = 32
      "0100000" when "01110111100100111", -- t[61223] = 32
      "0100000" when "01110111100101000", -- t[61224] = 32
      "0100000" when "01110111100101001", -- t[61225] = 32
      "0100000" when "01110111100101010", -- t[61226] = 32
      "0100000" when "01110111100101011", -- t[61227] = 32
      "0100000" when "01110111100101100", -- t[61228] = 32
      "0100000" when "01110111100101101", -- t[61229] = 32
      "0100000" when "01110111100101110", -- t[61230] = 32
      "0100000" when "01110111100101111", -- t[61231] = 32
      "0100000" when "01110111100110000", -- t[61232] = 32
      "0100000" when "01110111100110001", -- t[61233] = 32
      "0100000" when "01110111100110010", -- t[61234] = 32
      "0100000" when "01110111100110011", -- t[61235] = 32
      "0100000" when "01110111100110100", -- t[61236] = 32
      "0100000" when "01110111100110101", -- t[61237] = 32
      "0100000" when "01110111100110110", -- t[61238] = 32
      "0100000" when "01110111100110111", -- t[61239] = 32
      "0100000" when "01110111100111000", -- t[61240] = 32
      "0100000" when "01110111100111001", -- t[61241] = 32
      "0100000" when "01110111100111010", -- t[61242] = 32
      "0100000" when "01110111100111011", -- t[61243] = 32
      "0100000" when "01110111100111100", -- t[61244] = 32
      "0100000" when "01110111100111101", -- t[61245] = 32
      "0100000" when "01110111100111110", -- t[61246] = 32
      "0100000" when "01110111100111111", -- t[61247] = 32
      "0100000" when "01110111101000000", -- t[61248] = 32
      "0100000" when "01110111101000001", -- t[61249] = 32
      "0100000" when "01110111101000010", -- t[61250] = 32
      "0100000" when "01110111101000011", -- t[61251] = 32
      "0100000" when "01110111101000100", -- t[61252] = 32
      "0100000" when "01110111101000101", -- t[61253] = 32
      "0100000" when "01110111101000110", -- t[61254] = 32
      "0100000" when "01110111101000111", -- t[61255] = 32
      "0100000" when "01110111101001000", -- t[61256] = 32
      "0100000" when "01110111101001001", -- t[61257] = 32
      "0100000" when "01110111101001010", -- t[61258] = 32
      "0100000" when "01110111101001011", -- t[61259] = 32
      "0100000" when "01110111101001100", -- t[61260] = 32
      "0100000" when "01110111101001101", -- t[61261] = 32
      "0100000" when "01110111101001110", -- t[61262] = 32
      "0100000" when "01110111101001111", -- t[61263] = 32
      "0100000" when "01110111101010000", -- t[61264] = 32
      "0100000" when "01110111101010001", -- t[61265] = 32
      "0100000" when "01110111101010010", -- t[61266] = 32
      "0100000" when "01110111101010011", -- t[61267] = 32
      "0100000" when "01110111101010100", -- t[61268] = 32
      "0100000" when "01110111101010101", -- t[61269] = 32
      "0100000" when "01110111101010110", -- t[61270] = 32
      "0100000" when "01110111101010111", -- t[61271] = 32
      "0100000" when "01110111101011000", -- t[61272] = 32
      "0100000" when "01110111101011001", -- t[61273] = 32
      "0100000" when "01110111101011010", -- t[61274] = 32
      "0100000" when "01110111101011011", -- t[61275] = 32
      "0100000" when "01110111101011100", -- t[61276] = 32
      "0100000" when "01110111101011101", -- t[61277] = 32
      "0100000" when "01110111101011110", -- t[61278] = 32
      "0100000" when "01110111101011111", -- t[61279] = 32
      "0100000" when "01110111101100000", -- t[61280] = 32
      "0100000" when "01110111101100001", -- t[61281] = 32
      "0100000" when "01110111101100010", -- t[61282] = 32
      "0100000" when "01110111101100011", -- t[61283] = 32
      "0100000" when "01110111101100100", -- t[61284] = 32
      "0100000" when "01110111101100101", -- t[61285] = 32
      "0100000" when "01110111101100110", -- t[61286] = 32
      "0100000" when "01110111101100111", -- t[61287] = 32
      "0100000" when "01110111101101000", -- t[61288] = 32
      "0100000" when "01110111101101001", -- t[61289] = 32
      "0100000" when "01110111101101010", -- t[61290] = 32
      "0100000" when "01110111101101011", -- t[61291] = 32
      "0100000" when "01110111101101100", -- t[61292] = 32
      "0100000" when "01110111101101101", -- t[61293] = 32
      "0100000" when "01110111101101110", -- t[61294] = 32
      "0100000" when "01110111101101111", -- t[61295] = 32
      "0100000" when "01110111101110000", -- t[61296] = 32
      "0100000" when "01110111101110001", -- t[61297] = 32
      "0100000" when "01110111101110010", -- t[61298] = 32
      "0100000" when "01110111101110011", -- t[61299] = 32
      "0100000" when "01110111101110100", -- t[61300] = 32
      "0100000" when "01110111101110101", -- t[61301] = 32
      "0100000" when "01110111101110110", -- t[61302] = 32
      "0100000" when "01110111101110111", -- t[61303] = 32
      "0100000" when "01110111101111000", -- t[61304] = 32
      "0100000" when "01110111101111001", -- t[61305] = 32
      "0100000" when "01110111101111010", -- t[61306] = 32
      "0100000" when "01110111101111011", -- t[61307] = 32
      "0100000" when "01110111101111100", -- t[61308] = 32
      "0100000" when "01110111101111101", -- t[61309] = 32
      "0100000" when "01110111101111110", -- t[61310] = 32
      "0100000" when "01110111101111111", -- t[61311] = 32
      "0100000" when "01110111110000000", -- t[61312] = 32
      "0100000" when "01110111110000001", -- t[61313] = 32
      "0100000" when "01110111110000010", -- t[61314] = 32
      "0100000" when "01110111110000011", -- t[61315] = 32
      "0100000" when "01110111110000100", -- t[61316] = 32
      "0100000" when "01110111110000101", -- t[61317] = 32
      "0100000" when "01110111110000110", -- t[61318] = 32
      "0100000" when "01110111110000111", -- t[61319] = 32
      "0100000" when "01110111110001000", -- t[61320] = 32
      "0100000" when "01110111110001001", -- t[61321] = 32
      "0100000" when "01110111110001010", -- t[61322] = 32
      "0100000" when "01110111110001011", -- t[61323] = 32
      "0100000" when "01110111110001100", -- t[61324] = 32
      "0100000" when "01110111110001101", -- t[61325] = 32
      "0100000" when "01110111110001110", -- t[61326] = 32
      "0100000" when "01110111110001111", -- t[61327] = 32
      "0100000" when "01110111110010000", -- t[61328] = 32
      "0100000" when "01110111110010001", -- t[61329] = 32
      "0100000" when "01110111110010010", -- t[61330] = 32
      "0100000" when "01110111110010011", -- t[61331] = 32
      "0100000" when "01110111110010100", -- t[61332] = 32
      "0100000" when "01110111110010101", -- t[61333] = 32
      "0100000" when "01110111110010110", -- t[61334] = 32
      "0100000" when "01110111110010111", -- t[61335] = 32
      "0100000" when "01110111110011000", -- t[61336] = 32
      "0100000" when "01110111110011001", -- t[61337] = 32
      "0100000" when "01110111110011010", -- t[61338] = 32
      "0100000" when "01110111110011011", -- t[61339] = 32
      "0100000" when "01110111110011100", -- t[61340] = 32
      "0100000" when "01110111110011101", -- t[61341] = 32
      "0100000" when "01110111110011110", -- t[61342] = 32
      "0100000" when "01110111110011111", -- t[61343] = 32
      "0100000" when "01110111110100000", -- t[61344] = 32
      "0100000" when "01110111110100001", -- t[61345] = 32
      "0100000" when "01110111110100010", -- t[61346] = 32
      "0100000" when "01110111110100011", -- t[61347] = 32
      "0100000" when "01110111110100100", -- t[61348] = 32
      "0100000" when "01110111110100101", -- t[61349] = 32
      "0100000" when "01110111110100110", -- t[61350] = 32
      "0100000" when "01110111110100111", -- t[61351] = 32
      "0100000" when "01110111110101000", -- t[61352] = 32
      "0100000" when "01110111110101001", -- t[61353] = 32
      "0100000" when "01110111110101010", -- t[61354] = 32
      "0100000" when "01110111110101011", -- t[61355] = 32
      "0100000" when "01110111110101100", -- t[61356] = 32
      "0100000" when "01110111110101101", -- t[61357] = 32
      "0100000" when "01110111110101110", -- t[61358] = 32
      "0100000" when "01110111110101111", -- t[61359] = 32
      "0100000" when "01110111110110000", -- t[61360] = 32
      "0100000" when "01110111110110001", -- t[61361] = 32
      "0100000" when "01110111110110010", -- t[61362] = 32
      "0100000" when "01110111110110011", -- t[61363] = 32
      "0100000" when "01110111110110100", -- t[61364] = 32
      "0100000" when "01110111110110101", -- t[61365] = 32
      "0100000" when "01110111110110110", -- t[61366] = 32
      "0100000" when "01110111110110111", -- t[61367] = 32
      "0100000" when "01110111110111000", -- t[61368] = 32
      "0100000" when "01110111110111001", -- t[61369] = 32
      "0100000" when "01110111110111010", -- t[61370] = 32
      "0100000" when "01110111110111011", -- t[61371] = 32
      "0100001" when "01110111110111100", -- t[61372] = 33
      "0100001" when "01110111110111101", -- t[61373] = 33
      "0100001" when "01110111110111110", -- t[61374] = 33
      "0100001" when "01110111110111111", -- t[61375] = 33
      "0100001" when "01110111111000000", -- t[61376] = 33
      "0100001" when "01110111111000001", -- t[61377] = 33
      "0100001" when "01110111111000010", -- t[61378] = 33
      "0100001" when "01110111111000011", -- t[61379] = 33
      "0100001" when "01110111111000100", -- t[61380] = 33
      "0100001" when "01110111111000101", -- t[61381] = 33
      "0100001" when "01110111111000110", -- t[61382] = 33
      "0100001" when "01110111111000111", -- t[61383] = 33
      "0100001" when "01110111111001000", -- t[61384] = 33
      "0100001" when "01110111111001001", -- t[61385] = 33
      "0100001" when "01110111111001010", -- t[61386] = 33
      "0100001" when "01110111111001011", -- t[61387] = 33
      "0100001" when "01110111111001100", -- t[61388] = 33
      "0100001" when "01110111111001101", -- t[61389] = 33
      "0100001" when "01110111111001110", -- t[61390] = 33
      "0100001" when "01110111111001111", -- t[61391] = 33
      "0100001" when "01110111111010000", -- t[61392] = 33
      "0100001" when "01110111111010001", -- t[61393] = 33
      "0100001" when "01110111111010010", -- t[61394] = 33
      "0100001" when "01110111111010011", -- t[61395] = 33
      "0100001" when "01110111111010100", -- t[61396] = 33
      "0100001" when "01110111111010101", -- t[61397] = 33
      "0100001" when "01110111111010110", -- t[61398] = 33
      "0100001" when "01110111111010111", -- t[61399] = 33
      "0100001" when "01110111111011000", -- t[61400] = 33
      "0100001" when "01110111111011001", -- t[61401] = 33
      "0100001" when "01110111111011010", -- t[61402] = 33
      "0100001" when "01110111111011011", -- t[61403] = 33
      "0100001" when "01110111111011100", -- t[61404] = 33
      "0100001" when "01110111111011101", -- t[61405] = 33
      "0100001" when "01110111111011110", -- t[61406] = 33
      "0100001" when "01110111111011111", -- t[61407] = 33
      "0100001" when "01110111111100000", -- t[61408] = 33
      "0100001" when "01110111111100001", -- t[61409] = 33
      "0100001" when "01110111111100010", -- t[61410] = 33
      "0100001" when "01110111111100011", -- t[61411] = 33
      "0100001" when "01110111111100100", -- t[61412] = 33
      "0100001" when "01110111111100101", -- t[61413] = 33
      "0100001" when "01110111111100110", -- t[61414] = 33
      "0100001" when "01110111111100111", -- t[61415] = 33
      "0100001" when "01110111111101000", -- t[61416] = 33
      "0100001" when "01110111111101001", -- t[61417] = 33
      "0100001" when "01110111111101010", -- t[61418] = 33
      "0100001" when "01110111111101011", -- t[61419] = 33
      "0100001" when "01110111111101100", -- t[61420] = 33
      "0100001" when "01110111111101101", -- t[61421] = 33
      "0100001" when "01110111111101110", -- t[61422] = 33
      "0100001" when "01110111111101111", -- t[61423] = 33
      "0100001" when "01110111111110000", -- t[61424] = 33
      "0100001" when "01110111111110001", -- t[61425] = 33
      "0100001" when "01110111111110010", -- t[61426] = 33
      "0100001" when "01110111111110011", -- t[61427] = 33
      "0100001" when "01110111111110100", -- t[61428] = 33
      "0100001" when "01110111111110101", -- t[61429] = 33
      "0100001" when "01110111111110110", -- t[61430] = 33
      "0100001" when "01110111111110111", -- t[61431] = 33
      "0100001" when "01110111111111000", -- t[61432] = 33
      "0100001" when "01110111111111001", -- t[61433] = 33
      "0100001" when "01110111111111010", -- t[61434] = 33
      "0100001" when "01110111111111011", -- t[61435] = 33
      "0100001" when "01110111111111100", -- t[61436] = 33
      "0100001" when "01110111111111101", -- t[61437] = 33
      "0100001" when "01110111111111110", -- t[61438] = 33
      "0100001" when "01110111111111111", -- t[61439] = 33
      "0100001" when "01111000000000000", -- t[61440] = 33
      "0100001" when "01111000000000001", -- t[61441] = 33
      "0100001" when "01111000000000010", -- t[61442] = 33
      "0100001" when "01111000000000011", -- t[61443] = 33
      "0100001" when "01111000000000100", -- t[61444] = 33
      "0100001" when "01111000000000101", -- t[61445] = 33
      "0100001" when "01111000000000110", -- t[61446] = 33
      "0100001" when "01111000000000111", -- t[61447] = 33
      "0100001" when "01111000000001000", -- t[61448] = 33
      "0100001" when "01111000000001001", -- t[61449] = 33
      "0100001" when "01111000000001010", -- t[61450] = 33
      "0100001" when "01111000000001011", -- t[61451] = 33
      "0100001" when "01111000000001100", -- t[61452] = 33
      "0100001" when "01111000000001101", -- t[61453] = 33
      "0100001" when "01111000000001110", -- t[61454] = 33
      "0100001" when "01111000000001111", -- t[61455] = 33
      "0100001" when "01111000000010000", -- t[61456] = 33
      "0100001" when "01111000000010001", -- t[61457] = 33
      "0100001" when "01111000000010010", -- t[61458] = 33
      "0100001" when "01111000000010011", -- t[61459] = 33
      "0100001" when "01111000000010100", -- t[61460] = 33
      "0100001" when "01111000000010101", -- t[61461] = 33
      "0100001" when "01111000000010110", -- t[61462] = 33
      "0100001" when "01111000000010111", -- t[61463] = 33
      "0100001" when "01111000000011000", -- t[61464] = 33
      "0100001" when "01111000000011001", -- t[61465] = 33
      "0100001" when "01111000000011010", -- t[61466] = 33
      "0100001" when "01111000000011011", -- t[61467] = 33
      "0100001" when "01111000000011100", -- t[61468] = 33
      "0100001" when "01111000000011101", -- t[61469] = 33
      "0100001" when "01111000000011110", -- t[61470] = 33
      "0100001" when "01111000000011111", -- t[61471] = 33
      "0100001" when "01111000000100000", -- t[61472] = 33
      "0100001" when "01111000000100001", -- t[61473] = 33
      "0100001" when "01111000000100010", -- t[61474] = 33
      "0100001" when "01111000000100011", -- t[61475] = 33
      "0100001" when "01111000000100100", -- t[61476] = 33
      "0100001" when "01111000000100101", -- t[61477] = 33
      "0100001" when "01111000000100110", -- t[61478] = 33
      "0100001" when "01111000000100111", -- t[61479] = 33
      "0100001" when "01111000000101000", -- t[61480] = 33
      "0100001" when "01111000000101001", -- t[61481] = 33
      "0100001" when "01111000000101010", -- t[61482] = 33
      "0100001" when "01111000000101011", -- t[61483] = 33
      "0100001" when "01111000000101100", -- t[61484] = 33
      "0100001" when "01111000000101101", -- t[61485] = 33
      "0100001" when "01111000000101110", -- t[61486] = 33
      "0100001" when "01111000000101111", -- t[61487] = 33
      "0100001" when "01111000000110000", -- t[61488] = 33
      "0100001" when "01111000000110001", -- t[61489] = 33
      "0100001" when "01111000000110010", -- t[61490] = 33
      "0100001" when "01111000000110011", -- t[61491] = 33
      "0100001" when "01111000000110100", -- t[61492] = 33
      "0100001" when "01111000000110101", -- t[61493] = 33
      "0100001" when "01111000000110110", -- t[61494] = 33
      "0100001" when "01111000000110111", -- t[61495] = 33
      "0100001" when "01111000000111000", -- t[61496] = 33
      "0100001" when "01111000000111001", -- t[61497] = 33
      "0100001" when "01111000000111010", -- t[61498] = 33
      "0100001" when "01111000000111011", -- t[61499] = 33
      "0100001" when "01111000000111100", -- t[61500] = 33
      "0100001" when "01111000000111101", -- t[61501] = 33
      "0100001" when "01111000000111110", -- t[61502] = 33
      "0100001" when "01111000000111111", -- t[61503] = 33
      "0100001" when "01111000001000000", -- t[61504] = 33
      "0100001" when "01111000001000001", -- t[61505] = 33
      "0100001" when "01111000001000010", -- t[61506] = 33
      "0100001" when "01111000001000011", -- t[61507] = 33
      "0100001" when "01111000001000100", -- t[61508] = 33
      "0100001" when "01111000001000101", -- t[61509] = 33
      "0100001" when "01111000001000110", -- t[61510] = 33
      "0100001" when "01111000001000111", -- t[61511] = 33
      "0100001" when "01111000001001000", -- t[61512] = 33
      "0100001" when "01111000001001001", -- t[61513] = 33
      "0100001" when "01111000001001010", -- t[61514] = 33
      "0100001" when "01111000001001011", -- t[61515] = 33
      "0100001" when "01111000001001100", -- t[61516] = 33
      "0100001" when "01111000001001101", -- t[61517] = 33
      "0100001" when "01111000001001110", -- t[61518] = 33
      "0100001" when "01111000001001111", -- t[61519] = 33
      "0100001" when "01111000001010000", -- t[61520] = 33
      "0100001" when "01111000001010001", -- t[61521] = 33
      "0100001" when "01111000001010010", -- t[61522] = 33
      "0100001" when "01111000001010011", -- t[61523] = 33
      "0100001" when "01111000001010100", -- t[61524] = 33
      "0100001" when "01111000001010101", -- t[61525] = 33
      "0100001" when "01111000001010110", -- t[61526] = 33
      "0100001" when "01111000001010111", -- t[61527] = 33
      "0100001" when "01111000001011000", -- t[61528] = 33
      "0100001" when "01111000001011001", -- t[61529] = 33
      "0100001" when "01111000001011010", -- t[61530] = 33
      "0100001" when "01111000001011011", -- t[61531] = 33
      "0100001" when "01111000001011100", -- t[61532] = 33
      "0100001" when "01111000001011101", -- t[61533] = 33
      "0100001" when "01111000001011110", -- t[61534] = 33
      "0100001" when "01111000001011111", -- t[61535] = 33
      "0100001" when "01111000001100000", -- t[61536] = 33
      "0100001" when "01111000001100001", -- t[61537] = 33
      "0100001" when "01111000001100010", -- t[61538] = 33
      "0100001" when "01111000001100011", -- t[61539] = 33
      "0100001" when "01111000001100100", -- t[61540] = 33
      "0100001" when "01111000001100101", -- t[61541] = 33
      "0100001" when "01111000001100110", -- t[61542] = 33
      "0100001" when "01111000001100111", -- t[61543] = 33
      "0100001" when "01111000001101000", -- t[61544] = 33
      "0100001" when "01111000001101001", -- t[61545] = 33
      "0100001" when "01111000001101010", -- t[61546] = 33
      "0100001" when "01111000001101011", -- t[61547] = 33
      "0100001" when "01111000001101100", -- t[61548] = 33
      "0100001" when "01111000001101101", -- t[61549] = 33
      "0100001" when "01111000001101110", -- t[61550] = 33
      "0100001" when "01111000001101111", -- t[61551] = 33
      "0100001" when "01111000001110000", -- t[61552] = 33
      "0100001" when "01111000001110001", -- t[61553] = 33
      "0100001" when "01111000001110010", -- t[61554] = 33
      "0100001" when "01111000001110011", -- t[61555] = 33
      "0100001" when "01111000001110100", -- t[61556] = 33
      "0100001" when "01111000001110101", -- t[61557] = 33
      "0100001" when "01111000001110110", -- t[61558] = 33
      "0100001" when "01111000001110111", -- t[61559] = 33
      "0100001" when "01111000001111000", -- t[61560] = 33
      "0100001" when "01111000001111001", -- t[61561] = 33
      "0100001" when "01111000001111010", -- t[61562] = 33
      "0100001" when "01111000001111011", -- t[61563] = 33
      "0100001" when "01111000001111100", -- t[61564] = 33
      "0100001" when "01111000001111101", -- t[61565] = 33
      "0100001" when "01111000001111110", -- t[61566] = 33
      "0100001" when "01111000001111111", -- t[61567] = 33
      "0100001" when "01111000010000000", -- t[61568] = 33
      "0100001" when "01111000010000001", -- t[61569] = 33
      "0100001" when "01111000010000010", -- t[61570] = 33
      "0100001" when "01111000010000011", -- t[61571] = 33
      "0100001" when "01111000010000100", -- t[61572] = 33
      "0100001" when "01111000010000101", -- t[61573] = 33
      "0100001" when "01111000010000110", -- t[61574] = 33
      "0100001" when "01111000010000111", -- t[61575] = 33
      "0100001" when "01111000010001000", -- t[61576] = 33
      "0100001" when "01111000010001001", -- t[61577] = 33
      "0100001" when "01111000010001010", -- t[61578] = 33
      "0100001" when "01111000010001011", -- t[61579] = 33
      "0100001" when "01111000010001100", -- t[61580] = 33
      "0100001" when "01111000010001101", -- t[61581] = 33
      "0100001" when "01111000010001110", -- t[61582] = 33
      "0100001" when "01111000010001111", -- t[61583] = 33
      "0100001" when "01111000010010000", -- t[61584] = 33
      "0100001" when "01111000010010001", -- t[61585] = 33
      "0100001" when "01111000010010010", -- t[61586] = 33
      "0100001" when "01111000010010011", -- t[61587] = 33
      "0100001" when "01111000010010100", -- t[61588] = 33
      "0100001" when "01111000010010101", -- t[61589] = 33
      "0100001" when "01111000010010110", -- t[61590] = 33
      "0100001" when "01111000010010111", -- t[61591] = 33
      "0100001" when "01111000010011000", -- t[61592] = 33
      "0100001" when "01111000010011001", -- t[61593] = 33
      "0100001" when "01111000010011010", -- t[61594] = 33
      "0100001" when "01111000010011011", -- t[61595] = 33
      "0100001" when "01111000010011100", -- t[61596] = 33
      "0100001" when "01111000010011101", -- t[61597] = 33
      "0100001" when "01111000010011110", -- t[61598] = 33
      "0100001" when "01111000010011111", -- t[61599] = 33
      "0100001" when "01111000010100000", -- t[61600] = 33
      "0100001" when "01111000010100001", -- t[61601] = 33
      "0100001" when "01111000010100010", -- t[61602] = 33
      "0100001" when "01111000010100011", -- t[61603] = 33
      "0100001" when "01111000010100100", -- t[61604] = 33
      "0100001" when "01111000010100101", -- t[61605] = 33
      "0100001" when "01111000010100110", -- t[61606] = 33
      "0100001" when "01111000010100111", -- t[61607] = 33
      "0100001" when "01111000010101000", -- t[61608] = 33
      "0100001" when "01111000010101001", -- t[61609] = 33
      "0100001" when "01111000010101010", -- t[61610] = 33
      "0100001" when "01111000010101011", -- t[61611] = 33
      "0100001" when "01111000010101100", -- t[61612] = 33
      "0100001" when "01111000010101101", -- t[61613] = 33
      "0100001" when "01111000010101110", -- t[61614] = 33
      "0100001" when "01111000010101111", -- t[61615] = 33
      "0100001" when "01111000010110000", -- t[61616] = 33
      "0100001" when "01111000010110001", -- t[61617] = 33
      "0100001" when "01111000010110010", -- t[61618] = 33
      "0100001" when "01111000010110011", -- t[61619] = 33
      "0100001" when "01111000010110100", -- t[61620] = 33
      "0100001" when "01111000010110101", -- t[61621] = 33
      "0100001" when "01111000010110110", -- t[61622] = 33
      "0100001" when "01111000010110111", -- t[61623] = 33
      "0100001" when "01111000010111000", -- t[61624] = 33
      "0100001" when "01111000010111001", -- t[61625] = 33
      "0100001" when "01111000010111010", -- t[61626] = 33
      "0100001" when "01111000010111011", -- t[61627] = 33
      "0100001" when "01111000010111100", -- t[61628] = 33
      "0100001" when "01111000010111101", -- t[61629] = 33
      "0100001" when "01111000010111110", -- t[61630] = 33
      "0100001" when "01111000010111111", -- t[61631] = 33
      "0100001" when "01111000011000000", -- t[61632] = 33
      "0100001" when "01111000011000001", -- t[61633] = 33
      "0100001" when "01111000011000010", -- t[61634] = 33
      "0100001" when "01111000011000011", -- t[61635] = 33
      "0100001" when "01111000011000100", -- t[61636] = 33
      "0100001" when "01111000011000101", -- t[61637] = 33
      "0100001" when "01111000011000110", -- t[61638] = 33
      "0100001" when "01111000011000111", -- t[61639] = 33
      "0100001" when "01111000011001000", -- t[61640] = 33
      "0100001" when "01111000011001001", -- t[61641] = 33
      "0100001" when "01111000011001010", -- t[61642] = 33
      "0100001" when "01111000011001011", -- t[61643] = 33
      "0100001" when "01111000011001100", -- t[61644] = 33
      "0100001" when "01111000011001101", -- t[61645] = 33
      "0100001" when "01111000011001110", -- t[61646] = 33
      "0100001" when "01111000011001111", -- t[61647] = 33
      "0100001" when "01111000011010000", -- t[61648] = 33
      "0100001" when "01111000011010001", -- t[61649] = 33
      "0100001" when "01111000011010010", -- t[61650] = 33
      "0100001" when "01111000011010011", -- t[61651] = 33
      "0100001" when "01111000011010100", -- t[61652] = 33
      "0100001" when "01111000011010101", -- t[61653] = 33
      "0100001" when "01111000011010110", -- t[61654] = 33
      "0100001" when "01111000011010111", -- t[61655] = 33
      "0100001" when "01111000011011000", -- t[61656] = 33
      "0100001" when "01111000011011001", -- t[61657] = 33
      "0100001" when "01111000011011010", -- t[61658] = 33
      "0100001" when "01111000011011011", -- t[61659] = 33
      "0100001" when "01111000011011100", -- t[61660] = 33
      "0100001" when "01111000011011101", -- t[61661] = 33
      "0100001" when "01111000011011110", -- t[61662] = 33
      "0100001" when "01111000011011111", -- t[61663] = 33
      "0100001" when "01111000011100000", -- t[61664] = 33
      "0100001" when "01111000011100001", -- t[61665] = 33
      "0100001" when "01111000011100010", -- t[61666] = 33
      "0100001" when "01111000011100011", -- t[61667] = 33
      "0100001" when "01111000011100100", -- t[61668] = 33
      "0100001" when "01111000011100101", -- t[61669] = 33
      "0100001" when "01111000011100110", -- t[61670] = 33
      "0100001" when "01111000011100111", -- t[61671] = 33
      "0100001" when "01111000011101000", -- t[61672] = 33
      "0100001" when "01111000011101001", -- t[61673] = 33
      "0100001" when "01111000011101010", -- t[61674] = 33
      "0100001" when "01111000011101011", -- t[61675] = 33
      "0100001" when "01111000011101100", -- t[61676] = 33
      "0100001" when "01111000011101101", -- t[61677] = 33
      "0100001" when "01111000011101110", -- t[61678] = 33
      "0100001" when "01111000011101111", -- t[61679] = 33
      "0100001" when "01111000011110000", -- t[61680] = 33
      "0100001" when "01111000011110001", -- t[61681] = 33
      "0100001" when "01111000011110010", -- t[61682] = 33
      "0100001" when "01111000011110011", -- t[61683] = 33
      "0100001" when "01111000011110100", -- t[61684] = 33
      "0100001" when "01111000011110101", -- t[61685] = 33
      "0100001" when "01111000011110110", -- t[61686] = 33
      "0100001" when "01111000011110111", -- t[61687] = 33
      "0100001" when "01111000011111000", -- t[61688] = 33
      "0100001" when "01111000011111001", -- t[61689] = 33
      "0100001" when "01111000011111010", -- t[61690] = 33
      "0100001" when "01111000011111011", -- t[61691] = 33
      "0100001" when "01111000011111100", -- t[61692] = 33
      "0100001" when "01111000011111101", -- t[61693] = 33
      "0100001" when "01111000011111110", -- t[61694] = 33
      "0100001" when "01111000011111111", -- t[61695] = 33
      "0100001" when "01111000100000000", -- t[61696] = 33
      "0100001" when "01111000100000001", -- t[61697] = 33
      "0100001" when "01111000100000010", -- t[61698] = 33
      "0100001" when "01111000100000011", -- t[61699] = 33
      "0100001" when "01111000100000100", -- t[61700] = 33
      "0100001" when "01111000100000101", -- t[61701] = 33
      "0100001" when "01111000100000110", -- t[61702] = 33
      "0100001" when "01111000100000111", -- t[61703] = 33
      "0100001" when "01111000100001000", -- t[61704] = 33
      "0100001" when "01111000100001001", -- t[61705] = 33
      "0100001" when "01111000100001010", -- t[61706] = 33
      "0100001" when "01111000100001011", -- t[61707] = 33
      "0100001" when "01111000100001100", -- t[61708] = 33
      "0100001" when "01111000100001101", -- t[61709] = 33
      "0100001" when "01111000100001110", -- t[61710] = 33
      "0100001" when "01111000100001111", -- t[61711] = 33
      "0100001" when "01111000100010000", -- t[61712] = 33
      "0100001" when "01111000100010001", -- t[61713] = 33
      "0100001" when "01111000100010010", -- t[61714] = 33
      "0100001" when "01111000100010011", -- t[61715] = 33
      "0100001" when "01111000100010100", -- t[61716] = 33
      "0100001" when "01111000100010101", -- t[61717] = 33
      "0100001" when "01111000100010110", -- t[61718] = 33
      "0100001" when "01111000100010111", -- t[61719] = 33
      "0100001" when "01111000100011000", -- t[61720] = 33
      "0100001" when "01111000100011001", -- t[61721] = 33
      "0100001" when "01111000100011010", -- t[61722] = 33
      "0100001" when "01111000100011011", -- t[61723] = 33
      "0100001" when "01111000100011100", -- t[61724] = 33
      "0100001" when "01111000100011101", -- t[61725] = 33
      "0100001" when "01111000100011110", -- t[61726] = 33
      "0100001" when "01111000100011111", -- t[61727] = 33
      "0100001" when "01111000100100000", -- t[61728] = 33
      "0100001" when "01111000100100001", -- t[61729] = 33
      "0100010" when "01111000100100010", -- t[61730] = 34
      "0100010" when "01111000100100011", -- t[61731] = 34
      "0100010" when "01111000100100100", -- t[61732] = 34
      "0100010" when "01111000100100101", -- t[61733] = 34
      "0100010" when "01111000100100110", -- t[61734] = 34
      "0100010" when "01111000100100111", -- t[61735] = 34
      "0100010" when "01111000100101000", -- t[61736] = 34
      "0100010" when "01111000100101001", -- t[61737] = 34
      "0100010" when "01111000100101010", -- t[61738] = 34
      "0100010" when "01111000100101011", -- t[61739] = 34
      "0100010" when "01111000100101100", -- t[61740] = 34
      "0100010" when "01111000100101101", -- t[61741] = 34
      "0100010" when "01111000100101110", -- t[61742] = 34
      "0100010" when "01111000100101111", -- t[61743] = 34
      "0100010" when "01111000100110000", -- t[61744] = 34
      "0100010" when "01111000100110001", -- t[61745] = 34
      "0100010" when "01111000100110010", -- t[61746] = 34
      "0100010" when "01111000100110011", -- t[61747] = 34
      "0100010" when "01111000100110100", -- t[61748] = 34
      "0100010" when "01111000100110101", -- t[61749] = 34
      "0100010" when "01111000100110110", -- t[61750] = 34
      "0100010" when "01111000100110111", -- t[61751] = 34
      "0100010" when "01111000100111000", -- t[61752] = 34
      "0100010" when "01111000100111001", -- t[61753] = 34
      "0100010" when "01111000100111010", -- t[61754] = 34
      "0100010" when "01111000100111011", -- t[61755] = 34
      "0100010" when "01111000100111100", -- t[61756] = 34
      "0100010" when "01111000100111101", -- t[61757] = 34
      "0100010" when "01111000100111110", -- t[61758] = 34
      "0100010" when "01111000100111111", -- t[61759] = 34
      "0100010" when "01111000101000000", -- t[61760] = 34
      "0100010" when "01111000101000001", -- t[61761] = 34
      "0100010" when "01111000101000010", -- t[61762] = 34
      "0100010" when "01111000101000011", -- t[61763] = 34
      "0100010" when "01111000101000100", -- t[61764] = 34
      "0100010" when "01111000101000101", -- t[61765] = 34
      "0100010" when "01111000101000110", -- t[61766] = 34
      "0100010" when "01111000101000111", -- t[61767] = 34
      "0100010" when "01111000101001000", -- t[61768] = 34
      "0100010" when "01111000101001001", -- t[61769] = 34
      "0100010" when "01111000101001010", -- t[61770] = 34
      "0100010" when "01111000101001011", -- t[61771] = 34
      "0100010" when "01111000101001100", -- t[61772] = 34
      "0100010" when "01111000101001101", -- t[61773] = 34
      "0100010" when "01111000101001110", -- t[61774] = 34
      "0100010" when "01111000101001111", -- t[61775] = 34
      "0100010" when "01111000101010000", -- t[61776] = 34
      "0100010" when "01111000101010001", -- t[61777] = 34
      "0100010" when "01111000101010010", -- t[61778] = 34
      "0100010" when "01111000101010011", -- t[61779] = 34
      "0100010" when "01111000101010100", -- t[61780] = 34
      "0100010" when "01111000101010101", -- t[61781] = 34
      "0100010" when "01111000101010110", -- t[61782] = 34
      "0100010" when "01111000101010111", -- t[61783] = 34
      "0100010" when "01111000101011000", -- t[61784] = 34
      "0100010" when "01111000101011001", -- t[61785] = 34
      "0100010" when "01111000101011010", -- t[61786] = 34
      "0100010" when "01111000101011011", -- t[61787] = 34
      "0100010" when "01111000101011100", -- t[61788] = 34
      "0100010" when "01111000101011101", -- t[61789] = 34
      "0100010" when "01111000101011110", -- t[61790] = 34
      "0100010" when "01111000101011111", -- t[61791] = 34
      "0100010" when "01111000101100000", -- t[61792] = 34
      "0100010" when "01111000101100001", -- t[61793] = 34
      "0100010" when "01111000101100010", -- t[61794] = 34
      "0100010" when "01111000101100011", -- t[61795] = 34
      "0100010" when "01111000101100100", -- t[61796] = 34
      "0100010" when "01111000101100101", -- t[61797] = 34
      "0100010" when "01111000101100110", -- t[61798] = 34
      "0100010" when "01111000101100111", -- t[61799] = 34
      "0100010" when "01111000101101000", -- t[61800] = 34
      "0100010" when "01111000101101001", -- t[61801] = 34
      "0100010" when "01111000101101010", -- t[61802] = 34
      "0100010" when "01111000101101011", -- t[61803] = 34
      "0100010" when "01111000101101100", -- t[61804] = 34
      "0100010" when "01111000101101101", -- t[61805] = 34
      "0100010" when "01111000101101110", -- t[61806] = 34
      "0100010" when "01111000101101111", -- t[61807] = 34
      "0100010" when "01111000101110000", -- t[61808] = 34
      "0100010" when "01111000101110001", -- t[61809] = 34
      "0100010" when "01111000101110010", -- t[61810] = 34
      "0100010" when "01111000101110011", -- t[61811] = 34
      "0100010" when "01111000101110100", -- t[61812] = 34
      "0100010" when "01111000101110101", -- t[61813] = 34
      "0100010" when "01111000101110110", -- t[61814] = 34
      "0100010" when "01111000101110111", -- t[61815] = 34
      "0100010" when "01111000101111000", -- t[61816] = 34
      "0100010" when "01111000101111001", -- t[61817] = 34
      "0100010" when "01111000101111010", -- t[61818] = 34
      "0100010" when "01111000101111011", -- t[61819] = 34
      "0100010" when "01111000101111100", -- t[61820] = 34
      "0100010" when "01111000101111101", -- t[61821] = 34
      "0100010" when "01111000101111110", -- t[61822] = 34
      "0100010" when "01111000101111111", -- t[61823] = 34
      "0100010" when "01111000110000000", -- t[61824] = 34
      "0100010" when "01111000110000001", -- t[61825] = 34
      "0100010" when "01111000110000010", -- t[61826] = 34
      "0100010" when "01111000110000011", -- t[61827] = 34
      "0100010" when "01111000110000100", -- t[61828] = 34
      "0100010" when "01111000110000101", -- t[61829] = 34
      "0100010" when "01111000110000110", -- t[61830] = 34
      "0100010" when "01111000110000111", -- t[61831] = 34
      "0100010" when "01111000110001000", -- t[61832] = 34
      "0100010" when "01111000110001001", -- t[61833] = 34
      "0100010" when "01111000110001010", -- t[61834] = 34
      "0100010" when "01111000110001011", -- t[61835] = 34
      "0100010" when "01111000110001100", -- t[61836] = 34
      "0100010" when "01111000110001101", -- t[61837] = 34
      "0100010" when "01111000110001110", -- t[61838] = 34
      "0100010" when "01111000110001111", -- t[61839] = 34
      "0100010" when "01111000110010000", -- t[61840] = 34
      "0100010" when "01111000110010001", -- t[61841] = 34
      "0100010" when "01111000110010010", -- t[61842] = 34
      "0100010" when "01111000110010011", -- t[61843] = 34
      "0100010" when "01111000110010100", -- t[61844] = 34
      "0100010" when "01111000110010101", -- t[61845] = 34
      "0100010" when "01111000110010110", -- t[61846] = 34
      "0100010" when "01111000110010111", -- t[61847] = 34
      "0100010" when "01111000110011000", -- t[61848] = 34
      "0100010" when "01111000110011001", -- t[61849] = 34
      "0100010" when "01111000110011010", -- t[61850] = 34
      "0100010" when "01111000110011011", -- t[61851] = 34
      "0100010" when "01111000110011100", -- t[61852] = 34
      "0100010" when "01111000110011101", -- t[61853] = 34
      "0100010" when "01111000110011110", -- t[61854] = 34
      "0100010" when "01111000110011111", -- t[61855] = 34
      "0100010" when "01111000110100000", -- t[61856] = 34
      "0100010" when "01111000110100001", -- t[61857] = 34
      "0100010" when "01111000110100010", -- t[61858] = 34
      "0100010" when "01111000110100011", -- t[61859] = 34
      "0100010" when "01111000110100100", -- t[61860] = 34
      "0100010" when "01111000110100101", -- t[61861] = 34
      "0100010" when "01111000110100110", -- t[61862] = 34
      "0100010" when "01111000110100111", -- t[61863] = 34
      "0100010" when "01111000110101000", -- t[61864] = 34
      "0100010" when "01111000110101001", -- t[61865] = 34
      "0100010" when "01111000110101010", -- t[61866] = 34
      "0100010" when "01111000110101011", -- t[61867] = 34
      "0100010" when "01111000110101100", -- t[61868] = 34
      "0100010" when "01111000110101101", -- t[61869] = 34
      "0100010" when "01111000110101110", -- t[61870] = 34
      "0100010" when "01111000110101111", -- t[61871] = 34
      "0100010" when "01111000110110000", -- t[61872] = 34
      "0100010" when "01111000110110001", -- t[61873] = 34
      "0100010" when "01111000110110010", -- t[61874] = 34
      "0100010" when "01111000110110011", -- t[61875] = 34
      "0100010" when "01111000110110100", -- t[61876] = 34
      "0100010" when "01111000110110101", -- t[61877] = 34
      "0100010" when "01111000110110110", -- t[61878] = 34
      "0100010" when "01111000110110111", -- t[61879] = 34
      "0100010" when "01111000110111000", -- t[61880] = 34
      "0100010" when "01111000110111001", -- t[61881] = 34
      "0100010" when "01111000110111010", -- t[61882] = 34
      "0100010" when "01111000110111011", -- t[61883] = 34
      "0100010" when "01111000110111100", -- t[61884] = 34
      "0100010" when "01111000110111101", -- t[61885] = 34
      "0100010" when "01111000110111110", -- t[61886] = 34
      "0100010" when "01111000110111111", -- t[61887] = 34
      "0100010" when "01111000111000000", -- t[61888] = 34
      "0100010" when "01111000111000001", -- t[61889] = 34
      "0100010" when "01111000111000010", -- t[61890] = 34
      "0100010" when "01111000111000011", -- t[61891] = 34
      "0100010" when "01111000111000100", -- t[61892] = 34
      "0100010" when "01111000111000101", -- t[61893] = 34
      "0100010" when "01111000111000110", -- t[61894] = 34
      "0100010" when "01111000111000111", -- t[61895] = 34
      "0100010" when "01111000111001000", -- t[61896] = 34
      "0100010" when "01111000111001001", -- t[61897] = 34
      "0100010" when "01111000111001010", -- t[61898] = 34
      "0100010" when "01111000111001011", -- t[61899] = 34
      "0100010" when "01111000111001100", -- t[61900] = 34
      "0100010" when "01111000111001101", -- t[61901] = 34
      "0100010" when "01111000111001110", -- t[61902] = 34
      "0100010" when "01111000111001111", -- t[61903] = 34
      "0100010" when "01111000111010000", -- t[61904] = 34
      "0100010" when "01111000111010001", -- t[61905] = 34
      "0100010" when "01111000111010010", -- t[61906] = 34
      "0100010" when "01111000111010011", -- t[61907] = 34
      "0100010" when "01111000111010100", -- t[61908] = 34
      "0100010" when "01111000111010101", -- t[61909] = 34
      "0100010" when "01111000111010110", -- t[61910] = 34
      "0100010" when "01111000111010111", -- t[61911] = 34
      "0100010" when "01111000111011000", -- t[61912] = 34
      "0100010" when "01111000111011001", -- t[61913] = 34
      "0100010" when "01111000111011010", -- t[61914] = 34
      "0100010" when "01111000111011011", -- t[61915] = 34
      "0100010" when "01111000111011100", -- t[61916] = 34
      "0100010" when "01111000111011101", -- t[61917] = 34
      "0100010" when "01111000111011110", -- t[61918] = 34
      "0100010" when "01111000111011111", -- t[61919] = 34
      "0100010" when "01111000111100000", -- t[61920] = 34
      "0100010" when "01111000111100001", -- t[61921] = 34
      "0100010" when "01111000111100010", -- t[61922] = 34
      "0100010" when "01111000111100011", -- t[61923] = 34
      "0100010" when "01111000111100100", -- t[61924] = 34
      "0100010" when "01111000111100101", -- t[61925] = 34
      "0100010" when "01111000111100110", -- t[61926] = 34
      "0100010" when "01111000111100111", -- t[61927] = 34
      "0100010" when "01111000111101000", -- t[61928] = 34
      "0100010" when "01111000111101001", -- t[61929] = 34
      "0100010" when "01111000111101010", -- t[61930] = 34
      "0100010" when "01111000111101011", -- t[61931] = 34
      "0100010" when "01111000111101100", -- t[61932] = 34
      "0100010" when "01111000111101101", -- t[61933] = 34
      "0100010" when "01111000111101110", -- t[61934] = 34
      "0100010" when "01111000111101111", -- t[61935] = 34
      "0100010" when "01111000111110000", -- t[61936] = 34
      "0100010" when "01111000111110001", -- t[61937] = 34
      "0100010" when "01111000111110010", -- t[61938] = 34
      "0100010" when "01111000111110011", -- t[61939] = 34
      "0100010" when "01111000111110100", -- t[61940] = 34
      "0100010" when "01111000111110101", -- t[61941] = 34
      "0100010" when "01111000111110110", -- t[61942] = 34
      "0100010" when "01111000111110111", -- t[61943] = 34
      "0100010" when "01111000111111000", -- t[61944] = 34
      "0100010" when "01111000111111001", -- t[61945] = 34
      "0100010" when "01111000111111010", -- t[61946] = 34
      "0100010" when "01111000111111011", -- t[61947] = 34
      "0100010" when "01111000111111100", -- t[61948] = 34
      "0100010" when "01111000111111101", -- t[61949] = 34
      "0100010" when "01111000111111110", -- t[61950] = 34
      "0100010" when "01111000111111111", -- t[61951] = 34
      "0100010" when "01111001000000000", -- t[61952] = 34
      "0100010" when "01111001000000001", -- t[61953] = 34
      "0100010" when "01111001000000010", -- t[61954] = 34
      "0100010" when "01111001000000011", -- t[61955] = 34
      "0100010" when "01111001000000100", -- t[61956] = 34
      "0100010" when "01111001000000101", -- t[61957] = 34
      "0100010" when "01111001000000110", -- t[61958] = 34
      "0100010" when "01111001000000111", -- t[61959] = 34
      "0100010" when "01111001000001000", -- t[61960] = 34
      "0100010" when "01111001000001001", -- t[61961] = 34
      "0100010" when "01111001000001010", -- t[61962] = 34
      "0100010" when "01111001000001011", -- t[61963] = 34
      "0100010" when "01111001000001100", -- t[61964] = 34
      "0100010" when "01111001000001101", -- t[61965] = 34
      "0100010" when "01111001000001110", -- t[61966] = 34
      "0100010" when "01111001000001111", -- t[61967] = 34
      "0100010" when "01111001000010000", -- t[61968] = 34
      "0100010" when "01111001000010001", -- t[61969] = 34
      "0100010" when "01111001000010010", -- t[61970] = 34
      "0100010" when "01111001000010011", -- t[61971] = 34
      "0100010" when "01111001000010100", -- t[61972] = 34
      "0100010" when "01111001000010101", -- t[61973] = 34
      "0100010" when "01111001000010110", -- t[61974] = 34
      "0100010" when "01111001000010111", -- t[61975] = 34
      "0100010" when "01111001000011000", -- t[61976] = 34
      "0100010" when "01111001000011001", -- t[61977] = 34
      "0100010" when "01111001000011010", -- t[61978] = 34
      "0100010" when "01111001000011011", -- t[61979] = 34
      "0100010" when "01111001000011100", -- t[61980] = 34
      "0100010" when "01111001000011101", -- t[61981] = 34
      "0100010" when "01111001000011110", -- t[61982] = 34
      "0100010" when "01111001000011111", -- t[61983] = 34
      "0100010" when "01111001000100000", -- t[61984] = 34
      "0100010" when "01111001000100001", -- t[61985] = 34
      "0100010" when "01111001000100010", -- t[61986] = 34
      "0100010" when "01111001000100011", -- t[61987] = 34
      "0100010" when "01111001000100100", -- t[61988] = 34
      "0100010" when "01111001000100101", -- t[61989] = 34
      "0100010" when "01111001000100110", -- t[61990] = 34
      "0100010" when "01111001000100111", -- t[61991] = 34
      "0100010" when "01111001000101000", -- t[61992] = 34
      "0100010" when "01111001000101001", -- t[61993] = 34
      "0100010" when "01111001000101010", -- t[61994] = 34
      "0100010" when "01111001000101011", -- t[61995] = 34
      "0100010" when "01111001000101100", -- t[61996] = 34
      "0100010" when "01111001000101101", -- t[61997] = 34
      "0100010" when "01111001000101110", -- t[61998] = 34
      "0100010" when "01111001000101111", -- t[61999] = 34
      "0100010" when "01111001000110000", -- t[62000] = 34
      "0100010" when "01111001000110001", -- t[62001] = 34
      "0100010" when "01111001000110010", -- t[62002] = 34
      "0100010" when "01111001000110011", -- t[62003] = 34
      "0100010" when "01111001000110100", -- t[62004] = 34
      "0100010" when "01111001000110101", -- t[62005] = 34
      "0100010" when "01111001000110110", -- t[62006] = 34
      "0100010" when "01111001000110111", -- t[62007] = 34
      "0100010" when "01111001000111000", -- t[62008] = 34
      "0100010" when "01111001000111001", -- t[62009] = 34
      "0100010" when "01111001000111010", -- t[62010] = 34
      "0100010" when "01111001000111011", -- t[62011] = 34
      "0100010" when "01111001000111100", -- t[62012] = 34
      "0100010" when "01111001000111101", -- t[62013] = 34
      "0100010" when "01111001000111110", -- t[62014] = 34
      "0100010" when "01111001000111111", -- t[62015] = 34
      "0100010" when "01111001001000000", -- t[62016] = 34
      "0100010" when "01111001001000001", -- t[62017] = 34
      "0100010" when "01111001001000010", -- t[62018] = 34
      "0100010" when "01111001001000011", -- t[62019] = 34
      "0100010" when "01111001001000100", -- t[62020] = 34
      "0100010" when "01111001001000101", -- t[62021] = 34
      "0100010" when "01111001001000110", -- t[62022] = 34
      "0100010" when "01111001001000111", -- t[62023] = 34
      "0100010" when "01111001001001000", -- t[62024] = 34
      "0100010" when "01111001001001001", -- t[62025] = 34
      "0100010" when "01111001001001010", -- t[62026] = 34
      "0100010" when "01111001001001011", -- t[62027] = 34
      "0100010" when "01111001001001100", -- t[62028] = 34
      "0100010" when "01111001001001101", -- t[62029] = 34
      "0100010" when "01111001001001110", -- t[62030] = 34
      "0100010" when "01111001001001111", -- t[62031] = 34
      "0100010" when "01111001001010000", -- t[62032] = 34
      "0100010" when "01111001001010001", -- t[62033] = 34
      "0100010" when "01111001001010010", -- t[62034] = 34
      "0100010" when "01111001001010011", -- t[62035] = 34
      "0100010" when "01111001001010100", -- t[62036] = 34
      "0100010" when "01111001001010101", -- t[62037] = 34
      "0100010" when "01111001001010110", -- t[62038] = 34
      "0100010" when "01111001001010111", -- t[62039] = 34
      "0100010" when "01111001001011000", -- t[62040] = 34
      "0100010" when "01111001001011001", -- t[62041] = 34
      "0100010" when "01111001001011010", -- t[62042] = 34
      "0100010" when "01111001001011011", -- t[62043] = 34
      "0100010" when "01111001001011100", -- t[62044] = 34
      "0100010" when "01111001001011101", -- t[62045] = 34
      "0100010" when "01111001001011110", -- t[62046] = 34
      "0100010" when "01111001001011111", -- t[62047] = 34
      "0100010" when "01111001001100000", -- t[62048] = 34
      "0100010" when "01111001001100001", -- t[62049] = 34
      "0100010" when "01111001001100010", -- t[62050] = 34
      "0100010" when "01111001001100011", -- t[62051] = 34
      "0100010" when "01111001001100100", -- t[62052] = 34
      "0100010" when "01111001001100101", -- t[62053] = 34
      "0100010" when "01111001001100110", -- t[62054] = 34
      "0100010" when "01111001001100111", -- t[62055] = 34
      "0100010" when "01111001001101000", -- t[62056] = 34
      "0100010" when "01111001001101001", -- t[62057] = 34
      "0100010" when "01111001001101010", -- t[62058] = 34
      "0100010" when "01111001001101011", -- t[62059] = 34
      "0100010" when "01111001001101100", -- t[62060] = 34
      "0100010" when "01111001001101101", -- t[62061] = 34
      "0100010" when "01111001001101110", -- t[62062] = 34
      "0100010" when "01111001001101111", -- t[62063] = 34
      "0100010" when "01111001001110000", -- t[62064] = 34
      "0100010" when "01111001001110001", -- t[62065] = 34
      "0100010" when "01111001001110010", -- t[62066] = 34
      "0100010" when "01111001001110011", -- t[62067] = 34
      "0100010" when "01111001001110100", -- t[62068] = 34
      "0100010" when "01111001001110101", -- t[62069] = 34
      "0100010" when "01111001001110110", -- t[62070] = 34
      "0100010" when "01111001001110111", -- t[62071] = 34
      "0100010" when "01111001001111000", -- t[62072] = 34
      "0100010" when "01111001001111001", -- t[62073] = 34
      "0100010" when "01111001001111010", -- t[62074] = 34
      "0100010" when "01111001001111011", -- t[62075] = 34
      "0100010" when "01111001001111100", -- t[62076] = 34
      "0100011" when "01111001001111101", -- t[62077] = 35
      "0100011" when "01111001001111110", -- t[62078] = 35
      "0100011" when "01111001001111111", -- t[62079] = 35
      "0100011" when "01111001010000000", -- t[62080] = 35
      "0100011" when "01111001010000001", -- t[62081] = 35
      "0100011" when "01111001010000010", -- t[62082] = 35
      "0100011" when "01111001010000011", -- t[62083] = 35
      "0100011" when "01111001010000100", -- t[62084] = 35
      "0100011" when "01111001010000101", -- t[62085] = 35
      "0100011" when "01111001010000110", -- t[62086] = 35
      "0100011" when "01111001010000111", -- t[62087] = 35
      "0100011" when "01111001010001000", -- t[62088] = 35
      "0100011" when "01111001010001001", -- t[62089] = 35
      "0100011" when "01111001010001010", -- t[62090] = 35
      "0100011" when "01111001010001011", -- t[62091] = 35
      "0100011" when "01111001010001100", -- t[62092] = 35
      "0100011" when "01111001010001101", -- t[62093] = 35
      "0100011" when "01111001010001110", -- t[62094] = 35
      "0100011" when "01111001010001111", -- t[62095] = 35
      "0100011" when "01111001010010000", -- t[62096] = 35
      "0100011" when "01111001010010001", -- t[62097] = 35
      "0100011" when "01111001010010010", -- t[62098] = 35
      "0100011" when "01111001010010011", -- t[62099] = 35
      "0100011" when "01111001010010100", -- t[62100] = 35
      "0100011" when "01111001010010101", -- t[62101] = 35
      "0100011" when "01111001010010110", -- t[62102] = 35
      "0100011" when "01111001010010111", -- t[62103] = 35
      "0100011" when "01111001010011000", -- t[62104] = 35
      "0100011" when "01111001010011001", -- t[62105] = 35
      "0100011" when "01111001010011010", -- t[62106] = 35
      "0100011" when "01111001010011011", -- t[62107] = 35
      "0100011" when "01111001010011100", -- t[62108] = 35
      "0100011" when "01111001010011101", -- t[62109] = 35
      "0100011" when "01111001010011110", -- t[62110] = 35
      "0100011" when "01111001010011111", -- t[62111] = 35
      "0100011" when "01111001010100000", -- t[62112] = 35
      "0100011" when "01111001010100001", -- t[62113] = 35
      "0100011" when "01111001010100010", -- t[62114] = 35
      "0100011" when "01111001010100011", -- t[62115] = 35
      "0100011" when "01111001010100100", -- t[62116] = 35
      "0100011" when "01111001010100101", -- t[62117] = 35
      "0100011" when "01111001010100110", -- t[62118] = 35
      "0100011" when "01111001010100111", -- t[62119] = 35
      "0100011" when "01111001010101000", -- t[62120] = 35
      "0100011" when "01111001010101001", -- t[62121] = 35
      "0100011" when "01111001010101010", -- t[62122] = 35
      "0100011" when "01111001010101011", -- t[62123] = 35
      "0100011" when "01111001010101100", -- t[62124] = 35
      "0100011" when "01111001010101101", -- t[62125] = 35
      "0100011" when "01111001010101110", -- t[62126] = 35
      "0100011" when "01111001010101111", -- t[62127] = 35
      "0100011" when "01111001010110000", -- t[62128] = 35
      "0100011" when "01111001010110001", -- t[62129] = 35
      "0100011" when "01111001010110010", -- t[62130] = 35
      "0100011" when "01111001010110011", -- t[62131] = 35
      "0100011" when "01111001010110100", -- t[62132] = 35
      "0100011" when "01111001010110101", -- t[62133] = 35
      "0100011" when "01111001010110110", -- t[62134] = 35
      "0100011" when "01111001010110111", -- t[62135] = 35
      "0100011" when "01111001010111000", -- t[62136] = 35
      "0100011" when "01111001010111001", -- t[62137] = 35
      "0100011" when "01111001010111010", -- t[62138] = 35
      "0100011" when "01111001010111011", -- t[62139] = 35
      "0100011" when "01111001010111100", -- t[62140] = 35
      "0100011" when "01111001010111101", -- t[62141] = 35
      "0100011" when "01111001010111110", -- t[62142] = 35
      "0100011" when "01111001010111111", -- t[62143] = 35
      "0100011" when "01111001011000000", -- t[62144] = 35
      "0100011" when "01111001011000001", -- t[62145] = 35
      "0100011" when "01111001011000010", -- t[62146] = 35
      "0100011" when "01111001011000011", -- t[62147] = 35
      "0100011" when "01111001011000100", -- t[62148] = 35
      "0100011" when "01111001011000101", -- t[62149] = 35
      "0100011" when "01111001011000110", -- t[62150] = 35
      "0100011" when "01111001011000111", -- t[62151] = 35
      "0100011" when "01111001011001000", -- t[62152] = 35
      "0100011" when "01111001011001001", -- t[62153] = 35
      "0100011" when "01111001011001010", -- t[62154] = 35
      "0100011" when "01111001011001011", -- t[62155] = 35
      "0100011" when "01111001011001100", -- t[62156] = 35
      "0100011" when "01111001011001101", -- t[62157] = 35
      "0100011" when "01111001011001110", -- t[62158] = 35
      "0100011" when "01111001011001111", -- t[62159] = 35
      "0100011" when "01111001011010000", -- t[62160] = 35
      "0100011" when "01111001011010001", -- t[62161] = 35
      "0100011" when "01111001011010010", -- t[62162] = 35
      "0100011" when "01111001011010011", -- t[62163] = 35
      "0100011" when "01111001011010100", -- t[62164] = 35
      "0100011" when "01111001011010101", -- t[62165] = 35
      "0100011" when "01111001011010110", -- t[62166] = 35
      "0100011" when "01111001011010111", -- t[62167] = 35
      "0100011" when "01111001011011000", -- t[62168] = 35
      "0100011" when "01111001011011001", -- t[62169] = 35
      "0100011" when "01111001011011010", -- t[62170] = 35
      "0100011" when "01111001011011011", -- t[62171] = 35
      "0100011" when "01111001011011100", -- t[62172] = 35
      "0100011" when "01111001011011101", -- t[62173] = 35
      "0100011" when "01111001011011110", -- t[62174] = 35
      "0100011" when "01111001011011111", -- t[62175] = 35
      "0100011" when "01111001011100000", -- t[62176] = 35
      "0100011" when "01111001011100001", -- t[62177] = 35
      "0100011" when "01111001011100010", -- t[62178] = 35
      "0100011" when "01111001011100011", -- t[62179] = 35
      "0100011" when "01111001011100100", -- t[62180] = 35
      "0100011" when "01111001011100101", -- t[62181] = 35
      "0100011" when "01111001011100110", -- t[62182] = 35
      "0100011" when "01111001011100111", -- t[62183] = 35
      "0100011" when "01111001011101000", -- t[62184] = 35
      "0100011" when "01111001011101001", -- t[62185] = 35
      "0100011" when "01111001011101010", -- t[62186] = 35
      "0100011" when "01111001011101011", -- t[62187] = 35
      "0100011" when "01111001011101100", -- t[62188] = 35
      "0100011" when "01111001011101101", -- t[62189] = 35
      "0100011" when "01111001011101110", -- t[62190] = 35
      "0100011" when "01111001011101111", -- t[62191] = 35
      "0100011" when "01111001011110000", -- t[62192] = 35
      "0100011" when "01111001011110001", -- t[62193] = 35
      "0100011" when "01111001011110010", -- t[62194] = 35
      "0100011" when "01111001011110011", -- t[62195] = 35
      "0100011" when "01111001011110100", -- t[62196] = 35
      "0100011" when "01111001011110101", -- t[62197] = 35
      "0100011" when "01111001011110110", -- t[62198] = 35
      "0100011" when "01111001011110111", -- t[62199] = 35
      "0100011" when "01111001011111000", -- t[62200] = 35
      "0100011" when "01111001011111001", -- t[62201] = 35
      "0100011" when "01111001011111010", -- t[62202] = 35
      "0100011" when "01111001011111011", -- t[62203] = 35
      "0100011" when "01111001011111100", -- t[62204] = 35
      "0100011" when "01111001011111101", -- t[62205] = 35
      "0100011" when "01111001011111110", -- t[62206] = 35
      "0100011" when "01111001011111111", -- t[62207] = 35
      "0100011" when "01111001100000000", -- t[62208] = 35
      "0100011" when "01111001100000001", -- t[62209] = 35
      "0100011" when "01111001100000010", -- t[62210] = 35
      "0100011" when "01111001100000011", -- t[62211] = 35
      "0100011" when "01111001100000100", -- t[62212] = 35
      "0100011" when "01111001100000101", -- t[62213] = 35
      "0100011" when "01111001100000110", -- t[62214] = 35
      "0100011" when "01111001100000111", -- t[62215] = 35
      "0100011" when "01111001100001000", -- t[62216] = 35
      "0100011" when "01111001100001001", -- t[62217] = 35
      "0100011" when "01111001100001010", -- t[62218] = 35
      "0100011" when "01111001100001011", -- t[62219] = 35
      "0100011" when "01111001100001100", -- t[62220] = 35
      "0100011" when "01111001100001101", -- t[62221] = 35
      "0100011" when "01111001100001110", -- t[62222] = 35
      "0100011" when "01111001100001111", -- t[62223] = 35
      "0100011" when "01111001100010000", -- t[62224] = 35
      "0100011" when "01111001100010001", -- t[62225] = 35
      "0100011" when "01111001100010010", -- t[62226] = 35
      "0100011" when "01111001100010011", -- t[62227] = 35
      "0100011" when "01111001100010100", -- t[62228] = 35
      "0100011" when "01111001100010101", -- t[62229] = 35
      "0100011" when "01111001100010110", -- t[62230] = 35
      "0100011" when "01111001100010111", -- t[62231] = 35
      "0100011" when "01111001100011000", -- t[62232] = 35
      "0100011" when "01111001100011001", -- t[62233] = 35
      "0100011" when "01111001100011010", -- t[62234] = 35
      "0100011" when "01111001100011011", -- t[62235] = 35
      "0100011" when "01111001100011100", -- t[62236] = 35
      "0100011" when "01111001100011101", -- t[62237] = 35
      "0100011" when "01111001100011110", -- t[62238] = 35
      "0100011" when "01111001100011111", -- t[62239] = 35
      "0100011" when "01111001100100000", -- t[62240] = 35
      "0100011" when "01111001100100001", -- t[62241] = 35
      "0100011" when "01111001100100010", -- t[62242] = 35
      "0100011" when "01111001100100011", -- t[62243] = 35
      "0100011" when "01111001100100100", -- t[62244] = 35
      "0100011" when "01111001100100101", -- t[62245] = 35
      "0100011" when "01111001100100110", -- t[62246] = 35
      "0100011" when "01111001100100111", -- t[62247] = 35
      "0100011" when "01111001100101000", -- t[62248] = 35
      "0100011" when "01111001100101001", -- t[62249] = 35
      "0100011" when "01111001100101010", -- t[62250] = 35
      "0100011" when "01111001100101011", -- t[62251] = 35
      "0100011" when "01111001100101100", -- t[62252] = 35
      "0100011" when "01111001100101101", -- t[62253] = 35
      "0100011" when "01111001100101110", -- t[62254] = 35
      "0100011" when "01111001100101111", -- t[62255] = 35
      "0100011" when "01111001100110000", -- t[62256] = 35
      "0100011" when "01111001100110001", -- t[62257] = 35
      "0100011" when "01111001100110010", -- t[62258] = 35
      "0100011" when "01111001100110011", -- t[62259] = 35
      "0100011" when "01111001100110100", -- t[62260] = 35
      "0100011" when "01111001100110101", -- t[62261] = 35
      "0100011" when "01111001100110110", -- t[62262] = 35
      "0100011" when "01111001100110111", -- t[62263] = 35
      "0100011" when "01111001100111000", -- t[62264] = 35
      "0100011" when "01111001100111001", -- t[62265] = 35
      "0100011" when "01111001100111010", -- t[62266] = 35
      "0100011" when "01111001100111011", -- t[62267] = 35
      "0100011" when "01111001100111100", -- t[62268] = 35
      "0100011" when "01111001100111101", -- t[62269] = 35
      "0100011" when "01111001100111110", -- t[62270] = 35
      "0100011" when "01111001100111111", -- t[62271] = 35
      "0100011" when "01111001101000000", -- t[62272] = 35
      "0100011" when "01111001101000001", -- t[62273] = 35
      "0100011" when "01111001101000010", -- t[62274] = 35
      "0100011" when "01111001101000011", -- t[62275] = 35
      "0100011" when "01111001101000100", -- t[62276] = 35
      "0100011" when "01111001101000101", -- t[62277] = 35
      "0100011" when "01111001101000110", -- t[62278] = 35
      "0100011" when "01111001101000111", -- t[62279] = 35
      "0100011" when "01111001101001000", -- t[62280] = 35
      "0100011" when "01111001101001001", -- t[62281] = 35
      "0100011" when "01111001101001010", -- t[62282] = 35
      "0100011" when "01111001101001011", -- t[62283] = 35
      "0100011" when "01111001101001100", -- t[62284] = 35
      "0100011" when "01111001101001101", -- t[62285] = 35
      "0100011" when "01111001101001110", -- t[62286] = 35
      "0100011" when "01111001101001111", -- t[62287] = 35
      "0100011" when "01111001101010000", -- t[62288] = 35
      "0100011" when "01111001101010001", -- t[62289] = 35
      "0100011" when "01111001101010010", -- t[62290] = 35
      "0100011" when "01111001101010011", -- t[62291] = 35
      "0100011" when "01111001101010100", -- t[62292] = 35
      "0100011" when "01111001101010101", -- t[62293] = 35
      "0100011" when "01111001101010110", -- t[62294] = 35
      "0100011" when "01111001101010111", -- t[62295] = 35
      "0100011" when "01111001101011000", -- t[62296] = 35
      "0100011" when "01111001101011001", -- t[62297] = 35
      "0100011" when "01111001101011010", -- t[62298] = 35
      "0100011" when "01111001101011011", -- t[62299] = 35
      "0100011" when "01111001101011100", -- t[62300] = 35
      "0100011" when "01111001101011101", -- t[62301] = 35
      "0100011" when "01111001101011110", -- t[62302] = 35
      "0100011" when "01111001101011111", -- t[62303] = 35
      "0100011" when "01111001101100000", -- t[62304] = 35
      "0100011" when "01111001101100001", -- t[62305] = 35
      "0100011" when "01111001101100010", -- t[62306] = 35
      "0100011" when "01111001101100011", -- t[62307] = 35
      "0100011" when "01111001101100100", -- t[62308] = 35
      "0100011" when "01111001101100101", -- t[62309] = 35
      "0100011" when "01111001101100110", -- t[62310] = 35
      "0100011" when "01111001101100111", -- t[62311] = 35
      "0100011" when "01111001101101000", -- t[62312] = 35
      "0100011" when "01111001101101001", -- t[62313] = 35
      "0100011" when "01111001101101010", -- t[62314] = 35
      "0100011" when "01111001101101011", -- t[62315] = 35
      "0100011" when "01111001101101100", -- t[62316] = 35
      "0100011" when "01111001101101101", -- t[62317] = 35
      "0100011" when "01111001101101110", -- t[62318] = 35
      "0100011" when "01111001101101111", -- t[62319] = 35
      "0100011" when "01111001101110000", -- t[62320] = 35
      "0100011" when "01111001101110001", -- t[62321] = 35
      "0100011" when "01111001101110010", -- t[62322] = 35
      "0100011" when "01111001101110011", -- t[62323] = 35
      "0100011" when "01111001101110100", -- t[62324] = 35
      "0100011" when "01111001101110101", -- t[62325] = 35
      "0100011" when "01111001101110110", -- t[62326] = 35
      "0100011" when "01111001101110111", -- t[62327] = 35
      "0100011" when "01111001101111000", -- t[62328] = 35
      "0100011" when "01111001101111001", -- t[62329] = 35
      "0100011" when "01111001101111010", -- t[62330] = 35
      "0100011" when "01111001101111011", -- t[62331] = 35
      "0100011" when "01111001101111100", -- t[62332] = 35
      "0100011" when "01111001101111101", -- t[62333] = 35
      "0100011" when "01111001101111110", -- t[62334] = 35
      "0100011" when "01111001101111111", -- t[62335] = 35
      "0100011" when "01111001110000000", -- t[62336] = 35
      "0100011" when "01111001110000001", -- t[62337] = 35
      "0100011" when "01111001110000010", -- t[62338] = 35
      "0100011" when "01111001110000011", -- t[62339] = 35
      "0100011" when "01111001110000100", -- t[62340] = 35
      "0100011" when "01111001110000101", -- t[62341] = 35
      "0100011" when "01111001110000110", -- t[62342] = 35
      "0100011" when "01111001110000111", -- t[62343] = 35
      "0100011" when "01111001110001000", -- t[62344] = 35
      "0100011" when "01111001110001001", -- t[62345] = 35
      "0100011" when "01111001110001010", -- t[62346] = 35
      "0100011" when "01111001110001011", -- t[62347] = 35
      "0100011" when "01111001110001100", -- t[62348] = 35
      "0100011" when "01111001110001101", -- t[62349] = 35
      "0100011" when "01111001110001110", -- t[62350] = 35
      "0100011" when "01111001110001111", -- t[62351] = 35
      "0100011" when "01111001110010000", -- t[62352] = 35
      "0100011" when "01111001110010001", -- t[62353] = 35
      "0100011" when "01111001110010010", -- t[62354] = 35
      "0100011" when "01111001110010011", -- t[62355] = 35
      "0100011" when "01111001110010100", -- t[62356] = 35
      "0100011" when "01111001110010101", -- t[62357] = 35
      "0100011" when "01111001110010110", -- t[62358] = 35
      "0100011" when "01111001110010111", -- t[62359] = 35
      "0100011" when "01111001110011000", -- t[62360] = 35
      "0100011" when "01111001110011001", -- t[62361] = 35
      "0100011" when "01111001110011010", -- t[62362] = 35
      "0100011" when "01111001110011011", -- t[62363] = 35
      "0100011" when "01111001110011100", -- t[62364] = 35
      "0100011" when "01111001110011101", -- t[62365] = 35
      "0100011" when "01111001110011110", -- t[62366] = 35
      "0100011" when "01111001110011111", -- t[62367] = 35
      "0100011" when "01111001110100000", -- t[62368] = 35
      "0100011" when "01111001110100001", -- t[62369] = 35
      "0100011" when "01111001110100010", -- t[62370] = 35
      "0100011" when "01111001110100011", -- t[62371] = 35
      "0100011" when "01111001110100100", -- t[62372] = 35
      "0100011" when "01111001110100101", -- t[62373] = 35
      "0100011" when "01111001110100110", -- t[62374] = 35
      "0100011" when "01111001110100111", -- t[62375] = 35
      "0100011" when "01111001110101000", -- t[62376] = 35
      "0100011" when "01111001110101001", -- t[62377] = 35
      "0100011" when "01111001110101010", -- t[62378] = 35
      "0100011" when "01111001110101011", -- t[62379] = 35
      "0100011" when "01111001110101100", -- t[62380] = 35
      "0100011" when "01111001110101101", -- t[62381] = 35
      "0100011" when "01111001110101110", -- t[62382] = 35
      "0100011" when "01111001110101111", -- t[62383] = 35
      "0100011" when "01111001110110000", -- t[62384] = 35
      "0100011" when "01111001110110001", -- t[62385] = 35
      "0100011" when "01111001110110010", -- t[62386] = 35
      "0100011" when "01111001110110011", -- t[62387] = 35
      "0100011" when "01111001110110100", -- t[62388] = 35
      "0100011" when "01111001110110101", -- t[62389] = 35
      "0100011" when "01111001110110110", -- t[62390] = 35
      "0100011" when "01111001110110111", -- t[62391] = 35
      "0100011" when "01111001110111000", -- t[62392] = 35
      "0100011" when "01111001110111001", -- t[62393] = 35
      "0100011" when "01111001110111010", -- t[62394] = 35
      "0100011" when "01111001110111011", -- t[62395] = 35
      "0100011" when "01111001110111100", -- t[62396] = 35
      "0100011" when "01111001110111101", -- t[62397] = 35
      "0100011" when "01111001110111110", -- t[62398] = 35
      "0100011" when "01111001110111111", -- t[62399] = 35
      "0100011" when "01111001111000000", -- t[62400] = 35
      "0100011" when "01111001111000001", -- t[62401] = 35
      "0100011" when "01111001111000010", -- t[62402] = 35
      "0100011" when "01111001111000011", -- t[62403] = 35
      "0100011" when "01111001111000100", -- t[62404] = 35
      "0100011" when "01111001111000101", -- t[62405] = 35
      "0100011" when "01111001111000110", -- t[62406] = 35
      "0100011" when "01111001111000111", -- t[62407] = 35
      "0100011" when "01111001111001000", -- t[62408] = 35
      "0100011" when "01111001111001001", -- t[62409] = 35
      "0100011" when "01111001111001010", -- t[62410] = 35
      "0100011" when "01111001111001011", -- t[62411] = 35
      "0100011" when "01111001111001100", -- t[62412] = 35
      "0100011" when "01111001111001101", -- t[62413] = 35
      "0100100" when "01111001111001110", -- t[62414] = 36
      "0100100" when "01111001111001111", -- t[62415] = 36
      "0100100" when "01111001111010000", -- t[62416] = 36
      "0100100" when "01111001111010001", -- t[62417] = 36
      "0100100" when "01111001111010010", -- t[62418] = 36
      "0100100" when "01111001111010011", -- t[62419] = 36
      "0100100" when "01111001111010100", -- t[62420] = 36
      "0100100" when "01111001111010101", -- t[62421] = 36
      "0100100" when "01111001111010110", -- t[62422] = 36
      "0100100" when "01111001111010111", -- t[62423] = 36
      "0100100" when "01111001111011000", -- t[62424] = 36
      "0100100" when "01111001111011001", -- t[62425] = 36
      "0100100" when "01111001111011010", -- t[62426] = 36
      "0100100" when "01111001111011011", -- t[62427] = 36
      "0100100" when "01111001111011100", -- t[62428] = 36
      "0100100" when "01111001111011101", -- t[62429] = 36
      "0100100" when "01111001111011110", -- t[62430] = 36
      "0100100" when "01111001111011111", -- t[62431] = 36
      "0100100" when "01111001111100000", -- t[62432] = 36
      "0100100" when "01111001111100001", -- t[62433] = 36
      "0100100" when "01111001111100010", -- t[62434] = 36
      "0100100" when "01111001111100011", -- t[62435] = 36
      "0100100" when "01111001111100100", -- t[62436] = 36
      "0100100" when "01111001111100101", -- t[62437] = 36
      "0100100" when "01111001111100110", -- t[62438] = 36
      "0100100" when "01111001111100111", -- t[62439] = 36
      "0100100" when "01111001111101000", -- t[62440] = 36
      "0100100" when "01111001111101001", -- t[62441] = 36
      "0100100" when "01111001111101010", -- t[62442] = 36
      "0100100" when "01111001111101011", -- t[62443] = 36
      "0100100" when "01111001111101100", -- t[62444] = 36
      "0100100" when "01111001111101101", -- t[62445] = 36
      "0100100" when "01111001111101110", -- t[62446] = 36
      "0100100" when "01111001111101111", -- t[62447] = 36
      "0100100" when "01111001111110000", -- t[62448] = 36
      "0100100" when "01111001111110001", -- t[62449] = 36
      "0100100" when "01111001111110010", -- t[62450] = 36
      "0100100" when "01111001111110011", -- t[62451] = 36
      "0100100" when "01111001111110100", -- t[62452] = 36
      "0100100" when "01111001111110101", -- t[62453] = 36
      "0100100" when "01111001111110110", -- t[62454] = 36
      "0100100" when "01111001111110111", -- t[62455] = 36
      "0100100" when "01111001111111000", -- t[62456] = 36
      "0100100" when "01111001111111001", -- t[62457] = 36
      "0100100" when "01111001111111010", -- t[62458] = 36
      "0100100" when "01111001111111011", -- t[62459] = 36
      "0100100" when "01111001111111100", -- t[62460] = 36
      "0100100" when "01111001111111101", -- t[62461] = 36
      "0100100" when "01111001111111110", -- t[62462] = 36
      "0100100" when "01111001111111111", -- t[62463] = 36
      "0100100" when "01111010000000000", -- t[62464] = 36
      "0100100" when "01111010000000001", -- t[62465] = 36
      "0100100" when "01111010000000010", -- t[62466] = 36
      "0100100" when "01111010000000011", -- t[62467] = 36
      "0100100" when "01111010000000100", -- t[62468] = 36
      "0100100" when "01111010000000101", -- t[62469] = 36
      "0100100" when "01111010000000110", -- t[62470] = 36
      "0100100" when "01111010000000111", -- t[62471] = 36
      "0100100" when "01111010000001000", -- t[62472] = 36
      "0100100" when "01111010000001001", -- t[62473] = 36
      "0100100" when "01111010000001010", -- t[62474] = 36
      "0100100" when "01111010000001011", -- t[62475] = 36
      "0100100" when "01111010000001100", -- t[62476] = 36
      "0100100" when "01111010000001101", -- t[62477] = 36
      "0100100" when "01111010000001110", -- t[62478] = 36
      "0100100" when "01111010000001111", -- t[62479] = 36
      "0100100" when "01111010000010000", -- t[62480] = 36
      "0100100" when "01111010000010001", -- t[62481] = 36
      "0100100" when "01111010000010010", -- t[62482] = 36
      "0100100" when "01111010000010011", -- t[62483] = 36
      "0100100" when "01111010000010100", -- t[62484] = 36
      "0100100" when "01111010000010101", -- t[62485] = 36
      "0100100" when "01111010000010110", -- t[62486] = 36
      "0100100" when "01111010000010111", -- t[62487] = 36
      "0100100" when "01111010000011000", -- t[62488] = 36
      "0100100" when "01111010000011001", -- t[62489] = 36
      "0100100" when "01111010000011010", -- t[62490] = 36
      "0100100" when "01111010000011011", -- t[62491] = 36
      "0100100" when "01111010000011100", -- t[62492] = 36
      "0100100" when "01111010000011101", -- t[62493] = 36
      "0100100" when "01111010000011110", -- t[62494] = 36
      "0100100" when "01111010000011111", -- t[62495] = 36
      "0100100" when "01111010000100000", -- t[62496] = 36
      "0100100" when "01111010000100001", -- t[62497] = 36
      "0100100" when "01111010000100010", -- t[62498] = 36
      "0100100" when "01111010000100011", -- t[62499] = 36
      "0100100" when "01111010000100100", -- t[62500] = 36
      "0100100" when "01111010000100101", -- t[62501] = 36
      "0100100" when "01111010000100110", -- t[62502] = 36
      "0100100" when "01111010000100111", -- t[62503] = 36
      "0100100" when "01111010000101000", -- t[62504] = 36
      "0100100" when "01111010000101001", -- t[62505] = 36
      "0100100" when "01111010000101010", -- t[62506] = 36
      "0100100" when "01111010000101011", -- t[62507] = 36
      "0100100" when "01111010000101100", -- t[62508] = 36
      "0100100" when "01111010000101101", -- t[62509] = 36
      "0100100" when "01111010000101110", -- t[62510] = 36
      "0100100" when "01111010000101111", -- t[62511] = 36
      "0100100" when "01111010000110000", -- t[62512] = 36
      "0100100" when "01111010000110001", -- t[62513] = 36
      "0100100" when "01111010000110010", -- t[62514] = 36
      "0100100" when "01111010000110011", -- t[62515] = 36
      "0100100" when "01111010000110100", -- t[62516] = 36
      "0100100" when "01111010000110101", -- t[62517] = 36
      "0100100" when "01111010000110110", -- t[62518] = 36
      "0100100" when "01111010000110111", -- t[62519] = 36
      "0100100" when "01111010000111000", -- t[62520] = 36
      "0100100" when "01111010000111001", -- t[62521] = 36
      "0100100" when "01111010000111010", -- t[62522] = 36
      "0100100" when "01111010000111011", -- t[62523] = 36
      "0100100" when "01111010000111100", -- t[62524] = 36
      "0100100" when "01111010000111101", -- t[62525] = 36
      "0100100" when "01111010000111110", -- t[62526] = 36
      "0100100" when "01111010000111111", -- t[62527] = 36
      "0100100" when "01111010001000000", -- t[62528] = 36
      "0100100" when "01111010001000001", -- t[62529] = 36
      "0100100" when "01111010001000010", -- t[62530] = 36
      "0100100" when "01111010001000011", -- t[62531] = 36
      "0100100" when "01111010001000100", -- t[62532] = 36
      "0100100" when "01111010001000101", -- t[62533] = 36
      "0100100" when "01111010001000110", -- t[62534] = 36
      "0100100" when "01111010001000111", -- t[62535] = 36
      "0100100" when "01111010001001000", -- t[62536] = 36
      "0100100" when "01111010001001001", -- t[62537] = 36
      "0100100" when "01111010001001010", -- t[62538] = 36
      "0100100" when "01111010001001011", -- t[62539] = 36
      "0100100" when "01111010001001100", -- t[62540] = 36
      "0100100" when "01111010001001101", -- t[62541] = 36
      "0100100" when "01111010001001110", -- t[62542] = 36
      "0100100" when "01111010001001111", -- t[62543] = 36
      "0100100" when "01111010001010000", -- t[62544] = 36
      "0100100" when "01111010001010001", -- t[62545] = 36
      "0100100" when "01111010001010010", -- t[62546] = 36
      "0100100" when "01111010001010011", -- t[62547] = 36
      "0100100" when "01111010001010100", -- t[62548] = 36
      "0100100" when "01111010001010101", -- t[62549] = 36
      "0100100" when "01111010001010110", -- t[62550] = 36
      "0100100" when "01111010001010111", -- t[62551] = 36
      "0100100" when "01111010001011000", -- t[62552] = 36
      "0100100" when "01111010001011001", -- t[62553] = 36
      "0100100" when "01111010001011010", -- t[62554] = 36
      "0100100" when "01111010001011011", -- t[62555] = 36
      "0100100" when "01111010001011100", -- t[62556] = 36
      "0100100" when "01111010001011101", -- t[62557] = 36
      "0100100" when "01111010001011110", -- t[62558] = 36
      "0100100" when "01111010001011111", -- t[62559] = 36
      "0100100" when "01111010001100000", -- t[62560] = 36
      "0100100" when "01111010001100001", -- t[62561] = 36
      "0100100" when "01111010001100010", -- t[62562] = 36
      "0100100" when "01111010001100011", -- t[62563] = 36
      "0100100" when "01111010001100100", -- t[62564] = 36
      "0100100" when "01111010001100101", -- t[62565] = 36
      "0100100" when "01111010001100110", -- t[62566] = 36
      "0100100" when "01111010001100111", -- t[62567] = 36
      "0100100" when "01111010001101000", -- t[62568] = 36
      "0100100" when "01111010001101001", -- t[62569] = 36
      "0100100" when "01111010001101010", -- t[62570] = 36
      "0100100" when "01111010001101011", -- t[62571] = 36
      "0100100" when "01111010001101100", -- t[62572] = 36
      "0100100" when "01111010001101101", -- t[62573] = 36
      "0100100" when "01111010001101110", -- t[62574] = 36
      "0100100" when "01111010001101111", -- t[62575] = 36
      "0100100" when "01111010001110000", -- t[62576] = 36
      "0100100" when "01111010001110001", -- t[62577] = 36
      "0100100" when "01111010001110010", -- t[62578] = 36
      "0100100" when "01111010001110011", -- t[62579] = 36
      "0100100" when "01111010001110100", -- t[62580] = 36
      "0100100" when "01111010001110101", -- t[62581] = 36
      "0100100" when "01111010001110110", -- t[62582] = 36
      "0100100" when "01111010001110111", -- t[62583] = 36
      "0100100" when "01111010001111000", -- t[62584] = 36
      "0100100" when "01111010001111001", -- t[62585] = 36
      "0100100" when "01111010001111010", -- t[62586] = 36
      "0100100" when "01111010001111011", -- t[62587] = 36
      "0100100" when "01111010001111100", -- t[62588] = 36
      "0100100" when "01111010001111101", -- t[62589] = 36
      "0100100" when "01111010001111110", -- t[62590] = 36
      "0100100" when "01111010001111111", -- t[62591] = 36
      "0100100" when "01111010010000000", -- t[62592] = 36
      "0100100" when "01111010010000001", -- t[62593] = 36
      "0100100" when "01111010010000010", -- t[62594] = 36
      "0100100" when "01111010010000011", -- t[62595] = 36
      "0100100" when "01111010010000100", -- t[62596] = 36
      "0100100" when "01111010010000101", -- t[62597] = 36
      "0100100" when "01111010010000110", -- t[62598] = 36
      "0100100" when "01111010010000111", -- t[62599] = 36
      "0100100" when "01111010010001000", -- t[62600] = 36
      "0100100" when "01111010010001001", -- t[62601] = 36
      "0100100" when "01111010010001010", -- t[62602] = 36
      "0100100" when "01111010010001011", -- t[62603] = 36
      "0100100" when "01111010010001100", -- t[62604] = 36
      "0100100" when "01111010010001101", -- t[62605] = 36
      "0100100" when "01111010010001110", -- t[62606] = 36
      "0100100" when "01111010010001111", -- t[62607] = 36
      "0100100" when "01111010010010000", -- t[62608] = 36
      "0100100" when "01111010010010001", -- t[62609] = 36
      "0100100" when "01111010010010010", -- t[62610] = 36
      "0100100" when "01111010010010011", -- t[62611] = 36
      "0100100" when "01111010010010100", -- t[62612] = 36
      "0100100" when "01111010010010101", -- t[62613] = 36
      "0100100" when "01111010010010110", -- t[62614] = 36
      "0100100" when "01111010010010111", -- t[62615] = 36
      "0100100" when "01111010010011000", -- t[62616] = 36
      "0100100" when "01111010010011001", -- t[62617] = 36
      "0100100" when "01111010010011010", -- t[62618] = 36
      "0100100" when "01111010010011011", -- t[62619] = 36
      "0100100" when "01111010010011100", -- t[62620] = 36
      "0100100" when "01111010010011101", -- t[62621] = 36
      "0100100" when "01111010010011110", -- t[62622] = 36
      "0100100" when "01111010010011111", -- t[62623] = 36
      "0100100" when "01111010010100000", -- t[62624] = 36
      "0100100" when "01111010010100001", -- t[62625] = 36
      "0100100" when "01111010010100010", -- t[62626] = 36
      "0100100" when "01111010010100011", -- t[62627] = 36
      "0100100" when "01111010010100100", -- t[62628] = 36
      "0100100" when "01111010010100101", -- t[62629] = 36
      "0100100" when "01111010010100110", -- t[62630] = 36
      "0100100" when "01111010010100111", -- t[62631] = 36
      "0100100" when "01111010010101000", -- t[62632] = 36
      "0100100" when "01111010010101001", -- t[62633] = 36
      "0100100" when "01111010010101010", -- t[62634] = 36
      "0100100" when "01111010010101011", -- t[62635] = 36
      "0100100" when "01111010010101100", -- t[62636] = 36
      "0100100" when "01111010010101101", -- t[62637] = 36
      "0100100" when "01111010010101110", -- t[62638] = 36
      "0100100" when "01111010010101111", -- t[62639] = 36
      "0100100" when "01111010010110000", -- t[62640] = 36
      "0100100" when "01111010010110001", -- t[62641] = 36
      "0100100" when "01111010010110010", -- t[62642] = 36
      "0100100" when "01111010010110011", -- t[62643] = 36
      "0100100" when "01111010010110100", -- t[62644] = 36
      "0100100" when "01111010010110101", -- t[62645] = 36
      "0100100" when "01111010010110110", -- t[62646] = 36
      "0100100" when "01111010010110111", -- t[62647] = 36
      "0100100" when "01111010010111000", -- t[62648] = 36
      "0100100" when "01111010010111001", -- t[62649] = 36
      "0100100" when "01111010010111010", -- t[62650] = 36
      "0100100" when "01111010010111011", -- t[62651] = 36
      "0100100" when "01111010010111100", -- t[62652] = 36
      "0100100" when "01111010010111101", -- t[62653] = 36
      "0100100" when "01111010010111110", -- t[62654] = 36
      "0100100" when "01111010010111111", -- t[62655] = 36
      "0100100" when "01111010011000000", -- t[62656] = 36
      "0100100" when "01111010011000001", -- t[62657] = 36
      "0100100" when "01111010011000010", -- t[62658] = 36
      "0100100" when "01111010011000011", -- t[62659] = 36
      "0100100" when "01111010011000100", -- t[62660] = 36
      "0100100" when "01111010011000101", -- t[62661] = 36
      "0100100" when "01111010011000110", -- t[62662] = 36
      "0100100" when "01111010011000111", -- t[62663] = 36
      "0100100" when "01111010011001000", -- t[62664] = 36
      "0100100" when "01111010011001001", -- t[62665] = 36
      "0100100" when "01111010011001010", -- t[62666] = 36
      "0100100" when "01111010011001011", -- t[62667] = 36
      "0100100" when "01111010011001100", -- t[62668] = 36
      "0100100" when "01111010011001101", -- t[62669] = 36
      "0100100" when "01111010011001110", -- t[62670] = 36
      "0100100" when "01111010011001111", -- t[62671] = 36
      "0100100" when "01111010011010000", -- t[62672] = 36
      "0100100" when "01111010011010001", -- t[62673] = 36
      "0100100" when "01111010011010010", -- t[62674] = 36
      "0100100" when "01111010011010011", -- t[62675] = 36
      "0100100" when "01111010011010100", -- t[62676] = 36
      "0100100" when "01111010011010101", -- t[62677] = 36
      "0100100" when "01111010011010110", -- t[62678] = 36
      "0100100" when "01111010011010111", -- t[62679] = 36
      "0100100" when "01111010011011000", -- t[62680] = 36
      "0100100" when "01111010011011001", -- t[62681] = 36
      "0100100" when "01111010011011010", -- t[62682] = 36
      "0100100" when "01111010011011011", -- t[62683] = 36
      "0100100" when "01111010011011100", -- t[62684] = 36
      "0100100" when "01111010011011101", -- t[62685] = 36
      "0100100" when "01111010011011110", -- t[62686] = 36
      "0100100" when "01111010011011111", -- t[62687] = 36
      "0100100" when "01111010011100000", -- t[62688] = 36
      "0100100" when "01111010011100001", -- t[62689] = 36
      "0100100" when "01111010011100010", -- t[62690] = 36
      "0100100" when "01111010011100011", -- t[62691] = 36
      "0100100" when "01111010011100100", -- t[62692] = 36
      "0100100" when "01111010011100101", -- t[62693] = 36
      "0100100" when "01111010011100110", -- t[62694] = 36
      "0100100" when "01111010011100111", -- t[62695] = 36
      "0100100" when "01111010011101000", -- t[62696] = 36
      "0100100" when "01111010011101001", -- t[62697] = 36
      "0100100" when "01111010011101010", -- t[62698] = 36
      "0100100" when "01111010011101011", -- t[62699] = 36
      "0100100" when "01111010011101100", -- t[62700] = 36
      "0100100" when "01111010011101101", -- t[62701] = 36
      "0100100" when "01111010011101110", -- t[62702] = 36
      "0100100" when "01111010011101111", -- t[62703] = 36
      "0100100" when "01111010011110000", -- t[62704] = 36
      "0100100" when "01111010011110001", -- t[62705] = 36
      "0100100" when "01111010011110010", -- t[62706] = 36
      "0100100" when "01111010011110011", -- t[62707] = 36
      "0100100" when "01111010011110100", -- t[62708] = 36
      "0100100" when "01111010011110101", -- t[62709] = 36
      "0100100" when "01111010011110110", -- t[62710] = 36
      "0100100" when "01111010011110111", -- t[62711] = 36
      "0100100" when "01111010011111000", -- t[62712] = 36
      "0100100" when "01111010011111001", -- t[62713] = 36
      "0100100" when "01111010011111010", -- t[62714] = 36
      "0100100" when "01111010011111011", -- t[62715] = 36
      "0100100" when "01111010011111100", -- t[62716] = 36
      "0100100" when "01111010011111101", -- t[62717] = 36
      "0100100" when "01111010011111110", -- t[62718] = 36
      "0100100" when "01111010011111111", -- t[62719] = 36
      "0100100" when "01111010100000000", -- t[62720] = 36
      "0100100" when "01111010100000001", -- t[62721] = 36
      "0100100" when "01111010100000010", -- t[62722] = 36
      "0100100" when "01111010100000011", -- t[62723] = 36
      "0100100" when "01111010100000100", -- t[62724] = 36
      "0100100" when "01111010100000101", -- t[62725] = 36
      "0100100" when "01111010100000110", -- t[62726] = 36
      "0100100" when "01111010100000111", -- t[62727] = 36
      "0100100" when "01111010100001000", -- t[62728] = 36
      "0100100" when "01111010100001001", -- t[62729] = 36
      "0100100" when "01111010100001010", -- t[62730] = 36
      "0100100" when "01111010100001011", -- t[62731] = 36
      "0100100" when "01111010100001100", -- t[62732] = 36
      "0100100" when "01111010100001101", -- t[62733] = 36
      "0100100" when "01111010100001110", -- t[62734] = 36
      "0100100" when "01111010100001111", -- t[62735] = 36
      "0100100" when "01111010100010000", -- t[62736] = 36
      "0100100" when "01111010100010001", -- t[62737] = 36
      "0100100" when "01111010100010010", -- t[62738] = 36
      "0100100" when "01111010100010011", -- t[62739] = 36
      "0100100" when "01111010100010100", -- t[62740] = 36
      "0100100" when "01111010100010101", -- t[62741] = 36
      "0100101" when "01111010100010110", -- t[62742] = 37
      "0100101" when "01111010100010111", -- t[62743] = 37
      "0100101" when "01111010100011000", -- t[62744] = 37
      "0100101" when "01111010100011001", -- t[62745] = 37
      "0100101" when "01111010100011010", -- t[62746] = 37
      "0100101" when "01111010100011011", -- t[62747] = 37
      "0100101" when "01111010100011100", -- t[62748] = 37
      "0100101" when "01111010100011101", -- t[62749] = 37
      "0100101" when "01111010100011110", -- t[62750] = 37
      "0100101" when "01111010100011111", -- t[62751] = 37
      "0100101" when "01111010100100000", -- t[62752] = 37
      "0100101" when "01111010100100001", -- t[62753] = 37
      "0100101" when "01111010100100010", -- t[62754] = 37
      "0100101" when "01111010100100011", -- t[62755] = 37
      "0100101" when "01111010100100100", -- t[62756] = 37
      "0100101" when "01111010100100101", -- t[62757] = 37
      "0100101" when "01111010100100110", -- t[62758] = 37
      "0100101" when "01111010100100111", -- t[62759] = 37
      "0100101" when "01111010100101000", -- t[62760] = 37
      "0100101" when "01111010100101001", -- t[62761] = 37
      "0100101" when "01111010100101010", -- t[62762] = 37
      "0100101" when "01111010100101011", -- t[62763] = 37
      "0100101" when "01111010100101100", -- t[62764] = 37
      "0100101" when "01111010100101101", -- t[62765] = 37
      "0100101" when "01111010100101110", -- t[62766] = 37
      "0100101" when "01111010100101111", -- t[62767] = 37
      "0100101" when "01111010100110000", -- t[62768] = 37
      "0100101" when "01111010100110001", -- t[62769] = 37
      "0100101" when "01111010100110010", -- t[62770] = 37
      "0100101" when "01111010100110011", -- t[62771] = 37
      "0100101" when "01111010100110100", -- t[62772] = 37
      "0100101" when "01111010100110101", -- t[62773] = 37
      "0100101" when "01111010100110110", -- t[62774] = 37
      "0100101" when "01111010100110111", -- t[62775] = 37
      "0100101" when "01111010100111000", -- t[62776] = 37
      "0100101" when "01111010100111001", -- t[62777] = 37
      "0100101" when "01111010100111010", -- t[62778] = 37
      "0100101" when "01111010100111011", -- t[62779] = 37
      "0100101" when "01111010100111100", -- t[62780] = 37
      "0100101" when "01111010100111101", -- t[62781] = 37
      "0100101" when "01111010100111110", -- t[62782] = 37
      "0100101" when "01111010100111111", -- t[62783] = 37
      "0100101" when "01111010101000000", -- t[62784] = 37
      "0100101" when "01111010101000001", -- t[62785] = 37
      "0100101" when "01111010101000010", -- t[62786] = 37
      "0100101" when "01111010101000011", -- t[62787] = 37
      "0100101" when "01111010101000100", -- t[62788] = 37
      "0100101" when "01111010101000101", -- t[62789] = 37
      "0100101" when "01111010101000110", -- t[62790] = 37
      "0100101" when "01111010101000111", -- t[62791] = 37
      "0100101" when "01111010101001000", -- t[62792] = 37
      "0100101" when "01111010101001001", -- t[62793] = 37
      "0100101" when "01111010101001010", -- t[62794] = 37
      "0100101" when "01111010101001011", -- t[62795] = 37
      "0100101" when "01111010101001100", -- t[62796] = 37
      "0100101" when "01111010101001101", -- t[62797] = 37
      "0100101" when "01111010101001110", -- t[62798] = 37
      "0100101" when "01111010101001111", -- t[62799] = 37
      "0100101" when "01111010101010000", -- t[62800] = 37
      "0100101" when "01111010101010001", -- t[62801] = 37
      "0100101" when "01111010101010010", -- t[62802] = 37
      "0100101" when "01111010101010011", -- t[62803] = 37
      "0100101" when "01111010101010100", -- t[62804] = 37
      "0100101" when "01111010101010101", -- t[62805] = 37
      "0100101" when "01111010101010110", -- t[62806] = 37
      "0100101" when "01111010101010111", -- t[62807] = 37
      "0100101" when "01111010101011000", -- t[62808] = 37
      "0100101" when "01111010101011001", -- t[62809] = 37
      "0100101" when "01111010101011010", -- t[62810] = 37
      "0100101" when "01111010101011011", -- t[62811] = 37
      "0100101" when "01111010101011100", -- t[62812] = 37
      "0100101" when "01111010101011101", -- t[62813] = 37
      "0100101" when "01111010101011110", -- t[62814] = 37
      "0100101" when "01111010101011111", -- t[62815] = 37
      "0100101" when "01111010101100000", -- t[62816] = 37
      "0100101" when "01111010101100001", -- t[62817] = 37
      "0100101" when "01111010101100010", -- t[62818] = 37
      "0100101" when "01111010101100011", -- t[62819] = 37
      "0100101" when "01111010101100100", -- t[62820] = 37
      "0100101" when "01111010101100101", -- t[62821] = 37
      "0100101" when "01111010101100110", -- t[62822] = 37
      "0100101" when "01111010101100111", -- t[62823] = 37
      "0100101" when "01111010101101000", -- t[62824] = 37
      "0100101" when "01111010101101001", -- t[62825] = 37
      "0100101" when "01111010101101010", -- t[62826] = 37
      "0100101" when "01111010101101011", -- t[62827] = 37
      "0100101" when "01111010101101100", -- t[62828] = 37
      "0100101" when "01111010101101101", -- t[62829] = 37
      "0100101" when "01111010101101110", -- t[62830] = 37
      "0100101" when "01111010101101111", -- t[62831] = 37
      "0100101" when "01111010101110000", -- t[62832] = 37
      "0100101" when "01111010101110001", -- t[62833] = 37
      "0100101" when "01111010101110010", -- t[62834] = 37
      "0100101" when "01111010101110011", -- t[62835] = 37
      "0100101" when "01111010101110100", -- t[62836] = 37
      "0100101" when "01111010101110101", -- t[62837] = 37
      "0100101" when "01111010101110110", -- t[62838] = 37
      "0100101" when "01111010101110111", -- t[62839] = 37
      "0100101" when "01111010101111000", -- t[62840] = 37
      "0100101" when "01111010101111001", -- t[62841] = 37
      "0100101" when "01111010101111010", -- t[62842] = 37
      "0100101" when "01111010101111011", -- t[62843] = 37
      "0100101" when "01111010101111100", -- t[62844] = 37
      "0100101" when "01111010101111101", -- t[62845] = 37
      "0100101" when "01111010101111110", -- t[62846] = 37
      "0100101" when "01111010101111111", -- t[62847] = 37
      "0100101" when "01111010110000000", -- t[62848] = 37
      "0100101" when "01111010110000001", -- t[62849] = 37
      "0100101" when "01111010110000010", -- t[62850] = 37
      "0100101" when "01111010110000011", -- t[62851] = 37
      "0100101" when "01111010110000100", -- t[62852] = 37
      "0100101" when "01111010110000101", -- t[62853] = 37
      "0100101" when "01111010110000110", -- t[62854] = 37
      "0100101" when "01111010110000111", -- t[62855] = 37
      "0100101" when "01111010110001000", -- t[62856] = 37
      "0100101" when "01111010110001001", -- t[62857] = 37
      "0100101" when "01111010110001010", -- t[62858] = 37
      "0100101" when "01111010110001011", -- t[62859] = 37
      "0100101" when "01111010110001100", -- t[62860] = 37
      "0100101" when "01111010110001101", -- t[62861] = 37
      "0100101" when "01111010110001110", -- t[62862] = 37
      "0100101" when "01111010110001111", -- t[62863] = 37
      "0100101" when "01111010110010000", -- t[62864] = 37
      "0100101" when "01111010110010001", -- t[62865] = 37
      "0100101" when "01111010110010010", -- t[62866] = 37
      "0100101" when "01111010110010011", -- t[62867] = 37
      "0100101" when "01111010110010100", -- t[62868] = 37
      "0100101" when "01111010110010101", -- t[62869] = 37
      "0100101" when "01111010110010110", -- t[62870] = 37
      "0100101" when "01111010110010111", -- t[62871] = 37
      "0100101" when "01111010110011000", -- t[62872] = 37
      "0100101" when "01111010110011001", -- t[62873] = 37
      "0100101" when "01111010110011010", -- t[62874] = 37
      "0100101" when "01111010110011011", -- t[62875] = 37
      "0100101" when "01111010110011100", -- t[62876] = 37
      "0100101" when "01111010110011101", -- t[62877] = 37
      "0100101" when "01111010110011110", -- t[62878] = 37
      "0100101" when "01111010110011111", -- t[62879] = 37
      "0100101" when "01111010110100000", -- t[62880] = 37
      "0100101" when "01111010110100001", -- t[62881] = 37
      "0100101" when "01111010110100010", -- t[62882] = 37
      "0100101" when "01111010110100011", -- t[62883] = 37
      "0100101" when "01111010110100100", -- t[62884] = 37
      "0100101" when "01111010110100101", -- t[62885] = 37
      "0100101" when "01111010110100110", -- t[62886] = 37
      "0100101" when "01111010110100111", -- t[62887] = 37
      "0100101" when "01111010110101000", -- t[62888] = 37
      "0100101" when "01111010110101001", -- t[62889] = 37
      "0100101" when "01111010110101010", -- t[62890] = 37
      "0100101" when "01111010110101011", -- t[62891] = 37
      "0100101" when "01111010110101100", -- t[62892] = 37
      "0100101" when "01111010110101101", -- t[62893] = 37
      "0100101" when "01111010110101110", -- t[62894] = 37
      "0100101" when "01111010110101111", -- t[62895] = 37
      "0100101" when "01111010110110000", -- t[62896] = 37
      "0100101" when "01111010110110001", -- t[62897] = 37
      "0100101" when "01111010110110010", -- t[62898] = 37
      "0100101" when "01111010110110011", -- t[62899] = 37
      "0100101" when "01111010110110100", -- t[62900] = 37
      "0100101" when "01111010110110101", -- t[62901] = 37
      "0100101" when "01111010110110110", -- t[62902] = 37
      "0100101" when "01111010110110111", -- t[62903] = 37
      "0100101" when "01111010110111000", -- t[62904] = 37
      "0100101" when "01111010110111001", -- t[62905] = 37
      "0100101" when "01111010110111010", -- t[62906] = 37
      "0100101" when "01111010110111011", -- t[62907] = 37
      "0100101" when "01111010110111100", -- t[62908] = 37
      "0100101" when "01111010110111101", -- t[62909] = 37
      "0100101" when "01111010110111110", -- t[62910] = 37
      "0100101" when "01111010110111111", -- t[62911] = 37
      "0100101" when "01111010111000000", -- t[62912] = 37
      "0100101" when "01111010111000001", -- t[62913] = 37
      "0100101" when "01111010111000010", -- t[62914] = 37
      "0100101" when "01111010111000011", -- t[62915] = 37
      "0100101" when "01111010111000100", -- t[62916] = 37
      "0100101" when "01111010111000101", -- t[62917] = 37
      "0100101" when "01111010111000110", -- t[62918] = 37
      "0100101" when "01111010111000111", -- t[62919] = 37
      "0100101" when "01111010111001000", -- t[62920] = 37
      "0100101" when "01111010111001001", -- t[62921] = 37
      "0100101" when "01111010111001010", -- t[62922] = 37
      "0100101" when "01111010111001011", -- t[62923] = 37
      "0100101" when "01111010111001100", -- t[62924] = 37
      "0100101" when "01111010111001101", -- t[62925] = 37
      "0100101" when "01111010111001110", -- t[62926] = 37
      "0100101" when "01111010111001111", -- t[62927] = 37
      "0100101" when "01111010111010000", -- t[62928] = 37
      "0100101" when "01111010111010001", -- t[62929] = 37
      "0100101" when "01111010111010010", -- t[62930] = 37
      "0100101" when "01111010111010011", -- t[62931] = 37
      "0100101" when "01111010111010100", -- t[62932] = 37
      "0100101" when "01111010111010101", -- t[62933] = 37
      "0100101" when "01111010111010110", -- t[62934] = 37
      "0100101" when "01111010111010111", -- t[62935] = 37
      "0100101" when "01111010111011000", -- t[62936] = 37
      "0100101" when "01111010111011001", -- t[62937] = 37
      "0100101" when "01111010111011010", -- t[62938] = 37
      "0100101" when "01111010111011011", -- t[62939] = 37
      "0100101" when "01111010111011100", -- t[62940] = 37
      "0100101" when "01111010111011101", -- t[62941] = 37
      "0100101" when "01111010111011110", -- t[62942] = 37
      "0100101" when "01111010111011111", -- t[62943] = 37
      "0100101" when "01111010111100000", -- t[62944] = 37
      "0100101" when "01111010111100001", -- t[62945] = 37
      "0100101" when "01111010111100010", -- t[62946] = 37
      "0100101" when "01111010111100011", -- t[62947] = 37
      "0100101" when "01111010111100100", -- t[62948] = 37
      "0100101" when "01111010111100101", -- t[62949] = 37
      "0100101" when "01111010111100110", -- t[62950] = 37
      "0100101" when "01111010111100111", -- t[62951] = 37
      "0100101" when "01111010111101000", -- t[62952] = 37
      "0100101" when "01111010111101001", -- t[62953] = 37
      "0100101" when "01111010111101010", -- t[62954] = 37
      "0100101" when "01111010111101011", -- t[62955] = 37
      "0100101" when "01111010111101100", -- t[62956] = 37
      "0100101" when "01111010111101101", -- t[62957] = 37
      "0100101" when "01111010111101110", -- t[62958] = 37
      "0100101" when "01111010111101111", -- t[62959] = 37
      "0100101" when "01111010111110000", -- t[62960] = 37
      "0100101" when "01111010111110001", -- t[62961] = 37
      "0100101" when "01111010111110010", -- t[62962] = 37
      "0100101" when "01111010111110011", -- t[62963] = 37
      "0100101" when "01111010111110100", -- t[62964] = 37
      "0100101" when "01111010111110101", -- t[62965] = 37
      "0100101" when "01111010111110110", -- t[62966] = 37
      "0100101" when "01111010111110111", -- t[62967] = 37
      "0100101" when "01111010111111000", -- t[62968] = 37
      "0100101" when "01111010111111001", -- t[62969] = 37
      "0100101" when "01111010111111010", -- t[62970] = 37
      "0100101" when "01111010111111011", -- t[62971] = 37
      "0100101" when "01111010111111100", -- t[62972] = 37
      "0100101" when "01111010111111101", -- t[62973] = 37
      "0100101" when "01111010111111110", -- t[62974] = 37
      "0100101" when "01111010111111111", -- t[62975] = 37
      "0100101" when "01111011000000000", -- t[62976] = 37
      "0100101" when "01111011000000001", -- t[62977] = 37
      "0100101" when "01111011000000010", -- t[62978] = 37
      "0100101" when "01111011000000011", -- t[62979] = 37
      "0100101" when "01111011000000100", -- t[62980] = 37
      "0100101" when "01111011000000101", -- t[62981] = 37
      "0100101" when "01111011000000110", -- t[62982] = 37
      "0100101" when "01111011000000111", -- t[62983] = 37
      "0100101" when "01111011000001000", -- t[62984] = 37
      "0100101" when "01111011000001001", -- t[62985] = 37
      "0100101" when "01111011000001010", -- t[62986] = 37
      "0100101" when "01111011000001011", -- t[62987] = 37
      "0100101" when "01111011000001100", -- t[62988] = 37
      "0100101" when "01111011000001101", -- t[62989] = 37
      "0100101" when "01111011000001110", -- t[62990] = 37
      "0100101" when "01111011000001111", -- t[62991] = 37
      "0100101" when "01111011000010000", -- t[62992] = 37
      "0100101" when "01111011000010001", -- t[62993] = 37
      "0100101" when "01111011000010010", -- t[62994] = 37
      "0100101" when "01111011000010011", -- t[62995] = 37
      "0100101" when "01111011000010100", -- t[62996] = 37
      "0100101" when "01111011000010101", -- t[62997] = 37
      "0100101" when "01111011000010110", -- t[62998] = 37
      "0100101" when "01111011000010111", -- t[62999] = 37
      "0100101" when "01111011000011000", -- t[63000] = 37
      "0100101" when "01111011000011001", -- t[63001] = 37
      "0100101" when "01111011000011010", -- t[63002] = 37
      "0100101" when "01111011000011011", -- t[63003] = 37
      "0100101" when "01111011000011100", -- t[63004] = 37
      "0100101" when "01111011000011101", -- t[63005] = 37
      "0100101" when "01111011000011110", -- t[63006] = 37
      "0100101" when "01111011000011111", -- t[63007] = 37
      "0100101" when "01111011000100000", -- t[63008] = 37
      "0100101" when "01111011000100001", -- t[63009] = 37
      "0100101" when "01111011000100010", -- t[63010] = 37
      "0100101" when "01111011000100011", -- t[63011] = 37
      "0100101" when "01111011000100100", -- t[63012] = 37
      "0100101" when "01111011000100101", -- t[63013] = 37
      "0100101" when "01111011000100110", -- t[63014] = 37
      "0100101" when "01111011000100111", -- t[63015] = 37
      "0100101" when "01111011000101000", -- t[63016] = 37
      "0100101" when "01111011000101001", -- t[63017] = 37
      "0100101" when "01111011000101010", -- t[63018] = 37
      "0100101" when "01111011000101011", -- t[63019] = 37
      "0100101" when "01111011000101100", -- t[63020] = 37
      "0100101" when "01111011000101101", -- t[63021] = 37
      "0100101" when "01111011000101110", -- t[63022] = 37
      "0100101" when "01111011000101111", -- t[63023] = 37
      "0100101" when "01111011000110000", -- t[63024] = 37
      "0100101" when "01111011000110001", -- t[63025] = 37
      "0100101" when "01111011000110010", -- t[63026] = 37
      "0100101" when "01111011000110011", -- t[63027] = 37
      "0100101" when "01111011000110100", -- t[63028] = 37
      "0100101" when "01111011000110101", -- t[63029] = 37
      "0100101" when "01111011000110110", -- t[63030] = 37
      "0100101" when "01111011000110111", -- t[63031] = 37
      "0100101" when "01111011000111000", -- t[63032] = 37
      "0100101" when "01111011000111001", -- t[63033] = 37
      "0100101" when "01111011000111010", -- t[63034] = 37
      "0100101" when "01111011000111011", -- t[63035] = 37
      "0100101" when "01111011000111100", -- t[63036] = 37
      "0100101" when "01111011000111101", -- t[63037] = 37
      "0100101" when "01111011000111110", -- t[63038] = 37
      "0100101" when "01111011000111111", -- t[63039] = 37
      "0100101" when "01111011001000000", -- t[63040] = 37
      "0100101" when "01111011001000001", -- t[63041] = 37
      "0100101" when "01111011001000010", -- t[63042] = 37
      "0100101" when "01111011001000011", -- t[63043] = 37
      "0100101" when "01111011001000100", -- t[63044] = 37
      "0100101" when "01111011001000101", -- t[63045] = 37
      "0100101" when "01111011001000110", -- t[63046] = 37
      "0100101" when "01111011001000111", -- t[63047] = 37
      "0100101" when "01111011001001000", -- t[63048] = 37
      "0100101" when "01111011001001001", -- t[63049] = 37
      "0100101" when "01111011001001010", -- t[63050] = 37
      "0100101" when "01111011001001011", -- t[63051] = 37
      "0100101" when "01111011001001100", -- t[63052] = 37
      "0100101" when "01111011001001101", -- t[63053] = 37
      "0100101" when "01111011001001110", -- t[63054] = 37
      "0100101" when "01111011001001111", -- t[63055] = 37
      "0100101" when "01111011001010000", -- t[63056] = 37
      "0100101" when "01111011001010001", -- t[63057] = 37
      "0100101" when "01111011001010010", -- t[63058] = 37
      "0100101" when "01111011001010011", -- t[63059] = 37
      "0100101" when "01111011001010100", -- t[63060] = 37
      "0100110" when "01111011001010101", -- t[63061] = 38
      "0100110" when "01111011001010110", -- t[63062] = 38
      "0100110" when "01111011001010111", -- t[63063] = 38
      "0100110" when "01111011001011000", -- t[63064] = 38
      "0100110" when "01111011001011001", -- t[63065] = 38
      "0100110" when "01111011001011010", -- t[63066] = 38
      "0100110" when "01111011001011011", -- t[63067] = 38
      "0100110" when "01111011001011100", -- t[63068] = 38
      "0100110" when "01111011001011101", -- t[63069] = 38
      "0100110" when "01111011001011110", -- t[63070] = 38
      "0100110" when "01111011001011111", -- t[63071] = 38
      "0100110" when "01111011001100000", -- t[63072] = 38
      "0100110" when "01111011001100001", -- t[63073] = 38
      "0100110" when "01111011001100010", -- t[63074] = 38
      "0100110" when "01111011001100011", -- t[63075] = 38
      "0100110" when "01111011001100100", -- t[63076] = 38
      "0100110" when "01111011001100101", -- t[63077] = 38
      "0100110" when "01111011001100110", -- t[63078] = 38
      "0100110" when "01111011001100111", -- t[63079] = 38
      "0100110" when "01111011001101000", -- t[63080] = 38
      "0100110" when "01111011001101001", -- t[63081] = 38
      "0100110" when "01111011001101010", -- t[63082] = 38
      "0100110" when "01111011001101011", -- t[63083] = 38
      "0100110" when "01111011001101100", -- t[63084] = 38
      "0100110" when "01111011001101101", -- t[63085] = 38
      "0100110" when "01111011001101110", -- t[63086] = 38
      "0100110" when "01111011001101111", -- t[63087] = 38
      "0100110" when "01111011001110000", -- t[63088] = 38
      "0100110" when "01111011001110001", -- t[63089] = 38
      "0100110" when "01111011001110010", -- t[63090] = 38
      "0100110" when "01111011001110011", -- t[63091] = 38
      "0100110" when "01111011001110100", -- t[63092] = 38
      "0100110" when "01111011001110101", -- t[63093] = 38
      "0100110" when "01111011001110110", -- t[63094] = 38
      "0100110" when "01111011001110111", -- t[63095] = 38
      "0100110" when "01111011001111000", -- t[63096] = 38
      "0100110" when "01111011001111001", -- t[63097] = 38
      "0100110" when "01111011001111010", -- t[63098] = 38
      "0100110" when "01111011001111011", -- t[63099] = 38
      "0100110" when "01111011001111100", -- t[63100] = 38
      "0100110" when "01111011001111101", -- t[63101] = 38
      "0100110" when "01111011001111110", -- t[63102] = 38
      "0100110" when "01111011001111111", -- t[63103] = 38
      "0100110" when "01111011010000000", -- t[63104] = 38
      "0100110" when "01111011010000001", -- t[63105] = 38
      "0100110" when "01111011010000010", -- t[63106] = 38
      "0100110" when "01111011010000011", -- t[63107] = 38
      "0100110" when "01111011010000100", -- t[63108] = 38
      "0100110" when "01111011010000101", -- t[63109] = 38
      "0100110" when "01111011010000110", -- t[63110] = 38
      "0100110" when "01111011010000111", -- t[63111] = 38
      "0100110" when "01111011010001000", -- t[63112] = 38
      "0100110" when "01111011010001001", -- t[63113] = 38
      "0100110" when "01111011010001010", -- t[63114] = 38
      "0100110" when "01111011010001011", -- t[63115] = 38
      "0100110" when "01111011010001100", -- t[63116] = 38
      "0100110" when "01111011010001101", -- t[63117] = 38
      "0100110" when "01111011010001110", -- t[63118] = 38
      "0100110" when "01111011010001111", -- t[63119] = 38
      "0100110" when "01111011010010000", -- t[63120] = 38
      "0100110" when "01111011010010001", -- t[63121] = 38
      "0100110" when "01111011010010010", -- t[63122] = 38
      "0100110" when "01111011010010011", -- t[63123] = 38
      "0100110" when "01111011010010100", -- t[63124] = 38
      "0100110" when "01111011010010101", -- t[63125] = 38
      "0100110" when "01111011010010110", -- t[63126] = 38
      "0100110" when "01111011010010111", -- t[63127] = 38
      "0100110" when "01111011010011000", -- t[63128] = 38
      "0100110" when "01111011010011001", -- t[63129] = 38
      "0100110" when "01111011010011010", -- t[63130] = 38
      "0100110" when "01111011010011011", -- t[63131] = 38
      "0100110" when "01111011010011100", -- t[63132] = 38
      "0100110" when "01111011010011101", -- t[63133] = 38
      "0100110" when "01111011010011110", -- t[63134] = 38
      "0100110" when "01111011010011111", -- t[63135] = 38
      "0100110" when "01111011010100000", -- t[63136] = 38
      "0100110" when "01111011010100001", -- t[63137] = 38
      "0100110" when "01111011010100010", -- t[63138] = 38
      "0100110" when "01111011010100011", -- t[63139] = 38
      "0100110" when "01111011010100100", -- t[63140] = 38
      "0100110" when "01111011010100101", -- t[63141] = 38
      "0100110" when "01111011010100110", -- t[63142] = 38
      "0100110" when "01111011010100111", -- t[63143] = 38
      "0100110" when "01111011010101000", -- t[63144] = 38
      "0100110" when "01111011010101001", -- t[63145] = 38
      "0100110" when "01111011010101010", -- t[63146] = 38
      "0100110" when "01111011010101011", -- t[63147] = 38
      "0100110" when "01111011010101100", -- t[63148] = 38
      "0100110" when "01111011010101101", -- t[63149] = 38
      "0100110" when "01111011010101110", -- t[63150] = 38
      "0100110" when "01111011010101111", -- t[63151] = 38
      "0100110" when "01111011010110000", -- t[63152] = 38
      "0100110" when "01111011010110001", -- t[63153] = 38
      "0100110" when "01111011010110010", -- t[63154] = 38
      "0100110" when "01111011010110011", -- t[63155] = 38
      "0100110" when "01111011010110100", -- t[63156] = 38
      "0100110" when "01111011010110101", -- t[63157] = 38
      "0100110" when "01111011010110110", -- t[63158] = 38
      "0100110" when "01111011010110111", -- t[63159] = 38
      "0100110" when "01111011010111000", -- t[63160] = 38
      "0100110" when "01111011010111001", -- t[63161] = 38
      "0100110" when "01111011010111010", -- t[63162] = 38
      "0100110" when "01111011010111011", -- t[63163] = 38
      "0100110" when "01111011010111100", -- t[63164] = 38
      "0100110" when "01111011010111101", -- t[63165] = 38
      "0100110" when "01111011010111110", -- t[63166] = 38
      "0100110" when "01111011010111111", -- t[63167] = 38
      "0100110" when "01111011011000000", -- t[63168] = 38
      "0100110" when "01111011011000001", -- t[63169] = 38
      "0100110" when "01111011011000010", -- t[63170] = 38
      "0100110" when "01111011011000011", -- t[63171] = 38
      "0100110" when "01111011011000100", -- t[63172] = 38
      "0100110" when "01111011011000101", -- t[63173] = 38
      "0100110" when "01111011011000110", -- t[63174] = 38
      "0100110" when "01111011011000111", -- t[63175] = 38
      "0100110" when "01111011011001000", -- t[63176] = 38
      "0100110" when "01111011011001001", -- t[63177] = 38
      "0100110" when "01111011011001010", -- t[63178] = 38
      "0100110" when "01111011011001011", -- t[63179] = 38
      "0100110" when "01111011011001100", -- t[63180] = 38
      "0100110" when "01111011011001101", -- t[63181] = 38
      "0100110" when "01111011011001110", -- t[63182] = 38
      "0100110" when "01111011011001111", -- t[63183] = 38
      "0100110" when "01111011011010000", -- t[63184] = 38
      "0100110" when "01111011011010001", -- t[63185] = 38
      "0100110" when "01111011011010010", -- t[63186] = 38
      "0100110" when "01111011011010011", -- t[63187] = 38
      "0100110" when "01111011011010100", -- t[63188] = 38
      "0100110" when "01111011011010101", -- t[63189] = 38
      "0100110" when "01111011011010110", -- t[63190] = 38
      "0100110" when "01111011011010111", -- t[63191] = 38
      "0100110" when "01111011011011000", -- t[63192] = 38
      "0100110" when "01111011011011001", -- t[63193] = 38
      "0100110" when "01111011011011010", -- t[63194] = 38
      "0100110" when "01111011011011011", -- t[63195] = 38
      "0100110" when "01111011011011100", -- t[63196] = 38
      "0100110" when "01111011011011101", -- t[63197] = 38
      "0100110" when "01111011011011110", -- t[63198] = 38
      "0100110" when "01111011011011111", -- t[63199] = 38
      "0100110" when "01111011011100000", -- t[63200] = 38
      "0100110" when "01111011011100001", -- t[63201] = 38
      "0100110" when "01111011011100010", -- t[63202] = 38
      "0100110" when "01111011011100011", -- t[63203] = 38
      "0100110" when "01111011011100100", -- t[63204] = 38
      "0100110" when "01111011011100101", -- t[63205] = 38
      "0100110" when "01111011011100110", -- t[63206] = 38
      "0100110" when "01111011011100111", -- t[63207] = 38
      "0100110" when "01111011011101000", -- t[63208] = 38
      "0100110" when "01111011011101001", -- t[63209] = 38
      "0100110" when "01111011011101010", -- t[63210] = 38
      "0100110" when "01111011011101011", -- t[63211] = 38
      "0100110" when "01111011011101100", -- t[63212] = 38
      "0100110" when "01111011011101101", -- t[63213] = 38
      "0100110" when "01111011011101110", -- t[63214] = 38
      "0100110" when "01111011011101111", -- t[63215] = 38
      "0100110" when "01111011011110000", -- t[63216] = 38
      "0100110" when "01111011011110001", -- t[63217] = 38
      "0100110" when "01111011011110010", -- t[63218] = 38
      "0100110" when "01111011011110011", -- t[63219] = 38
      "0100110" when "01111011011110100", -- t[63220] = 38
      "0100110" when "01111011011110101", -- t[63221] = 38
      "0100110" when "01111011011110110", -- t[63222] = 38
      "0100110" when "01111011011110111", -- t[63223] = 38
      "0100110" when "01111011011111000", -- t[63224] = 38
      "0100110" when "01111011011111001", -- t[63225] = 38
      "0100110" when "01111011011111010", -- t[63226] = 38
      "0100110" when "01111011011111011", -- t[63227] = 38
      "0100110" when "01111011011111100", -- t[63228] = 38
      "0100110" when "01111011011111101", -- t[63229] = 38
      "0100110" when "01111011011111110", -- t[63230] = 38
      "0100110" when "01111011011111111", -- t[63231] = 38
      "0100110" when "01111011100000000", -- t[63232] = 38
      "0100110" when "01111011100000001", -- t[63233] = 38
      "0100110" when "01111011100000010", -- t[63234] = 38
      "0100110" when "01111011100000011", -- t[63235] = 38
      "0100110" when "01111011100000100", -- t[63236] = 38
      "0100110" when "01111011100000101", -- t[63237] = 38
      "0100110" when "01111011100000110", -- t[63238] = 38
      "0100110" when "01111011100000111", -- t[63239] = 38
      "0100110" when "01111011100001000", -- t[63240] = 38
      "0100110" when "01111011100001001", -- t[63241] = 38
      "0100110" when "01111011100001010", -- t[63242] = 38
      "0100110" when "01111011100001011", -- t[63243] = 38
      "0100110" when "01111011100001100", -- t[63244] = 38
      "0100110" when "01111011100001101", -- t[63245] = 38
      "0100110" when "01111011100001110", -- t[63246] = 38
      "0100110" when "01111011100001111", -- t[63247] = 38
      "0100110" when "01111011100010000", -- t[63248] = 38
      "0100110" when "01111011100010001", -- t[63249] = 38
      "0100110" when "01111011100010010", -- t[63250] = 38
      "0100110" when "01111011100010011", -- t[63251] = 38
      "0100110" when "01111011100010100", -- t[63252] = 38
      "0100110" when "01111011100010101", -- t[63253] = 38
      "0100110" when "01111011100010110", -- t[63254] = 38
      "0100110" when "01111011100010111", -- t[63255] = 38
      "0100110" when "01111011100011000", -- t[63256] = 38
      "0100110" when "01111011100011001", -- t[63257] = 38
      "0100110" when "01111011100011010", -- t[63258] = 38
      "0100110" when "01111011100011011", -- t[63259] = 38
      "0100110" when "01111011100011100", -- t[63260] = 38
      "0100110" when "01111011100011101", -- t[63261] = 38
      "0100110" when "01111011100011110", -- t[63262] = 38
      "0100110" when "01111011100011111", -- t[63263] = 38
      "0100110" when "01111011100100000", -- t[63264] = 38
      "0100110" when "01111011100100001", -- t[63265] = 38
      "0100110" when "01111011100100010", -- t[63266] = 38
      "0100110" when "01111011100100011", -- t[63267] = 38
      "0100110" when "01111011100100100", -- t[63268] = 38
      "0100110" when "01111011100100101", -- t[63269] = 38
      "0100110" when "01111011100100110", -- t[63270] = 38
      "0100110" when "01111011100100111", -- t[63271] = 38
      "0100110" when "01111011100101000", -- t[63272] = 38
      "0100110" when "01111011100101001", -- t[63273] = 38
      "0100110" when "01111011100101010", -- t[63274] = 38
      "0100110" when "01111011100101011", -- t[63275] = 38
      "0100110" when "01111011100101100", -- t[63276] = 38
      "0100110" when "01111011100101101", -- t[63277] = 38
      "0100110" when "01111011100101110", -- t[63278] = 38
      "0100110" when "01111011100101111", -- t[63279] = 38
      "0100110" when "01111011100110000", -- t[63280] = 38
      "0100110" when "01111011100110001", -- t[63281] = 38
      "0100110" when "01111011100110010", -- t[63282] = 38
      "0100110" when "01111011100110011", -- t[63283] = 38
      "0100110" when "01111011100110100", -- t[63284] = 38
      "0100110" when "01111011100110101", -- t[63285] = 38
      "0100110" when "01111011100110110", -- t[63286] = 38
      "0100110" when "01111011100110111", -- t[63287] = 38
      "0100110" when "01111011100111000", -- t[63288] = 38
      "0100110" when "01111011100111001", -- t[63289] = 38
      "0100110" when "01111011100111010", -- t[63290] = 38
      "0100110" when "01111011100111011", -- t[63291] = 38
      "0100110" when "01111011100111100", -- t[63292] = 38
      "0100110" when "01111011100111101", -- t[63293] = 38
      "0100110" when "01111011100111110", -- t[63294] = 38
      "0100110" when "01111011100111111", -- t[63295] = 38
      "0100110" when "01111011101000000", -- t[63296] = 38
      "0100110" when "01111011101000001", -- t[63297] = 38
      "0100110" when "01111011101000010", -- t[63298] = 38
      "0100110" when "01111011101000011", -- t[63299] = 38
      "0100110" when "01111011101000100", -- t[63300] = 38
      "0100110" when "01111011101000101", -- t[63301] = 38
      "0100110" when "01111011101000110", -- t[63302] = 38
      "0100110" when "01111011101000111", -- t[63303] = 38
      "0100110" when "01111011101001000", -- t[63304] = 38
      "0100110" when "01111011101001001", -- t[63305] = 38
      "0100110" when "01111011101001010", -- t[63306] = 38
      "0100110" when "01111011101001011", -- t[63307] = 38
      "0100110" when "01111011101001100", -- t[63308] = 38
      "0100110" when "01111011101001101", -- t[63309] = 38
      "0100110" when "01111011101001110", -- t[63310] = 38
      "0100110" when "01111011101001111", -- t[63311] = 38
      "0100110" when "01111011101010000", -- t[63312] = 38
      "0100110" when "01111011101010001", -- t[63313] = 38
      "0100110" when "01111011101010010", -- t[63314] = 38
      "0100110" when "01111011101010011", -- t[63315] = 38
      "0100110" when "01111011101010100", -- t[63316] = 38
      "0100110" when "01111011101010101", -- t[63317] = 38
      "0100110" when "01111011101010110", -- t[63318] = 38
      "0100110" when "01111011101010111", -- t[63319] = 38
      "0100110" when "01111011101011000", -- t[63320] = 38
      "0100110" when "01111011101011001", -- t[63321] = 38
      "0100110" when "01111011101011010", -- t[63322] = 38
      "0100110" when "01111011101011011", -- t[63323] = 38
      "0100110" when "01111011101011100", -- t[63324] = 38
      "0100110" when "01111011101011101", -- t[63325] = 38
      "0100110" when "01111011101011110", -- t[63326] = 38
      "0100110" when "01111011101011111", -- t[63327] = 38
      "0100110" when "01111011101100000", -- t[63328] = 38
      "0100110" when "01111011101100001", -- t[63329] = 38
      "0100110" when "01111011101100010", -- t[63330] = 38
      "0100110" when "01111011101100011", -- t[63331] = 38
      "0100110" when "01111011101100100", -- t[63332] = 38
      "0100110" when "01111011101100101", -- t[63333] = 38
      "0100110" when "01111011101100110", -- t[63334] = 38
      "0100110" when "01111011101100111", -- t[63335] = 38
      "0100110" when "01111011101101000", -- t[63336] = 38
      "0100110" when "01111011101101001", -- t[63337] = 38
      "0100110" when "01111011101101010", -- t[63338] = 38
      "0100110" when "01111011101101011", -- t[63339] = 38
      "0100110" when "01111011101101100", -- t[63340] = 38
      "0100110" when "01111011101101101", -- t[63341] = 38
      "0100110" when "01111011101101110", -- t[63342] = 38
      "0100110" when "01111011101101111", -- t[63343] = 38
      "0100110" when "01111011101110000", -- t[63344] = 38
      "0100110" when "01111011101110001", -- t[63345] = 38
      "0100110" when "01111011101110010", -- t[63346] = 38
      "0100110" when "01111011101110011", -- t[63347] = 38
      "0100110" when "01111011101110100", -- t[63348] = 38
      "0100110" when "01111011101110101", -- t[63349] = 38
      "0100110" when "01111011101110110", -- t[63350] = 38
      "0100110" when "01111011101110111", -- t[63351] = 38
      "0100110" when "01111011101111000", -- t[63352] = 38
      "0100110" when "01111011101111001", -- t[63353] = 38
      "0100110" when "01111011101111010", -- t[63354] = 38
      "0100110" when "01111011101111011", -- t[63355] = 38
      "0100110" when "01111011101111100", -- t[63356] = 38
      "0100110" when "01111011101111101", -- t[63357] = 38
      "0100110" when "01111011101111110", -- t[63358] = 38
      "0100110" when "01111011101111111", -- t[63359] = 38
      "0100110" when "01111011110000000", -- t[63360] = 38
      "0100110" when "01111011110000001", -- t[63361] = 38
      "0100110" when "01111011110000010", -- t[63362] = 38
      "0100110" when "01111011110000011", -- t[63363] = 38
      "0100110" when "01111011110000100", -- t[63364] = 38
      "0100110" when "01111011110000101", -- t[63365] = 38
      "0100110" when "01111011110000110", -- t[63366] = 38
      "0100110" when "01111011110000111", -- t[63367] = 38
      "0100110" when "01111011110001000", -- t[63368] = 38
      "0100110" when "01111011110001001", -- t[63369] = 38
      "0100110" when "01111011110001010", -- t[63370] = 38
      "0100111" when "01111011110001011", -- t[63371] = 39
      "0100111" when "01111011110001100", -- t[63372] = 39
      "0100111" when "01111011110001101", -- t[63373] = 39
      "0100111" when "01111011110001110", -- t[63374] = 39
      "0100111" when "01111011110001111", -- t[63375] = 39
      "0100111" when "01111011110010000", -- t[63376] = 39
      "0100111" when "01111011110010001", -- t[63377] = 39
      "0100111" when "01111011110010010", -- t[63378] = 39
      "0100111" when "01111011110010011", -- t[63379] = 39
      "0100111" when "01111011110010100", -- t[63380] = 39
      "0100111" when "01111011110010101", -- t[63381] = 39
      "0100111" when "01111011110010110", -- t[63382] = 39
      "0100111" when "01111011110010111", -- t[63383] = 39
      "0100111" when "01111011110011000", -- t[63384] = 39
      "0100111" when "01111011110011001", -- t[63385] = 39
      "0100111" when "01111011110011010", -- t[63386] = 39
      "0100111" when "01111011110011011", -- t[63387] = 39
      "0100111" when "01111011110011100", -- t[63388] = 39
      "0100111" when "01111011110011101", -- t[63389] = 39
      "0100111" when "01111011110011110", -- t[63390] = 39
      "0100111" when "01111011110011111", -- t[63391] = 39
      "0100111" when "01111011110100000", -- t[63392] = 39
      "0100111" when "01111011110100001", -- t[63393] = 39
      "0100111" when "01111011110100010", -- t[63394] = 39
      "0100111" when "01111011110100011", -- t[63395] = 39
      "0100111" when "01111011110100100", -- t[63396] = 39
      "0100111" when "01111011110100101", -- t[63397] = 39
      "0100111" when "01111011110100110", -- t[63398] = 39
      "0100111" when "01111011110100111", -- t[63399] = 39
      "0100111" when "01111011110101000", -- t[63400] = 39
      "0100111" when "01111011110101001", -- t[63401] = 39
      "0100111" when "01111011110101010", -- t[63402] = 39
      "0100111" when "01111011110101011", -- t[63403] = 39
      "0100111" when "01111011110101100", -- t[63404] = 39
      "0100111" when "01111011110101101", -- t[63405] = 39
      "0100111" when "01111011110101110", -- t[63406] = 39
      "0100111" when "01111011110101111", -- t[63407] = 39
      "0100111" when "01111011110110000", -- t[63408] = 39
      "0100111" when "01111011110110001", -- t[63409] = 39
      "0100111" when "01111011110110010", -- t[63410] = 39
      "0100111" when "01111011110110011", -- t[63411] = 39
      "0100111" when "01111011110110100", -- t[63412] = 39
      "0100111" when "01111011110110101", -- t[63413] = 39
      "0100111" when "01111011110110110", -- t[63414] = 39
      "0100111" when "01111011110110111", -- t[63415] = 39
      "0100111" when "01111011110111000", -- t[63416] = 39
      "0100111" when "01111011110111001", -- t[63417] = 39
      "0100111" when "01111011110111010", -- t[63418] = 39
      "0100111" when "01111011110111011", -- t[63419] = 39
      "0100111" when "01111011110111100", -- t[63420] = 39
      "0100111" when "01111011110111101", -- t[63421] = 39
      "0100111" when "01111011110111110", -- t[63422] = 39
      "0100111" when "01111011110111111", -- t[63423] = 39
      "0100111" when "01111011111000000", -- t[63424] = 39
      "0100111" when "01111011111000001", -- t[63425] = 39
      "0100111" when "01111011111000010", -- t[63426] = 39
      "0100111" when "01111011111000011", -- t[63427] = 39
      "0100111" when "01111011111000100", -- t[63428] = 39
      "0100111" when "01111011111000101", -- t[63429] = 39
      "0100111" when "01111011111000110", -- t[63430] = 39
      "0100111" when "01111011111000111", -- t[63431] = 39
      "0100111" when "01111011111001000", -- t[63432] = 39
      "0100111" when "01111011111001001", -- t[63433] = 39
      "0100111" when "01111011111001010", -- t[63434] = 39
      "0100111" when "01111011111001011", -- t[63435] = 39
      "0100111" when "01111011111001100", -- t[63436] = 39
      "0100111" when "01111011111001101", -- t[63437] = 39
      "0100111" when "01111011111001110", -- t[63438] = 39
      "0100111" when "01111011111001111", -- t[63439] = 39
      "0100111" when "01111011111010000", -- t[63440] = 39
      "0100111" when "01111011111010001", -- t[63441] = 39
      "0100111" when "01111011111010010", -- t[63442] = 39
      "0100111" when "01111011111010011", -- t[63443] = 39
      "0100111" when "01111011111010100", -- t[63444] = 39
      "0100111" when "01111011111010101", -- t[63445] = 39
      "0100111" when "01111011111010110", -- t[63446] = 39
      "0100111" when "01111011111010111", -- t[63447] = 39
      "0100111" when "01111011111011000", -- t[63448] = 39
      "0100111" when "01111011111011001", -- t[63449] = 39
      "0100111" when "01111011111011010", -- t[63450] = 39
      "0100111" when "01111011111011011", -- t[63451] = 39
      "0100111" when "01111011111011100", -- t[63452] = 39
      "0100111" when "01111011111011101", -- t[63453] = 39
      "0100111" when "01111011111011110", -- t[63454] = 39
      "0100111" when "01111011111011111", -- t[63455] = 39
      "0100111" when "01111011111100000", -- t[63456] = 39
      "0100111" when "01111011111100001", -- t[63457] = 39
      "0100111" when "01111011111100010", -- t[63458] = 39
      "0100111" when "01111011111100011", -- t[63459] = 39
      "0100111" when "01111011111100100", -- t[63460] = 39
      "0100111" when "01111011111100101", -- t[63461] = 39
      "0100111" when "01111011111100110", -- t[63462] = 39
      "0100111" when "01111011111100111", -- t[63463] = 39
      "0100111" when "01111011111101000", -- t[63464] = 39
      "0100111" when "01111011111101001", -- t[63465] = 39
      "0100111" when "01111011111101010", -- t[63466] = 39
      "0100111" when "01111011111101011", -- t[63467] = 39
      "0100111" when "01111011111101100", -- t[63468] = 39
      "0100111" when "01111011111101101", -- t[63469] = 39
      "0100111" when "01111011111101110", -- t[63470] = 39
      "0100111" when "01111011111101111", -- t[63471] = 39
      "0100111" when "01111011111110000", -- t[63472] = 39
      "0100111" when "01111011111110001", -- t[63473] = 39
      "0100111" when "01111011111110010", -- t[63474] = 39
      "0100111" when "01111011111110011", -- t[63475] = 39
      "0100111" when "01111011111110100", -- t[63476] = 39
      "0100111" when "01111011111110101", -- t[63477] = 39
      "0100111" when "01111011111110110", -- t[63478] = 39
      "0100111" when "01111011111110111", -- t[63479] = 39
      "0100111" when "01111011111111000", -- t[63480] = 39
      "0100111" when "01111011111111001", -- t[63481] = 39
      "0100111" when "01111011111111010", -- t[63482] = 39
      "0100111" when "01111011111111011", -- t[63483] = 39
      "0100111" when "01111011111111100", -- t[63484] = 39
      "0100111" when "01111011111111101", -- t[63485] = 39
      "0100111" when "01111011111111110", -- t[63486] = 39
      "0100111" when "01111011111111111", -- t[63487] = 39
      "0100111" when "01111100000000000", -- t[63488] = 39
      "0100111" when "01111100000000001", -- t[63489] = 39
      "0100111" when "01111100000000010", -- t[63490] = 39
      "0100111" when "01111100000000011", -- t[63491] = 39
      "0100111" when "01111100000000100", -- t[63492] = 39
      "0100111" when "01111100000000101", -- t[63493] = 39
      "0100111" when "01111100000000110", -- t[63494] = 39
      "0100111" when "01111100000000111", -- t[63495] = 39
      "0100111" when "01111100000001000", -- t[63496] = 39
      "0100111" when "01111100000001001", -- t[63497] = 39
      "0100111" when "01111100000001010", -- t[63498] = 39
      "0100111" when "01111100000001011", -- t[63499] = 39
      "0100111" when "01111100000001100", -- t[63500] = 39
      "0100111" when "01111100000001101", -- t[63501] = 39
      "0100111" when "01111100000001110", -- t[63502] = 39
      "0100111" when "01111100000001111", -- t[63503] = 39
      "0100111" when "01111100000010000", -- t[63504] = 39
      "0100111" when "01111100000010001", -- t[63505] = 39
      "0100111" when "01111100000010010", -- t[63506] = 39
      "0100111" when "01111100000010011", -- t[63507] = 39
      "0100111" when "01111100000010100", -- t[63508] = 39
      "0100111" when "01111100000010101", -- t[63509] = 39
      "0100111" when "01111100000010110", -- t[63510] = 39
      "0100111" when "01111100000010111", -- t[63511] = 39
      "0100111" when "01111100000011000", -- t[63512] = 39
      "0100111" when "01111100000011001", -- t[63513] = 39
      "0100111" when "01111100000011010", -- t[63514] = 39
      "0100111" when "01111100000011011", -- t[63515] = 39
      "0100111" when "01111100000011100", -- t[63516] = 39
      "0100111" when "01111100000011101", -- t[63517] = 39
      "0100111" when "01111100000011110", -- t[63518] = 39
      "0100111" when "01111100000011111", -- t[63519] = 39
      "0100111" when "01111100000100000", -- t[63520] = 39
      "0100111" when "01111100000100001", -- t[63521] = 39
      "0100111" when "01111100000100010", -- t[63522] = 39
      "0100111" when "01111100000100011", -- t[63523] = 39
      "0100111" when "01111100000100100", -- t[63524] = 39
      "0100111" when "01111100000100101", -- t[63525] = 39
      "0100111" when "01111100000100110", -- t[63526] = 39
      "0100111" when "01111100000100111", -- t[63527] = 39
      "0100111" when "01111100000101000", -- t[63528] = 39
      "0100111" when "01111100000101001", -- t[63529] = 39
      "0100111" when "01111100000101010", -- t[63530] = 39
      "0100111" when "01111100000101011", -- t[63531] = 39
      "0100111" when "01111100000101100", -- t[63532] = 39
      "0100111" when "01111100000101101", -- t[63533] = 39
      "0100111" when "01111100000101110", -- t[63534] = 39
      "0100111" when "01111100000101111", -- t[63535] = 39
      "0100111" when "01111100000110000", -- t[63536] = 39
      "0100111" when "01111100000110001", -- t[63537] = 39
      "0100111" when "01111100000110010", -- t[63538] = 39
      "0100111" when "01111100000110011", -- t[63539] = 39
      "0100111" when "01111100000110100", -- t[63540] = 39
      "0100111" when "01111100000110101", -- t[63541] = 39
      "0100111" when "01111100000110110", -- t[63542] = 39
      "0100111" when "01111100000110111", -- t[63543] = 39
      "0100111" when "01111100000111000", -- t[63544] = 39
      "0100111" when "01111100000111001", -- t[63545] = 39
      "0100111" when "01111100000111010", -- t[63546] = 39
      "0100111" when "01111100000111011", -- t[63547] = 39
      "0100111" when "01111100000111100", -- t[63548] = 39
      "0100111" when "01111100000111101", -- t[63549] = 39
      "0100111" when "01111100000111110", -- t[63550] = 39
      "0100111" when "01111100000111111", -- t[63551] = 39
      "0100111" when "01111100001000000", -- t[63552] = 39
      "0100111" when "01111100001000001", -- t[63553] = 39
      "0100111" when "01111100001000010", -- t[63554] = 39
      "0100111" when "01111100001000011", -- t[63555] = 39
      "0100111" when "01111100001000100", -- t[63556] = 39
      "0100111" when "01111100001000101", -- t[63557] = 39
      "0100111" when "01111100001000110", -- t[63558] = 39
      "0100111" when "01111100001000111", -- t[63559] = 39
      "0100111" when "01111100001001000", -- t[63560] = 39
      "0100111" when "01111100001001001", -- t[63561] = 39
      "0100111" when "01111100001001010", -- t[63562] = 39
      "0100111" when "01111100001001011", -- t[63563] = 39
      "0100111" when "01111100001001100", -- t[63564] = 39
      "0100111" when "01111100001001101", -- t[63565] = 39
      "0100111" when "01111100001001110", -- t[63566] = 39
      "0100111" when "01111100001001111", -- t[63567] = 39
      "0100111" when "01111100001010000", -- t[63568] = 39
      "0100111" when "01111100001010001", -- t[63569] = 39
      "0100111" when "01111100001010010", -- t[63570] = 39
      "0100111" when "01111100001010011", -- t[63571] = 39
      "0100111" when "01111100001010100", -- t[63572] = 39
      "0100111" when "01111100001010101", -- t[63573] = 39
      "0100111" when "01111100001010110", -- t[63574] = 39
      "0100111" when "01111100001010111", -- t[63575] = 39
      "0100111" when "01111100001011000", -- t[63576] = 39
      "0100111" when "01111100001011001", -- t[63577] = 39
      "0100111" when "01111100001011010", -- t[63578] = 39
      "0100111" when "01111100001011011", -- t[63579] = 39
      "0100111" when "01111100001011100", -- t[63580] = 39
      "0100111" when "01111100001011101", -- t[63581] = 39
      "0100111" when "01111100001011110", -- t[63582] = 39
      "0100111" when "01111100001011111", -- t[63583] = 39
      "0100111" when "01111100001100000", -- t[63584] = 39
      "0100111" when "01111100001100001", -- t[63585] = 39
      "0100111" when "01111100001100010", -- t[63586] = 39
      "0100111" when "01111100001100011", -- t[63587] = 39
      "0100111" when "01111100001100100", -- t[63588] = 39
      "0100111" when "01111100001100101", -- t[63589] = 39
      "0100111" when "01111100001100110", -- t[63590] = 39
      "0100111" when "01111100001100111", -- t[63591] = 39
      "0100111" when "01111100001101000", -- t[63592] = 39
      "0100111" when "01111100001101001", -- t[63593] = 39
      "0100111" when "01111100001101010", -- t[63594] = 39
      "0100111" when "01111100001101011", -- t[63595] = 39
      "0100111" when "01111100001101100", -- t[63596] = 39
      "0100111" when "01111100001101101", -- t[63597] = 39
      "0100111" when "01111100001101110", -- t[63598] = 39
      "0100111" when "01111100001101111", -- t[63599] = 39
      "0100111" when "01111100001110000", -- t[63600] = 39
      "0100111" when "01111100001110001", -- t[63601] = 39
      "0100111" when "01111100001110010", -- t[63602] = 39
      "0100111" when "01111100001110011", -- t[63603] = 39
      "0100111" when "01111100001110100", -- t[63604] = 39
      "0100111" when "01111100001110101", -- t[63605] = 39
      "0100111" when "01111100001110110", -- t[63606] = 39
      "0100111" when "01111100001110111", -- t[63607] = 39
      "0100111" when "01111100001111000", -- t[63608] = 39
      "0100111" when "01111100001111001", -- t[63609] = 39
      "0100111" when "01111100001111010", -- t[63610] = 39
      "0100111" when "01111100001111011", -- t[63611] = 39
      "0100111" when "01111100001111100", -- t[63612] = 39
      "0100111" when "01111100001111101", -- t[63613] = 39
      "0100111" when "01111100001111110", -- t[63614] = 39
      "0100111" when "01111100001111111", -- t[63615] = 39
      "0100111" when "01111100010000000", -- t[63616] = 39
      "0100111" when "01111100010000001", -- t[63617] = 39
      "0100111" when "01111100010000010", -- t[63618] = 39
      "0100111" when "01111100010000011", -- t[63619] = 39
      "0100111" when "01111100010000100", -- t[63620] = 39
      "0100111" when "01111100010000101", -- t[63621] = 39
      "0100111" when "01111100010000110", -- t[63622] = 39
      "0100111" when "01111100010000111", -- t[63623] = 39
      "0100111" when "01111100010001000", -- t[63624] = 39
      "0100111" when "01111100010001001", -- t[63625] = 39
      "0100111" when "01111100010001010", -- t[63626] = 39
      "0100111" when "01111100010001011", -- t[63627] = 39
      "0100111" when "01111100010001100", -- t[63628] = 39
      "0100111" when "01111100010001101", -- t[63629] = 39
      "0100111" when "01111100010001110", -- t[63630] = 39
      "0100111" when "01111100010001111", -- t[63631] = 39
      "0100111" when "01111100010010000", -- t[63632] = 39
      "0100111" when "01111100010010001", -- t[63633] = 39
      "0100111" when "01111100010010010", -- t[63634] = 39
      "0100111" when "01111100010010011", -- t[63635] = 39
      "0100111" when "01111100010010100", -- t[63636] = 39
      "0100111" when "01111100010010101", -- t[63637] = 39
      "0100111" when "01111100010010110", -- t[63638] = 39
      "0100111" when "01111100010010111", -- t[63639] = 39
      "0100111" when "01111100010011000", -- t[63640] = 39
      "0100111" when "01111100010011001", -- t[63641] = 39
      "0100111" when "01111100010011010", -- t[63642] = 39
      "0100111" when "01111100010011011", -- t[63643] = 39
      "0100111" when "01111100010011100", -- t[63644] = 39
      "0100111" when "01111100010011101", -- t[63645] = 39
      "0100111" when "01111100010011110", -- t[63646] = 39
      "0100111" when "01111100010011111", -- t[63647] = 39
      "0100111" when "01111100010100000", -- t[63648] = 39
      "0100111" when "01111100010100001", -- t[63649] = 39
      "0100111" when "01111100010100010", -- t[63650] = 39
      "0100111" when "01111100010100011", -- t[63651] = 39
      "0100111" when "01111100010100100", -- t[63652] = 39
      "0100111" when "01111100010100101", -- t[63653] = 39
      "0100111" when "01111100010100110", -- t[63654] = 39
      "0100111" when "01111100010100111", -- t[63655] = 39
      "0100111" when "01111100010101000", -- t[63656] = 39
      "0100111" when "01111100010101001", -- t[63657] = 39
      "0100111" when "01111100010101010", -- t[63658] = 39
      "0100111" when "01111100010101011", -- t[63659] = 39
      "0100111" when "01111100010101100", -- t[63660] = 39
      "0100111" when "01111100010101101", -- t[63661] = 39
      "0100111" when "01111100010101110", -- t[63662] = 39
      "0100111" when "01111100010101111", -- t[63663] = 39
      "0100111" when "01111100010110000", -- t[63664] = 39
      "0100111" when "01111100010110001", -- t[63665] = 39
      "0100111" when "01111100010110010", -- t[63666] = 39
      "0100111" when "01111100010110011", -- t[63667] = 39
      "0100111" when "01111100010110100", -- t[63668] = 39
      "0100111" when "01111100010110101", -- t[63669] = 39
      "0100111" when "01111100010110110", -- t[63670] = 39
      "0100111" when "01111100010110111", -- t[63671] = 39
      "0100111" when "01111100010111000", -- t[63672] = 39
      "0100111" when "01111100010111001", -- t[63673] = 39
      "0101000" when "01111100010111010", -- t[63674] = 40
      "0101000" when "01111100010111011", -- t[63675] = 40
      "0101000" when "01111100010111100", -- t[63676] = 40
      "0101000" when "01111100010111101", -- t[63677] = 40
      "0101000" when "01111100010111110", -- t[63678] = 40
      "0101000" when "01111100010111111", -- t[63679] = 40
      "0101000" when "01111100011000000", -- t[63680] = 40
      "0101000" when "01111100011000001", -- t[63681] = 40
      "0101000" when "01111100011000010", -- t[63682] = 40
      "0101000" when "01111100011000011", -- t[63683] = 40
      "0101000" when "01111100011000100", -- t[63684] = 40
      "0101000" when "01111100011000101", -- t[63685] = 40
      "0101000" when "01111100011000110", -- t[63686] = 40
      "0101000" when "01111100011000111", -- t[63687] = 40
      "0101000" when "01111100011001000", -- t[63688] = 40
      "0101000" when "01111100011001001", -- t[63689] = 40
      "0101000" when "01111100011001010", -- t[63690] = 40
      "0101000" when "01111100011001011", -- t[63691] = 40
      "0101000" when "01111100011001100", -- t[63692] = 40
      "0101000" when "01111100011001101", -- t[63693] = 40
      "0101000" when "01111100011001110", -- t[63694] = 40
      "0101000" when "01111100011001111", -- t[63695] = 40
      "0101000" when "01111100011010000", -- t[63696] = 40
      "0101000" when "01111100011010001", -- t[63697] = 40
      "0101000" when "01111100011010010", -- t[63698] = 40
      "0101000" when "01111100011010011", -- t[63699] = 40
      "0101000" when "01111100011010100", -- t[63700] = 40
      "0101000" when "01111100011010101", -- t[63701] = 40
      "0101000" when "01111100011010110", -- t[63702] = 40
      "0101000" when "01111100011010111", -- t[63703] = 40
      "0101000" when "01111100011011000", -- t[63704] = 40
      "0101000" when "01111100011011001", -- t[63705] = 40
      "0101000" when "01111100011011010", -- t[63706] = 40
      "0101000" when "01111100011011011", -- t[63707] = 40
      "0101000" when "01111100011011100", -- t[63708] = 40
      "0101000" when "01111100011011101", -- t[63709] = 40
      "0101000" when "01111100011011110", -- t[63710] = 40
      "0101000" when "01111100011011111", -- t[63711] = 40
      "0101000" when "01111100011100000", -- t[63712] = 40
      "0101000" when "01111100011100001", -- t[63713] = 40
      "0101000" when "01111100011100010", -- t[63714] = 40
      "0101000" when "01111100011100011", -- t[63715] = 40
      "0101000" when "01111100011100100", -- t[63716] = 40
      "0101000" when "01111100011100101", -- t[63717] = 40
      "0101000" when "01111100011100110", -- t[63718] = 40
      "0101000" when "01111100011100111", -- t[63719] = 40
      "0101000" when "01111100011101000", -- t[63720] = 40
      "0101000" when "01111100011101001", -- t[63721] = 40
      "0101000" when "01111100011101010", -- t[63722] = 40
      "0101000" when "01111100011101011", -- t[63723] = 40
      "0101000" when "01111100011101100", -- t[63724] = 40
      "0101000" when "01111100011101101", -- t[63725] = 40
      "0101000" when "01111100011101110", -- t[63726] = 40
      "0101000" when "01111100011101111", -- t[63727] = 40
      "0101000" when "01111100011110000", -- t[63728] = 40
      "0101000" when "01111100011110001", -- t[63729] = 40
      "0101000" when "01111100011110010", -- t[63730] = 40
      "0101000" when "01111100011110011", -- t[63731] = 40
      "0101000" when "01111100011110100", -- t[63732] = 40
      "0101000" when "01111100011110101", -- t[63733] = 40
      "0101000" when "01111100011110110", -- t[63734] = 40
      "0101000" when "01111100011110111", -- t[63735] = 40
      "0101000" when "01111100011111000", -- t[63736] = 40
      "0101000" when "01111100011111001", -- t[63737] = 40
      "0101000" when "01111100011111010", -- t[63738] = 40
      "0101000" when "01111100011111011", -- t[63739] = 40
      "0101000" when "01111100011111100", -- t[63740] = 40
      "0101000" when "01111100011111101", -- t[63741] = 40
      "0101000" when "01111100011111110", -- t[63742] = 40
      "0101000" when "01111100011111111", -- t[63743] = 40
      "0101000" when "01111100100000000", -- t[63744] = 40
      "0101000" when "01111100100000001", -- t[63745] = 40
      "0101000" when "01111100100000010", -- t[63746] = 40
      "0101000" when "01111100100000011", -- t[63747] = 40
      "0101000" when "01111100100000100", -- t[63748] = 40
      "0101000" when "01111100100000101", -- t[63749] = 40
      "0101000" when "01111100100000110", -- t[63750] = 40
      "0101000" when "01111100100000111", -- t[63751] = 40
      "0101000" when "01111100100001000", -- t[63752] = 40
      "0101000" when "01111100100001001", -- t[63753] = 40
      "0101000" when "01111100100001010", -- t[63754] = 40
      "0101000" when "01111100100001011", -- t[63755] = 40
      "0101000" when "01111100100001100", -- t[63756] = 40
      "0101000" when "01111100100001101", -- t[63757] = 40
      "0101000" when "01111100100001110", -- t[63758] = 40
      "0101000" when "01111100100001111", -- t[63759] = 40
      "0101000" when "01111100100010000", -- t[63760] = 40
      "0101000" when "01111100100010001", -- t[63761] = 40
      "0101000" when "01111100100010010", -- t[63762] = 40
      "0101000" when "01111100100010011", -- t[63763] = 40
      "0101000" when "01111100100010100", -- t[63764] = 40
      "0101000" when "01111100100010101", -- t[63765] = 40
      "0101000" when "01111100100010110", -- t[63766] = 40
      "0101000" when "01111100100010111", -- t[63767] = 40
      "0101000" when "01111100100011000", -- t[63768] = 40
      "0101000" when "01111100100011001", -- t[63769] = 40
      "0101000" when "01111100100011010", -- t[63770] = 40
      "0101000" when "01111100100011011", -- t[63771] = 40
      "0101000" when "01111100100011100", -- t[63772] = 40
      "0101000" when "01111100100011101", -- t[63773] = 40
      "0101000" when "01111100100011110", -- t[63774] = 40
      "0101000" when "01111100100011111", -- t[63775] = 40
      "0101000" when "01111100100100000", -- t[63776] = 40
      "0101000" when "01111100100100001", -- t[63777] = 40
      "0101000" when "01111100100100010", -- t[63778] = 40
      "0101000" when "01111100100100011", -- t[63779] = 40
      "0101000" when "01111100100100100", -- t[63780] = 40
      "0101000" when "01111100100100101", -- t[63781] = 40
      "0101000" when "01111100100100110", -- t[63782] = 40
      "0101000" when "01111100100100111", -- t[63783] = 40
      "0101000" when "01111100100101000", -- t[63784] = 40
      "0101000" when "01111100100101001", -- t[63785] = 40
      "0101000" when "01111100100101010", -- t[63786] = 40
      "0101000" when "01111100100101011", -- t[63787] = 40
      "0101000" when "01111100100101100", -- t[63788] = 40
      "0101000" when "01111100100101101", -- t[63789] = 40
      "0101000" when "01111100100101110", -- t[63790] = 40
      "0101000" when "01111100100101111", -- t[63791] = 40
      "0101000" when "01111100100110000", -- t[63792] = 40
      "0101000" when "01111100100110001", -- t[63793] = 40
      "0101000" when "01111100100110010", -- t[63794] = 40
      "0101000" when "01111100100110011", -- t[63795] = 40
      "0101000" when "01111100100110100", -- t[63796] = 40
      "0101000" when "01111100100110101", -- t[63797] = 40
      "0101000" when "01111100100110110", -- t[63798] = 40
      "0101000" when "01111100100110111", -- t[63799] = 40
      "0101000" when "01111100100111000", -- t[63800] = 40
      "0101000" when "01111100100111001", -- t[63801] = 40
      "0101000" when "01111100100111010", -- t[63802] = 40
      "0101000" when "01111100100111011", -- t[63803] = 40
      "0101000" when "01111100100111100", -- t[63804] = 40
      "0101000" when "01111100100111101", -- t[63805] = 40
      "0101000" when "01111100100111110", -- t[63806] = 40
      "0101000" when "01111100100111111", -- t[63807] = 40
      "0101000" when "01111100101000000", -- t[63808] = 40
      "0101000" when "01111100101000001", -- t[63809] = 40
      "0101000" when "01111100101000010", -- t[63810] = 40
      "0101000" when "01111100101000011", -- t[63811] = 40
      "0101000" when "01111100101000100", -- t[63812] = 40
      "0101000" when "01111100101000101", -- t[63813] = 40
      "0101000" when "01111100101000110", -- t[63814] = 40
      "0101000" when "01111100101000111", -- t[63815] = 40
      "0101000" when "01111100101001000", -- t[63816] = 40
      "0101000" when "01111100101001001", -- t[63817] = 40
      "0101000" when "01111100101001010", -- t[63818] = 40
      "0101000" when "01111100101001011", -- t[63819] = 40
      "0101000" when "01111100101001100", -- t[63820] = 40
      "0101000" when "01111100101001101", -- t[63821] = 40
      "0101000" when "01111100101001110", -- t[63822] = 40
      "0101000" when "01111100101001111", -- t[63823] = 40
      "0101000" when "01111100101010000", -- t[63824] = 40
      "0101000" when "01111100101010001", -- t[63825] = 40
      "0101000" when "01111100101010010", -- t[63826] = 40
      "0101000" when "01111100101010011", -- t[63827] = 40
      "0101000" when "01111100101010100", -- t[63828] = 40
      "0101000" when "01111100101010101", -- t[63829] = 40
      "0101000" when "01111100101010110", -- t[63830] = 40
      "0101000" when "01111100101010111", -- t[63831] = 40
      "0101000" when "01111100101011000", -- t[63832] = 40
      "0101000" when "01111100101011001", -- t[63833] = 40
      "0101000" when "01111100101011010", -- t[63834] = 40
      "0101000" when "01111100101011011", -- t[63835] = 40
      "0101000" when "01111100101011100", -- t[63836] = 40
      "0101000" when "01111100101011101", -- t[63837] = 40
      "0101000" when "01111100101011110", -- t[63838] = 40
      "0101000" when "01111100101011111", -- t[63839] = 40
      "0101000" when "01111100101100000", -- t[63840] = 40
      "0101000" when "01111100101100001", -- t[63841] = 40
      "0101000" when "01111100101100010", -- t[63842] = 40
      "0101000" when "01111100101100011", -- t[63843] = 40
      "0101000" when "01111100101100100", -- t[63844] = 40
      "0101000" when "01111100101100101", -- t[63845] = 40
      "0101000" when "01111100101100110", -- t[63846] = 40
      "0101000" when "01111100101100111", -- t[63847] = 40
      "0101000" when "01111100101101000", -- t[63848] = 40
      "0101000" when "01111100101101001", -- t[63849] = 40
      "0101000" when "01111100101101010", -- t[63850] = 40
      "0101000" when "01111100101101011", -- t[63851] = 40
      "0101000" when "01111100101101100", -- t[63852] = 40
      "0101000" when "01111100101101101", -- t[63853] = 40
      "0101000" when "01111100101101110", -- t[63854] = 40
      "0101000" when "01111100101101111", -- t[63855] = 40
      "0101000" when "01111100101110000", -- t[63856] = 40
      "0101000" when "01111100101110001", -- t[63857] = 40
      "0101000" when "01111100101110010", -- t[63858] = 40
      "0101000" when "01111100101110011", -- t[63859] = 40
      "0101000" when "01111100101110100", -- t[63860] = 40
      "0101000" when "01111100101110101", -- t[63861] = 40
      "0101000" when "01111100101110110", -- t[63862] = 40
      "0101000" when "01111100101110111", -- t[63863] = 40
      "0101000" when "01111100101111000", -- t[63864] = 40
      "0101000" when "01111100101111001", -- t[63865] = 40
      "0101000" when "01111100101111010", -- t[63866] = 40
      "0101000" when "01111100101111011", -- t[63867] = 40
      "0101000" when "01111100101111100", -- t[63868] = 40
      "0101000" when "01111100101111101", -- t[63869] = 40
      "0101000" when "01111100101111110", -- t[63870] = 40
      "0101000" when "01111100101111111", -- t[63871] = 40
      "0101000" when "01111100110000000", -- t[63872] = 40
      "0101000" when "01111100110000001", -- t[63873] = 40
      "0101000" when "01111100110000010", -- t[63874] = 40
      "0101000" when "01111100110000011", -- t[63875] = 40
      "0101000" when "01111100110000100", -- t[63876] = 40
      "0101000" when "01111100110000101", -- t[63877] = 40
      "0101000" when "01111100110000110", -- t[63878] = 40
      "0101000" when "01111100110000111", -- t[63879] = 40
      "0101000" when "01111100110001000", -- t[63880] = 40
      "0101000" when "01111100110001001", -- t[63881] = 40
      "0101000" when "01111100110001010", -- t[63882] = 40
      "0101000" when "01111100110001011", -- t[63883] = 40
      "0101000" when "01111100110001100", -- t[63884] = 40
      "0101000" when "01111100110001101", -- t[63885] = 40
      "0101000" when "01111100110001110", -- t[63886] = 40
      "0101000" when "01111100110001111", -- t[63887] = 40
      "0101000" when "01111100110010000", -- t[63888] = 40
      "0101000" when "01111100110010001", -- t[63889] = 40
      "0101000" when "01111100110010010", -- t[63890] = 40
      "0101000" when "01111100110010011", -- t[63891] = 40
      "0101000" when "01111100110010100", -- t[63892] = 40
      "0101000" when "01111100110010101", -- t[63893] = 40
      "0101000" when "01111100110010110", -- t[63894] = 40
      "0101000" when "01111100110010111", -- t[63895] = 40
      "0101000" when "01111100110011000", -- t[63896] = 40
      "0101000" when "01111100110011001", -- t[63897] = 40
      "0101000" when "01111100110011010", -- t[63898] = 40
      "0101000" when "01111100110011011", -- t[63899] = 40
      "0101000" when "01111100110011100", -- t[63900] = 40
      "0101000" when "01111100110011101", -- t[63901] = 40
      "0101000" when "01111100110011110", -- t[63902] = 40
      "0101000" when "01111100110011111", -- t[63903] = 40
      "0101000" when "01111100110100000", -- t[63904] = 40
      "0101000" when "01111100110100001", -- t[63905] = 40
      "0101000" when "01111100110100010", -- t[63906] = 40
      "0101000" when "01111100110100011", -- t[63907] = 40
      "0101000" when "01111100110100100", -- t[63908] = 40
      "0101000" when "01111100110100101", -- t[63909] = 40
      "0101000" when "01111100110100110", -- t[63910] = 40
      "0101000" when "01111100110100111", -- t[63911] = 40
      "0101000" when "01111100110101000", -- t[63912] = 40
      "0101000" when "01111100110101001", -- t[63913] = 40
      "0101000" when "01111100110101010", -- t[63914] = 40
      "0101000" when "01111100110101011", -- t[63915] = 40
      "0101000" when "01111100110101100", -- t[63916] = 40
      "0101000" when "01111100110101101", -- t[63917] = 40
      "0101000" when "01111100110101110", -- t[63918] = 40
      "0101000" when "01111100110101111", -- t[63919] = 40
      "0101000" when "01111100110110000", -- t[63920] = 40
      "0101000" when "01111100110110001", -- t[63921] = 40
      "0101000" when "01111100110110010", -- t[63922] = 40
      "0101000" when "01111100110110011", -- t[63923] = 40
      "0101000" when "01111100110110100", -- t[63924] = 40
      "0101000" when "01111100110110101", -- t[63925] = 40
      "0101000" when "01111100110110110", -- t[63926] = 40
      "0101000" when "01111100110110111", -- t[63927] = 40
      "0101000" when "01111100110111000", -- t[63928] = 40
      "0101000" when "01111100110111001", -- t[63929] = 40
      "0101000" when "01111100110111010", -- t[63930] = 40
      "0101000" when "01111100110111011", -- t[63931] = 40
      "0101000" when "01111100110111100", -- t[63932] = 40
      "0101000" when "01111100110111101", -- t[63933] = 40
      "0101000" when "01111100110111110", -- t[63934] = 40
      "0101000" when "01111100110111111", -- t[63935] = 40
      "0101000" when "01111100111000000", -- t[63936] = 40
      "0101000" when "01111100111000001", -- t[63937] = 40
      "0101000" when "01111100111000010", -- t[63938] = 40
      "0101000" when "01111100111000011", -- t[63939] = 40
      "0101000" when "01111100111000100", -- t[63940] = 40
      "0101000" when "01111100111000101", -- t[63941] = 40
      "0101000" when "01111100111000110", -- t[63942] = 40
      "0101000" when "01111100111000111", -- t[63943] = 40
      "0101000" when "01111100111001000", -- t[63944] = 40
      "0101000" when "01111100111001001", -- t[63945] = 40
      "0101000" when "01111100111001010", -- t[63946] = 40
      "0101000" when "01111100111001011", -- t[63947] = 40
      "0101000" when "01111100111001100", -- t[63948] = 40
      "0101000" when "01111100111001101", -- t[63949] = 40
      "0101000" when "01111100111001110", -- t[63950] = 40
      "0101000" when "01111100111001111", -- t[63951] = 40
      "0101000" when "01111100111010000", -- t[63952] = 40
      "0101000" when "01111100111010001", -- t[63953] = 40
      "0101000" when "01111100111010010", -- t[63954] = 40
      "0101000" when "01111100111010011", -- t[63955] = 40
      "0101000" when "01111100111010100", -- t[63956] = 40
      "0101000" when "01111100111010101", -- t[63957] = 40
      "0101000" when "01111100111010110", -- t[63958] = 40
      "0101000" when "01111100111010111", -- t[63959] = 40
      "0101000" when "01111100111011000", -- t[63960] = 40
      "0101000" when "01111100111011001", -- t[63961] = 40
      "0101000" when "01111100111011010", -- t[63962] = 40
      "0101000" when "01111100111011011", -- t[63963] = 40
      "0101000" when "01111100111011100", -- t[63964] = 40
      "0101000" when "01111100111011101", -- t[63965] = 40
      "0101000" when "01111100111011110", -- t[63966] = 40
      "0101000" when "01111100111011111", -- t[63967] = 40
      "0101000" when "01111100111100000", -- t[63968] = 40
      "0101001" when "01111100111100001", -- t[63969] = 41
      "0101001" when "01111100111100010", -- t[63970] = 41
      "0101001" when "01111100111100011", -- t[63971] = 41
      "0101001" when "01111100111100100", -- t[63972] = 41
      "0101001" when "01111100111100101", -- t[63973] = 41
      "0101001" when "01111100111100110", -- t[63974] = 41
      "0101001" when "01111100111100111", -- t[63975] = 41
      "0101001" when "01111100111101000", -- t[63976] = 41
      "0101001" when "01111100111101001", -- t[63977] = 41
      "0101001" when "01111100111101010", -- t[63978] = 41
      "0101001" when "01111100111101011", -- t[63979] = 41
      "0101001" when "01111100111101100", -- t[63980] = 41
      "0101001" when "01111100111101101", -- t[63981] = 41
      "0101001" when "01111100111101110", -- t[63982] = 41
      "0101001" when "01111100111101111", -- t[63983] = 41
      "0101001" when "01111100111110000", -- t[63984] = 41
      "0101001" when "01111100111110001", -- t[63985] = 41
      "0101001" when "01111100111110010", -- t[63986] = 41
      "0101001" when "01111100111110011", -- t[63987] = 41
      "0101001" when "01111100111110100", -- t[63988] = 41
      "0101001" when "01111100111110101", -- t[63989] = 41
      "0101001" when "01111100111110110", -- t[63990] = 41
      "0101001" when "01111100111110111", -- t[63991] = 41
      "0101001" when "01111100111111000", -- t[63992] = 41
      "0101001" when "01111100111111001", -- t[63993] = 41
      "0101001" when "01111100111111010", -- t[63994] = 41
      "0101001" when "01111100111111011", -- t[63995] = 41
      "0101001" when "01111100111111100", -- t[63996] = 41
      "0101001" when "01111100111111101", -- t[63997] = 41
      "0101001" when "01111100111111110", -- t[63998] = 41
      "0101001" when "01111100111111111", -- t[63999] = 41
      "0101001" when "01111101000000000", -- t[64000] = 41
      "0101001" when "01111101000000001", -- t[64001] = 41
      "0101001" when "01111101000000010", -- t[64002] = 41
      "0101001" when "01111101000000011", -- t[64003] = 41
      "0101001" when "01111101000000100", -- t[64004] = 41
      "0101001" when "01111101000000101", -- t[64005] = 41
      "0101001" when "01111101000000110", -- t[64006] = 41
      "0101001" when "01111101000000111", -- t[64007] = 41
      "0101001" when "01111101000001000", -- t[64008] = 41
      "0101001" when "01111101000001001", -- t[64009] = 41
      "0101001" when "01111101000001010", -- t[64010] = 41
      "0101001" when "01111101000001011", -- t[64011] = 41
      "0101001" when "01111101000001100", -- t[64012] = 41
      "0101001" when "01111101000001101", -- t[64013] = 41
      "0101001" when "01111101000001110", -- t[64014] = 41
      "0101001" when "01111101000001111", -- t[64015] = 41
      "0101001" when "01111101000010000", -- t[64016] = 41
      "0101001" when "01111101000010001", -- t[64017] = 41
      "0101001" when "01111101000010010", -- t[64018] = 41
      "0101001" when "01111101000010011", -- t[64019] = 41
      "0101001" when "01111101000010100", -- t[64020] = 41
      "0101001" when "01111101000010101", -- t[64021] = 41
      "0101001" when "01111101000010110", -- t[64022] = 41
      "0101001" when "01111101000010111", -- t[64023] = 41
      "0101001" when "01111101000011000", -- t[64024] = 41
      "0101001" when "01111101000011001", -- t[64025] = 41
      "0101001" when "01111101000011010", -- t[64026] = 41
      "0101001" when "01111101000011011", -- t[64027] = 41
      "0101001" when "01111101000011100", -- t[64028] = 41
      "0101001" when "01111101000011101", -- t[64029] = 41
      "0101001" when "01111101000011110", -- t[64030] = 41
      "0101001" when "01111101000011111", -- t[64031] = 41
      "0101001" when "01111101000100000", -- t[64032] = 41
      "0101001" when "01111101000100001", -- t[64033] = 41
      "0101001" when "01111101000100010", -- t[64034] = 41
      "0101001" when "01111101000100011", -- t[64035] = 41
      "0101001" when "01111101000100100", -- t[64036] = 41
      "0101001" when "01111101000100101", -- t[64037] = 41
      "0101001" when "01111101000100110", -- t[64038] = 41
      "0101001" when "01111101000100111", -- t[64039] = 41
      "0101001" when "01111101000101000", -- t[64040] = 41
      "0101001" when "01111101000101001", -- t[64041] = 41
      "0101001" when "01111101000101010", -- t[64042] = 41
      "0101001" when "01111101000101011", -- t[64043] = 41
      "0101001" when "01111101000101100", -- t[64044] = 41
      "0101001" when "01111101000101101", -- t[64045] = 41
      "0101001" when "01111101000101110", -- t[64046] = 41
      "0101001" when "01111101000101111", -- t[64047] = 41
      "0101001" when "01111101000110000", -- t[64048] = 41
      "0101001" when "01111101000110001", -- t[64049] = 41
      "0101001" when "01111101000110010", -- t[64050] = 41
      "0101001" when "01111101000110011", -- t[64051] = 41
      "0101001" when "01111101000110100", -- t[64052] = 41
      "0101001" when "01111101000110101", -- t[64053] = 41
      "0101001" when "01111101000110110", -- t[64054] = 41
      "0101001" when "01111101000110111", -- t[64055] = 41
      "0101001" when "01111101000111000", -- t[64056] = 41
      "0101001" when "01111101000111001", -- t[64057] = 41
      "0101001" when "01111101000111010", -- t[64058] = 41
      "0101001" when "01111101000111011", -- t[64059] = 41
      "0101001" when "01111101000111100", -- t[64060] = 41
      "0101001" when "01111101000111101", -- t[64061] = 41
      "0101001" when "01111101000111110", -- t[64062] = 41
      "0101001" when "01111101000111111", -- t[64063] = 41
      "0101001" when "01111101001000000", -- t[64064] = 41
      "0101001" when "01111101001000001", -- t[64065] = 41
      "0101001" when "01111101001000010", -- t[64066] = 41
      "0101001" when "01111101001000011", -- t[64067] = 41
      "0101001" when "01111101001000100", -- t[64068] = 41
      "0101001" when "01111101001000101", -- t[64069] = 41
      "0101001" when "01111101001000110", -- t[64070] = 41
      "0101001" when "01111101001000111", -- t[64071] = 41
      "0101001" when "01111101001001000", -- t[64072] = 41
      "0101001" when "01111101001001001", -- t[64073] = 41
      "0101001" when "01111101001001010", -- t[64074] = 41
      "0101001" when "01111101001001011", -- t[64075] = 41
      "0101001" when "01111101001001100", -- t[64076] = 41
      "0101001" when "01111101001001101", -- t[64077] = 41
      "0101001" when "01111101001001110", -- t[64078] = 41
      "0101001" when "01111101001001111", -- t[64079] = 41
      "0101001" when "01111101001010000", -- t[64080] = 41
      "0101001" when "01111101001010001", -- t[64081] = 41
      "0101001" when "01111101001010010", -- t[64082] = 41
      "0101001" when "01111101001010011", -- t[64083] = 41
      "0101001" when "01111101001010100", -- t[64084] = 41
      "0101001" when "01111101001010101", -- t[64085] = 41
      "0101001" when "01111101001010110", -- t[64086] = 41
      "0101001" when "01111101001010111", -- t[64087] = 41
      "0101001" when "01111101001011000", -- t[64088] = 41
      "0101001" when "01111101001011001", -- t[64089] = 41
      "0101001" when "01111101001011010", -- t[64090] = 41
      "0101001" when "01111101001011011", -- t[64091] = 41
      "0101001" when "01111101001011100", -- t[64092] = 41
      "0101001" when "01111101001011101", -- t[64093] = 41
      "0101001" when "01111101001011110", -- t[64094] = 41
      "0101001" when "01111101001011111", -- t[64095] = 41
      "0101001" when "01111101001100000", -- t[64096] = 41
      "0101001" when "01111101001100001", -- t[64097] = 41
      "0101001" when "01111101001100010", -- t[64098] = 41
      "0101001" when "01111101001100011", -- t[64099] = 41
      "0101001" when "01111101001100100", -- t[64100] = 41
      "0101001" when "01111101001100101", -- t[64101] = 41
      "0101001" when "01111101001100110", -- t[64102] = 41
      "0101001" when "01111101001100111", -- t[64103] = 41
      "0101001" when "01111101001101000", -- t[64104] = 41
      "0101001" when "01111101001101001", -- t[64105] = 41
      "0101001" when "01111101001101010", -- t[64106] = 41
      "0101001" when "01111101001101011", -- t[64107] = 41
      "0101001" when "01111101001101100", -- t[64108] = 41
      "0101001" when "01111101001101101", -- t[64109] = 41
      "0101001" when "01111101001101110", -- t[64110] = 41
      "0101001" when "01111101001101111", -- t[64111] = 41
      "0101001" when "01111101001110000", -- t[64112] = 41
      "0101001" when "01111101001110001", -- t[64113] = 41
      "0101001" when "01111101001110010", -- t[64114] = 41
      "0101001" when "01111101001110011", -- t[64115] = 41
      "0101001" when "01111101001110100", -- t[64116] = 41
      "0101001" when "01111101001110101", -- t[64117] = 41
      "0101001" when "01111101001110110", -- t[64118] = 41
      "0101001" when "01111101001110111", -- t[64119] = 41
      "0101001" when "01111101001111000", -- t[64120] = 41
      "0101001" when "01111101001111001", -- t[64121] = 41
      "0101001" when "01111101001111010", -- t[64122] = 41
      "0101001" when "01111101001111011", -- t[64123] = 41
      "0101001" when "01111101001111100", -- t[64124] = 41
      "0101001" when "01111101001111101", -- t[64125] = 41
      "0101001" when "01111101001111110", -- t[64126] = 41
      "0101001" when "01111101001111111", -- t[64127] = 41
      "0101001" when "01111101010000000", -- t[64128] = 41
      "0101001" when "01111101010000001", -- t[64129] = 41
      "0101001" when "01111101010000010", -- t[64130] = 41
      "0101001" when "01111101010000011", -- t[64131] = 41
      "0101001" when "01111101010000100", -- t[64132] = 41
      "0101001" when "01111101010000101", -- t[64133] = 41
      "0101001" when "01111101010000110", -- t[64134] = 41
      "0101001" when "01111101010000111", -- t[64135] = 41
      "0101001" when "01111101010001000", -- t[64136] = 41
      "0101001" when "01111101010001001", -- t[64137] = 41
      "0101001" when "01111101010001010", -- t[64138] = 41
      "0101001" when "01111101010001011", -- t[64139] = 41
      "0101001" when "01111101010001100", -- t[64140] = 41
      "0101001" when "01111101010001101", -- t[64141] = 41
      "0101001" when "01111101010001110", -- t[64142] = 41
      "0101001" when "01111101010001111", -- t[64143] = 41
      "0101001" when "01111101010010000", -- t[64144] = 41
      "0101001" when "01111101010010001", -- t[64145] = 41
      "0101001" when "01111101010010010", -- t[64146] = 41
      "0101001" when "01111101010010011", -- t[64147] = 41
      "0101001" when "01111101010010100", -- t[64148] = 41
      "0101001" when "01111101010010101", -- t[64149] = 41
      "0101001" when "01111101010010110", -- t[64150] = 41
      "0101001" when "01111101010010111", -- t[64151] = 41
      "0101001" when "01111101010011000", -- t[64152] = 41
      "0101001" when "01111101010011001", -- t[64153] = 41
      "0101001" when "01111101010011010", -- t[64154] = 41
      "0101001" when "01111101010011011", -- t[64155] = 41
      "0101001" when "01111101010011100", -- t[64156] = 41
      "0101001" when "01111101010011101", -- t[64157] = 41
      "0101001" when "01111101010011110", -- t[64158] = 41
      "0101001" when "01111101010011111", -- t[64159] = 41
      "0101001" when "01111101010100000", -- t[64160] = 41
      "0101001" when "01111101010100001", -- t[64161] = 41
      "0101001" when "01111101010100010", -- t[64162] = 41
      "0101001" when "01111101010100011", -- t[64163] = 41
      "0101001" when "01111101010100100", -- t[64164] = 41
      "0101001" when "01111101010100101", -- t[64165] = 41
      "0101001" when "01111101010100110", -- t[64166] = 41
      "0101001" when "01111101010100111", -- t[64167] = 41
      "0101001" when "01111101010101000", -- t[64168] = 41
      "0101001" when "01111101010101001", -- t[64169] = 41
      "0101001" when "01111101010101010", -- t[64170] = 41
      "0101001" when "01111101010101011", -- t[64171] = 41
      "0101001" when "01111101010101100", -- t[64172] = 41
      "0101001" when "01111101010101101", -- t[64173] = 41
      "0101001" when "01111101010101110", -- t[64174] = 41
      "0101001" when "01111101010101111", -- t[64175] = 41
      "0101001" when "01111101010110000", -- t[64176] = 41
      "0101001" when "01111101010110001", -- t[64177] = 41
      "0101001" when "01111101010110010", -- t[64178] = 41
      "0101001" when "01111101010110011", -- t[64179] = 41
      "0101001" when "01111101010110100", -- t[64180] = 41
      "0101001" when "01111101010110101", -- t[64181] = 41
      "0101001" when "01111101010110110", -- t[64182] = 41
      "0101001" when "01111101010110111", -- t[64183] = 41
      "0101001" when "01111101010111000", -- t[64184] = 41
      "0101001" when "01111101010111001", -- t[64185] = 41
      "0101001" when "01111101010111010", -- t[64186] = 41
      "0101001" when "01111101010111011", -- t[64187] = 41
      "0101001" when "01111101010111100", -- t[64188] = 41
      "0101001" when "01111101010111101", -- t[64189] = 41
      "0101001" when "01111101010111110", -- t[64190] = 41
      "0101001" when "01111101010111111", -- t[64191] = 41
      "0101001" when "01111101011000000", -- t[64192] = 41
      "0101001" when "01111101011000001", -- t[64193] = 41
      "0101001" when "01111101011000010", -- t[64194] = 41
      "0101001" when "01111101011000011", -- t[64195] = 41
      "0101001" when "01111101011000100", -- t[64196] = 41
      "0101001" when "01111101011000101", -- t[64197] = 41
      "0101001" when "01111101011000110", -- t[64198] = 41
      "0101001" when "01111101011000111", -- t[64199] = 41
      "0101001" when "01111101011001000", -- t[64200] = 41
      "0101001" when "01111101011001001", -- t[64201] = 41
      "0101001" when "01111101011001010", -- t[64202] = 41
      "0101001" when "01111101011001011", -- t[64203] = 41
      "0101001" when "01111101011001100", -- t[64204] = 41
      "0101001" when "01111101011001101", -- t[64205] = 41
      "0101001" when "01111101011001110", -- t[64206] = 41
      "0101001" when "01111101011001111", -- t[64207] = 41
      "0101001" when "01111101011010000", -- t[64208] = 41
      "0101001" when "01111101011010001", -- t[64209] = 41
      "0101001" when "01111101011010010", -- t[64210] = 41
      "0101001" when "01111101011010011", -- t[64211] = 41
      "0101001" when "01111101011010100", -- t[64212] = 41
      "0101001" when "01111101011010101", -- t[64213] = 41
      "0101001" when "01111101011010110", -- t[64214] = 41
      "0101001" when "01111101011010111", -- t[64215] = 41
      "0101001" when "01111101011011000", -- t[64216] = 41
      "0101001" when "01111101011011001", -- t[64217] = 41
      "0101001" when "01111101011011010", -- t[64218] = 41
      "0101001" when "01111101011011011", -- t[64219] = 41
      "0101001" when "01111101011011100", -- t[64220] = 41
      "0101001" when "01111101011011101", -- t[64221] = 41
      "0101001" when "01111101011011110", -- t[64222] = 41
      "0101001" when "01111101011011111", -- t[64223] = 41
      "0101001" when "01111101011100000", -- t[64224] = 41
      "0101001" when "01111101011100001", -- t[64225] = 41
      "0101001" when "01111101011100010", -- t[64226] = 41
      "0101001" when "01111101011100011", -- t[64227] = 41
      "0101001" when "01111101011100100", -- t[64228] = 41
      "0101001" when "01111101011100101", -- t[64229] = 41
      "0101001" when "01111101011100110", -- t[64230] = 41
      "0101001" when "01111101011100111", -- t[64231] = 41
      "0101001" when "01111101011101000", -- t[64232] = 41
      "0101001" when "01111101011101001", -- t[64233] = 41
      "0101001" when "01111101011101010", -- t[64234] = 41
      "0101001" when "01111101011101011", -- t[64235] = 41
      "0101001" when "01111101011101100", -- t[64236] = 41
      "0101001" when "01111101011101101", -- t[64237] = 41
      "0101001" when "01111101011101110", -- t[64238] = 41
      "0101001" when "01111101011101111", -- t[64239] = 41
      "0101001" when "01111101011110000", -- t[64240] = 41
      "0101001" when "01111101011110001", -- t[64241] = 41
      "0101001" when "01111101011110010", -- t[64242] = 41
      "0101001" when "01111101011110011", -- t[64243] = 41
      "0101001" when "01111101011110100", -- t[64244] = 41
      "0101001" when "01111101011110101", -- t[64245] = 41
      "0101001" when "01111101011110110", -- t[64246] = 41
      "0101001" when "01111101011110111", -- t[64247] = 41
      "0101001" when "01111101011111000", -- t[64248] = 41
      "0101001" when "01111101011111001", -- t[64249] = 41
      "0101001" when "01111101011111010", -- t[64250] = 41
      "0101001" when "01111101011111011", -- t[64251] = 41
      "0101001" when "01111101011111100", -- t[64252] = 41
      "0101001" when "01111101011111101", -- t[64253] = 41
      "0101001" when "01111101011111110", -- t[64254] = 41
      "0101001" when "01111101011111111", -- t[64255] = 41
      "0101010" when "01111101100000000", -- t[64256] = 42
      "0101010" when "01111101100000001", -- t[64257] = 42
      "0101010" when "01111101100000010", -- t[64258] = 42
      "0101010" when "01111101100000011", -- t[64259] = 42
      "0101010" when "01111101100000100", -- t[64260] = 42
      "0101010" when "01111101100000101", -- t[64261] = 42
      "0101010" when "01111101100000110", -- t[64262] = 42
      "0101010" when "01111101100000111", -- t[64263] = 42
      "0101010" when "01111101100001000", -- t[64264] = 42
      "0101010" when "01111101100001001", -- t[64265] = 42
      "0101010" when "01111101100001010", -- t[64266] = 42
      "0101010" when "01111101100001011", -- t[64267] = 42
      "0101010" when "01111101100001100", -- t[64268] = 42
      "0101010" when "01111101100001101", -- t[64269] = 42
      "0101010" when "01111101100001110", -- t[64270] = 42
      "0101010" when "01111101100001111", -- t[64271] = 42
      "0101010" when "01111101100010000", -- t[64272] = 42
      "0101010" when "01111101100010001", -- t[64273] = 42
      "0101010" when "01111101100010010", -- t[64274] = 42
      "0101010" when "01111101100010011", -- t[64275] = 42
      "0101010" when "01111101100010100", -- t[64276] = 42
      "0101010" when "01111101100010101", -- t[64277] = 42
      "0101010" when "01111101100010110", -- t[64278] = 42
      "0101010" when "01111101100010111", -- t[64279] = 42
      "0101010" when "01111101100011000", -- t[64280] = 42
      "0101010" when "01111101100011001", -- t[64281] = 42
      "0101010" when "01111101100011010", -- t[64282] = 42
      "0101010" when "01111101100011011", -- t[64283] = 42
      "0101010" when "01111101100011100", -- t[64284] = 42
      "0101010" when "01111101100011101", -- t[64285] = 42
      "0101010" when "01111101100011110", -- t[64286] = 42
      "0101010" when "01111101100011111", -- t[64287] = 42
      "0101010" when "01111101100100000", -- t[64288] = 42
      "0101010" when "01111101100100001", -- t[64289] = 42
      "0101010" when "01111101100100010", -- t[64290] = 42
      "0101010" when "01111101100100011", -- t[64291] = 42
      "0101010" when "01111101100100100", -- t[64292] = 42
      "0101010" when "01111101100100101", -- t[64293] = 42
      "0101010" when "01111101100100110", -- t[64294] = 42
      "0101010" when "01111101100100111", -- t[64295] = 42
      "0101010" when "01111101100101000", -- t[64296] = 42
      "0101010" when "01111101100101001", -- t[64297] = 42
      "0101010" when "01111101100101010", -- t[64298] = 42
      "0101010" when "01111101100101011", -- t[64299] = 42
      "0101010" when "01111101100101100", -- t[64300] = 42
      "0101010" when "01111101100101101", -- t[64301] = 42
      "0101010" when "01111101100101110", -- t[64302] = 42
      "0101010" when "01111101100101111", -- t[64303] = 42
      "0101010" when "01111101100110000", -- t[64304] = 42
      "0101010" when "01111101100110001", -- t[64305] = 42
      "0101010" when "01111101100110010", -- t[64306] = 42
      "0101010" when "01111101100110011", -- t[64307] = 42
      "0101010" when "01111101100110100", -- t[64308] = 42
      "0101010" when "01111101100110101", -- t[64309] = 42
      "0101010" when "01111101100110110", -- t[64310] = 42
      "0101010" when "01111101100110111", -- t[64311] = 42
      "0101010" when "01111101100111000", -- t[64312] = 42
      "0101010" when "01111101100111001", -- t[64313] = 42
      "0101010" when "01111101100111010", -- t[64314] = 42
      "0101010" when "01111101100111011", -- t[64315] = 42
      "0101010" when "01111101100111100", -- t[64316] = 42
      "0101010" when "01111101100111101", -- t[64317] = 42
      "0101010" when "01111101100111110", -- t[64318] = 42
      "0101010" when "01111101100111111", -- t[64319] = 42
      "0101010" when "01111101101000000", -- t[64320] = 42
      "0101010" when "01111101101000001", -- t[64321] = 42
      "0101010" when "01111101101000010", -- t[64322] = 42
      "0101010" when "01111101101000011", -- t[64323] = 42
      "0101010" when "01111101101000100", -- t[64324] = 42
      "0101010" when "01111101101000101", -- t[64325] = 42
      "0101010" when "01111101101000110", -- t[64326] = 42
      "0101010" when "01111101101000111", -- t[64327] = 42
      "0101010" when "01111101101001000", -- t[64328] = 42
      "0101010" when "01111101101001001", -- t[64329] = 42
      "0101010" when "01111101101001010", -- t[64330] = 42
      "0101010" when "01111101101001011", -- t[64331] = 42
      "0101010" when "01111101101001100", -- t[64332] = 42
      "0101010" when "01111101101001101", -- t[64333] = 42
      "0101010" when "01111101101001110", -- t[64334] = 42
      "0101010" when "01111101101001111", -- t[64335] = 42
      "0101010" when "01111101101010000", -- t[64336] = 42
      "0101010" when "01111101101010001", -- t[64337] = 42
      "0101010" when "01111101101010010", -- t[64338] = 42
      "0101010" when "01111101101010011", -- t[64339] = 42
      "0101010" when "01111101101010100", -- t[64340] = 42
      "0101010" when "01111101101010101", -- t[64341] = 42
      "0101010" when "01111101101010110", -- t[64342] = 42
      "0101010" when "01111101101010111", -- t[64343] = 42
      "0101010" when "01111101101011000", -- t[64344] = 42
      "0101010" when "01111101101011001", -- t[64345] = 42
      "0101010" when "01111101101011010", -- t[64346] = 42
      "0101010" when "01111101101011011", -- t[64347] = 42
      "0101010" when "01111101101011100", -- t[64348] = 42
      "0101010" when "01111101101011101", -- t[64349] = 42
      "0101010" when "01111101101011110", -- t[64350] = 42
      "0101010" when "01111101101011111", -- t[64351] = 42
      "0101010" when "01111101101100000", -- t[64352] = 42
      "0101010" when "01111101101100001", -- t[64353] = 42
      "0101010" when "01111101101100010", -- t[64354] = 42
      "0101010" when "01111101101100011", -- t[64355] = 42
      "0101010" when "01111101101100100", -- t[64356] = 42
      "0101010" when "01111101101100101", -- t[64357] = 42
      "0101010" when "01111101101100110", -- t[64358] = 42
      "0101010" when "01111101101100111", -- t[64359] = 42
      "0101010" when "01111101101101000", -- t[64360] = 42
      "0101010" when "01111101101101001", -- t[64361] = 42
      "0101010" when "01111101101101010", -- t[64362] = 42
      "0101010" when "01111101101101011", -- t[64363] = 42
      "0101010" when "01111101101101100", -- t[64364] = 42
      "0101010" when "01111101101101101", -- t[64365] = 42
      "0101010" when "01111101101101110", -- t[64366] = 42
      "0101010" when "01111101101101111", -- t[64367] = 42
      "0101010" when "01111101101110000", -- t[64368] = 42
      "0101010" when "01111101101110001", -- t[64369] = 42
      "0101010" when "01111101101110010", -- t[64370] = 42
      "0101010" when "01111101101110011", -- t[64371] = 42
      "0101010" when "01111101101110100", -- t[64372] = 42
      "0101010" when "01111101101110101", -- t[64373] = 42
      "0101010" when "01111101101110110", -- t[64374] = 42
      "0101010" when "01111101101110111", -- t[64375] = 42
      "0101010" when "01111101101111000", -- t[64376] = 42
      "0101010" when "01111101101111001", -- t[64377] = 42
      "0101010" when "01111101101111010", -- t[64378] = 42
      "0101010" when "01111101101111011", -- t[64379] = 42
      "0101010" when "01111101101111100", -- t[64380] = 42
      "0101010" when "01111101101111101", -- t[64381] = 42
      "0101010" when "01111101101111110", -- t[64382] = 42
      "0101010" when "01111101101111111", -- t[64383] = 42
      "0101010" when "01111101110000000", -- t[64384] = 42
      "0101010" when "01111101110000001", -- t[64385] = 42
      "0101010" when "01111101110000010", -- t[64386] = 42
      "0101010" when "01111101110000011", -- t[64387] = 42
      "0101010" when "01111101110000100", -- t[64388] = 42
      "0101010" when "01111101110000101", -- t[64389] = 42
      "0101010" when "01111101110000110", -- t[64390] = 42
      "0101010" when "01111101110000111", -- t[64391] = 42
      "0101010" when "01111101110001000", -- t[64392] = 42
      "0101010" when "01111101110001001", -- t[64393] = 42
      "0101010" when "01111101110001010", -- t[64394] = 42
      "0101010" when "01111101110001011", -- t[64395] = 42
      "0101010" when "01111101110001100", -- t[64396] = 42
      "0101010" when "01111101110001101", -- t[64397] = 42
      "0101010" when "01111101110001110", -- t[64398] = 42
      "0101010" when "01111101110001111", -- t[64399] = 42
      "0101010" when "01111101110010000", -- t[64400] = 42
      "0101010" when "01111101110010001", -- t[64401] = 42
      "0101010" when "01111101110010010", -- t[64402] = 42
      "0101010" when "01111101110010011", -- t[64403] = 42
      "0101010" when "01111101110010100", -- t[64404] = 42
      "0101010" when "01111101110010101", -- t[64405] = 42
      "0101010" when "01111101110010110", -- t[64406] = 42
      "0101010" when "01111101110010111", -- t[64407] = 42
      "0101010" when "01111101110011000", -- t[64408] = 42
      "0101010" when "01111101110011001", -- t[64409] = 42
      "0101010" when "01111101110011010", -- t[64410] = 42
      "0101010" when "01111101110011011", -- t[64411] = 42
      "0101010" when "01111101110011100", -- t[64412] = 42
      "0101010" when "01111101110011101", -- t[64413] = 42
      "0101010" when "01111101110011110", -- t[64414] = 42
      "0101010" when "01111101110011111", -- t[64415] = 42
      "0101010" when "01111101110100000", -- t[64416] = 42
      "0101010" when "01111101110100001", -- t[64417] = 42
      "0101010" when "01111101110100010", -- t[64418] = 42
      "0101010" when "01111101110100011", -- t[64419] = 42
      "0101010" when "01111101110100100", -- t[64420] = 42
      "0101010" when "01111101110100101", -- t[64421] = 42
      "0101010" when "01111101110100110", -- t[64422] = 42
      "0101010" when "01111101110100111", -- t[64423] = 42
      "0101010" when "01111101110101000", -- t[64424] = 42
      "0101010" when "01111101110101001", -- t[64425] = 42
      "0101010" when "01111101110101010", -- t[64426] = 42
      "0101010" when "01111101110101011", -- t[64427] = 42
      "0101010" when "01111101110101100", -- t[64428] = 42
      "0101010" when "01111101110101101", -- t[64429] = 42
      "0101010" when "01111101110101110", -- t[64430] = 42
      "0101010" when "01111101110101111", -- t[64431] = 42
      "0101010" when "01111101110110000", -- t[64432] = 42
      "0101010" when "01111101110110001", -- t[64433] = 42
      "0101010" when "01111101110110010", -- t[64434] = 42
      "0101010" when "01111101110110011", -- t[64435] = 42
      "0101010" when "01111101110110100", -- t[64436] = 42
      "0101010" when "01111101110110101", -- t[64437] = 42
      "0101010" when "01111101110110110", -- t[64438] = 42
      "0101010" when "01111101110110111", -- t[64439] = 42
      "0101010" when "01111101110111000", -- t[64440] = 42
      "0101010" when "01111101110111001", -- t[64441] = 42
      "0101010" when "01111101110111010", -- t[64442] = 42
      "0101010" when "01111101110111011", -- t[64443] = 42
      "0101010" when "01111101110111100", -- t[64444] = 42
      "0101010" when "01111101110111101", -- t[64445] = 42
      "0101010" when "01111101110111110", -- t[64446] = 42
      "0101010" when "01111101110111111", -- t[64447] = 42
      "0101010" when "01111101111000000", -- t[64448] = 42
      "0101010" when "01111101111000001", -- t[64449] = 42
      "0101010" when "01111101111000010", -- t[64450] = 42
      "0101010" when "01111101111000011", -- t[64451] = 42
      "0101010" when "01111101111000100", -- t[64452] = 42
      "0101010" when "01111101111000101", -- t[64453] = 42
      "0101010" when "01111101111000110", -- t[64454] = 42
      "0101010" when "01111101111000111", -- t[64455] = 42
      "0101010" when "01111101111001000", -- t[64456] = 42
      "0101010" when "01111101111001001", -- t[64457] = 42
      "0101010" when "01111101111001010", -- t[64458] = 42
      "0101010" when "01111101111001011", -- t[64459] = 42
      "0101010" when "01111101111001100", -- t[64460] = 42
      "0101010" when "01111101111001101", -- t[64461] = 42
      "0101010" when "01111101111001110", -- t[64462] = 42
      "0101010" when "01111101111001111", -- t[64463] = 42
      "0101010" when "01111101111010000", -- t[64464] = 42
      "0101010" when "01111101111010001", -- t[64465] = 42
      "0101010" when "01111101111010010", -- t[64466] = 42
      "0101010" when "01111101111010011", -- t[64467] = 42
      "0101010" when "01111101111010100", -- t[64468] = 42
      "0101010" when "01111101111010101", -- t[64469] = 42
      "0101010" when "01111101111010110", -- t[64470] = 42
      "0101010" when "01111101111010111", -- t[64471] = 42
      "0101010" when "01111101111011000", -- t[64472] = 42
      "0101010" when "01111101111011001", -- t[64473] = 42
      "0101010" when "01111101111011010", -- t[64474] = 42
      "0101010" when "01111101111011011", -- t[64475] = 42
      "0101010" when "01111101111011100", -- t[64476] = 42
      "0101010" when "01111101111011101", -- t[64477] = 42
      "0101010" when "01111101111011110", -- t[64478] = 42
      "0101010" when "01111101111011111", -- t[64479] = 42
      "0101010" when "01111101111100000", -- t[64480] = 42
      "0101010" when "01111101111100001", -- t[64481] = 42
      "0101010" when "01111101111100010", -- t[64482] = 42
      "0101010" when "01111101111100011", -- t[64483] = 42
      "0101010" when "01111101111100100", -- t[64484] = 42
      "0101010" when "01111101111100101", -- t[64485] = 42
      "0101010" when "01111101111100110", -- t[64486] = 42
      "0101010" when "01111101111100111", -- t[64487] = 42
      "0101010" when "01111101111101000", -- t[64488] = 42
      "0101010" when "01111101111101001", -- t[64489] = 42
      "0101010" when "01111101111101010", -- t[64490] = 42
      "0101010" when "01111101111101011", -- t[64491] = 42
      "0101010" when "01111101111101100", -- t[64492] = 42
      "0101010" when "01111101111101101", -- t[64493] = 42
      "0101010" when "01111101111101110", -- t[64494] = 42
      "0101010" when "01111101111101111", -- t[64495] = 42
      "0101010" when "01111101111110000", -- t[64496] = 42
      "0101010" when "01111101111110001", -- t[64497] = 42
      "0101010" when "01111101111110010", -- t[64498] = 42
      "0101010" when "01111101111110011", -- t[64499] = 42
      "0101010" when "01111101111110100", -- t[64500] = 42
      "0101010" when "01111101111110101", -- t[64501] = 42
      "0101010" when "01111101111110110", -- t[64502] = 42
      "0101010" when "01111101111110111", -- t[64503] = 42
      "0101010" when "01111101111111000", -- t[64504] = 42
      "0101010" when "01111101111111001", -- t[64505] = 42
      "0101010" when "01111101111111010", -- t[64506] = 42
      "0101010" when "01111101111111011", -- t[64507] = 42
      "0101010" when "01111101111111100", -- t[64508] = 42
      "0101010" when "01111101111111101", -- t[64509] = 42
      "0101010" when "01111101111111110", -- t[64510] = 42
      "0101010" when "01111101111111111", -- t[64511] = 42
      "0101010" when "01111110000000000", -- t[64512] = 42
      "0101010" when "01111110000000001", -- t[64513] = 42
      "0101010" when "01111110000000010", -- t[64514] = 42
      "0101010" when "01111110000000011", -- t[64515] = 42
      "0101010" when "01111110000000100", -- t[64516] = 42
      "0101010" when "01111110000000101", -- t[64517] = 42
      "0101010" when "01111110000000110", -- t[64518] = 42
      "0101010" when "01111110000000111", -- t[64519] = 42
      "0101010" when "01111110000001000", -- t[64520] = 42
      "0101010" when "01111110000001001", -- t[64521] = 42
      "0101010" when "01111110000001010", -- t[64522] = 42
      "0101010" when "01111110000001011", -- t[64523] = 42
      "0101010" when "01111110000001100", -- t[64524] = 42
      "0101010" when "01111110000001101", -- t[64525] = 42
      "0101010" when "01111110000001110", -- t[64526] = 42
      "0101010" when "01111110000001111", -- t[64527] = 42
      "0101010" when "01111110000010000", -- t[64528] = 42
      "0101010" when "01111110000010001", -- t[64529] = 42
      "0101010" when "01111110000010010", -- t[64530] = 42
      "0101010" when "01111110000010011", -- t[64531] = 42
      "0101010" when "01111110000010100", -- t[64532] = 42
      "0101010" when "01111110000010101", -- t[64533] = 42
      "0101010" when "01111110000010110", -- t[64534] = 42
      "0101010" when "01111110000010111", -- t[64535] = 42
      "0101010" when "01111110000011000", -- t[64536] = 42
      "0101011" when "01111110000011001", -- t[64537] = 43
      "0101011" when "01111110000011010", -- t[64538] = 43
      "0101011" when "01111110000011011", -- t[64539] = 43
      "0101011" when "01111110000011100", -- t[64540] = 43
      "0101011" when "01111110000011101", -- t[64541] = 43
      "0101011" when "01111110000011110", -- t[64542] = 43
      "0101011" when "01111110000011111", -- t[64543] = 43
      "0101011" when "01111110000100000", -- t[64544] = 43
      "0101011" when "01111110000100001", -- t[64545] = 43
      "0101011" when "01111110000100010", -- t[64546] = 43
      "0101011" when "01111110000100011", -- t[64547] = 43
      "0101011" when "01111110000100100", -- t[64548] = 43
      "0101011" when "01111110000100101", -- t[64549] = 43
      "0101011" when "01111110000100110", -- t[64550] = 43
      "0101011" when "01111110000100111", -- t[64551] = 43
      "0101011" when "01111110000101000", -- t[64552] = 43
      "0101011" when "01111110000101001", -- t[64553] = 43
      "0101011" when "01111110000101010", -- t[64554] = 43
      "0101011" when "01111110000101011", -- t[64555] = 43
      "0101011" when "01111110000101100", -- t[64556] = 43
      "0101011" when "01111110000101101", -- t[64557] = 43
      "0101011" when "01111110000101110", -- t[64558] = 43
      "0101011" when "01111110000101111", -- t[64559] = 43
      "0101011" when "01111110000110000", -- t[64560] = 43
      "0101011" when "01111110000110001", -- t[64561] = 43
      "0101011" when "01111110000110010", -- t[64562] = 43
      "0101011" when "01111110000110011", -- t[64563] = 43
      "0101011" when "01111110000110100", -- t[64564] = 43
      "0101011" when "01111110000110101", -- t[64565] = 43
      "0101011" when "01111110000110110", -- t[64566] = 43
      "0101011" when "01111110000110111", -- t[64567] = 43
      "0101011" when "01111110000111000", -- t[64568] = 43
      "0101011" when "01111110000111001", -- t[64569] = 43
      "0101011" when "01111110000111010", -- t[64570] = 43
      "0101011" when "01111110000111011", -- t[64571] = 43
      "0101011" when "01111110000111100", -- t[64572] = 43
      "0101011" when "01111110000111101", -- t[64573] = 43
      "0101011" when "01111110000111110", -- t[64574] = 43
      "0101011" when "01111110000111111", -- t[64575] = 43
      "0101011" when "01111110001000000", -- t[64576] = 43
      "0101011" when "01111110001000001", -- t[64577] = 43
      "0101011" when "01111110001000010", -- t[64578] = 43
      "0101011" when "01111110001000011", -- t[64579] = 43
      "0101011" when "01111110001000100", -- t[64580] = 43
      "0101011" when "01111110001000101", -- t[64581] = 43
      "0101011" when "01111110001000110", -- t[64582] = 43
      "0101011" when "01111110001000111", -- t[64583] = 43
      "0101011" when "01111110001001000", -- t[64584] = 43
      "0101011" when "01111110001001001", -- t[64585] = 43
      "0101011" when "01111110001001010", -- t[64586] = 43
      "0101011" when "01111110001001011", -- t[64587] = 43
      "0101011" when "01111110001001100", -- t[64588] = 43
      "0101011" when "01111110001001101", -- t[64589] = 43
      "0101011" when "01111110001001110", -- t[64590] = 43
      "0101011" when "01111110001001111", -- t[64591] = 43
      "0101011" when "01111110001010000", -- t[64592] = 43
      "0101011" when "01111110001010001", -- t[64593] = 43
      "0101011" when "01111110001010010", -- t[64594] = 43
      "0101011" when "01111110001010011", -- t[64595] = 43
      "0101011" when "01111110001010100", -- t[64596] = 43
      "0101011" when "01111110001010101", -- t[64597] = 43
      "0101011" when "01111110001010110", -- t[64598] = 43
      "0101011" when "01111110001010111", -- t[64599] = 43
      "0101011" when "01111110001011000", -- t[64600] = 43
      "0101011" when "01111110001011001", -- t[64601] = 43
      "0101011" when "01111110001011010", -- t[64602] = 43
      "0101011" when "01111110001011011", -- t[64603] = 43
      "0101011" when "01111110001011100", -- t[64604] = 43
      "0101011" when "01111110001011101", -- t[64605] = 43
      "0101011" when "01111110001011110", -- t[64606] = 43
      "0101011" when "01111110001011111", -- t[64607] = 43
      "0101011" when "01111110001100000", -- t[64608] = 43
      "0101011" when "01111110001100001", -- t[64609] = 43
      "0101011" when "01111110001100010", -- t[64610] = 43
      "0101011" when "01111110001100011", -- t[64611] = 43
      "0101011" when "01111110001100100", -- t[64612] = 43
      "0101011" when "01111110001100101", -- t[64613] = 43
      "0101011" when "01111110001100110", -- t[64614] = 43
      "0101011" when "01111110001100111", -- t[64615] = 43
      "0101011" when "01111110001101000", -- t[64616] = 43
      "0101011" when "01111110001101001", -- t[64617] = 43
      "0101011" when "01111110001101010", -- t[64618] = 43
      "0101011" when "01111110001101011", -- t[64619] = 43
      "0101011" when "01111110001101100", -- t[64620] = 43
      "0101011" when "01111110001101101", -- t[64621] = 43
      "0101011" when "01111110001101110", -- t[64622] = 43
      "0101011" when "01111110001101111", -- t[64623] = 43
      "0101011" when "01111110001110000", -- t[64624] = 43
      "0101011" when "01111110001110001", -- t[64625] = 43
      "0101011" when "01111110001110010", -- t[64626] = 43
      "0101011" when "01111110001110011", -- t[64627] = 43
      "0101011" when "01111110001110100", -- t[64628] = 43
      "0101011" when "01111110001110101", -- t[64629] = 43
      "0101011" when "01111110001110110", -- t[64630] = 43
      "0101011" when "01111110001110111", -- t[64631] = 43
      "0101011" when "01111110001111000", -- t[64632] = 43
      "0101011" when "01111110001111001", -- t[64633] = 43
      "0101011" when "01111110001111010", -- t[64634] = 43
      "0101011" when "01111110001111011", -- t[64635] = 43
      "0101011" when "01111110001111100", -- t[64636] = 43
      "0101011" when "01111110001111101", -- t[64637] = 43
      "0101011" when "01111110001111110", -- t[64638] = 43
      "0101011" when "01111110001111111", -- t[64639] = 43
      "0101011" when "01111110010000000", -- t[64640] = 43
      "0101011" when "01111110010000001", -- t[64641] = 43
      "0101011" when "01111110010000010", -- t[64642] = 43
      "0101011" when "01111110010000011", -- t[64643] = 43
      "0101011" when "01111110010000100", -- t[64644] = 43
      "0101011" when "01111110010000101", -- t[64645] = 43
      "0101011" when "01111110010000110", -- t[64646] = 43
      "0101011" when "01111110010000111", -- t[64647] = 43
      "0101011" when "01111110010001000", -- t[64648] = 43
      "0101011" when "01111110010001001", -- t[64649] = 43
      "0101011" when "01111110010001010", -- t[64650] = 43
      "0101011" when "01111110010001011", -- t[64651] = 43
      "0101011" when "01111110010001100", -- t[64652] = 43
      "0101011" when "01111110010001101", -- t[64653] = 43
      "0101011" when "01111110010001110", -- t[64654] = 43
      "0101011" when "01111110010001111", -- t[64655] = 43
      "0101011" when "01111110010010000", -- t[64656] = 43
      "0101011" when "01111110010010001", -- t[64657] = 43
      "0101011" when "01111110010010010", -- t[64658] = 43
      "0101011" when "01111110010010011", -- t[64659] = 43
      "0101011" when "01111110010010100", -- t[64660] = 43
      "0101011" when "01111110010010101", -- t[64661] = 43
      "0101011" when "01111110010010110", -- t[64662] = 43
      "0101011" when "01111110010010111", -- t[64663] = 43
      "0101011" when "01111110010011000", -- t[64664] = 43
      "0101011" when "01111110010011001", -- t[64665] = 43
      "0101011" when "01111110010011010", -- t[64666] = 43
      "0101011" when "01111110010011011", -- t[64667] = 43
      "0101011" when "01111110010011100", -- t[64668] = 43
      "0101011" when "01111110010011101", -- t[64669] = 43
      "0101011" when "01111110010011110", -- t[64670] = 43
      "0101011" when "01111110010011111", -- t[64671] = 43
      "0101011" when "01111110010100000", -- t[64672] = 43
      "0101011" when "01111110010100001", -- t[64673] = 43
      "0101011" when "01111110010100010", -- t[64674] = 43
      "0101011" when "01111110010100011", -- t[64675] = 43
      "0101011" when "01111110010100100", -- t[64676] = 43
      "0101011" when "01111110010100101", -- t[64677] = 43
      "0101011" when "01111110010100110", -- t[64678] = 43
      "0101011" when "01111110010100111", -- t[64679] = 43
      "0101011" when "01111110010101000", -- t[64680] = 43
      "0101011" when "01111110010101001", -- t[64681] = 43
      "0101011" when "01111110010101010", -- t[64682] = 43
      "0101011" when "01111110010101011", -- t[64683] = 43
      "0101011" when "01111110010101100", -- t[64684] = 43
      "0101011" when "01111110010101101", -- t[64685] = 43
      "0101011" when "01111110010101110", -- t[64686] = 43
      "0101011" when "01111110010101111", -- t[64687] = 43
      "0101011" when "01111110010110000", -- t[64688] = 43
      "0101011" when "01111110010110001", -- t[64689] = 43
      "0101011" when "01111110010110010", -- t[64690] = 43
      "0101011" when "01111110010110011", -- t[64691] = 43
      "0101011" when "01111110010110100", -- t[64692] = 43
      "0101011" when "01111110010110101", -- t[64693] = 43
      "0101011" when "01111110010110110", -- t[64694] = 43
      "0101011" when "01111110010110111", -- t[64695] = 43
      "0101011" when "01111110010111000", -- t[64696] = 43
      "0101011" when "01111110010111001", -- t[64697] = 43
      "0101011" when "01111110010111010", -- t[64698] = 43
      "0101011" when "01111110010111011", -- t[64699] = 43
      "0101011" when "01111110010111100", -- t[64700] = 43
      "0101011" when "01111110010111101", -- t[64701] = 43
      "0101011" when "01111110010111110", -- t[64702] = 43
      "0101011" when "01111110010111111", -- t[64703] = 43
      "0101011" when "01111110011000000", -- t[64704] = 43
      "0101011" when "01111110011000001", -- t[64705] = 43
      "0101011" when "01111110011000010", -- t[64706] = 43
      "0101011" when "01111110011000011", -- t[64707] = 43
      "0101011" when "01111110011000100", -- t[64708] = 43
      "0101011" when "01111110011000101", -- t[64709] = 43
      "0101011" when "01111110011000110", -- t[64710] = 43
      "0101011" when "01111110011000111", -- t[64711] = 43
      "0101011" when "01111110011001000", -- t[64712] = 43
      "0101011" when "01111110011001001", -- t[64713] = 43
      "0101011" when "01111110011001010", -- t[64714] = 43
      "0101011" when "01111110011001011", -- t[64715] = 43
      "0101011" when "01111110011001100", -- t[64716] = 43
      "0101011" when "01111110011001101", -- t[64717] = 43
      "0101011" when "01111110011001110", -- t[64718] = 43
      "0101011" when "01111110011001111", -- t[64719] = 43
      "0101011" when "01111110011010000", -- t[64720] = 43
      "0101011" when "01111110011010001", -- t[64721] = 43
      "0101011" when "01111110011010010", -- t[64722] = 43
      "0101011" when "01111110011010011", -- t[64723] = 43
      "0101011" when "01111110011010100", -- t[64724] = 43
      "0101011" when "01111110011010101", -- t[64725] = 43
      "0101011" when "01111110011010110", -- t[64726] = 43
      "0101011" when "01111110011010111", -- t[64727] = 43
      "0101011" when "01111110011011000", -- t[64728] = 43
      "0101011" when "01111110011011001", -- t[64729] = 43
      "0101011" when "01111110011011010", -- t[64730] = 43
      "0101011" when "01111110011011011", -- t[64731] = 43
      "0101011" when "01111110011011100", -- t[64732] = 43
      "0101011" when "01111110011011101", -- t[64733] = 43
      "0101011" when "01111110011011110", -- t[64734] = 43
      "0101011" when "01111110011011111", -- t[64735] = 43
      "0101011" when "01111110011100000", -- t[64736] = 43
      "0101011" when "01111110011100001", -- t[64737] = 43
      "0101011" when "01111110011100010", -- t[64738] = 43
      "0101011" when "01111110011100011", -- t[64739] = 43
      "0101011" when "01111110011100100", -- t[64740] = 43
      "0101011" when "01111110011100101", -- t[64741] = 43
      "0101011" when "01111110011100110", -- t[64742] = 43
      "0101011" when "01111110011100111", -- t[64743] = 43
      "0101011" when "01111110011101000", -- t[64744] = 43
      "0101011" when "01111110011101001", -- t[64745] = 43
      "0101011" when "01111110011101010", -- t[64746] = 43
      "0101011" when "01111110011101011", -- t[64747] = 43
      "0101011" when "01111110011101100", -- t[64748] = 43
      "0101011" when "01111110011101101", -- t[64749] = 43
      "0101011" when "01111110011101110", -- t[64750] = 43
      "0101011" when "01111110011101111", -- t[64751] = 43
      "0101011" when "01111110011110000", -- t[64752] = 43
      "0101011" when "01111110011110001", -- t[64753] = 43
      "0101011" when "01111110011110010", -- t[64754] = 43
      "0101011" when "01111110011110011", -- t[64755] = 43
      "0101011" when "01111110011110100", -- t[64756] = 43
      "0101011" when "01111110011110101", -- t[64757] = 43
      "0101011" when "01111110011110110", -- t[64758] = 43
      "0101011" when "01111110011110111", -- t[64759] = 43
      "0101011" when "01111110011111000", -- t[64760] = 43
      "0101011" when "01111110011111001", -- t[64761] = 43
      "0101011" when "01111110011111010", -- t[64762] = 43
      "0101011" when "01111110011111011", -- t[64763] = 43
      "0101011" when "01111110011111100", -- t[64764] = 43
      "0101011" when "01111110011111101", -- t[64765] = 43
      "0101011" when "01111110011111110", -- t[64766] = 43
      "0101011" when "01111110011111111", -- t[64767] = 43
      "0101011" when "01111110100000000", -- t[64768] = 43
      "0101011" when "01111110100000001", -- t[64769] = 43
      "0101011" when "01111110100000010", -- t[64770] = 43
      "0101011" when "01111110100000011", -- t[64771] = 43
      "0101011" when "01111110100000100", -- t[64772] = 43
      "0101011" when "01111110100000101", -- t[64773] = 43
      "0101011" when "01111110100000110", -- t[64774] = 43
      "0101011" when "01111110100000111", -- t[64775] = 43
      "0101011" when "01111110100001000", -- t[64776] = 43
      "0101011" when "01111110100001001", -- t[64777] = 43
      "0101011" when "01111110100001010", -- t[64778] = 43
      "0101011" when "01111110100001011", -- t[64779] = 43
      "0101011" when "01111110100001100", -- t[64780] = 43
      "0101011" when "01111110100001101", -- t[64781] = 43
      "0101011" when "01111110100001110", -- t[64782] = 43
      "0101011" when "01111110100001111", -- t[64783] = 43
      "0101011" when "01111110100010000", -- t[64784] = 43
      "0101011" when "01111110100010001", -- t[64785] = 43
      "0101011" when "01111110100010010", -- t[64786] = 43
      "0101011" when "01111110100010011", -- t[64787] = 43
      "0101011" when "01111110100010100", -- t[64788] = 43
      "0101011" when "01111110100010101", -- t[64789] = 43
      "0101011" when "01111110100010110", -- t[64790] = 43
      "0101011" when "01111110100010111", -- t[64791] = 43
      "0101011" when "01111110100011000", -- t[64792] = 43
      "0101011" when "01111110100011001", -- t[64793] = 43
      "0101011" when "01111110100011010", -- t[64794] = 43
      "0101011" when "01111110100011011", -- t[64795] = 43
      "0101011" when "01111110100011100", -- t[64796] = 43
      "0101011" when "01111110100011101", -- t[64797] = 43
      "0101011" when "01111110100011110", -- t[64798] = 43
      "0101011" when "01111110100011111", -- t[64799] = 43
      "0101011" when "01111110100100000", -- t[64800] = 43
      "0101011" when "01111110100100001", -- t[64801] = 43
      "0101011" when "01111110100100010", -- t[64802] = 43
      "0101011" when "01111110100100011", -- t[64803] = 43
      "0101011" when "01111110100100100", -- t[64804] = 43
      "0101011" when "01111110100100101", -- t[64805] = 43
      "0101011" when "01111110100100110", -- t[64806] = 43
      "0101011" when "01111110100100111", -- t[64807] = 43
      "0101011" when "01111110100101000", -- t[64808] = 43
      "0101011" when "01111110100101001", -- t[64809] = 43
      "0101011" when "01111110100101010", -- t[64810] = 43
      "0101011" when "01111110100101011", -- t[64811] = 43
      "0101100" when "01111110100101100", -- t[64812] = 44
      "0101100" when "01111110100101101", -- t[64813] = 44
      "0101100" when "01111110100101110", -- t[64814] = 44
      "0101100" when "01111110100101111", -- t[64815] = 44
      "0101100" when "01111110100110000", -- t[64816] = 44
      "0101100" when "01111110100110001", -- t[64817] = 44
      "0101100" when "01111110100110010", -- t[64818] = 44
      "0101100" when "01111110100110011", -- t[64819] = 44
      "0101100" when "01111110100110100", -- t[64820] = 44
      "0101100" when "01111110100110101", -- t[64821] = 44
      "0101100" when "01111110100110110", -- t[64822] = 44
      "0101100" when "01111110100110111", -- t[64823] = 44
      "0101100" when "01111110100111000", -- t[64824] = 44
      "0101100" when "01111110100111001", -- t[64825] = 44
      "0101100" when "01111110100111010", -- t[64826] = 44
      "0101100" when "01111110100111011", -- t[64827] = 44
      "0101100" when "01111110100111100", -- t[64828] = 44
      "0101100" when "01111110100111101", -- t[64829] = 44
      "0101100" when "01111110100111110", -- t[64830] = 44
      "0101100" when "01111110100111111", -- t[64831] = 44
      "0101100" when "01111110101000000", -- t[64832] = 44
      "0101100" when "01111110101000001", -- t[64833] = 44
      "0101100" when "01111110101000010", -- t[64834] = 44
      "0101100" when "01111110101000011", -- t[64835] = 44
      "0101100" when "01111110101000100", -- t[64836] = 44
      "0101100" when "01111110101000101", -- t[64837] = 44
      "0101100" when "01111110101000110", -- t[64838] = 44
      "0101100" when "01111110101000111", -- t[64839] = 44
      "0101100" when "01111110101001000", -- t[64840] = 44
      "0101100" when "01111110101001001", -- t[64841] = 44
      "0101100" when "01111110101001010", -- t[64842] = 44
      "0101100" when "01111110101001011", -- t[64843] = 44
      "0101100" when "01111110101001100", -- t[64844] = 44
      "0101100" when "01111110101001101", -- t[64845] = 44
      "0101100" when "01111110101001110", -- t[64846] = 44
      "0101100" when "01111110101001111", -- t[64847] = 44
      "0101100" when "01111110101010000", -- t[64848] = 44
      "0101100" when "01111110101010001", -- t[64849] = 44
      "0101100" when "01111110101010010", -- t[64850] = 44
      "0101100" when "01111110101010011", -- t[64851] = 44
      "0101100" when "01111110101010100", -- t[64852] = 44
      "0101100" when "01111110101010101", -- t[64853] = 44
      "0101100" when "01111110101010110", -- t[64854] = 44
      "0101100" when "01111110101010111", -- t[64855] = 44
      "0101100" when "01111110101011000", -- t[64856] = 44
      "0101100" when "01111110101011001", -- t[64857] = 44
      "0101100" when "01111110101011010", -- t[64858] = 44
      "0101100" when "01111110101011011", -- t[64859] = 44
      "0101100" when "01111110101011100", -- t[64860] = 44
      "0101100" when "01111110101011101", -- t[64861] = 44
      "0101100" when "01111110101011110", -- t[64862] = 44
      "0101100" when "01111110101011111", -- t[64863] = 44
      "0101100" when "01111110101100000", -- t[64864] = 44
      "0101100" when "01111110101100001", -- t[64865] = 44
      "0101100" when "01111110101100010", -- t[64866] = 44
      "0101100" when "01111110101100011", -- t[64867] = 44
      "0101100" when "01111110101100100", -- t[64868] = 44
      "0101100" when "01111110101100101", -- t[64869] = 44
      "0101100" when "01111110101100110", -- t[64870] = 44
      "0101100" when "01111110101100111", -- t[64871] = 44
      "0101100" when "01111110101101000", -- t[64872] = 44
      "0101100" when "01111110101101001", -- t[64873] = 44
      "0101100" when "01111110101101010", -- t[64874] = 44
      "0101100" when "01111110101101011", -- t[64875] = 44
      "0101100" when "01111110101101100", -- t[64876] = 44
      "0101100" when "01111110101101101", -- t[64877] = 44
      "0101100" when "01111110101101110", -- t[64878] = 44
      "0101100" when "01111110101101111", -- t[64879] = 44
      "0101100" when "01111110101110000", -- t[64880] = 44
      "0101100" when "01111110101110001", -- t[64881] = 44
      "0101100" when "01111110101110010", -- t[64882] = 44
      "0101100" when "01111110101110011", -- t[64883] = 44
      "0101100" when "01111110101110100", -- t[64884] = 44
      "0101100" when "01111110101110101", -- t[64885] = 44
      "0101100" when "01111110101110110", -- t[64886] = 44
      "0101100" when "01111110101110111", -- t[64887] = 44
      "0101100" when "01111110101111000", -- t[64888] = 44
      "0101100" when "01111110101111001", -- t[64889] = 44
      "0101100" when "01111110101111010", -- t[64890] = 44
      "0101100" when "01111110101111011", -- t[64891] = 44
      "0101100" when "01111110101111100", -- t[64892] = 44
      "0101100" when "01111110101111101", -- t[64893] = 44
      "0101100" when "01111110101111110", -- t[64894] = 44
      "0101100" when "01111110101111111", -- t[64895] = 44
      "0101100" when "01111110110000000", -- t[64896] = 44
      "0101100" when "01111110110000001", -- t[64897] = 44
      "0101100" when "01111110110000010", -- t[64898] = 44
      "0101100" when "01111110110000011", -- t[64899] = 44
      "0101100" when "01111110110000100", -- t[64900] = 44
      "0101100" when "01111110110000101", -- t[64901] = 44
      "0101100" when "01111110110000110", -- t[64902] = 44
      "0101100" when "01111110110000111", -- t[64903] = 44
      "0101100" when "01111110110001000", -- t[64904] = 44
      "0101100" when "01111110110001001", -- t[64905] = 44
      "0101100" when "01111110110001010", -- t[64906] = 44
      "0101100" when "01111110110001011", -- t[64907] = 44
      "0101100" when "01111110110001100", -- t[64908] = 44
      "0101100" when "01111110110001101", -- t[64909] = 44
      "0101100" when "01111110110001110", -- t[64910] = 44
      "0101100" when "01111110110001111", -- t[64911] = 44
      "0101100" when "01111110110010000", -- t[64912] = 44
      "0101100" when "01111110110010001", -- t[64913] = 44
      "0101100" when "01111110110010010", -- t[64914] = 44
      "0101100" when "01111110110010011", -- t[64915] = 44
      "0101100" when "01111110110010100", -- t[64916] = 44
      "0101100" when "01111110110010101", -- t[64917] = 44
      "0101100" when "01111110110010110", -- t[64918] = 44
      "0101100" when "01111110110010111", -- t[64919] = 44
      "0101100" when "01111110110011000", -- t[64920] = 44
      "0101100" when "01111110110011001", -- t[64921] = 44
      "0101100" when "01111110110011010", -- t[64922] = 44
      "0101100" when "01111110110011011", -- t[64923] = 44
      "0101100" when "01111110110011100", -- t[64924] = 44
      "0101100" when "01111110110011101", -- t[64925] = 44
      "0101100" when "01111110110011110", -- t[64926] = 44
      "0101100" when "01111110110011111", -- t[64927] = 44
      "0101100" when "01111110110100000", -- t[64928] = 44
      "0101100" when "01111110110100001", -- t[64929] = 44
      "0101100" when "01111110110100010", -- t[64930] = 44
      "0101100" when "01111110110100011", -- t[64931] = 44
      "0101100" when "01111110110100100", -- t[64932] = 44
      "0101100" when "01111110110100101", -- t[64933] = 44
      "0101100" when "01111110110100110", -- t[64934] = 44
      "0101100" when "01111110110100111", -- t[64935] = 44
      "0101100" when "01111110110101000", -- t[64936] = 44
      "0101100" when "01111110110101001", -- t[64937] = 44
      "0101100" when "01111110110101010", -- t[64938] = 44
      "0101100" when "01111110110101011", -- t[64939] = 44
      "0101100" when "01111110110101100", -- t[64940] = 44
      "0101100" when "01111110110101101", -- t[64941] = 44
      "0101100" when "01111110110101110", -- t[64942] = 44
      "0101100" when "01111110110101111", -- t[64943] = 44
      "0101100" when "01111110110110000", -- t[64944] = 44
      "0101100" when "01111110110110001", -- t[64945] = 44
      "0101100" when "01111110110110010", -- t[64946] = 44
      "0101100" when "01111110110110011", -- t[64947] = 44
      "0101100" when "01111110110110100", -- t[64948] = 44
      "0101100" when "01111110110110101", -- t[64949] = 44
      "0101100" when "01111110110110110", -- t[64950] = 44
      "0101100" when "01111110110110111", -- t[64951] = 44
      "0101100" when "01111110110111000", -- t[64952] = 44
      "0101100" when "01111110110111001", -- t[64953] = 44
      "0101100" when "01111110110111010", -- t[64954] = 44
      "0101100" when "01111110110111011", -- t[64955] = 44
      "0101100" when "01111110110111100", -- t[64956] = 44
      "0101100" when "01111110110111101", -- t[64957] = 44
      "0101100" when "01111110110111110", -- t[64958] = 44
      "0101100" when "01111110110111111", -- t[64959] = 44
      "0101100" when "01111110111000000", -- t[64960] = 44
      "0101100" when "01111110111000001", -- t[64961] = 44
      "0101100" when "01111110111000010", -- t[64962] = 44
      "0101100" when "01111110111000011", -- t[64963] = 44
      "0101100" when "01111110111000100", -- t[64964] = 44
      "0101100" when "01111110111000101", -- t[64965] = 44
      "0101100" when "01111110111000110", -- t[64966] = 44
      "0101100" when "01111110111000111", -- t[64967] = 44
      "0101100" when "01111110111001000", -- t[64968] = 44
      "0101100" when "01111110111001001", -- t[64969] = 44
      "0101100" when "01111110111001010", -- t[64970] = 44
      "0101100" when "01111110111001011", -- t[64971] = 44
      "0101100" when "01111110111001100", -- t[64972] = 44
      "0101100" when "01111110111001101", -- t[64973] = 44
      "0101100" when "01111110111001110", -- t[64974] = 44
      "0101100" when "01111110111001111", -- t[64975] = 44
      "0101100" when "01111110111010000", -- t[64976] = 44
      "0101100" when "01111110111010001", -- t[64977] = 44
      "0101100" when "01111110111010010", -- t[64978] = 44
      "0101100" when "01111110111010011", -- t[64979] = 44
      "0101100" when "01111110111010100", -- t[64980] = 44
      "0101100" when "01111110111010101", -- t[64981] = 44
      "0101100" when "01111110111010110", -- t[64982] = 44
      "0101100" when "01111110111010111", -- t[64983] = 44
      "0101100" when "01111110111011000", -- t[64984] = 44
      "0101100" when "01111110111011001", -- t[64985] = 44
      "0101100" when "01111110111011010", -- t[64986] = 44
      "0101100" when "01111110111011011", -- t[64987] = 44
      "0101100" when "01111110111011100", -- t[64988] = 44
      "0101100" when "01111110111011101", -- t[64989] = 44
      "0101100" when "01111110111011110", -- t[64990] = 44
      "0101100" when "01111110111011111", -- t[64991] = 44
      "0101100" when "01111110111100000", -- t[64992] = 44
      "0101100" when "01111110111100001", -- t[64993] = 44
      "0101100" when "01111110111100010", -- t[64994] = 44
      "0101100" when "01111110111100011", -- t[64995] = 44
      "0101100" when "01111110111100100", -- t[64996] = 44
      "0101100" when "01111110111100101", -- t[64997] = 44
      "0101100" when "01111110111100110", -- t[64998] = 44
      "0101100" when "01111110111100111", -- t[64999] = 44
      "0101100" when "01111110111101000", -- t[65000] = 44
      "0101100" when "01111110111101001", -- t[65001] = 44
      "0101100" when "01111110111101010", -- t[65002] = 44
      "0101100" when "01111110111101011", -- t[65003] = 44
      "0101100" when "01111110111101100", -- t[65004] = 44
      "0101100" when "01111110111101101", -- t[65005] = 44
      "0101100" when "01111110111101110", -- t[65006] = 44
      "0101100" when "01111110111101111", -- t[65007] = 44
      "0101100" when "01111110111110000", -- t[65008] = 44
      "0101100" when "01111110111110001", -- t[65009] = 44
      "0101100" when "01111110111110010", -- t[65010] = 44
      "0101100" when "01111110111110011", -- t[65011] = 44
      "0101100" when "01111110111110100", -- t[65012] = 44
      "0101100" when "01111110111110101", -- t[65013] = 44
      "0101100" when "01111110111110110", -- t[65014] = 44
      "0101100" when "01111110111110111", -- t[65015] = 44
      "0101100" when "01111110111111000", -- t[65016] = 44
      "0101100" when "01111110111111001", -- t[65017] = 44
      "0101100" when "01111110111111010", -- t[65018] = 44
      "0101100" when "01111110111111011", -- t[65019] = 44
      "0101100" when "01111110111111100", -- t[65020] = 44
      "0101100" when "01111110111111101", -- t[65021] = 44
      "0101100" when "01111110111111110", -- t[65022] = 44
      "0101100" when "01111110111111111", -- t[65023] = 44
      "0101100" when "01111111000000000", -- t[65024] = 44
      "0101100" when "01111111000000001", -- t[65025] = 44
      "0101100" when "01111111000000010", -- t[65026] = 44
      "0101100" when "01111111000000011", -- t[65027] = 44
      "0101100" when "01111111000000100", -- t[65028] = 44
      "0101100" when "01111111000000101", -- t[65029] = 44
      "0101100" when "01111111000000110", -- t[65030] = 44
      "0101100" when "01111111000000111", -- t[65031] = 44
      "0101100" when "01111111000001000", -- t[65032] = 44
      "0101100" when "01111111000001001", -- t[65033] = 44
      "0101100" when "01111111000001010", -- t[65034] = 44
      "0101100" when "01111111000001011", -- t[65035] = 44
      "0101100" when "01111111000001100", -- t[65036] = 44
      "0101100" when "01111111000001101", -- t[65037] = 44
      "0101100" when "01111111000001110", -- t[65038] = 44
      "0101100" when "01111111000001111", -- t[65039] = 44
      "0101100" when "01111111000010000", -- t[65040] = 44
      "0101100" when "01111111000010001", -- t[65041] = 44
      "0101100" when "01111111000010010", -- t[65042] = 44
      "0101100" when "01111111000010011", -- t[65043] = 44
      "0101100" when "01111111000010100", -- t[65044] = 44
      "0101100" when "01111111000010101", -- t[65045] = 44
      "0101100" when "01111111000010110", -- t[65046] = 44
      "0101100" when "01111111000010111", -- t[65047] = 44
      "0101100" when "01111111000011000", -- t[65048] = 44
      "0101100" when "01111111000011001", -- t[65049] = 44
      "0101100" when "01111111000011010", -- t[65050] = 44
      "0101100" when "01111111000011011", -- t[65051] = 44
      "0101100" when "01111111000011100", -- t[65052] = 44
      "0101100" when "01111111000011101", -- t[65053] = 44
      "0101100" when "01111111000011110", -- t[65054] = 44
      "0101100" when "01111111000011111", -- t[65055] = 44
      "0101100" when "01111111000100000", -- t[65056] = 44
      "0101100" when "01111111000100001", -- t[65057] = 44
      "0101100" when "01111111000100010", -- t[65058] = 44
      "0101100" when "01111111000100011", -- t[65059] = 44
      "0101100" when "01111111000100100", -- t[65060] = 44
      "0101100" when "01111111000100101", -- t[65061] = 44
      "0101100" when "01111111000100110", -- t[65062] = 44
      "0101100" when "01111111000100111", -- t[65063] = 44
      "0101100" when "01111111000101000", -- t[65064] = 44
      "0101100" when "01111111000101001", -- t[65065] = 44
      "0101100" when "01111111000101010", -- t[65066] = 44
      "0101100" when "01111111000101011", -- t[65067] = 44
      "0101100" when "01111111000101100", -- t[65068] = 44
      "0101100" when "01111111000101101", -- t[65069] = 44
      "0101100" when "01111111000101110", -- t[65070] = 44
      "0101100" when "01111111000101111", -- t[65071] = 44
      "0101100" when "01111111000110000", -- t[65072] = 44
      "0101100" when "01111111000110001", -- t[65073] = 44
      "0101100" when "01111111000110010", -- t[65074] = 44
      "0101100" when "01111111000110011", -- t[65075] = 44
      "0101100" when "01111111000110100", -- t[65076] = 44
      "0101100" when "01111111000110101", -- t[65077] = 44
      "0101100" when "01111111000110110", -- t[65078] = 44
      "0101100" when "01111111000110111", -- t[65079] = 44
      "0101101" when "01111111000111000", -- t[65080] = 45
      "0101101" when "01111111000111001", -- t[65081] = 45
      "0101101" when "01111111000111010", -- t[65082] = 45
      "0101101" when "01111111000111011", -- t[65083] = 45
      "0101101" when "01111111000111100", -- t[65084] = 45
      "0101101" when "01111111000111101", -- t[65085] = 45
      "0101101" when "01111111000111110", -- t[65086] = 45
      "0101101" when "01111111000111111", -- t[65087] = 45
      "0101101" when "01111111001000000", -- t[65088] = 45
      "0101101" when "01111111001000001", -- t[65089] = 45
      "0101101" when "01111111001000010", -- t[65090] = 45
      "0101101" when "01111111001000011", -- t[65091] = 45
      "0101101" when "01111111001000100", -- t[65092] = 45
      "0101101" when "01111111001000101", -- t[65093] = 45
      "0101101" when "01111111001000110", -- t[65094] = 45
      "0101101" when "01111111001000111", -- t[65095] = 45
      "0101101" when "01111111001001000", -- t[65096] = 45
      "0101101" when "01111111001001001", -- t[65097] = 45
      "0101101" when "01111111001001010", -- t[65098] = 45
      "0101101" when "01111111001001011", -- t[65099] = 45
      "0101101" when "01111111001001100", -- t[65100] = 45
      "0101101" when "01111111001001101", -- t[65101] = 45
      "0101101" when "01111111001001110", -- t[65102] = 45
      "0101101" when "01111111001001111", -- t[65103] = 45
      "0101101" when "01111111001010000", -- t[65104] = 45
      "0101101" when "01111111001010001", -- t[65105] = 45
      "0101101" when "01111111001010010", -- t[65106] = 45
      "0101101" when "01111111001010011", -- t[65107] = 45
      "0101101" when "01111111001010100", -- t[65108] = 45
      "0101101" when "01111111001010101", -- t[65109] = 45
      "0101101" when "01111111001010110", -- t[65110] = 45
      "0101101" when "01111111001010111", -- t[65111] = 45
      "0101101" when "01111111001011000", -- t[65112] = 45
      "0101101" when "01111111001011001", -- t[65113] = 45
      "0101101" when "01111111001011010", -- t[65114] = 45
      "0101101" when "01111111001011011", -- t[65115] = 45
      "0101101" when "01111111001011100", -- t[65116] = 45
      "0101101" when "01111111001011101", -- t[65117] = 45
      "0101101" when "01111111001011110", -- t[65118] = 45
      "0101101" when "01111111001011111", -- t[65119] = 45
      "0101101" when "01111111001100000", -- t[65120] = 45
      "0101101" when "01111111001100001", -- t[65121] = 45
      "0101101" when "01111111001100010", -- t[65122] = 45
      "0101101" when "01111111001100011", -- t[65123] = 45
      "0101101" when "01111111001100100", -- t[65124] = 45
      "0101101" when "01111111001100101", -- t[65125] = 45
      "0101101" when "01111111001100110", -- t[65126] = 45
      "0101101" when "01111111001100111", -- t[65127] = 45
      "0101101" when "01111111001101000", -- t[65128] = 45
      "0101101" when "01111111001101001", -- t[65129] = 45
      "0101101" when "01111111001101010", -- t[65130] = 45
      "0101101" when "01111111001101011", -- t[65131] = 45
      "0101101" when "01111111001101100", -- t[65132] = 45
      "0101101" when "01111111001101101", -- t[65133] = 45
      "0101101" when "01111111001101110", -- t[65134] = 45
      "0101101" when "01111111001101111", -- t[65135] = 45
      "0101101" when "01111111001110000", -- t[65136] = 45
      "0101101" when "01111111001110001", -- t[65137] = 45
      "0101101" when "01111111001110010", -- t[65138] = 45
      "0101101" when "01111111001110011", -- t[65139] = 45
      "0101101" when "01111111001110100", -- t[65140] = 45
      "0101101" when "01111111001110101", -- t[65141] = 45
      "0101101" when "01111111001110110", -- t[65142] = 45
      "0101101" when "01111111001110111", -- t[65143] = 45
      "0101101" when "01111111001111000", -- t[65144] = 45
      "0101101" when "01111111001111001", -- t[65145] = 45
      "0101101" when "01111111001111010", -- t[65146] = 45
      "0101101" when "01111111001111011", -- t[65147] = 45
      "0101101" when "01111111001111100", -- t[65148] = 45
      "0101101" when "01111111001111101", -- t[65149] = 45
      "0101101" when "01111111001111110", -- t[65150] = 45
      "0101101" when "01111111001111111", -- t[65151] = 45
      "0101101" when "01111111010000000", -- t[65152] = 45
      "0101101" when "01111111010000001", -- t[65153] = 45
      "0101101" when "01111111010000010", -- t[65154] = 45
      "0101101" when "01111111010000011", -- t[65155] = 45
      "0101101" when "01111111010000100", -- t[65156] = 45
      "0101101" when "01111111010000101", -- t[65157] = 45
      "0101101" when "01111111010000110", -- t[65158] = 45
      "0101101" when "01111111010000111", -- t[65159] = 45
      "0101101" when "01111111010001000", -- t[65160] = 45
      "0101101" when "01111111010001001", -- t[65161] = 45
      "0101101" when "01111111010001010", -- t[65162] = 45
      "0101101" when "01111111010001011", -- t[65163] = 45
      "0101101" when "01111111010001100", -- t[65164] = 45
      "0101101" when "01111111010001101", -- t[65165] = 45
      "0101101" when "01111111010001110", -- t[65166] = 45
      "0101101" when "01111111010001111", -- t[65167] = 45
      "0101101" when "01111111010010000", -- t[65168] = 45
      "0101101" when "01111111010010001", -- t[65169] = 45
      "0101101" when "01111111010010010", -- t[65170] = 45
      "0101101" when "01111111010010011", -- t[65171] = 45
      "0101101" when "01111111010010100", -- t[65172] = 45
      "0101101" when "01111111010010101", -- t[65173] = 45
      "0101101" when "01111111010010110", -- t[65174] = 45
      "0101101" when "01111111010010111", -- t[65175] = 45
      "0101101" when "01111111010011000", -- t[65176] = 45
      "0101101" when "01111111010011001", -- t[65177] = 45
      "0101101" when "01111111010011010", -- t[65178] = 45
      "0101101" when "01111111010011011", -- t[65179] = 45
      "0101101" when "01111111010011100", -- t[65180] = 45
      "0101101" when "01111111010011101", -- t[65181] = 45
      "0101101" when "01111111010011110", -- t[65182] = 45
      "0101101" when "01111111010011111", -- t[65183] = 45
      "0101101" when "01111111010100000", -- t[65184] = 45
      "0101101" when "01111111010100001", -- t[65185] = 45
      "0101101" when "01111111010100010", -- t[65186] = 45
      "0101101" when "01111111010100011", -- t[65187] = 45
      "0101101" when "01111111010100100", -- t[65188] = 45
      "0101101" when "01111111010100101", -- t[65189] = 45
      "0101101" when "01111111010100110", -- t[65190] = 45
      "0101101" when "01111111010100111", -- t[65191] = 45
      "0101101" when "01111111010101000", -- t[65192] = 45
      "0101101" when "01111111010101001", -- t[65193] = 45
      "0101101" when "01111111010101010", -- t[65194] = 45
      "0101101" when "01111111010101011", -- t[65195] = 45
      "0101101" when "01111111010101100", -- t[65196] = 45
      "0101101" when "01111111010101101", -- t[65197] = 45
      "0101101" when "01111111010101110", -- t[65198] = 45
      "0101101" when "01111111010101111", -- t[65199] = 45
      "0101101" when "01111111010110000", -- t[65200] = 45
      "0101101" when "01111111010110001", -- t[65201] = 45
      "0101101" when "01111111010110010", -- t[65202] = 45
      "0101101" when "01111111010110011", -- t[65203] = 45
      "0101101" when "01111111010110100", -- t[65204] = 45
      "0101101" when "01111111010110101", -- t[65205] = 45
      "0101101" when "01111111010110110", -- t[65206] = 45
      "0101101" when "01111111010110111", -- t[65207] = 45
      "0101101" when "01111111010111000", -- t[65208] = 45
      "0101101" when "01111111010111001", -- t[65209] = 45
      "0101101" when "01111111010111010", -- t[65210] = 45
      "0101101" when "01111111010111011", -- t[65211] = 45
      "0101101" when "01111111010111100", -- t[65212] = 45
      "0101101" when "01111111010111101", -- t[65213] = 45
      "0101101" when "01111111010111110", -- t[65214] = 45
      "0101101" when "01111111010111111", -- t[65215] = 45
      "0101101" when "01111111011000000", -- t[65216] = 45
      "0101101" when "01111111011000001", -- t[65217] = 45
      "0101101" when "01111111011000010", -- t[65218] = 45
      "0101101" when "01111111011000011", -- t[65219] = 45
      "0101101" when "01111111011000100", -- t[65220] = 45
      "0101101" when "01111111011000101", -- t[65221] = 45
      "0101101" when "01111111011000110", -- t[65222] = 45
      "0101101" when "01111111011000111", -- t[65223] = 45
      "0101101" when "01111111011001000", -- t[65224] = 45
      "0101101" when "01111111011001001", -- t[65225] = 45
      "0101101" when "01111111011001010", -- t[65226] = 45
      "0101101" when "01111111011001011", -- t[65227] = 45
      "0101101" when "01111111011001100", -- t[65228] = 45
      "0101101" when "01111111011001101", -- t[65229] = 45
      "0101101" when "01111111011001110", -- t[65230] = 45
      "0101101" when "01111111011001111", -- t[65231] = 45
      "0101101" when "01111111011010000", -- t[65232] = 45
      "0101101" when "01111111011010001", -- t[65233] = 45
      "0101101" when "01111111011010010", -- t[65234] = 45
      "0101101" when "01111111011010011", -- t[65235] = 45
      "0101101" when "01111111011010100", -- t[65236] = 45
      "0101101" when "01111111011010101", -- t[65237] = 45
      "0101101" when "01111111011010110", -- t[65238] = 45
      "0101101" when "01111111011010111", -- t[65239] = 45
      "0101101" when "01111111011011000", -- t[65240] = 45
      "0101101" when "01111111011011001", -- t[65241] = 45
      "0101101" when "01111111011011010", -- t[65242] = 45
      "0101101" when "01111111011011011", -- t[65243] = 45
      "0101101" when "01111111011011100", -- t[65244] = 45
      "0101101" when "01111111011011101", -- t[65245] = 45
      "0101101" when "01111111011011110", -- t[65246] = 45
      "0101101" when "01111111011011111", -- t[65247] = 45
      "0101101" when "01111111011100000", -- t[65248] = 45
      "0101101" when "01111111011100001", -- t[65249] = 45
      "0101101" when "01111111011100010", -- t[65250] = 45
      "0101101" when "01111111011100011", -- t[65251] = 45
      "0101101" when "01111111011100100", -- t[65252] = 45
      "0101101" when "01111111011100101", -- t[65253] = 45
      "0101101" when "01111111011100110", -- t[65254] = 45
      "0101101" when "01111111011100111", -- t[65255] = 45
      "0101101" when "01111111011101000", -- t[65256] = 45
      "0101101" when "01111111011101001", -- t[65257] = 45
      "0101101" when "01111111011101010", -- t[65258] = 45
      "0101101" when "01111111011101011", -- t[65259] = 45
      "0101101" when "01111111011101100", -- t[65260] = 45
      "0101101" when "01111111011101101", -- t[65261] = 45
      "0101101" when "01111111011101110", -- t[65262] = 45
      "0101101" when "01111111011101111", -- t[65263] = 45
      "0101101" when "01111111011110000", -- t[65264] = 45
      "0101101" when "01111111011110001", -- t[65265] = 45
      "0101101" when "01111111011110010", -- t[65266] = 45
      "0101101" when "01111111011110011", -- t[65267] = 45
      "0101101" when "01111111011110100", -- t[65268] = 45
      "0101101" when "01111111011110101", -- t[65269] = 45
      "0101101" when "01111111011110110", -- t[65270] = 45
      "0101101" when "01111111011110111", -- t[65271] = 45
      "0101101" when "01111111011111000", -- t[65272] = 45
      "0101101" when "01111111011111001", -- t[65273] = 45
      "0101101" when "01111111011111010", -- t[65274] = 45
      "0101101" when "01111111011111011", -- t[65275] = 45
      "0101101" when "01111111011111100", -- t[65276] = 45
      "0101101" when "01111111011111101", -- t[65277] = 45
      "0101101" when "01111111011111110", -- t[65278] = 45
      "0101101" when "01111111011111111", -- t[65279] = 45
      "0101101" when "01111111100000000", -- t[65280] = 45
      "0101101" when "01111111100000001", -- t[65281] = 45
      "0101101" when "01111111100000010", -- t[65282] = 45
      "0101101" when "01111111100000011", -- t[65283] = 45
      "0101101" when "01111111100000100", -- t[65284] = 45
      "0101101" when "01111111100000101", -- t[65285] = 45
      "0101101" when "01111111100000110", -- t[65286] = 45
      "0101101" when "01111111100000111", -- t[65287] = 45
      "0101101" when "01111111100001000", -- t[65288] = 45
      "0101101" when "01111111100001001", -- t[65289] = 45
      "0101101" when "01111111100001010", -- t[65290] = 45
      "0101101" when "01111111100001011", -- t[65291] = 45
      "0101101" when "01111111100001100", -- t[65292] = 45
      "0101101" when "01111111100001101", -- t[65293] = 45
      "0101101" when "01111111100001110", -- t[65294] = 45
      "0101101" when "01111111100001111", -- t[65295] = 45
      "0101101" when "01111111100010000", -- t[65296] = 45
      "0101101" when "01111111100010001", -- t[65297] = 45
      "0101101" when "01111111100010010", -- t[65298] = 45
      "0101101" when "01111111100010011", -- t[65299] = 45
      "0101101" when "01111111100010100", -- t[65300] = 45
      "0101101" when "01111111100010101", -- t[65301] = 45
      "0101101" when "01111111100010110", -- t[65302] = 45
      "0101101" when "01111111100010111", -- t[65303] = 45
      "0101101" when "01111111100011000", -- t[65304] = 45
      "0101101" when "01111111100011001", -- t[65305] = 45
      "0101101" when "01111111100011010", -- t[65306] = 45
      "0101101" when "01111111100011011", -- t[65307] = 45
      "0101101" when "01111111100011100", -- t[65308] = 45
      "0101101" when "01111111100011101", -- t[65309] = 45
      "0101101" when "01111111100011110", -- t[65310] = 45
      "0101101" when "01111111100011111", -- t[65311] = 45
      "0101101" when "01111111100100000", -- t[65312] = 45
      "0101101" when "01111111100100001", -- t[65313] = 45
      "0101101" when "01111111100100010", -- t[65314] = 45
      "0101101" when "01111111100100011", -- t[65315] = 45
      "0101101" when "01111111100100100", -- t[65316] = 45
      "0101101" when "01111111100100101", -- t[65317] = 45
      "0101101" when "01111111100100110", -- t[65318] = 45
      "0101101" when "01111111100100111", -- t[65319] = 45
      "0101101" when "01111111100101000", -- t[65320] = 45
      "0101101" when "01111111100101001", -- t[65321] = 45
      "0101101" when "01111111100101010", -- t[65322] = 45
      "0101101" when "01111111100101011", -- t[65323] = 45
      "0101101" when "01111111100101100", -- t[65324] = 45
      "0101101" when "01111111100101101", -- t[65325] = 45
      "0101101" when "01111111100101110", -- t[65326] = 45
      "0101101" when "01111111100101111", -- t[65327] = 45
      "0101101" when "01111111100110000", -- t[65328] = 45
      "0101101" when "01111111100110001", -- t[65329] = 45
      "0101101" when "01111111100110010", -- t[65330] = 45
      "0101101" when "01111111100110011", -- t[65331] = 45
      "0101101" when "01111111100110100", -- t[65332] = 45
      "0101101" when "01111111100110101", -- t[65333] = 45
      "0101101" when "01111111100110110", -- t[65334] = 45
      "0101101" when "01111111100110111", -- t[65335] = 45
      "0101101" when "01111111100111000", -- t[65336] = 45
      "0101101" when "01111111100111001", -- t[65337] = 45
      "0101101" when "01111111100111010", -- t[65338] = 45
      "0101101" when "01111111100111011", -- t[65339] = 45
      "0101101" when "01111111100111100", -- t[65340] = 45
      "0101101" when "01111111100111101", -- t[65341] = 45
      "0101110" when "01111111100111110", -- t[65342] = 46
      "0101110" when "01111111100111111", -- t[65343] = 46
      "0101110" when "01111111101000000", -- t[65344] = 46
      "0101110" when "01111111101000001", -- t[65345] = 46
      "0101110" when "01111111101000010", -- t[65346] = 46
      "0101110" when "01111111101000011", -- t[65347] = 46
      "0101110" when "01111111101000100", -- t[65348] = 46
      "0101110" when "01111111101000101", -- t[65349] = 46
      "0101110" when "01111111101000110", -- t[65350] = 46
      "0101110" when "01111111101000111", -- t[65351] = 46
      "0101110" when "01111111101001000", -- t[65352] = 46
      "0101110" when "01111111101001001", -- t[65353] = 46
      "0101110" when "01111111101001010", -- t[65354] = 46
      "0101110" when "01111111101001011", -- t[65355] = 46
      "0101110" when "01111111101001100", -- t[65356] = 46
      "0101110" when "01111111101001101", -- t[65357] = 46
      "0101110" when "01111111101001110", -- t[65358] = 46
      "0101110" when "01111111101001111", -- t[65359] = 46
      "0101110" when "01111111101010000", -- t[65360] = 46
      "0101110" when "01111111101010001", -- t[65361] = 46
      "0101110" when "01111111101010010", -- t[65362] = 46
      "0101110" when "01111111101010011", -- t[65363] = 46
      "0101110" when "01111111101010100", -- t[65364] = 46
      "0101110" when "01111111101010101", -- t[65365] = 46
      "0101110" when "01111111101010110", -- t[65366] = 46
      "0101110" when "01111111101010111", -- t[65367] = 46
      "0101110" when "01111111101011000", -- t[65368] = 46
      "0101110" when "01111111101011001", -- t[65369] = 46
      "0101110" when "01111111101011010", -- t[65370] = 46
      "0101110" when "01111111101011011", -- t[65371] = 46
      "0101110" when "01111111101011100", -- t[65372] = 46
      "0101110" when "01111111101011101", -- t[65373] = 46
      "0101110" when "01111111101011110", -- t[65374] = 46
      "0101110" when "01111111101011111", -- t[65375] = 46
      "0101110" when "01111111101100000", -- t[65376] = 46
      "0101110" when "01111111101100001", -- t[65377] = 46
      "0101110" when "01111111101100010", -- t[65378] = 46
      "0101110" when "01111111101100011", -- t[65379] = 46
      "0101110" when "01111111101100100", -- t[65380] = 46
      "0101110" when "01111111101100101", -- t[65381] = 46
      "0101110" when "01111111101100110", -- t[65382] = 46
      "0101110" when "01111111101100111", -- t[65383] = 46
      "0101110" when "01111111101101000", -- t[65384] = 46
      "0101110" when "01111111101101001", -- t[65385] = 46
      "0101110" when "01111111101101010", -- t[65386] = 46
      "0101110" when "01111111101101011", -- t[65387] = 46
      "0101110" when "01111111101101100", -- t[65388] = 46
      "0101110" when "01111111101101101", -- t[65389] = 46
      "0101110" when "01111111101101110", -- t[65390] = 46
      "0101110" when "01111111101101111", -- t[65391] = 46
      "0101110" when "01111111101110000", -- t[65392] = 46
      "0101110" when "01111111101110001", -- t[65393] = 46
      "0101110" when "01111111101110010", -- t[65394] = 46
      "0101110" when "01111111101110011", -- t[65395] = 46
      "0101110" when "01111111101110100", -- t[65396] = 46
      "0101110" when "01111111101110101", -- t[65397] = 46
      "0101110" when "01111111101110110", -- t[65398] = 46
      "0101110" when "01111111101110111", -- t[65399] = 46
      "0101110" when "01111111101111000", -- t[65400] = 46
      "0101110" when "01111111101111001", -- t[65401] = 46
      "0101110" when "01111111101111010", -- t[65402] = 46
      "0101110" when "01111111101111011", -- t[65403] = 46
      "0101110" when "01111111101111100", -- t[65404] = 46
      "0101110" when "01111111101111101", -- t[65405] = 46
      "0101110" when "01111111101111110", -- t[65406] = 46
      "0101110" when "01111111101111111", -- t[65407] = 46
      "0101110" when "01111111110000000", -- t[65408] = 46
      "0101110" when "01111111110000001", -- t[65409] = 46
      "0101110" when "01111111110000010", -- t[65410] = 46
      "0101110" when "01111111110000011", -- t[65411] = 46
      "0101110" when "01111111110000100", -- t[65412] = 46
      "0101110" when "01111111110000101", -- t[65413] = 46
      "0101110" when "01111111110000110", -- t[65414] = 46
      "0101110" when "01111111110000111", -- t[65415] = 46
      "0101110" when "01111111110001000", -- t[65416] = 46
      "0101110" when "01111111110001001", -- t[65417] = 46
      "0101110" when "01111111110001010", -- t[65418] = 46
      "0101110" when "01111111110001011", -- t[65419] = 46
      "0101110" when "01111111110001100", -- t[65420] = 46
      "0101110" when "01111111110001101", -- t[65421] = 46
      "0101110" when "01111111110001110", -- t[65422] = 46
      "0101110" when "01111111110001111", -- t[65423] = 46
      "0101110" when "01111111110010000", -- t[65424] = 46
      "0101110" when "01111111110010001", -- t[65425] = 46
      "0101110" when "01111111110010010", -- t[65426] = 46
      "0101110" when "01111111110010011", -- t[65427] = 46
      "0101110" when "01111111110010100", -- t[65428] = 46
      "0101110" when "01111111110010101", -- t[65429] = 46
      "0101110" when "01111111110010110", -- t[65430] = 46
      "0101110" when "01111111110010111", -- t[65431] = 46
      "0101110" when "01111111110011000", -- t[65432] = 46
      "0101110" when "01111111110011001", -- t[65433] = 46
      "0101110" when "01111111110011010", -- t[65434] = 46
      "0101110" when "01111111110011011", -- t[65435] = 46
      "0101110" when "01111111110011100", -- t[65436] = 46
      "0101110" when "01111111110011101", -- t[65437] = 46
      "0101110" when "01111111110011110", -- t[65438] = 46
      "0101110" when "01111111110011111", -- t[65439] = 46
      "0101110" when "01111111110100000", -- t[65440] = 46
      "0101110" when "01111111110100001", -- t[65441] = 46
      "0101110" when "01111111110100010", -- t[65442] = 46
      "0101110" when "01111111110100011", -- t[65443] = 46
      "0101110" when "01111111110100100", -- t[65444] = 46
      "0101110" when "01111111110100101", -- t[65445] = 46
      "0101110" when "01111111110100110", -- t[65446] = 46
      "0101110" when "01111111110100111", -- t[65447] = 46
      "0101110" when "01111111110101000", -- t[65448] = 46
      "0101110" when "01111111110101001", -- t[65449] = 46
      "0101110" when "01111111110101010", -- t[65450] = 46
      "0101110" when "01111111110101011", -- t[65451] = 46
      "0101110" when "01111111110101100", -- t[65452] = 46
      "0101110" when "01111111110101101", -- t[65453] = 46
      "0101110" when "01111111110101110", -- t[65454] = 46
      "0101110" when "01111111110101111", -- t[65455] = 46
      "0101110" when "01111111110110000", -- t[65456] = 46
      "0101110" when "01111111110110001", -- t[65457] = 46
      "0101110" when "01111111110110010", -- t[65458] = 46
      "0101110" when "01111111110110011", -- t[65459] = 46
      "0101110" when "01111111110110100", -- t[65460] = 46
      "0101110" when "01111111110110101", -- t[65461] = 46
      "0101110" when "01111111110110110", -- t[65462] = 46
      "0101110" when "01111111110110111", -- t[65463] = 46
      "0101110" when "01111111110111000", -- t[65464] = 46
      "0101110" when "01111111110111001", -- t[65465] = 46
      "0101110" when "01111111110111010", -- t[65466] = 46
      "0101110" when "01111111110111011", -- t[65467] = 46
      "0101110" when "01111111110111100", -- t[65468] = 46
      "0101110" when "01111111110111101", -- t[65469] = 46
      "0101110" when "01111111110111110", -- t[65470] = 46
      "0101110" when "01111111110111111", -- t[65471] = 46
      "0101110" when "01111111111000000", -- t[65472] = 46
      "0101110" when "01111111111000001", -- t[65473] = 46
      "0101110" when "01111111111000010", -- t[65474] = 46
      "0101110" when "01111111111000011", -- t[65475] = 46
      "0101110" when "01111111111000100", -- t[65476] = 46
      "0101110" when "01111111111000101", -- t[65477] = 46
      "0101110" when "01111111111000110", -- t[65478] = 46
      "0101110" when "01111111111000111", -- t[65479] = 46
      "0101110" when "01111111111001000", -- t[65480] = 46
      "0101110" when "01111111111001001", -- t[65481] = 46
      "0101110" when "01111111111001010", -- t[65482] = 46
      "0101110" when "01111111111001011", -- t[65483] = 46
      "0101110" when "01111111111001100", -- t[65484] = 46
      "0101110" when "01111111111001101", -- t[65485] = 46
      "0101110" when "01111111111001110", -- t[65486] = 46
      "0101110" when "01111111111001111", -- t[65487] = 46
      "0101110" when "01111111111010000", -- t[65488] = 46
      "0101110" when "01111111111010001", -- t[65489] = 46
      "0101110" when "01111111111010010", -- t[65490] = 46
      "0101110" when "01111111111010011", -- t[65491] = 46
      "0101110" when "01111111111010100", -- t[65492] = 46
      "0101110" when "01111111111010101", -- t[65493] = 46
      "0101110" when "01111111111010110", -- t[65494] = 46
      "0101110" when "01111111111010111", -- t[65495] = 46
      "0101110" when "01111111111011000", -- t[65496] = 46
      "0101110" when "01111111111011001", -- t[65497] = 46
      "0101110" when "01111111111011010", -- t[65498] = 46
      "0101110" when "01111111111011011", -- t[65499] = 46
      "0101110" when "01111111111011100", -- t[65500] = 46
      "0101110" when "01111111111011101", -- t[65501] = 46
      "0101110" when "01111111111011110", -- t[65502] = 46
      "0101110" when "01111111111011111", -- t[65503] = 46
      "0101110" when "01111111111100000", -- t[65504] = 46
      "0101110" when "01111111111100001", -- t[65505] = 46
      "0101110" when "01111111111100010", -- t[65506] = 46
      "0101110" when "01111111111100011", -- t[65507] = 46
      "0101110" when "01111111111100100", -- t[65508] = 46
      "0101110" when "01111111111100101", -- t[65509] = 46
      "0101110" when "01111111111100110", -- t[65510] = 46
      "0101110" when "01111111111100111", -- t[65511] = 46
      "0101110" when "01111111111101000", -- t[65512] = 46
      "0101110" when "01111111111101001", -- t[65513] = 46
      "0101110" when "01111111111101010", -- t[65514] = 46
      "0101110" when "01111111111101011", -- t[65515] = 46
      "0101110" when "01111111111101100", -- t[65516] = 46
      "0101110" when "01111111111101101", -- t[65517] = 46
      "0101110" when "01111111111101110", -- t[65518] = 46
      "0101110" when "01111111111101111", -- t[65519] = 46
      "0101110" when "01111111111110000", -- t[65520] = 46
      "0101110" when "01111111111110001", -- t[65521] = 46
      "0101110" when "01111111111110010", -- t[65522] = 46
      "0101110" when "01111111111110011", -- t[65523] = 46
      "0101110" when "01111111111110100", -- t[65524] = 46
      "0101110" when "01111111111110101", -- t[65525] = 46
      "0101110" when "01111111111110110", -- t[65526] = 46
      "0101110" when "01111111111110111", -- t[65527] = 46
      "0101110" when "01111111111111000", -- t[65528] = 46
      "0101110" when "01111111111111001", -- t[65529] = 46
      "0101110" when "01111111111111010", -- t[65530] = 46
      "0101110" when "01111111111111011", -- t[65531] = 46
      "0101110" when "01111111111111100", -- t[65532] = 46
      "0101110" when "01111111111111101", -- t[65533] = 46
      "0101110" when "01111111111111110", -- t[65534] = 46
      "0101110" when "01111111111111111", -- t[65535] = 46
      "-------" when others;
end architecture;


-- MultiPartite: LNS subtraction function: [-7.999999999999998 -4.0[ -> [0.0 0.12500000000000003[
-- wI = 15 bits
-- wO = 10 bits
-- Decomposition: 9, 6 / 7, 6, 3 / 2, 2, 2
-- Guard bits: 3
-- Size: 7952 = 13.2^9 + 4.2^8 + 2.2^7 + 1.2^4

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T1_13 is
  component LNSSub_MPT_T1_13_tiv is
    port( x : in  std_logic_vector(8 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to2 is
    port( x : in  std_logic_vector(7 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to1 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to0 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to2_xor is
    port( a : in  std_logic_vector(6 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to1_xor is
    port( a : in  std_logic_vector(5 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T1_13_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_13_tiv is
  port( x : in  std_logic_vector(8 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_tiv is
begin
  with x select
    r <=
      "0000101111000" when "000000000", -- t[0] = 376
      "0000101111010" when "000000001", -- t[1] = 378
      "0000101111100" when "000000010", -- t[2] = 380
      "0000101111110" when "000000011", -- t[3] = 382
      "0000110000000" when "000000100", -- t[4] = 384
      "0000110000010" when "000000101", -- t[5] = 386
      "0000110000100" when "000000110", -- t[6] = 388
      "0000110000110" when "000000111", -- t[7] = 390
      "0000110001001" when "000001000", -- t[8] = 393
      "0000110001011" when "000001001", -- t[9] = 395
      "0000110001101" when "000001010", -- t[10] = 397
      "0000110001111" when "000001011", -- t[11] = 399
      "0000110010001" when "000001100", -- t[12] = 401
      "0000110010011" when "000001101", -- t[13] = 403
      "0000110010101" when "000001110", -- t[14] = 405
      "0000110011000" when "000001111", -- t[15] = 408
      "0000110011010" when "000010000", -- t[16] = 410
      "0000110011100" when "000010001", -- t[17] = 412
      "0000110011110" when "000010010", -- t[18] = 414
      "0000110100000" when "000010011", -- t[19] = 416
      "0000110100011" when "000010100", -- t[20] = 419
      "0000110100101" when "000010101", -- t[21] = 421
      "0000110100111" when "000010110", -- t[22] = 423
      "0000110101001" when "000010111", -- t[23] = 425
      "0000110101100" when "000011000", -- t[24] = 428
      "0000110101110" when "000011001", -- t[25] = 430
      "0000110110000" when "000011010", -- t[26] = 432
      "0000110110011" when "000011011", -- t[27] = 435
      "0000110110101" when "000011100", -- t[28] = 437
      "0000110110111" when "000011101", -- t[29] = 439
      "0000110111010" when "000011110", -- t[30] = 442
      "0000110111100" when "000011111", -- t[31] = 444
      "0000110111110" when "000100000", -- t[32] = 446
      "0000111000001" when "000100001", -- t[33] = 449
      "0000111000011" when "000100010", -- t[34] = 451
      "0000111000110" when "000100011", -- t[35] = 454
      "0000111001000" when "000100100", -- t[36] = 456
      "0000111001011" when "000100101", -- t[37] = 459
      "0000111001101" when "000100110", -- t[38] = 461
      "0000111010000" when "000100111", -- t[39] = 464
      "0000111010010" when "000101000", -- t[40] = 466
      "0000111010101" when "000101001", -- t[41] = 469
      "0000111010111" when "000101010", -- t[42] = 471
      "0000111011010" when "000101011", -- t[43] = 474
      "0000111011100" when "000101100", -- t[44] = 476
      "0000111011111" when "000101101", -- t[45] = 479
      "0000111100001" when "000101110", -- t[46] = 481
      "0000111100100" when "000101111", -- t[47] = 484
      "0000111100110" when "000110000", -- t[48] = 486
      "0000111101001" when "000110001", -- t[49] = 489
      "0000111101100" when "000110010", -- t[50] = 492
      "0000111101110" when "000110011", -- t[51] = 494
      "0000111110001" when "000110100", -- t[52] = 497
      "0000111110100" when "000110101", -- t[53] = 500
      "0000111110110" when "000110110", -- t[54] = 502
      "0000111111001" when "000110111", -- t[55] = 505
      "0000111111100" when "000111000", -- t[56] = 508
      "0000111111111" when "000111001", -- t[57] = 511
      "0001000000001" when "000111010", -- t[58] = 513
      "0001000000100" when "000111011", -- t[59] = 516
      "0001000000111" when "000111100", -- t[60] = 519
      "0001000001010" when "000111101", -- t[61] = 522
      "0001000001100" when "000111110", -- t[62] = 524
      "0001000001111" when "000111111", -- t[63] = 527
      "0001000010010" when "001000000", -- t[64] = 530
      "0001000010101" when "001000001", -- t[65] = 533
      "0001000011000" when "001000010", -- t[66] = 536
      "0001000011011" when "001000011", -- t[67] = 539
      "0001000011110" when "001000100", -- t[68] = 542
      "0001000100001" when "001000101", -- t[69] = 545
      "0001000100100" when "001000110", -- t[70] = 548
      "0001000100111" when "001000111", -- t[71] = 551
      "0001000101001" when "001001000", -- t[72] = 553
      "0001000101100" when "001001001", -- t[73] = 556
      "0001000101111" when "001001010", -- t[74] = 559
      "0001000110010" when "001001011", -- t[75] = 562
      "0001000110110" when "001001100", -- t[76] = 566
      "0001000111001" when "001001101", -- t[77] = 569
      "0001000111100" when "001001110", -- t[78] = 572
      "0001000111111" when "001001111", -- t[79] = 575
      "0001001000010" when "001010000", -- t[80] = 578
      "0001001000101" when "001010001", -- t[81] = 581
      "0001001001000" when "001010010", -- t[82] = 584
      "0001001001011" when "001010011", -- t[83] = 587
      "0001001001110" when "001010100", -- t[84] = 590
      "0001001010010" when "001010101", -- t[85] = 594
      "0001001010101" when "001010110", -- t[86] = 597
      "0001001011000" when "001010111", -- t[87] = 600
      "0001001011011" when "001011000", -- t[88] = 603
      "0001001011111" when "001011001", -- t[89] = 607
      "0001001100010" when "001011010", -- t[90] = 610
      "0001001100101" when "001011011", -- t[91] = 613
      "0001001101000" when "001011100", -- t[92] = 616
      "0001001101100" when "001011101", -- t[93] = 620
      "0001001101111" when "001011110", -- t[94] = 623
      "0001001110010" when "001011111", -- t[95] = 626
      "0001001110110" when "001100000", -- t[96] = 630
      "0001001111001" when "001100001", -- t[97] = 633
      "0001001111101" when "001100010", -- t[98] = 637
      "0001010000000" when "001100011", -- t[99] = 640
      "0001010000100" when "001100100", -- t[100] = 644
      "0001010000111" when "001100101", -- t[101] = 647
      "0001010001011" when "001100110", -- t[102] = 651
      "0001010001110" when "001100111", -- t[103] = 654
      "0001010010010" when "001101000", -- t[104] = 658
      "0001010010101" when "001101001", -- t[105] = 661
      "0001010011001" when "001101010", -- t[106] = 665
      "0001010011100" when "001101011", -- t[107] = 668
      "0001010100000" when "001101100", -- t[108] = 672
      "0001010100100" when "001101101", -- t[109] = 676
      "0001010100111" when "001101110", -- t[110] = 679
      "0001010101011" when "001101111", -- t[111] = 683
      "0001010101111" when "001110000", -- t[112] = 687
      "0001010110010" when "001110001", -- t[113] = 690
      "0001010110110" when "001110010", -- t[114] = 694
      "0001010111010" when "001110011", -- t[115] = 698
      "0001010111110" when "001110100", -- t[116] = 702
      "0001011000001" when "001110101", -- t[117] = 705
      "0001011000101" when "001110110", -- t[118] = 709
      "0001011001001" when "001110111", -- t[119] = 713
      "0001011001101" when "001111000", -- t[120] = 717
      "0001011010001" when "001111001", -- t[121] = 721
      "0001011010101" when "001111010", -- t[122] = 725
      "0001011011001" when "001111011", -- t[123] = 729
      "0001011011101" when "001111100", -- t[124] = 733
      "0001011100001" when "001111101", -- t[125] = 737
      "0001011100101" when "001111110", -- t[126] = 741
      "0001011101001" when "001111111", -- t[127] = 745
      "0001011101101" when "010000000", -- t[128] = 749
      "0001011110001" when "010000001", -- t[129] = 753
      "0001011110101" when "010000010", -- t[130] = 757
      "0001011111001" when "010000011", -- t[131] = 761
      "0001011111101" when "010000100", -- t[132] = 765
      "0001100000001" when "010000101", -- t[133] = 769
      "0001100000101" when "010000110", -- t[134] = 773
      "0001100001001" when "010000111", -- t[135] = 777
      "0001100001110" when "010001000", -- t[136] = 782
      "0001100010010" when "010001001", -- t[137] = 786
      "0001100010110" when "010001010", -- t[138] = 790
      "0001100011010" when "010001011", -- t[139] = 794
      "0001100011111" when "010001100", -- t[140] = 799
      "0001100100011" when "010001101", -- t[141] = 803
      "0001100100111" when "010001110", -- t[142] = 807
      "0001100101100" when "010001111", -- t[143] = 812
      "0001100110000" when "010010000", -- t[144] = 816
      "0001100110101" when "010010001", -- t[145] = 821
      "0001100111001" when "010010010", -- t[146] = 825
      "0001100111101" when "010010011", -- t[147] = 829
      "0001101000010" when "010010100", -- t[148] = 834
      "0001101000110" when "010010101", -- t[149] = 838
      "0001101001011" when "010010110", -- t[150] = 843
      "0001101010000" when "010010111", -- t[151] = 848
      "0001101010100" when "010011000", -- t[152] = 852
      "0001101011001" when "010011001", -- t[153] = 857
      "0001101011101" when "010011010", -- t[154] = 861
      "0001101100010" when "010011011", -- t[155] = 866
      "0001101100111" when "010011100", -- t[156] = 871
      "0001101101100" when "010011101", -- t[157] = 876
      "0001101110000" when "010011110", -- t[158] = 880
      "0001101110101" when "010011111", -- t[159] = 885
      "0001101111010" when "010100000", -- t[160] = 890
      "0001101111111" when "010100001", -- t[161] = 895
      "0001110000100" when "010100010", -- t[162] = 900
      "0001110001000" when "010100011", -- t[163] = 904
      "0001110001101" when "010100100", -- t[164] = 909
      "0001110010010" when "010100101", -- t[165] = 914
      "0001110010111" when "010100110", -- t[166] = 919
      "0001110011100" when "010100111", -- t[167] = 924
      "0001110100001" when "010101000", -- t[168] = 929
      "0001110100110" when "010101001", -- t[169] = 934
      "0001110101011" when "010101010", -- t[170] = 939
      "0001110110000" when "010101011", -- t[171] = 944
      "0001110110110" when "010101100", -- t[172] = 950
      "0001110111011" when "010101101", -- t[173] = 955
      "0001111000000" when "010101110", -- t[174] = 960
      "0001111000101" when "010101111", -- t[175] = 965
      "0001111001010" when "010110000", -- t[176] = 970
      "0001111010000" when "010110001", -- t[177] = 976
      "0001111010101" when "010110010", -- t[178] = 981
      "0001111011010" when "010110011", -- t[179] = 986
      "0001111100000" when "010110100", -- t[180] = 992
      "0001111100101" when "010110101", -- t[181] = 997
      "0001111101010" when "010110110", -- t[182] = 1002
      "0001111110000" when "010110111", -- t[183] = 1008
      "0001111110101" when "010111000", -- t[184] = 1013
      "0001111111011" when "010111001", -- t[185] = 1019
      "0010000000000" when "010111010", -- t[186] = 1024
      "0010000000110" when "010111011", -- t[187] = 1030
      "0010000001100" when "010111100", -- t[188] = 1036
      "0010000010001" when "010111101", -- t[189] = 1041
      "0010000010111" when "010111110", -- t[190] = 1047
      "0010000011101" when "010111111", -- t[191] = 1053
      "0010000100010" when "011000000", -- t[192] = 1058
      "0010000101000" when "011000001", -- t[193] = 1064
      "0010000101110" when "011000010", -- t[194] = 1070
      "0010000110100" when "011000011", -- t[195] = 1076
      "0010000111001" when "011000100", -- t[196] = 1081
      "0010000111111" when "011000101", -- t[197] = 1087
      "0010001000101" when "011000110", -- t[198] = 1093
      "0010001001011" when "011000111", -- t[199] = 1099
      "0010001010001" when "011001000", -- t[200] = 1105
      "0010001010111" when "011001001", -- t[201] = 1111
      "0010001011101" when "011001010", -- t[202] = 1117
      "0010001100011" when "011001011", -- t[203] = 1123
      "0010001101001" when "011001100", -- t[204] = 1129
      "0010001110000" when "011001101", -- t[205] = 1136
      "0010001110110" when "011001110", -- t[206] = 1142
      "0010001111100" when "011001111", -- t[207] = 1148
      "0010010000010" when "011010000", -- t[208] = 1154
      "0010010001000" when "011010001", -- t[209] = 1160
      "0010010001111" when "011010010", -- t[210] = 1167
      "0010010010101" when "011010011", -- t[211] = 1173
      "0010010011011" when "011010100", -- t[212] = 1179
      "0010010100010" when "011010101", -- t[213] = 1186
      "0010010101000" when "011010110", -- t[214] = 1192
      "0010010101111" when "011010111", -- t[215] = 1199
      "0010010110101" when "011011000", -- t[216] = 1205
      "0010010111100" when "011011001", -- t[217] = 1212
      "0010011000011" when "011011010", -- t[218] = 1219
      "0010011001001" when "011011011", -- t[219] = 1225
      "0010011010000" when "011011100", -- t[220] = 1232
      "0010011010111" when "011011101", -- t[221] = 1239
      "0010011011101" when "011011110", -- t[222] = 1245
      "0010011100100" when "011011111", -- t[223] = 1252
      "0010011101011" when "011100000", -- t[224] = 1259
      "0010011110010" when "011100001", -- t[225] = 1266
      "0010011111001" when "011100010", -- t[226] = 1273
      "0010100000000" when "011100011", -- t[227] = 1280
      "0010100000111" when "011100100", -- t[228] = 1287
      "0010100001110" when "011100101", -- t[229] = 1294
      "0010100010101" when "011100110", -- t[230] = 1301
      "0010100011100" when "011100111", -- t[231] = 1308
      "0010100100011" when "011101000", -- t[232] = 1315
      "0010100101010" when "011101001", -- t[233] = 1322
      "0010100110001" when "011101010", -- t[234] = 1329
      "0010100111000" when "011101011", -- t[235] = 1336
      "0010101000000" when "011101100", -- t[236] = 1344
      "0010101000111" when "011101101", -- t[237] = 1351
      "0010101001110" when "011101110", -- t[238] = 1358
      "0010101010110" when "011101111", -- t[239] = 1366
      "0010101011101" when "011110000", -- t[240] = 1373
      "0010101100101" when "011110001", -- t[241] = 1381
      "0010101101100" when "011110010", -- t[242] = 1388
      "0010101110100" when "011110011", -- t[243] = 1396
      "0010101111011" when "011110100", -- t[244] = 1403
      "0010110000011" when "011110101", -- t[245] = 1411
      "0010110001011" when "011110110", -- t[246] = 1419
      "0010110010010" when "011110111", -- t[247] = 1426
      "0010110011010" when "011111000", -- t[248] = 1434
      "0010110100010" when "011111001", -- t[249] = 1442
      "0010110101010" when "011111010", -- t[250] = 1450
      "0010110110010" when "011111011", -- t[251] = 1458
      "0010110111010" when "011111100", -- t[252] = 1466
      "0010111000010" when "011111101", -- t[253] = 1474
      "0010111001010" when "011111110", -- t[254] = 1482
      "0010111010010" when "011111111", -- t[255] = 1490
      "0010111011010" when "100000000", -- t[256] = 1498
      "0010111100010" when "100000001", -- t[257] = 1506
      "0010111101010" when "100000010", -- t[258] = 1514
      "0010111110011" when "100000011", -- t[259] = 1523
      "0010111111011" when "100000100", -- t[260] = 1531
      "0011000000011" when "100000101", -- t[261] = 1539
      "0011000001100" when "100000110", -- t[262] = 1548
      "0011000010100" when "100000111", -- t[263] = 1556
      "0011000011101" when "100001000", -- t[264] = 1565
      "0011000100101" when "100001001", -- t[265] = 1573
      "0011000101110" when "100001010", -- t[266] = 1582
      "0011000110110" when "100001011", -- t[267] = 1590
      "0011000111111" when "100001100", -- t[268] = 1599
      "0011001001000" when "100001101", -- t[269] = 1608
      "0011001010001" when "100001110", -- t[270] = 1617
      "0011001011001" when "100001111", -- t[271] = 1625
      "0011001100010" when "100010000", -- t[272] = 1634
      "0011001101011" when "100010001", -- t[273] = 1643
      "0011001110100" when "100010010", -- t[274] = 1652
      "0011001111101" when "100010011", -- t[275] = 1661
      "0011010000110" when "100010100", -- t[276] = 1670
      "0011010001111" when "100010101", -- t[277] = 1679
      "0011010011001" when "100010110", -- t[278] = 1689
      "0011010100010" when "100010111", -- t[279] = 1698
      "0011010101011" when "100011000", -- t[280] = 1707
      "0011010110100" when "100011001", -- t[281] = 1716
      "0011010111110" when "100011010", -- t[282] = 1726
      "0011011000111" when "100011011", -- t[283] = 1735
      "0011011010001" when "100011100", -- t[284] = 1745
      "0011011011010" when "100011101", -- t[285] = 1754
      "0011011100100" when "100011110", -- t[286] = 1764
      "0011011101101" when "100011111", -- t[287] = 1773
      "0011011110111" when "100100000", -- t[288] = 1783
      "0011100000001" when "100100001", -- t[289] = 1793
      "0011100001011" when "100100010", -- t[290] = 1803
      "0011100010101" when "100100011", -- t[291] = 1813
      "0011100011110" when "100100100", -- t[292] = 1822
      "0011100101000" when "100100101", -- t[293] = 1832
      "0011100110010" when "100100110", -- t[294] = 1842
      "0011100111101" when "100100111", -- t[295] = 1853
      "0011101000111" when "100101000", -- t[296] = 1863
      "0011101010001" when "100101001", -- t[297] = 1873
      "0011101011011" when "100101010", -- t[298] = 1883
      "0011101100101" when "100101011", -- t[299] = 1893
      "0011101110000" when "100101100", -- t[300] = 1904
      "0011101111010" when "100101101", -- t[301] = 1914
      "0011110000101" when "100101110", -- t[302] = 1925
      "0011110001111" when "100101111", -- t[303] = 1935
      "0011110011010" when "100110000", -- t[304] = 1946
      "0011110100100" when "100110001", -- t[305] = 1956
      "0011110101111" when "100110010", -- t[306] = 1967
      "0011110111010" when "100110011", -- t[307] = 1978
      "0011111000101" when "100110100", -- t[308] = 1989
      "0011111010000" when "100110101", -- t[309] = 2000
      "0011111011011" when "100110110", -- t[310] = 2011
      "0011111100110" when "100110111", -- t[311] = 2022
      "0011111110001" when "100111000", -- t[312] = 2033
      "0011111111100" when "100111001", -- t[313] = 2044
      "0100000000111" when "100111010", -- t[314] = 2055
      "0100000010010" when "100111011", -- t[315] = 2066
      "0100000011101" when "100111100", -- t[316] = 2077
      "0100000101001" when "100111101", -- t[317] = 2089
      "0100000110100" when "100111110", -- t[318] = 2100
      "0100001000000" when "100111111", -- t[319] = 2112
      "0100001001011" when "101000000", -- t[320] = 2123
      "0100001010111" when "101000001", -- t[321] = 2135
      "0100001100011" when "101000010", -- t[322] = 2147
      "0100001101110" when "101000011", -- t[323] = 2158
      "0100001111010" when "101000100", -- t[324] = 2170
      "0100010000110" when "101000101", -- t[325] = 2182
      "0100010010010" when "101000110", -- t[326] = 2194
      "0100010011110" when "101000111", -- t[327] = 2206
      "0100010101010" when "101001000", -- t[328] = 2218
      "0100010110110" when "101001001", -- t[329] = 2230
      "0100011000011" when "101001010", -- t[330] = 2243
      "0100011001111" when "101001011", -- t[331] = 2255
      "0100011011011" when "101001100", -- t[332] = 2267
      "0100011101000" when "101001101", -- t[333] = 2280
      "0100011110100" when "101001110", -- t[334] = 2292
      "0100100000001" when "101001111", -- t[335] = 2305
      "0100100001101" when "101010000", -- t[336] = 2317
      "0100100011010" when "101010001", -- t[337] = 2330
      "0100100100111" when "101010010", -- t[338] = 2343
      "0100100110100" when "101010011", -- t[339] = 2356
      "0100101000001" when "101010100", -- t[340] = 2369
      "0100101001110" when "101010101", -- t[341] = 2382
      "0100101011011" when "101010110", -- t[342] = 2395
      "0100101101000" when "101010111", -- t[343] = 2408
      "0100101110101" when "101011000", -- t[344] = 2421
      "0100110000010" when "101011001", -- t[345] = 2434
      "0100110010000" when "101011010", -- t[346] = 2448
      "0100110011101" when "101011011", -- t[347] = 2461
      "0100110101011" when "101011100", -- t[348] = 2475
      "0100110111000" when "101011101", -- t[349] = 2488
      "0100111000110" when "101011110", -- t[350] = 2502
      "0100111010100" when "101011111", -- t[351] = 2516
      "0100111100010" when "101100000", -- t[352] = 2530
      "0100111101111" when "101100001", -- t[353] = 2543
      "0100111111101" when "101100010", -- t[354] = 2557
      "0101000001100" when "101100011", -- t[355] = 2572
      "0101000011010" when "101100100", -- t[356] = 2586
      "0101000101000" when "101100101", -- t[357] = 2600
      "0101000110110" when "101100110", -- t[358] = 2614
      "0101001000100" when "101100111", -- t[359] = 2628
      "0101001010011" when "101101000", -- t[360] = 2643
      "0101001100001" when "101101001", -- t[361] = 2657
      "0101001110000" when "101101010", -- t[362] = 2672
      "0101001111111" when "101101011", -- t[363] = 2687
      "0101010001110" when "101101100", -- t[364] = 2702
      "0101010011100" when "101101101", -- t[365] = 2716
      "0101010101011" when "101101110", -- t[366] = 2731
      "0101010111010" when "101101111", -- t[367] = 2746
      "0101011001001" when "101110000", -- t[368] = 2761
      "0101011011001" when "101110001", -- t[369] = 2777
      "0101011101000" when "101110010", -- t[370] = 2792
      "0101011110111" when "101110011", -- t[371] = 2807
      "0101100000111" when "101110100", -- t[372] = 2823
      "0101100010110" when "101110101", -- t[373] = 2838
      "0101100100110" when "101110110", -- t[374] = 2854
      "0101100110110" when "101110111", -- t[375] = 2870
      "0101101000101" when "101111000", -- t[376] = 2885
      "0101101010101" when "101111001", -- t[377] = 2901
      "0101101100101" when "101111010", -- t[378] = 2917
      "0101101110101" when "101111011", -- t[379] = 2933
      "0101110000101" when "101111100", -- t[380] = 2949
      "0101110010110" when "101111101", -- t[381] = 2966
      "0101110100110" when "101111110", -- t[382] = 2982
      "0101110110110" when "101111111", -- t[383] = 2998
      "0101111000111" when "110000000", -- t[384] = 3015
      "0101111011000" when "110000001", -- t[385] = 3032
      "0101111101000" when "110000010", -- t[386] = 3048
      "0101111111001" when "110000011", -- t[387] = 3065
      "0110000001010" when "110000100", -- t[388] = 3082
      "0110000011011" when "110000101", -- t[389] = 3099
      "0110000101100" when "110000110", -- t[390] = 3116
      "0110000111101" when "110000111", -- t[391] = 3133
      "0110001001110" when "110001000", -- t[392] = 3150
      "0110001100000" when "110001001", -- t[393] = 3168
      "0110001110001" when "110001010", -- t[394] = 3185
      "0110010000011" when "110001011", -- t[395] = 3203
      "0110010010101" when "110001100", -- t[396] = 3221
      "0110010100110" when "110001101", -- t[397] = 3238
      "0110010111000" when "110001110", -- t[398] = 3256
      "0110011001010" when "110001111", -- t[399] = 3274
      "0110011011100" when "110010000", -- t[400] = 3292
      "0110011101110" when "110010001", -- t[401] = 3310
      "0110100000001" when "110010010", -- t[402] = 3329
      "0110100010011" when "110010011", -- t[403] = 3347
      "0110100100101" when "110010100", -- t[404] = 3365
      "0110100111000" when "110010101", -- t[405] = 3384
      "0110101001011" when "110010110", -- t[406] = 3403
      "0110101011101" when "110010111", -- t[407] = 3421
      "0110101110000" when "110011000", -- t[408] = 3440
      "0110110000011" when "110011001", -- t[409] = 3459
      "0110110010110" when "110011010", -- t[410] = 3478
      "0110110101010" when "110011011", -- t[411] = 3498
      "0110110111101" when "110011100", -- t[412] = 3517
      "0110111010000" when "110011101", -- t[413] = 3536
      "0110111100100" when "110011110", -- t[414] = 3556
      "0110111111000" when "110011111", -- t[415] = 3576
      "0111000001011" when "110100000", -- t[416] = 3595
      "0111000011111" when "110100001", -- t[417] = 3615
      "0111000110011" when "110100010", -- t[418] = 3635
      "0111001000111" when "110100011", -- t[419] = 3655
      "0111001011100" when "110100100", -- t[420] = 3676
      "0111001110000" when "110100101", -- t[421] = 3696
      "0111010000100" when "110100110", -- t[422] = 3716
      "0111010011001" when "110100111", -- t[423] = 3737
      "0111010101110" when "110101000", -- t[424] = 3758
      "0111011000010" when "110101001", -- t[425] = 3778
      "0111011010111" when "110101010", -- t[426] = 3799
      "0111011101100" when "110101011", -- t[427] = 3820
      "0111100000001" when "110101100", -- t[428] = 3841
      "0111100010111" when "110101101", -- t[429] = 3863
      "0111100101100" when "110101110", -- t[430] = 3884
      "0111101000010" when "110101111", -- t[431] = 3906
      "0111101010111" when "110110000", -- t[432] = 3927
      "0111101101101" when "110110001", -- t[433] = 3949
      "0111110000011" when "110110010", -- t[434] = 3971
      "0111110011001" when "110110011", -- t[435] = 3993
      "0111110101111" when "110110100", -- t[436] = 4015
      "0111111000101" when "110110101", -- t[437] = 4037
      "0111111011100" when "110110110", -- t[438] = 4060
      "0111111110010" when "110110111", -- t[439] = 4082
      "1000000001001" when "110111000", -- t[440] = 4105
      "1000000011111" when "110111001", -- t[441] = 4127
      "1000000110110" when "110111010", -- t[442] = 4150
      "1000001001101" when "110111011", -- t[443] = 4173
      "1000001100100" when "110111100", -- t[444] = 4196
      "1000001111100" when "110111101", -- t[445] = 4220
      "1000010010011" when "110111110", -- t[446] = 4243
      "1000010101011" when "110111111", -- t[447] = 4267
      "1000011000010" when "111000000", -- t[448] = 4290
      "1000011011010" when "111000001", -- t[449] = 4314
      "1000011110010" when "111000010", -- t[450] = 4338
      "1000100001010" when "111000011", -- t[451] = 4362
      "1000100100010" when "111000100", -- t[452] = 4386
      "1000100111011" when "111000101", -- t[453] = 4411
      "1000101010011" when "111000110", -- t[454] = 4435
      "1000101101100" when "111000111", -- t[455] = 4460
      "1000110000101" when "111001000", -- t[456] = 4485
      "1000110011110" when "111001001", -- t[457] = 4510
      "1000110110111" when "111001010", -- t[458] = 4535
      "1000111010000" when "111001011", -- t[459] = 4560
      "1000111101001" when "111001100", -- t[460] = 4585
      "1001000000011" when "111001101", -- t[461] = 4611
      "1001000011100" when "111001110", -- t[462] = 4636
      "1001000110110" when "111001111", -- t[463] = 4662
      "1001001010000" when "111010000", -- t[464] = 4688
      "1001001101010" when "111010001", -- t[465] = 4714
      "1001010000100" when "111010010", -- t[466] = 4740
      "1001010011111" when "111010011", -- t[467] = 4767
      "1001010111001" when "111010100", -- t[468] = 4793
      "1001011010100" when "111010101", -- t[469] = 4820
      "1001011101111" when "111010110", -- t[470] = 4847
      "1001100001010" when "111010111", -- t[471] = 4874
      "1001100100101" when "111011000", -- t[472] = 4901
      "1001101000000" when "111011001", -- t[473] = 4928
      "1001101011011" when "111011010", -- t[474] = 4955
      "1001101110111" when "111011011", -- t[475] = 4983
      "1001110010011" when "111011100", -- t[476] = 5011
      "1001110101111" when "111011101", -- t[477] = 5039
      "1001111001011" when "111011110", -- t[478] = 5067
      "1001111100111" when "111011111", -- t[479] = 5095
      "1010000000011" when "111100000", -- t[480] = 5123
      "1010000100000" when "111100001", -- t[481] = 5152
      "1010000111101" when "111100010", -- t[482] = 5181
      "1010001011010" when "111100011", -- t[483] = 5210
      "1010001110111" when "111100100", -- t[484] = 5239
      "1010010010100" when "111100101", -- t[485] = 5268
      "1010010110001" when "111100110", -- t[486] = 5297
      "1010011001111" when "111100111", -- t[487] = 5327
      "1010011101101" when "111101000", -- t[488] = 5357
      "1010100001010" when "111101001", -- t[489] = 5386
      "1010100101001" when "111101010", -- t[490] = 5417
      "1010101000111" when "111101011", -- t[491] = 5447
      "1010101100101" when "111101100", -- t[492] = 5477
      "1010110000100" when "111101101", -- t[493] = 5508
      "1010110100011" when "111101110", -- t[494] = 5539
      "1010111000010" when "111101111", -- t[495] = 5570
      "1010111100001" when "111110000", -- t[496] = 5601
      "1011000000000" when "111110001", -- t[497] = 5632
      "1011000011111" when "111110010", -- t[498] = 5663
      "1011000111111" when "111110011", -- t[499] = 5695
      "1011001011111" when "111110100", -- t[500] = 5727
      "1011001111111" when "111110101", -- t[501] = 5759
      "1011010011111" when "111110110", -- t[502] = 5791
      "1011011000000" when "111110111", -- t[503] = 5824
      "1011011100000" when "111111000", -- t[504] = 5856
      "1011100000001" when "111111001", -- t[505] = 5889
      "1011100100010" when "111111010", -- t[506] = 5922
      "1011101000011" when "111111011", -- t[507] = 5955
      "1011101100101" when "111111100", -- t[508] = 5989
      "1011110000110" when "111111101", -- t[509] = 6022
      "1011110101000" when "111111110", -- t[510] = 6056
      "1011111001010" when "111111111", -- t[511] = 6090
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_13_to2 is
  port( x : in  std_logic_vector(7 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to2 is
begin
  with x select
    r <=
      "0000" when "00000000", -- t[0] = 0
      "0000" when "00000001", -- t[1] = 0
      "0000" when "00000010", -- t[2] = 0
      "0000" when "00000011", -- t[3] = 0
      "0000" when "00000100", -- t[4] = 0
      "0000" when "00000101", -- t[5] = 0
      "0000" when "00000110", -- t[6] = 0
      "0000" when "00000111", -- t[7] = 0
      "0000" when "00001000", -- t[8] = 0
      "0000" when "00001001", -- t[9] = 0
      "0000" when "00001010", -- t[10] = 0
      "0000" when "00001011", -- t[11] = 0
      "0000" when "00001100", -- t[12] = 0
      "0000" when "00001101", -- t[13] = 0
      "0000" when "00001110", -- t[14] = 0
      "0000" when "00001111", -- t[15] = 0
      "0000" when "00010000", -- t[16] = 0
      "0000" when "00010001", -- t[17] = 0
      "0000" when "00010010", -- t[18] = 0
      "0000" when "00010011", -- t[19] = 0
      "0000" when "00010100", -- t[20] = 0
      "0000" when "00010101", -- t[21] = 0
      "0000" when "00010110", -- t[22] = 0
      "0000" when "00010111", -- t[23] = 0
      "0000" when "00011000", -- t[24] = 0
      "0000" when "00011001", -- t[25] = 0
      "0000" when "00011010", -- t[26] = 0
      "0001" when "00011011", -- t[27] = 1
      "0000" when "00011100", -- t[28] = 0
      "0001" when "00011101", -- t[29] = 1
      "0000" when "00011110", -- t[30] = 0
      "0001" when "00011111", -- t[31] = 1
      "0000" when "00100000", -- t[32] = 0
      "0001" when "00100001", -- t[33] = 1
      "0000" when "00100010", -- t[34] = 0
      "0001" when "00100011", -- t[35] = 1
      "0000" when "00100100", -- t[36] = 0
      "0001" when "00100101", -- t[37] = 1
      "0000" when "00100110", -- t[38] = 0
      "0001" when "00100111", -- t[39] = 1
      "0000" when "00101000", -- t[40] = 0
      "0001" when "00101001", -- t[41] = 1
      "0000" when "00101010", -- t[42] = 0
      "0001" when "00101011", -- t[43] = 1
      "0000" when "00101100", -- t[44] = 0
      "0001" when "00101101", -- t[45] = 1
      "0000" when "00101110", -- t[46] = 0
      "0001" when "00101111", -- t[47] = 1
      "0000" when "00110000", -- t[48] = 0
      "0001" when "00110001", -- t[49] = 1
      "0000" when "00110010", -- t[50] = 0
      "0001" when "00110011", -- t[51] = 1
      "0000" when "00110100", -- t[52] = 0
      "0001" when "00110101", -- t[53] = 1
      "0000" when "00110110", -- t[54] = 0
      "0001" when "00110111", -- t[55] = 1
      "0000" when "00111000", -- t[56] = 0
      "0001" when "00111001", -- t[57] = 1
      "0000" when "00111010", -- t[58] = 0
      "0001" when "00111011", -- t[59] = 1
      "0000" when "00111100", -- t[60] = 0
      "0001" when "00111101", -- t[61] = 1
      "0000" when "00111110", -- t[62] = 0
      "0001" when "00111111", -- t[63] = 1
      "0000" when "01000000", -- t[64] = 0
      "0001" when "01000001", -- t[65] = 1
      "0000" when "01000010", -- t[66] = 0
      "0001" when "01000011", -- t[67] = 1
      "0000" when "01000100", -- t[68] = 0
      "0001" when "01000101", -- t[69] = 1
      "0000" when "01000110", -- t[70] = 0
      "0001" when "01000111", -- t[71] = 1
      "0000" when "01001000", -- t[72] = 0
      "0001" when "01001001", -- t[73] = 1
      "0000" when "01001010", -- t[74] = 0
      "0001" when "01001011", -- t[75] = 1
      "0000" when "01001100", -- t[76] = 0
      "0001" when "01001101", -- t[77] = 1
      "0000" when "01001110", -- t[78] = 0
      "0001" when "01001111", -- t[79] = 1
      "0000" when "01010000", -- t[80] = 0
      "0001" when "01010001", -- t[81] = 1
      "0000" when "01010010", -- t[82] = 0
      "0001" when "01010011", -- t[83] = 1
      "0000" when "01010100", -- t[84] = 0
      "0001" when "01010101", -- t[85] = 1
      "0000" when "01010110", -- t[86] = 0
      "0001" when "01010111", -- t[87] = 1
      "0000" when "01011000", -- t[88] = 0
      "0001" when "01011001", -- t[89] = 1
      "0000" when "01011010", -- t[90] = 0
      "0010" when "01011011", -- t[91] = 2
      "0000" when "01011100", -- t[92] = 0
      "0010" when "01011101", -- t[93] = 2
      "0000" when "01011110", -- t[94] = 0
      "0010" when "01011111", -- t[95] = 2
      "0000" when "01100000", -- t[96] = 0
      "0010" when "01100001", -- t[97] = 2
      "0000" when "01100010", -- t[98] = 0
      "0010" when "01100011", -- t[99] = 2
      "0000" when "01100100", -- t[100] = 0
      "0010" when "01100101", -- t[101] = 2
      "0000" when "01100110", -- t[102] = 0
      "0010" when "01100111", -- t[103] = 2
      "0000" when "01101000", -- t[104] = 0
      "0010" when "01101001", -- t[105] = 2
      "0000" when "01101010", -- t[106] = 0
      "0010" when "01101011", -- t[107] = 2
      "0000" when "01101100", -- t[108] = 0
      "0010" when "01101101", -- t[109] = 2
      "0000" when "01101110", -- t[110] = 0
      "0010" when "01101111", -- t[111] = 2
      "0000" when "01110000", -- t[112] = 0
      "0010" when "01110001", -- t[113] = 2
      "0000" when "01110010", -- t[114] = 0
      "0010" when "01110011", -- t[115] = 2
      "0000" when "01110100", -- t[116] = 0
      "0010" when "01110101", -- t[117] = 2
      "0000" when "01110110", -- t[118] = 0
      "0010" when "01110111", -- t[119] = 2
      "0000" when "01111000", -- t[120] = 0
      "0010" when "01111001", -- t[121] = 2
      "0000" when "01111010", -- t[122] = 0
      "0010" when "01111011", -- t[123] = 2
      "0000" when "01111100", -- t[124] = 0
      "0010" when "01111101", -- t[125] = 2
      "0001" when "01111110", -- t[126] = 1
      "0011" when "01111111", -- t[127] = 3
      "0001" when "10000000", -- t[128] = 1
      "0011" when "10000001", -- t[129] = 3
      "0001" when "10000010", -- t[130] = 1
      "0011" when "10000011", -- t[131] = 3
      "0001" when "10000100", -- t[132] = 1
      "0011" when "10000101", -- t[133] = 3
      "0001" when "10000110", -- t[134] = 1
      "0011" when "10000111", -- t[135] = 3
      "0001" when "10001000", -- t[136] = 1
      "0011" when "10001001", -- t[137] = 3
      "0001" when "10001010", -- t[138] = 1
      "0011" when "10001011", -- t[139] = 3
      "0001" when "10001100", -- t[140] = 1
      "0011" when "10001101", -- t[141] = 3
      "0001" when "10001110", -- t[142] = 1
      "0011" when "10001111", -- t[143] = 3
      "0001" when "10010000", -- t[144] = 1
      "0011" when "10010001", -- t[145] = 3
      "0001" when "10010010", -- t[146] = 1
      "0011" when "10010011", -- t[147] = 3
      "0001" when "10010100", -- t[148] = 1
      "0011" when "10010101", -- t[149] = 3
      "0001" when "10010110", -- t[150] = 1
      "0011" when "10010111", -- t[151] = 3
      "0001" when "10011000", -- t[152] = 1
      "0100" when "10011001", -- t[153] = 4
      "0001" when "10011010", -- t[154] = 1
      "0100" when "10011011", -- t[155] = 4
      "0001" when "10011100", -- t[156] = 1
      "0100" when "10011101", -- t[157] = 4
      "0001" when "10011110", -- t[158] = 1
      "0100" when "10011111", -- t[159] = 4
      "0001" when "10100000", -- t[160] = 1
      "0100" when "10100001", -- t[161] = 4
      "0001" when "10100010", -- t[162] = 1
      "0100" when "10100011", -- t[163] = 4
      "0001" when "10100100", -- t[164] = 1
      "0100" when "10100101", -- t[165] = 4
      "0001" when "10100110", -- t[166] = 1
      "0100" when "10100111", -- t[167] = 4
      "0001" when "10101000", -- t[168] = 1
      "0100" when "10101001", -- t[169] = 4
      "0001" when "10101010", -- t[170] = 1
      "0100" when "10101011", -- t[171] = 4
      "0001" when "10101100", -- t[172] = 1
      "0101" when "10101101", -- t[173] = 5
      "0001" when "10101110", -- t[174] = 1
      "0101" when "10101111", -- t[175] = 5
      "0001" when "10110000", -- t[176] = 1
      "0101" when "10110001", -- t[177] = 5
      "0001" when "10110010", -- t[178] = 1
      "0101" when "10110011", -- t[179] = 5
      "0001" when "10110100", -- t[180] = 1
      "0101" when "10110101", -- t[181] = 5
      "0001" when "10110110", -- t[182] = 1
      "0101" when "10110111", -- t[183] = 5
      "0001" when "10111000", -- t[184] = 1
      "0101" when "10111001", -- t[185] = 5
      "0001" when "10111010", -- t[186] = 1
      "0101" when "10111011", -- t[187] = 5
      "0001" when "10111100", -- t[188] = 1
      "0101" when "10111101", -- t[189] = 5
      "0010" when "10111110", -- t[190] = 2
      "0110" when "10111111", -- t[191] = 6
      "0010" when "11000000", -- t[192] = 2
      "0110" when "11000001", -- t[193] = 6
      "0010" when "11000010", -- t[194] = 2
      "0110" when "11000011", -- t[195] = 6
      "0010" when "11000100", -- t[196] = 2
      "0110" when "11000101", -- t[197] = 6
      "0010" when "11000110", -- t[198] = 2
      "0110" when "11000111", -- t[199] = 6
      "0010" when "11001000", -- t[200] = 2
      "0110" when "11001001", -- t[201] = 6
      "0010" when "11001010", -- t[202] = 2
      "0111" when "11001011", -- t[203] = 7
      "0010" when "11001100", -- t[204] = 2
      "0111" when "11001101", -- t[205] = 7
      "0010" when "11001110", -- t[206] = 2
      "0111" when "11001111", -- t[207] = 7
      "0010" when "11010000", -- t[208] = 2
      "0111" when "11010001", -- t[209] = 7
      "0010" when "11010010", -- t[210] = 2
      "0111" when "11010011", -- t[211] = 7
      "0010" when "11010100", -- t[212] = 2
      "0111" when "11010101", -- t[213] = 7
      "0010" when "11010110", -- t[214] = 2
      "1000" when "11010111", -- t[215] = 8
      "0010" when "11011000", -- t[216] = 2
      "1000" when "11011001", -- t[217] = 8
      "0010" when "11011010", -- t[218] = 2
      "1000" when "11011011", -- t[219] = 8
      "0010" when "11011100", -- t[220] = 2
      "1000" when "11011101", -- t[221] = 8
      "0010" when "11011110", -- t[222] = 2
      "1000" when "11011111", -- t[223] = 8
      "0010" when "11100000", -- t[224] = 2
      "1000" when "11100001", -- t[225] = 8
      "0011" when "11100010", -- t[226] = 3
      "1001" when "11100011", -- t[227] = 9
      "0011" when "11100100", -- t[228] = 3
      "1001" when "11100101", -- t[229] = 9
      "0011" when "11100110", -- t[230] = 3
      "1001" when "11100111", -- t[231] = 9
      "0011" when "11101000", -- t[232] = 3
      "1001" when "11101001", -- t[233] = 9
      "0011" when "11101010", -- t[234] = 3
      "1010" when "11101011", -- t[235] = 10
      "0011" when "11101100", -- t[236] = 3
      "1010" when "11101101", -- t[237] = 10
      "0011" when "11101110", -- t[238] = 3
      "1010" when "11101111", -- t[239] = 10
      "0011" when "11110000", -- t[240] = 3
      "1010" when "11110001", -- t[241] = 10
      "0011" when "11110010", -- t[242] = 3
      "1011" when "11110011", -- t[243] = 11
      "0011" when "11110100", -- t[244] = 3
      "1011" when "11110101", -- t[245] = 11
      "0011" when "11110110", -- t[246] = 3
      "1011" when "11110111", -- t[247] = 11
      "0011" when "11111000", -- t[248] = 3
      "1011" when "11111001", -- t[249] = 11
      "0100" when "11111010", -- t[250] = 4
      "1100" when "11111011", -- t[251] = 12
      "0100" when "11111100", -- t[252] = 4
      "1100" when "11111101", -- t[253] = 12
      "0100" when "11111110", -- t[254] = 4
      "1100" when "11111111", -- t[255] = 12
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_13_to1 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to1 is
begin
  with x select
    r <=
      "00" when "0000000", -- t[0] = 0
      "00" when "0000001", -- t[1] = 0
      "00" when "0000010", -- t[2] = 0
      "00" when "0000011", -- t[3] = 0
      "00" when "0000100", -- t[4] = 0
      "00" when "0000101", -- t[5] = 0
      "00" when "0000110", -- t[6] = 0
      "00" when "0000111", -- t[7] = 0
      "00" when "0001000", -- t[8] = 0
      "00" when "0001001", -- t[9] = 0
      "00" when "0001010", -- t[10] = 0
      "00" when "0001011", -- t[11] = 0
      "00" when "0001100", -- t[12] = 0
      "00" when "0001101", -- t[13] = 0
      "00" when "0001110", -- t[14] = 0
      "00" when "0001111", -- t[15] = 0
      "00" when "0010000", -- t[16] = 0
      "00" when "0010001", -- t[17] = 0
      "00" when "0010010", -- t[18] = 0
      "00" when "0010011", -- t[19] = 0
      "00" when "0010100", -- t[20] = 0
      "00" when "0010101", -- t[21] = 0
      "00" when "0010110", -- t[22] = 0
      "00" when "0010111", -- t[23] = 0
      "00" when "0011000", -- t[24] = 0
      "00" when "0011001", -- t[25] = 0
      "00" when "0011010", -- t[26] = 0
      "00" when "0011011", -- t[27] = 0
      "00" when "0011100", -- t[28] = 0
      "00" when "0011101", -- t[29] = 0
      "00" when "0011110", -- t[30] = 0
      "00" when "0011111", -- t[31] = 0
      "00" when "0100000", -- t[32] = 0
      "00" when "0100001", -- t[33] = 0
      "00" when "0100010", -- t[34] = 0
      "00" when "0100011", -- t[35] = 0
      "00" when "0100100", -- t[36] = 0
      "00" when "0100101", -- t[37] = 0
      "00" when "0100110", -- t[38] = 0
      "00" when "0100111", -- t[39] = 0
      "00" when "0101000", -- t[40] = 0
      "00" when "0101001", -- t[41] = 0
      "00" when "0101010", -- t[42] = 0
      "00" when "0101011", -- t[43] = 0
      "00" when "0101100", -- t[44] = 0
      "00" when "0101101", -- t[45] = 0
      "00" when "0101110", -- t[46] = 0
      "00" when "0101111", -- t[47] = 0
      "00" when "0110000", -- t[48] = 0
      "00" when "0110001", -- t[49] = 0
      "00" when "0110010", -- t[50] = 0
      "00" when "0110011", -- t[51] = 0
      "00" when "0110100", -- t[52] = 0
      "00" when "0110101", -- t[53] = 0
      "00" when "0110110", -- t[54] = 0
      "00" when "0110111", -- t[55] = 0
      "00" when "0111000", -- t[56] = 0
      "00" when "0111001", -- t[57] = 0
      "00" when "0111010", -- t[58] = 0
      "00" when "0111011", -- t[59] = 0
      "00" when "0111100", -- t[60] = 0
      "00" when "0111101", -- t[61] = 0
      "00" when "0111110", -- t[62] = 0
      "00" when "0111111", -- t[63] = 0
      "00" when "1000000", -- t[64] = 0
      "00" when "1000001", -- t[65] = 0
      "00" when "1000010", -- t[66] = 0
      "00" when "1000011", -- t[67] = 0
      "00" when "1000100", -- t[68] = 0
      "00" when "1000101", -- t[69] = 0
      "00" when "1000110", -- t[70] = 0
      "00" when "1000111", -- t[71] = 0
      "00" when "1001000", -- t[72] = 0
      "00" when "1001001", -- t[73] = 0
      "00" when "1001010", -- t[74] = 0
      "00" when "1001011", -- t[75] = 0
      "00" when "1001100", -- t[76] = 0
      "01" when "1001101", -- t[77] = 1
      "00" when "1001110", -- t[78] = 0
      "01" when "1001111", -- t[79] = 1
      "00" when "1010000", -- t[80] = 0
      "01" when "1010001", -- t[81] = 1
      "00" when "1010010", -- t[82] = 0
      "01" when "1010011", -- t[83] = 1
      "00" when "1010100", -- t[84] = 0
      "01" when "1010101", -- t[85] = 1
      "00" when "1010110", -- t[86] = 0
      "01" when "1010111", -- t[87] = 1
      "00" when "1011000", -- t[88] = 0
      "01" when "1011001", -- t[89] = 1
      "00" when "1011010", -- t[90] = 0
      "01" when "1011011", -- t[91] = 1
      "00" when "1011100", -- t[92] = 0
      "01" when "1011101", -- t[93] = 1
      "00" when "1011110", -- t[94] = 0
      "01" when "1011111", -- t[95] = 1
      "00" when "1100000", -- t[96] = 0
      "01" when "1100001", -- t[97] = 1
      "00" when "1100010", -- t[98] = 0
      "01" when "1100011", -- t[99] = 1
      "00" when "1100100", -- t[100] = 0
      "01" when "1100101", -- t[101] = 1
      "00" when "1100110", -- t[102] = 0
      "01" when "1100111", -- t[103] = 1
      "00" when "1101000", -- t[104] = 0
      "01" when "1101001", -- t[105] = 1
      "00" when "1101010", -- t[106] = 0
      "01" when "1101011", -- t[107] = 1
      "00" when "1101100", -- t[108] = 0
      "10" when "1101101", -- t[109] = 2
      "00" when "1101110", -- t[110] = 0
      "10" when "1101111", -- t[111] = 2
      "00" when "1110000", -- t[112] = 0
      "10" when "1110001", -- t[113] = 2
      "00" when "1110010", -- t[114] = 0
      "10" when "1110011", -- t[115] = 2
      "00" when "1110100", -- t[116] = 0
      "10" when "1110101", -- t[117] = 2
      "00" when "1110110", -- t[118] = 0
      "10" when "1110111", -- t[119] = 2
      "00" when "1111000", -- t[120] = 0
      "10" when "1111001", -- t[121] = 2
      "00" when "1111010", -- t[122] = 0
      "10" when "1111011", -- t[123] = 2
      "00" when "1111100", -- t[124] = 0
      "10" when "1111101", -- t[125] = 2
      "01" when "1111110", -- t[126] = 1
      "11" when "1111111", -- t[127] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_13_to0 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to0 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "0" when "1101", -- t[13] = 0
      "0" when "1110", -- t[14] = 0
      "0" when "1111", -- t[15] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_13.all;

entity LNSSub_MPT_T1_13_to2_xor is
  port( a : in  std_logic_vector(6 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(7 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(7 downto 1) <= a(6 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T1_13_to2
    port map( x => in_t,
              r => out_t );

  r(12 downto 4) <= (12 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_13.all;

entity LNSSub_MPT_T1_13_to1_xor is
  port( a : in  std_logic_vector(5 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(6 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(6 downto 1) <= a(5 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T1_13_to1
    port map( x => in_t,
              r => out_t );

  r(12 downto 2) <= (12 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_13.all;

entity LNSSub_MPT_T1_13_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T1_13_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 1) <= (12 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_13.all;

entity LNSSub_MPT_T1_13 is
  port( x : in  std_logic_vector(14 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_13 is
  signal in_tiv  : std_logic_vector(8 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a2      : std_logic_vector(6 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(12 downto 0);
  signal a1      : std_logic_vector(5 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(14 downto 6);
  inst_tiv : LNSSub_MPT_T1_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(14 downto 8);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T1_13_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(14 downto 9);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T1_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(14 downto 12);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T1_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(12 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T1_13_Clk is
  port( x   : in  std_logic_vector(14 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T1_13_Clk is
  signal in_tiv_1  : std_logic_vector(8 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a2_1      : std_logic_vector(6 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(12 downto 0);
  signal out2_2    : std_logic_vector(12 downto 0);
  signal a1_1      : std_logic_vector(5 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(12 downto 0);
  signal out1_2    : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(14 downto 6);
  inst_tiv : LNSSub_MPT_T1_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(14 downto 8);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T1_13_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(14 downto 9);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T1_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(14 downto 12);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T1_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-4.0 -2.0[ -> [0.0 0.5[
-- wI = 14 bits
-- wO = 12 bits
-- Decomposition: 7, 7 / 6, 5, 2 / 2, 3, 2
-- Guard bits: 2
-- Size: 3208 = 14.2^7 + 6.2^7 + 5.2^7 + 1.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T2_13 is
  component LNSSub_MPT_T2_13_tiv is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to2 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to1 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to2_xor is
    port( a : in  std_logic_vector(5 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to1_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MPT_T2_13_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(13 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_13_tiv is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_tiv is
begin
  with x select
    r <=
      "00101111111111" when "0000000", -- t[0] = 3071
      "00110000100010" when "0000001", -- t[1] = 3106
      "00110001000101" when "0000010", -- t[2] = 3141
      "00110001101000" when "0000011", -- t[3] = 3176
      "00110010001100" when "0000100", -- t[4] = 3212
      "00110010110000" when "0000101", -- t[5] = 3248
      "00110011010100" when "0000110", -- t[6] = 3284
      "00110011111001" when "0000111", -- t[7] = 3321
      "00110100011111" when "0001000", -- t[8] = 3359
      "00110101000101" when "0001001", -- t[9] = 3397
      "00110101101011" when "0001010", -- t[10] = 3435
      "00110110010010" when "0001011", -- t[11] = 3474
      "00110110111001" when "0001100", -- t[12] = 3513
      "00110111100001" when "0001101", -- t[13] = 3553
      "00111000001001" when "0001110", -- t[14] = 3593
      "00111000110010" when "0001111", -- t[15] = 3634
      "00111001011011" when "0010000", -- t[16] = 3675
      "00111010000100" when "0010001", -- t[17] = 3716
      "00111010101110" when "0010010", -- t[18] = 3758
      "00111011011001" when "0010011", -- t[19] = 3801
      "00111100000100" when "0010100", -- t[20] = 3844
      "00111100110000" when "0010101", -- t[21] = 3888
      "00111101011100" when "0010110", -- t[22] = 3932
      "00111110001000" when "0010111", -- t[23] = 3976
      "00111110110101" when "0011000", -- t[24] = 4021
      "00111111100011" when "0011001", -- t[25] = 4067
      "01000000010001" when "0011010", -- t[26] = 4113
      "01000001000000" when "0011011", -- t[27] = 4160
      "01000001110000" when "0011100", -- t[28] = 4208
      "01000010011111" when "0011101", -- t[29] = 4255
      "01000011010000" when "0011110", -- t[30] = 4304
      "01000100000001" when "0011111", -- t[31] = 4353
      "01000100110011" when "0100000", -- t[32] = 4403
      "01000101100101" when "0100001", -- t[33] = 4453
      "01000110011000" when "0100010", -- t[34] = 4504
      "01000111001011" when "0100011", -- t[35] = 4555
      "01000111111111" when "0100100", -- t[36] = 4607
      "01001000110100" when "0100101", -- t[37] = 4660
      "01001001101001" when "0100110", -- t[38] = 4713
      "01001010011111" when "0100111", -- t[39] = 4767
      "01001011010110" when "0101000", -- t[40] = 4822
      "01001100001101" when "0101001", -- t[41] = 4877
      "01001101000101" when "0101010", -- t[42] = 4933
      "01001101111110" when "0101011", -- t[43] = 4990
      "01001110110111" when "0101100", -- t[44] = 5047
      "01001111110001" when "0101101", -- t[45] = 5105
      "01010000101100" when "0101110", -- t[46] = 5164
      "01010001100111" when "0101111", -- t[47] = 5223
      "01010010100011" when "0110000", -- t[48] = 5283
      "01010011100000" when "0110001", -- t[49] = 5344
      "01010100011110" when "0110010", -- t[50] = 5406
      "01010101011100" when "0110011", -- t[51] = 5468
      "01010110011011" when "0110100", -- t[52] = 5531
      "01010111011011" when "0110101", -- t[53] = 5595
      "01011000011100" when "0110110", -- t[54] = 5660
      "01011001011101" when "0110111", -- t[55] = 5725
      "01011010011111" when "0111000", -- t[56] = 5791
      "01011011100011" when "0111001", -- t[57] = 5859
      "01011100100110" when "0111010", -- t[58] = 5926
      "01011101101011" when "0111011", -- t[59] = 5995
      "01011110110001" when "0111100", -- t[60] = 6065
      "01011111110111" when "0111101", -- t[61] = 6135
      "01100000111111" when "0111110", -- t[62] = 6207
      "01100010000111" when "0111111", -- t[63] = 6279
      "01100011010000" when "1000000", -- t[64] = 6352
      "01100100011010" when "1000001", -- t[65] = 6426
      "01100101100101" when "1000010", -- t[66] = 6501
      "01100110110001" when "1000011", -- t[67] = 6577
      "01100111111110" when "1000100", -- t[68] = 6654
      "01101001001100" when "1000101", -- t[69] = 6732
      "01101010011011" when "1000110", -- t[70] = 6811
      "01101011101010" when "1000111", -- t[71] = 6890
      "01101100111011" when "1001000", -- t[72] = 6971
      "01101110001101" when "1001001", -- t[73] = 7053
      "01101111100000" when "1001010", -- t[74] = 7136
      "01110000110100" when "1001011", -- t[75] = 7220
      "01110010001001" when "1001100", -- t[76] = 7305
      "01110011011111" when "1001101", -- t[77] = 7391
      "01110100110110" when "1001110", -- t[78] = 7478
      "01110110001110" when "1001111", -- t[79] = 7566
      "01110111101000" when "1010000", -- t[80] = 7656
      "01111001000010" when "1010001", -- t[81] = 7746
      "01111010011110" when "1010010", -- t[82] = 7838
      "01111011111011" when "1010011", -- t[83] = 7931
      "01111101011001" when "1010100", -- t[84] = 8025
      "01111110111000" when "1010101", -- t[85] = 8120
      "10000000011001" when "1010110", -- t[86] = 8217
      "10000001111010" when "1010111", -- t[87] = 8314
      "10000011011101" when "1011000", -- t[88] = 8413
      "10000101000010" when "1011001", -- t[89] = 8514
      "10000110100111" when "1011010", -- t[90] = 8615
      "10001000001110" when "1011011", -- t[91] = 8718
      "10001001110111" when "1011100", -- t[92] = 8823
      "10001011100001" when "1011101", -- t[93] = 8929
      "10001101001100" when "1011110", -- t[94] = 9036
      "10001110111000" when "1011111", -- t[95] = 9144
      "10010000100110" when "1100000", -- t[96] = 9254
      "10010010010101" when "1100001", -- t[97] = 9365
      "10010100000110" when "1100010", -- t[98] = 9478
      "10010101111001" when "1100011", -- t[99] = 9593
      "10010111101101" when "1100100", -- t[100] = 9709
      "10011001100010" when "1100101", -- t[101] = 9826
      "10011011011001" when "1100110", -- t[102] = 9945
      "10011101010010" when "1100111", -- t[103] = 10066
      "10011111001100" when "1101000", -- t[104] = 10188
      "10100001001000" when "1101001", -- t[105] = 10312
      "10100011000110" when "1101010", -- t[106] = 10438
      "10100101000101" when "1101011", -- t[107] = 10565
      "10100111000110" when "1101100", -- t[108] = 10694
      "10101001001001" when "1101101", -- t[109] = 10825
      "10101011001101" when "1101110", -- t[110] = 10957
      "10101101010100" when "1101111", -- t[111] = 11092
      "10101111011100" when "1110000", -- t[112] = 11228
      "10110001100110" when "1110001", -- t[113] = 11366
      "10110011110010" when "1110010", -- t[114] = 11506
      "10110110000000" when "1110011", -- t[115] = 11648
      "10111000010000" when "1110100", -- t[116] = 11792
      "10111010100010" when "1110101", -- t[117] = 11938
      "10111100110110" when "1110110", -- t[118] = 12086
      "10111111001101" when "1110111", -- t[119] = 12237
      "11000001100101" when "1111000", -- t[120] = 12389
      "11000011111111" when "1111001", -- t[121] = 12543
      "11000110011100" when "1111010", -- t[122] = 12700
      "11001000111011" when "1111011", -- t[123] = 12859
      "11001011011100" when "1111100", -- t[124] = 13020
      "11001110000000" when "1111101", -- t[125] = 13184
      "11010000100101" when "1111110", -- t[126] = 13349
      "11010011001110" when "1111111", -- t[127] = 13518
      "--------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_13_to2 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to2 is
begin
  with x select
    r <=
      "000100" when "0000000", -- t[0] = 4
      "001100" when "0000001", -- t[1] = 12
      "000100" when "0000010", -- t[2] = 4
      "001101" when "0000011", -- t[3] = 13
      "000100" when "0000100", -- t[4] = 4
      "001101" when "0000101", -- t[5] = 13
      "000100" when "0000110", -- t[6] = 4
      "001101" when "0000111", -- t[7] = 13
      "000100" when "0001000", -- t[8] = 4
      "001110" when "0001001", -- t[9] = 14
      "000100" when "0001010", -- t[10] = 4
      "001110" when "0001011", -- t[11] = 14
      "000100" when "0001100", -- t[12] = 4
      "001110" when "0001101", -- t[13] = 14
      "000101" when "0001110", -- t[14] = 5
      "001111" when "0001111", -- t[15] = 15
      "000101" when "0010000", -- t[16] = 5
      "001111" when "0010001", -- t[17] = 15
      "000101" when "0010010", -- t[18] = 5
      "001111" when "0010011", -- t[19] = 15
      "000101" when "0010100", -- t[20] = 5
      "010000" when "0010101", -- t[21] = 16
      "000101" when "0010110", -- t[22] = 5
      "010000" when "0010111", -- t[23] = 16
      "000101" when "0011000", -- t[24] = 5
      "010001" when "0011001", -- t[25] = 17
      "000101" when "0011010", -- t[26] = 5
      "010001" when "0011011", -- t[27] = 17
      "000101" when "0011100", -- t[28] = 5
      "010001" when "0011101", -- t[29] = 17
      "000110" when "0011110", -- t[30] = 6
      "010010" when "0011111", -- t[31] = 18
      "000110" when "0100000", -- t[32] = 6
      "010010" when "0100001", -- t[33] = 18
      "000110" when "0100010", -- t[34] = 6
      "010011" when "0100011", -- t[35] = 19
      "000110" when "0100100", -- t[36] = 6
      "010011" when "0100101", -- t[37] = 19
      "000110" when "0100110", -- t[38] = 6
      "010100" when "0100111", -- t[39] = 20
      "000110" when "0101000", -- t[40] = 6
      "010100" when "0101001", -- t[41] = 20
      "000111" when "0101010", -- t[42] = 7
      "010101" when "0101011", -- t[43] = 21
      "000111" when "0101100", -- t[44] = 7
      "010101" when "0101101", -- t[45] = 21
      "000111" when "0101110", -- t[46] = 7
      "010110" when "0101111", -- t[47] = 22
      "000111" when "0110000", -- t[48] = 7
      "010110" when "0110001", -- t[49] = 22
      "000111" when "0110010", -- t[50] = 7
      "010111" when "0110011", -- t[51] = 23
      "000111" when "0110100", -- t[52] = 7
      "010111" when "0110101", -- t[53] = 23
      "001000" when "0110110", -- t[54] = 8
      "011000" when "0110111", -- t[55] = 24
      "001000" when "0111000", -- t[56] = 8
      "011001" when "0111001", -- t[57] = 25
      "001000" when "0111010", -- t[58] = 8
      "011001" when "0111011", -- t[59] = 25
      "001000" when "0111100", -- t[60] = 8
      "011010" when "0111101", -- t[61] = 26
      "001001" when "0111110", -- t[62] = 9
      "011011" when "0111111", -- t[63] = 27
      "001001" when "1000000", -- t[64] = 9
      "011011" when "1000001", -- t[65] = 27
      "001001" when "1000010", -- t[66] = 9
      "011100" when "1000011", -- t[67] = 28
      "001001" when "1000100", -- t[68] = 9
      "011101" when "1000101", -- t[69] = 29
      "001001" when "1000110", -- t[70] = 9
      "011101" when "1000111", -- t[71] = 29
      "001010" when "1001000", -- t[72] = 10
      "011110" when "1001001", -- t[73] = 30
      "001010" when "1001010", -- t[74] = 10
      "011111" when "1001011", -- t[75] = 31
      "001010" when "1001100", -- t[76] = 10
      "100000" when "1001101", -- t[77] = 32
      "001011" when "1001110", -- t[78] = 11
      "100001" when "1001111", -- t[79] = 33
      "001011" when "1010000", -- t[80] = 11
      "100001" when "1010001", -- t[81] = 33
      "001011" when "1010010", -- t[82] = 11
      "100010" when "1010011", -- t[83] = 34
      "001011" when "1010100", -- t[84] = 11
      "100011" when "1010101", -- t[85] = 35
      "001100" when "1010110", -- t[86] = 12
      "100100" when "1010111", -- t[87] = 36
      "001100" when "1011000", -- t[88] = 12
      "100101" when "1011001", -- t[89] = 37
      "001100" when "1011010", -- t[90] = 12
      "100110" when "1011011", -- t[91] = 38
      "001101" when "1011100", -- t[92] = 13
      "100111" when "1011101", -- t[93] = 39
      "001101" when "1011110", -- t[94] = 13
      "101000" when "1011111", -- t[95] = 40
      "001101" when "1100000", -- t[96] = 13
      "101001" when "1100001", -- t[97] = 41
      "001110" when "1100010", -- t[98] = 14
      "101010" when "1100011", -- t[99] = 42
      "001110" when "1100100", -- t[100] = 14
      "101011" when "1100101", -- t[101] = 43
      "001111" when "1100110", -- t[102] = 15
      "101101" when "1100111", -- t[103] = 45
      "001111" when "1101000", -- t[104] = 15
      "101110" when "1101001", -- t[105] = 46
      "001111" when "1101010", -- t[106] = 15
      "101111" when "1101011", -- t[107] = 47
      "010000" when "1101100", -- t[108] = 16
      "110000" when "1101101", -- t[109] = 48
      "010000" when "1101110", -- t[110] = 16
      "110010" when "1101111", -- t[111] = 50
      "010001" when "1110000", -- t[112] = 17
      "110011" when "1110001", -- t[113] = 51
      "010001" when "1110010", -- t[114] = 17
      "110101" when "1110011", -- t[115] = 53
      "010010" when "1110100", -- t[116] = 18
      "110110" when "1110101", -- t[117] = 54
      "010010" when "1110110", -- t[118] = 18
      "111000" when "1110111", -- t[119] = 56
      "010011" when "1111000", -- t[120] = 19
      "111001" when "1111001", -- t[121] = 57
      "010011" when "1111010", -- t[122] = 19
      "111011" when "1111011", -- t[123] = 59
      "010100" when "1111100", -- t[124] = 20
      "111101" when "1111101", -- t[125] = 61
      "010100" when "1111110", -- t[126] = 20
      "111110" when "1111111", -- t[127] = 62
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_13_to1 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to1 is
begin
  with x select
    r <=
      "00000" when "0000000", -- t[0] = 0
      "00001" when "0000001", -- t[1] = 1
      "00010" when "0000010", -- t[2] = 2
      "00011" when "0000011", -- t[3] = 3
      "00000" when "0000100", -- t[4] = 0
      "00001" when "0000101", -- t[5] = 1
      "00010" when "0000110", -- t[6] = 2
      "00100" when "0000111", -- t[7] = 4
      "00000" when "0001000", -- t[8] = 0
      "00001" when "0001001", -- t[9] = 1
      "00010" when "0001010", -- t[10] = 2
      "00100" when "0001011", -- t[11] = 4
      "00000" when "0001100", -- t[12] = 0
      "00001" when "0001101", -- t[13] = 1
      "00011" when "0001110", -- t[14] = 3
      "00100" when "0001111", -- t[15] = 4
      "00000" when "0010000", -- t[16] = 0
      "00001" when "0010001", -- t[17] = 1
      "00011" when "0010010", -- t[18] = 3
      "00100" when "0010011", -- t[19] = 4
      "00000" when "0010100", -- t[20] = 0
      "00010" when "0010101", -- t[21] = 2
      "00011" when "0010110", -- t[22] = 3
      "00100" when "0010111", -- t[23] = 4
      "00000" when "0011000", -- t[24] = 0
      "00010" when "0011001", -- t[25] = 2
      "00011" when "0011010", -- t[26] = 3
      "00101" when "0011011", -- t[27] = 5
      "00000" when "0011100", -- t[28] = 0
      "00010" when "0011101", -- t[29] = 2
      "00011" when "0011110", -- t[30] = 3
      "00101" when "0011111", -- t[31] = 5
      "00000" when "0100000", -- t[32] = 0
      "00010" when "0100001", -- t[33] = 2
      "00011" when "0100010", -- t[34] = 3
      "00101" when "0100011", -- t[35] = 5
      "00000" when "0100100", -- t[36] = 0
      "00010" when "0100101", -- t[37] = 2
      "00100" when "0100110", -- t[38] = 4
      "00101" when "0100111", -- t[39] = 5
      "00000" when "0101000", -- t[40] = 0
      "00010" when "0101001", -- t[41] = 2
      "00100" when "0101010", -- t[42] = 4
      "00110" when "0101011", -- t[43] = 6
      "00000" when "0101100", -- t[44] = 0
      "00010" when "0101101", -- t[45] = 2
      "00100" when "0101110", -- t[46] = 4
      "00110" when "0101111", -- t[47] = 6
      "00000" when "0110000", -- t[48] = 0
      "00010" when "0110001", -- t[49] = 2
      "00100" when "0110010", -- t[50] = 4
      "00110" when "0110011", -- t[51] = 6
      "00001" when "0110100", -- t[52] = 1
      "00011" when "0110101", -- t[53] = 3
      "00101" when "0110110", -- t[54] = 5
      "00111" when "0110111", -- t[55] = 7
      "00001" when "0111000", -- t[56] = 1
      "00011" when "0111001", -- t[57] = 3
      "00101" when "0111010", -- t[58] = 5
      "00111" when "0111011", -- t[59] = 7
      "00001" when "0111100", -- t[60] = 1
      "00011" when "0111101", -- t[61] = 3
      "00101" when "0111110", -- t[62] = 5
      "00111" when "0111111", -- t[63] = 7
      "00001" when "1000000", -- t[64] = 1
      "00011" when "1000001", -- t[65] = 3
      "00101" when "1000010", -- t[66] = 5
      "01000" when "1000011", -- t[67] = 8
      "00001" when "1000100", -- t[68] = 1
      "00011" when "1000101", -- t[69] = 3
      "00110" when "1000110", -- t[70] = 6
      "01000" when "1000111", -- t[71] = 8
      "00001" when "1001000", -- t[72] = 1
      "00011" when "1001001", -- t[73] = 3
      "00110" when "1001010", -- t[74] = 6
      "01001" when "1001011", -- t[75] = 9
      "00001" when "1001100", -- t[76] = 1
      "00100" when "1001101", -- t[77] = 4
      "00110" when "1001110", -- t[78] = 6
      "01001" when "1001111", -- t[79] = 9
      "00001" when "1010000", -- t[80] = 1
      "00100" when "1010001", -- t[81] = 4
      "00111" when "1010010", -- t[82] = 7
      "01010" when "1010011", -- t[83] = 10
      "00001" when "1010100", -- t[84] = 1
      "00100" when "1010101", -- t[85] = 4
      "00111" when "1010110", -- t[86] = 7
      "01010" when "1010111", -- t[87] = 10
      "00001" when "1011000", -- t[88] = 1
      "00100" when "1011001", -- t[89] = 4
      "00111" when "1011010", -- t[90] = 7
      "01011" when "1011011", -- t[91] = 11
      "00001" when "1011100", -- t[92] = 1
      "00101" when "1011101", -- t[93] = 5
      "01000" when "1011110", -- t[94] = 8
      "01011" when "1011111", -- t[95] = 11
      "00001" when "1100000", -- t[96] = 1
      "00101" when "1100001", -- t[97] = 5
      "01000" when "1100010", -- t[98] = 8
      "01100" when "1100011", -- t[99] = 12
      "00001" when "1100100", -- t[100] = 1
      "00101" when "1100101", -- t[101] = 5
      "01001" when "1100110", -- t[102] = 9
      "01101" when "1100111", -- t[103] = 13
      "00001" when "1101000", -- t[104] = 1
      "00101" when "1101001", -- t[105] = 5
      "01001" when "1101010", -- t[106] = 9
      "01101" when "1101011", -- t[107] = 13
      "00010" when "1101100", -- t[108] = 2
      "00110" when "1101101", -- t[109] = 6
      "01010" when "1101110", -- t[110] = 10
      "01110" when "1101111", -- t[111] = 14
      "00010" when "1110000", -- t[112] = 2
      "00110" when "1110001", -- t[113] = 6
      "01010" when "1110010", -- t[114] = 10
      "01111" when "1110011", -- t[115] = 15
      "00010" when "1110100", -- t[116] = 2
      "00110" when "1110101", -- t[117] = 6
      "01011" when "1110110", -- t[118] = 11
      "10000" when "1110111", -- t[119] = 16
      "00010" when "1111000", -- t[120] = 2
      "00111" when "1111001", -- t[121] = 7
      "01100" when "1111010", -- t[122] = 12
      "10001" when "1111011", -- t[123] = 17
      "00010" when "1111100", -- t[124] = 2
      "00111" when "1111101", -- t[125] = 7
      "01100" when "1111110", -- t[126] = 12
      "10010" when "1111111", -- t[127] = 18
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_13_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to0 is
begin
  with x select
    r <=
      "0" when "000", -- t[0] = 0
      "0" when "001", -- t[1] = 0
      "0" when "010", -- t[2] = 0
      "0" when "011", -- t[3] = 0
      "0" when "100", -- t[4] = 0
      "1" when "101", -- t[5] = 1
      "0" when "110", -- t[6] = 0
      "1" when "111", -- t[7] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_13.all;

entity LNSSub_MPT_T2_13_to2_xor is
  port( a : in  std_logic_vector(5 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(6 downto 0);
  signal out_t : std_logic_vector(5 downto 0);
begin
  sign <= not b(1);
  in_t(6 downto 1) <= a(5 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T2_13_to2
    port map( x => in_t,
              r => out_t );

  r(13 downto 6) <= (13 downto 6 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_13.all;

entity LNSSub_MPT_T2_13_to1_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(6 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(2);
  in_t(6 downto 2) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to1 : LNSSub_MPT_T2_13_to1
    port map( x => in_t,
              r => out_t );

  r(13 downto 5) <= (13 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_13.all;

entity LNSSub_MPT_T2_13_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T2_13_to0
    port map( x => in_t,
              r => out_t );

  r(13 downto 1) <= (13 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_13.all;

entity LNSSub_MPT_T2_13 is
  port( x : in  std_logic_vector(13 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_13 is
  signal in_tiv  : std_logic_vector(6 downto 0);
  signal out_tiv : std_logic_vector(13 downto 0);
  signal a2      : std_logic_vector(5 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(13 downto 0);
  signal a1      : std_logic_vector(4 downto 0);
  signal b1      : std_logic_vector(2 downto 0);
  signal out1    : std_logic_vector(13 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(13 downto 0);
  signal sum     : std_logic_vector(13 downto 0);
begin
  in_tiv <= x(13 downto 7);
  inst_tiv : LNSSub_MPT_T2_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(13 downto 8);
  b2 <= x(6 downto 5);
  inst_to2_xor : LNSSub_MPT_T2_13_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(13 downto 9);
  b1 <= x(4 downto 2);
  inst_to1_xor : LNSSub_MPT_T2_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(13 downto 12);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T2_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(13 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T2_13_Clk is
  port( x   : in  std_logic_vector(13 downto 0);
        r   : out std_logic_vector(11 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T2_13_Clk is
  signal in_tiv_1  : std_logic_vector(6 downto 0);
  signal out_tiv_1 : std_logic_vector(13 downto 0);
  signal out_tiv_2 : std_logic_vector(13 downto 0);
  signal a2_1      : std_logic_vector(5 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(13 downto 0);
  signal out2_2    : std_logic_vector(13 downto 0);
  signal a1_1      : std_logic_vector(4 downto 0);
  signal b1_1      : std_logic_vector(2 downto 0);
  signal out1_1    : std_logic_vector(13 downto 0);
  signal out1_2    : std_logic_vector(13 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(13 downto 0);
  signal out0_2    : std_logic_vector(13 downto 0);
  signal psum1_2     : std_logic_vector(13 downto 0);
  signal psum1_3     : std_logic_vector(13 downto 0);
  signal psum2_2     : std_logic_vector(13 downto 0);
  signal psum2_3     : std_logic_vector(13 downto 0);
  signal sum_3     : std_logic_vector(13 downto 0);
begin
  in_tiv_1 <= x(13 downto 7);
  inst_tiv : LNSSub_MPT_T2_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(13 downto 8);
  b2_1 <= x(6 downto 5);
  inst_to2_xor : LNSSub_MPT_T2_13_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(13 downto 9);
  b1_1 <= x(4 downto 2);
  inst_to1_xor : LNSSub_MPT_T2_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(13 downto 12);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T2_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(13 downto 2);
end architecture;


-- MultiPartite: LNS subtraction function: [-2.0 -1.0[ -> [0.0 1.0[
-- wI = 13 bits
-- wO = 12 bits
-- Decomposition: 7, 6 / 5, 4, 2 / 2, 2, 2
-- Guard bits: 4
-- Size: 2784 = 16.2^7 + 8.2^6 + 6.2^5 + 4.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T3_13 is
  component LNSSub_MPT_T3_13_tiv is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to2 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to2_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T3_13_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_13_tiv is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_tiv is
begin
  with x select
    r <=
      "0110101010011101" when "0000000", -- t[0] = 27293
      "0110101101001001" when "0000001", -- t[1] = 27465
      "0110101111110110" when "0000010", -- t[2] = 27638
      "0110110010100101" when "0000011", -- t[3] = 27813
      "0110110101010100" when "0000100", -- t[4] = 27988
      "0110111000000101" when "0000101", -- t[5] = 28165
      "0110111010111000" when "0000110", -- t[6] = 28344
      "0110111101101011" when "0000111", -- t[7] = 28523
      "0111000000100000" when "0001000", -- t[8] = 28704
      "0111000011010110" when "0001001", -- t[9] = 28886
      "0111000110001110" when "0001010", -- t[10] = 29070
      "0111001001000111" when "0001011", -- t[11] = 29255
      "0111001100000001" when "0001100", -- t[12] = 29441
      "0111001110111101" when "0001101", -- t[13] = 29629
      "0111010001111010" when "0001110", -- t[14] = 29818
      "0111010100111000" when "0001111", -- t[15] = 30008
      "0111010111111000" when "0010000", -- t[16] = 30200
      "0111011010111001" when "0010001", -- t[17] = 30393
      "0111011101111100" when "0010010", -- t[18] = 30588
      "0111100001000000" when "0010011", -- t[19] = 30784
      "0111100100000110" when "0010100", -- t[20] = 30982
      "0111100111001101" when "0010101", -- t[21] = 31181
      "0111101010010110" when "0010110", -- t[22] = 31382
      "0111101101100000" when "0010111", -- t[23] = 31584
      "0111110000101100" when "0011000", -- t[24] = 31788
      "0111110011111001" when "0011001", -- t[25] = 31993
      "0111110111001000" when "0011010", -- t[26] = 32200
      "0111111010011001" when "0011011", -- t[27] = 32409
      "0111111101101011" when "0011100", -- t[28] = 32619
      "1000000000111110" when "0011101", -- t[29] = 32830
      "1000000100010100" when "0011110", -- t[30] = 33044
      "1000000111101011" when "0011111", -- t[31] = 33259
      "1000001011000011" when "0100000", -- t[32] = 33475
      "1000001110011110" when "0100001", -- t[33] = 33694
      "1000010001111010" when "0100010", -- t[34] = 33914
      "1000010101010111" when "0100011", -- t[35] = 34135
      "1000011000110111" when "0100100", -- t[36] = 34359
      "1000011100011000" when "0100101", -- t[37] = 34584
      "1000011111111011" when "0100110", -- t[38] = 34811
      "1000100011100000" when "0100111", -- t[39] = 35040
      "1000100111000110" when "0101000", -- t[40] = 35270
      "1000101010101110" when "0101001", -- t[41] = 35502
      "1000101110011001" when "0101010", -- t[42] = 35737
      "1000110010000101" when "0101011", -- t[43] = 35973
      "1000110101110011" when "0101100", -- t[44] = 36211
      "1000111001100010" when "0101101", -- t[45] = 36450
      "1000111101010100" when "0101110", -- t[46] = 36692
      "1001000001001000" when "0101111", -- t[47] = 36936
      "1001000100111101" when "0110000", -- t[48] = 37181
      "1001001000110101" when "0110001", -- t[49] = 37429
      "1001001100101111" when "0110010", -- t[50] = 37679
      "1001010000101010" when "0110011", -- t[51] = 37930
      "1001010100101000" when "0110100", -- t[52] = 38184
      "1001011000101000" when "0110101", -- t[53] = 38440
      "1001011100101001" when "0110110", -- t[54] = 38697
      "1001100000101101" when "0110111", -- t[55] = 38957
      "1001100100110011" when "0111000", -- t[56] = 39219
      "1001101000111100" when "0111001", -- t[57] = 39484
      "1001101101000110" when "0111010", -- t[58] = 39750
      "1001110001010011" when "0111011", -- t[59] = 40019
      "1001110101100001" when "0111100", -- t[60] = 40289
      "1001111001110010" when "0111101", -- t[61] = 40562
      "1001111110000110" when "0111110", -- t[62] = 40838
      "1010000010011100" when "0111111", -- t[63] = 41116
      "1010000110110100" when "1000000", -- t[64] = 41396
      "1010001011001110" when "1000001", -- t[65] = 41678
      "1010001111101011" when "1000010", -- t[66] = 41963
      "1010010100001010" when "1000011", -- t[67] = 42250
      "1010011000101011" when "1000100", -- t[68] = 42539
      "1010011101010000" when "1000101", -- t[69] = 42832
      "1010100001110110" when "1000110", -- t[70] = 43126
      "1010100110011111" when "1000111", -- t[71] = 43423
      "1010101011001011" when "1001000", -- t[72] = 43723
      "1010101111111001" when "1001001", -- t[73] = 44025
      "1010110100101010" when "1001010", -- t[74] = 44330
      "1010111001011101" when "1001011", -- t[75] = 44637
      "1010111110010100" when "1001100", -- t[76] = 44948
      "1011000011001101" when "1001101", -- t[77] = 45261
      "1011001000001000" when "1001110", -- t[78] = 45576
      "1011001101000111" when "1001111", -- t[79] = 45895
      "1011010010001000" when "1010000", -- t[80] = 46216
      "1011010111001100" when "1010001", -- t[81] = 46540
      "1011011100010011" when "1010010", -- t[82] = 46867
      "1011100001011101" when "1010011", -- t[83] = 47197
      "1011100110101010" when "1010100", -- t[84] = 47530
      "1011101011111010" when "1010101", -- t[85] = 47866
      "1011110001001101" when "1010110", -- t[86] = 48205
      "1011110110100010" when "1010111", -- t[87] = 48546
      "1011111011111100" when "1011000", -- t[88] = 48892
      "1100000001011000" when "1011001", -- t[89] = 49240
      "1100000110110111" when "1011010", -- t[90] = 49591
      "1100001100011010" when "1011011", -- t[91] = 49946
      "1100010010000000" when "1011100", -- t[92] = 50304
      "1100010111101001" when "1011101", -- t[93] = 50665
      "1100011101010101" when "1011110", -- t[94] = 51029
      "1100100011000101" when "1011111", -- t[95] = 51397
      "1100101000111001" when "1100000", -- t[96] = 51769
      "1100101110110000" when "1100001", -- t[97] = 52144
      "1100110100101010" when "1100010", -- t[98] = 52522
      "1100111010101000" when "1100011", -- t[99] = 52904
      "1101000000101010" when "1100100", -- t[100] = 53290
      "1101000110101111" when "1100101", -- t[101] = 53679
      "1101001100111000" when "1100110", -- t[102] = 54072
      "1101010011000101" when "1100111", -- t[103] = 54469
      "1101011001010110" when "1101000", -- t[104] = 54870
      "1101011111101011" when "1101001", -- t[105] = 55275
      "1101100110000011" when "1101010", -- t[106] = 55683
      "1101101100100000" when "1101011", -- t[107] = 56096
      "1101110011000001" when "1101100", -- t[108] = 56513
      "1101111001100101" when "1101101", -- t[109] = 56933
      "1110000000001110" when "1101110", -- t[110] = 57358
      "1110000110111011" when "1101111", -- t[111] = 57787
      "1110001101101101" when "1110000", -- t[112] = 58221
      "1110010100100011" when "1110001", -- t[113] = 58659
      "1110011011011101" when "1110010", -- t[114] = 59101
      "1110100010011100" when "1110011", -- t[115] = 59548
      "1110101001011111" when "1110100", -- t[116] = 59999
      "1110110000100111" when "1110101", -- t[117] = 60455
      "1110110111110100" when "1110110", -- t[118] = 60916
      "1110111111000101" when "1110111", -- t[119] = 61381
      "1111000110011100" when "1111000", -- t[120] = 61852
      "1111001101110111" when "1111001", -- t[121] = 62327
      "1111010101010111" when "1111010", -- t[122] = 62807
      "1111011100111101" when "1111011", -- t[123] = 63293
      "1111100100100111" when "1111100", -- t[124] = 63783
      "1111101100010111" when "1111101", -- t[125] = 64279
      "1111110100001100" when "1111110", -- t[126] = 64780
      "1111111100000110" when "1111111", -- t[127] = 65286
      "----------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_13_to2 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to2 is
begin
  with x select
    r <=
      "00010101" when "000000", -- t[0] = 21
      "01000000" when "000001", -- t[1] = 64
      "00010110" when "000010", -- t[2] = 22
      "01000010" when "000011", -- t[3] = 66
      "00010110" when "000100", -- t[4] = 22
      "01000100" when "000101", -- t[5] = 68
      "00010111" when "000110", -- t[6] = 23
      "01000110" when "000111", -- t[7] = 70
      "00011000" when "001000", -- t[8] = 24
      "01001000" when "001001", -- t[9] = 72
      "00011001" when "001010", -- t[10] = 25
      "01001011" when "001011", -- t[11] = 75
      "00011001" when "001100", -- t[12] = 25
      "01001101" when "001101", -- t[13] = 77
      "00011010" when "001110", -- t[14] = 26
      "01001111" when "001111", -- t[15] = 79
      "00011011" when "010000", -- t[16] = 27
      "01010010" when "010001", -- t[17] = 82
      "00011100" when "010010", -- t[18] = 28
      "01010101" when "010011", -- t[19] = 85
      "00011101" when "010100", -- t[20] = 29
      "01010111" when "010101", -- t[21] = 87
      "00011110" when "010110", -- t[22] = 30
      "01011010" when "010111", -- t[23] = 90
      "00011111" when "011000", -- t[24] = 31
      "01011101" when "011001", -- t[25] = 93
      "00100000" when "011010", -- t[26] = 32
      "01100000" when "011011", -- t[27] = 96
      "00100001" when "011100", -- t[28] = 33
      "01100011" when "011101", -- t[29] = 99
      "00100010" when "011110", -- t[30] = 34
      "01100111" when "011111", -- t[31] = 103
      "00100011" when "100000", -- t[32] = 35
      "01101010" when "100001", -- t[33] = 106
      "00100100" when "100010", -- t[34] = 36
      "01101110" when "100011", -- t[35] = 110
      "00100110" when "100100", -- t[36] = 38
      "01110010" when "100101", -- t[37] = 114
      "00100111" when "100110", -- t[38] = 39
      "01110110" when "100111", -- t[39] = 118
      "00101000" when "101000", -- t[40] = 40
      "01111010" when "101001", -- t[41] = 122
      "00101010" when "101010", -- t[42] = 42
      "01111110" when "101011", -- t[43] = 126
      "00101011" when "101100", -- t[44] = 43
      "10000011" when "101101", -- t[45] = 131
      "00101101" when "101110", -- t[46] = 45
      "10001000" when "101111", -- t[47] = 136
      "00101111" when "110000", -- t[48] = 47
      "10001101" when "110001", -- t[49] = 141
      "00110001" when "110010", -- t[50] = 49
      "10010011" when "110011", -- t[51] = 147
      "00110011" when "110100", -- t[52] = 51
      "10011001" when "110101", -- t[53] = 153
      "00110101" when "110110", -- t[54] = 53
      "10011111" when "110111", -- t[55] = 159
      "00110111" when "111000", -- t[56] = 55
      "10100101" when "111001", -- t[57] = 165
      "00111001" when "111010", -- t[58] = 57
      "10101100" when "111011", -- t[59] = 172
      "00111011" when "111100", -- t[60] = 59
      "10110011" when "111101", -- t[61] = 179
      "00111110" when "111110", -- t[62] = 62
      "10111011" when "111111", -- t[63] = 187
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_13_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to1 is
begin
  with x select
    r <=
      "000101" when "00000", -- t[0] = 5
      "010000" when "00001", -- t[1] = 16
      "000101" when "00010", -- t[2] = 5
      "010001" when "00011", -- t[3] = 17
      "000110" when "00100", -- t[4] = 6
      "010010" when "00101", -- t[5] = 18
      "000110" when "00110", -- t[6] = 6
      "010011" when "00111", -- t[7] = 19
      "000110" when "01000", -- t[8] = 6
      "010100" when "01001", -- t[9] = 20
      "000111" when "01010", -- t[10] = 7
      "010110" when "01011", -- t[11] = 22
      "000111" when "01100", -- t[12] = 7
      "010111" when "01101", -- t[13] = 23
      "001000" when "01110", -- t[14] = 8
      "011001" when "01111", -- t[15] = 25
      "001001" when "10000", -- t[16] = 9
      "011011" when "10001", -- t[17] = 27
      "001001" when "10010", -- t[18] = 9
      "011101" when "10011", -- t[19] = 29
      "001010" when "10100", -- t[20] = 10
      "011111" when "10101", -- t[21] = 31
      "001011" when "10110", -- t[22] = 11
      "100001" when "10111", -- t[23] = 33
      "001100" when "11000", -- t[24] = 12
      "100100" when "11001", -- t[25] = 36
      "001101" when "11010", -- t[26] = 13
      "100111" when "11011", -- t[27] = 39
      "001110" when "11100", -- t[28] = 14
      "101010" when "11101", -- t[29] = 42
      "001111" when "11110", -- t[30] = 15
      "101101" when "11111", -- t[31] = 45
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_13_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to0 is
begin
  with x select
    r <=
      "0001" when "000", -- t[0] = 1
      "0100" when "001", -- t[1] = 4
      "0001" when "010", -- t[2] = 1
      "0101" when "011", -- t[3] = 5
      "0010" when "100", -- t[4] = 2
      "0111" when "101", -- t[5] = 7
      "0011" when "110", -- t[6] = 3
      "1010" when "111", -- t[7] = 10
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_13.all;

entity LNSSub_MPT_T3_13_to2_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(7 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T3_13_to2
    port map( x => in_t,
              r => out_t );

  r(15 downto 8) <= (15 downto 8 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_13.all;

entity LNSSub_MPT_T3_13_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(5 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T3_13_to1
    port map( x => in_t,
              r => out_t );

  r(15 downto 6) <= (15 downto 6 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_13.all;

entity LNSSub_MPT_T3_13_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T3_13_to0
    port map( x => in_t,
              r => out_t );

  r(15 downto 4) <= (15 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_13.all;

entity LNSSub_MPT_T3_13 is
  port( x : in  std_logic_vector(12 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_13 is
  signal in_tiv  : std_logic_vector(6 downto 0);
  signal out_tiv : std_logic_vector(15 downto 0);
  signal a2      : std_logic_vector(4 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(15 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(15 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(15 downto 0);
  signal sum     : std_logic_vector(15 downto 0);
begin
  in_tiv <= x(12 downto 6);
  inst_tiv : LNSSub_MPT_T3_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(12 downto 8);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T3_13_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(12 downto 9);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T3_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(12 downto 11);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T3_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(15 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T3_13_Clk is
  port( x   : in  std_logic_vector(12 downto 0);
        r   : out std_logic_vector(11 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T3_13_Clk is
  signal in_tiv_1  : std_logic_vector(6 downto 0);
  signal out_tiv_1 : std_logic_vector(15 downto 0);
  signal out_tiv_2 : std_logic_vector(15 downto 0);
  signal a2_1      : std_logic_vector(4 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(15 downto 0);
  signal out2_2    : std_logic_vector(15 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(15 downto 0);
  signal out1_2    : std_logic_vector(15 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(15 downto 0);
  signal out0_2    : std_logic_vector(15 downto 0);
  signal psum1_2     : std_logic_vector(15 downto 0);
  signal psum1_3     : std_logic_vector(15 downto 0);
  signal psum2_2     : std_logic_vector(15 downto 0);
  signal psum2_3     : std_logic_vector(15 downto 0);
  signal sum_3     : std_logic_vector(15 downto 0);
begin
  in_tiv_1 <= x(12 downto 6);
  inst_tiv : LNSSub_MPT_T3_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(12 downto 8);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T3_13_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(12 downto 9);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T3_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(12 downto 11);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T3_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(15 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-1.0 -0.5[ -> [0.0 2.0[
-- wI = 12 bits
-- wO = 12 bits
-- Decomposition: 6, 6 / 5, 4, 3 / 2, 2, 2
-- Guard bits: 5
-- Size: 1968 = 17.2^6 + 9.2^6 + 7.2^5 + 5.2^4

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T4_13 is
  component LNSSub_MPT_T4_13_tiv is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to2 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to0 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to2_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T4_13_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_13_tiv is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_tiv is
begin
  with x select
    r <=
      "10000000100001110" when "000000", -- t[0] = 65806
      "10000001100010100" when "000001", -- t[1] = 66324
      "10000010100011111" when "000010", -- t[2] = 66847
      "10000011100110000" when "000011", -- t[3] = 67376
      "10000100101000111" when "000100", -- t[4] = 67911
      "10000101101100100" when "000101", -- t[5] = 68452
      "10000110110000111" when "000110", -- t[6] = 68999
      "10000111110110000" when "000111", -- t[7] = 69552
      "10001000111011111" when "001000", -- t[8] = 70111
      "10001010000010101" when "001001", -- t[9] = 70677
      "10001011001010010" when "001010", -- t[10] = 71250
      "10001100010010100" when "001011", -- t[11] = 71828
      "10001101011011110" when "001100", -- t[12] = 72414
      "10001110100101111" when "001101", -- t[13] = 73007
      "10001111110000110" when "001110", -- t[14] = 73606
      "10010000111100101" when "001111", -- t[15] = 74213
      "10010010001001011" when "010000", -- t[16] = 74827
      "10010011010111000" when "010001", -- t[17] = 75448
      "10010100100101101" when "010010", -- t[18] = 76077
      "10010101110101001" when "010011", -- t[19] = 76713
      "10010111000101101" when "010100", -- t[20] = 77357
      "10011000010111001" when "010101", -- t[21] = 78009
      "10011001101001110" when "010110", -- t[22] = 78670
      "10011010111101010" when "010111", -- t[23] = 79338
      "10011100010001111" when "011000", -- t[24] = 80015
      "10011101100111101" when "011001", -- t[25] = 80701
      "10011110111110011" when "011010", -- t[26] = 81395
      "10100000010110011" when "011011", -- t[27] = 82099
      "10100001101111011" when "011100", -- t[28] = 82811
      "10100011001001101" when "011101", -- t[29] = 83533
      "10100100100101000" when "011110", -- t[30] = 84264
      "10100110000001101" when "011111", -- t[31] = 85005
      "10100111011111100" when "100000", -- t[32] = 85756
      "10101000111110101" when "100001", -- t[33] = 86517
      "10101010011111000" when "100010", -- t[34] = 87288
      "10101100000000110" when "100011", -- t[35] = 88070
      "10101101100011111" when "100100", -- t[36] = 88863
      "10101111001000011" when "100101", -- t[37] = 89667
      "10110000101110010" when "100110", -- t[38] = 90482
      "10110010010101101" when "100111", -- t[39] = 91309
      "10110011111110100" when "101000", -- t[40] = 92148
      "10110101101000110" when "101001", -- t[41] = 92998
      "10110111010100110" when "101010", -- t[42] = 93862
      "10111001000010001" when "101011", -- t[43] = 94737
      "10111010110001010" when "101100", -- t[44] = 95626
      "10111100100010001" when "101101", -- t[45] = 96529
      "10111110010100100" when "101110", -- t[46] = 97444
      "11000000001000110" when "101111", -- t[47] = 98374
      "11000001111110110" when "110000", -- t[48] = 99318
      "11000011110110101" when "110001", -- t[49] = 100277
      "11000101110000011" when "110010", -- t[50] = 101251
      "11000111101100001" when "110011", -- t[51] = 102241
      "11001001101001111" when "110100", -- t[52] = 103247
      "11001011101001100" when "110101", -- t[53] = 104268
      "11001101101011011" when "110110", -- t[54] = 105307
      "11001111101111011" when "110111", -- t[55] = 106363
      "11010001110101101" when "111000", -- t[56] = 107437
      "11010011111110001" when "111001", -- t[57] = 108529
      "11010110001001000" when "111010", -- t[58] = 109640
      "11011000010110010" when "111011", -- t[59] = 110770
      "11011010100110000" when "111100", -- t[60] = 111920
      "11011100111000010" when "111101", -- t[61] = 113090
      "11011111001101010" when "111110", -- t[62] = 114282
      "11100001100100111" when "111111", -- t[63] = 115495
      "-----------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_13_to2 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to2 is
begin
  with x select
    r <=
      "001000000" when "000000", -- t[0] = 64
      "011000001" when "000001", -- t[1] = 193
      "001000010" when "000010", -- t[2] = 66
      "011000110" when "000011", -- t[3] = 198
      "001000011" when "000100", -- t[4] = 67
      "011001010" when "000101", -- t[5] = 202
      "001000101" when "000110", -- t[6] = 69
      "011001111" when "000111", -- t[7] = 207
      "001000110" when "001000", -- t[8] = 70
      "011010011" when "001001", -- t[9] = 211
      "001001000" when "001010", -- t[10] = 72
      "011011000" when "001011", -- t[11] = 216
      "001001001" when "001100", -- t[12] = 73
      "011011101" when "001101", -- t[13] = 221
      "001001011" when "001110", -- t[14] = 75
      "011100011" when "001111", -- t[15] = 227
      "001001101" when "010000", -- t[16] = 77
      "011101000" when "010001", -- t[17] = 232
      "001001111" when "010010", -- t[18] = 79
      "011101110" when "010011", -- t[19] = 238
      "001010001" when "010100", -- t[20] = 81
      "011110100" when "010101", -- t[21] = 244
      "001010011" when "010110", -- t[22] = 83
      "011111010" when "010111", -- t[23] = 250
      "001010101" when "011000", -- t[24] = 85
      "100000000" when "011001", -- t[25] = 256
      "001010111" when "011010", -- t[26] = 87
      "100000111" when "011011", -- t[27] = 263
      "001011010" when "011100", -- t[28] = 90
      "100001110" when "011101", -- t[29] = 270
      "001011100" when "011110", -- t[30] = 92
      "100010101" when "011111", -- t[31] = 277
      "001011110" when "100000", -- t[32] = 94
      "100011100" when "100001", -- t[33] = 284
      "001100001" when "100010", -- t[34] = 97
      "100100100" when "100011", -- t[35] = 292
      "001100100" when "100100", -- t[36] = 100
      "100101100" when "100101", -- t[37] = 300
      "001100111" when "100110", -- t[38] = 103
      "100110101" when "100111", -- t[39] = 309
      "001101010" when "101000", -- t[40] = 106
      "100111110" when "101001", -- t[41] = 318
      "001101101" when "101010", -- t[42] = 109
      "101000111" when "101011", -- t[43] = 327
      "001110000" when "101100", -- t[44] = 112
      "101010001" when "101101", -- t[45] = 337
      "001110100" when "101110", -- t[46] = 116
      "101011100" when "101111", -- t[47] = 348
      "001110111" when "110000", -- t[48] = 119
      "101100110" when "110001", -- t[49] = 358
      "001111011" when "110010", -- t[50] = 123
      "101110010" when "110011", -- t[51] = 370
      "001111111" when "110100", -- t[52] = 127
      "101111110" when "110101", -- t[53] = 382
      "010000011" when "110110", -- t[54] = 131
      "110001011" when "110111", -- t[55] = 395
      "010001000" when "111000", -- t[56] = 136
      "110011000" when "111001", -- t[57] = 408
      "010001100" when "111010", -- t[58] = 140
      "110100110" when "111011", -- t[59] = 422
      "010010010" when "111100", -- t[60] = 146
      "110110110" when "111101", -- t[61] = 438
      "010010111" when "111110", -- t[62] = 151
      "111000110" when "111111", -- t[63] = 454
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_13_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to1 is
begin
  with x select
    r <=
      "0010000" when "00000", -- t[0] = 16
      "0110001" when "00001", -- t[1] = 49
      "0010001" when "00010", -- t[2] = 17
      "0110011" when "00011", -- t[3] = 51
      "0010001" when "00100", -- t[4] = 17
      "0110101" when "00101", -- t[5] = 53
      "0010010" when "00110", -- t[6] = 18
      "0111000" when "00111", -- t[7] = 56
      "0010011" when "01000", -- t[8] = 19
      "0111010" when "01001", -- t[9] = 58
      "0010100" when "01010", -- t[10] = 20
      "0111101" when "01011", -- t[11] = 61
      "0010101" when "01100", -- t[12] = 21
      "1000001" when "01101", -- t[13] = 65
      "0010110" when "01110", -- t[14] = 22
      "1000100" when "01111", -- t[15] = 68
      "0011000" when "10000", -- t[16] = 24
      "1001000" when "10001", -- t[17] = 72
      "0011001" when "10010", -- t[18] = 25
      "1001100" when "10011", -- t[19] = 76
      "0011010" when "10100", -- t[20] = 26
      "1010000" when "10101", -- t[21] = 80
      "0011100" when "10110", -- t[22] = 28
      "1010101" when "10111", -- t[23] = 85
      "0011110" when "11000", -- t[24] = 30
      "1011011" when "11001", -- t[25] = 91
      "0100000" when "11010", -- t[26] = 32
      "1100001" when "11011", -- t[27] = 97
      "0100010" when "11100", -- t[28] = 34
      "1101000" when "11101", -- t[29] = 104
      "0100101" when "11110", -- t[30] = 37
      "1101111" when "11111", -- t[31] = 111
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_13_to0 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to0 is
begin
  with x select
    r <=
      "00100" when "0000", -- t[0] = 4
      "01100" when "0001", -- t[1] = 12
      "00100" when "0010", -- t[2] = 4
      "01101" when "0011", -- t[3] = 13
      "00101" when "0100", -- t[4] = 5
      "01111" when "0101", -- t[5] = 15
      "00101" when "0110", -- t[6] = 5
      "10000" when "0111", -- t[7] = 16
      "00110" when "1000", -- t[8] = 6
      "10010" when "1001", -- t[9] = 18
      "00110" when "1010", -- t[10] = 6
      "10100" when "1011", -- t[11] = 20
      "00111" when "1100", -- t[12] = 7
      "10111" when "1101", -- t[13] = 23
      "01000" when "1110", -- t[14] = 8
      "11010" when "1111", -- t[15] = 26
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_13.all;

entity LNSSub_MPT_T4_13_to2_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(8 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T4_13_to2
    port map( x => in_t,
              r => out_t );

  r(16 downto 9) <= (16 downto 9 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
  r(8) <= out_t(8) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_13.all;

entity LNSSub_MPT_T4_13_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(6 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T4_13_to1
    port map( x => in_t,
              r => out_t );

  r(16 downto 7) <= (16 downto 7 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_13.all;

entity LNSSub_MPT_T4_13_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T4_13_to0
    port map( x => in_t,
              r => out_t );

  r(16 downto 5) <= (16 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_13.all;

entity LNSSub_MPT_T4_13 is
  port( x : in  std_logic_vector(11 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_13 is
  signal in_tiv  : std_logic_vector(5 downto 0);
  signal out_tiv : std_logic_vector(16 downto 0);
  signal a2      : std_logic_vector(4 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(16 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(16 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(16 downto 0);
  signal sum     : std_logic_vector(16 downto 0);
begin
  in_tiv <= x(11 downto 6);
  inst_tiv : LNSSub_MPT_T4_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(11 downto 7);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T4_13_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(11 downto 8);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T4_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(11 downto 9);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T4_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(16 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T4_13_Clk is
  port( x   : in  std_logic_vector(11 downto 0);
        r   : out std_logic_vector(11 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T4_13_Clk is
  signal in_tiv_1  : std_logic_vector(5 downto 0);
  signal out_tiv_1 : std_logic_vector(16 downto 0);
  signal out_tiv_2 : std_logic_vector(16 downto 0);
  signal a2_1      : std_logic_vector(4 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(16 downto 0);
  signal out2_2    : std_logic_vector(16 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(16 downto 0);
  signal out1_2    : std_logic_vector(16 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(16 downto 0);
  signal out0_2    : std_logic_vector(16 downto 0);
  signal psum1_2     : std_logic_vector(16 downto 0);
  signal psum1_3     : std_logic_vector(16 downto 0);
  signal psum2_2     : std_logic_vector(16 downto 0);
  signal psum2_3     : std_logic_vector(16 downto 0);
  signal sum_3     : std_logic_vector(16 downto 0);
begin
  in_tiv_1 <= x(11 downto 6);
  inst_tiv : LNSSub_MPT_T4_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(11 downto 7);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T4_13_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(11 downto 8);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T4_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(11 downto 9);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T4_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(16 downto 5);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.5 -0.25[ -> [0.0 4.0[
-- wI = 11 bits
-- wO = 12 bits
-- Decomposition: 6, 5 / 5, 4 / 2, 3
-- Guard bits: 5
-- Size: 2048 = 17.2^6 + 8.2^6 + 7.2^6

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T5_13 is
  component LNSSub_MPT_T5_13_tiv is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T5_13_to1 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T5_13_to0 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T5_13_to1_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T5_13_to0_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_13_tiv is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13_tiv is
begin
  with x select
    r <=
      "01110001101101001" when "000000", -- t[0] = 58217
      "01110010010100001" when "000001", -- t[1] = 58529
      "01110010111011100" when "000010", -- t[2] = 58844
      "01110011100011010" when "000011", -- t[3] = 59162
      "01110100001011010" when "000100", -- t[4] = 59482
      "01110100110011110" when "000101", -- t[5] = 59806
      "01110101011100101" when "000110", -- t[6] = 60133
      "01110110000101111" when "000111", -- t[7] = 60463
      "01110110101111101" when "001000", -- t[8] = 60797
      "01110111011001101" when "001001", -- t[9] = 61133
      "01111000000100001" when "001010", -- t[10] = 61473
      "01111000101111001" when "001011", -- t[11] = 61817
      "01111001011010011" when "001100", -- t[12] = 62163
      "01111010000110010" when "001101", -- t[13] = 62514
      "01111010110010100" when "001110", -- t[14] = 62868
      "01111011011111001" when "001111", -- t[15] = 63225
      "01111100001100011" when "010000", -- t[16] = 63587
      "01111100111010000" when "010001", -- t[17] = 63952
      "01111101101000001" when "010010", -- t[18] = 64321
      "01111110010110101" when "010011", -- t[19] = 64693
      "01111111000101110" when "010100", -- t[20] = 65070
      "01111111110101011" when "010101", -- t[21] = 65451
      "10000000100101100" when "010110", -- t[22] = 65836
      "10000001010110001" when "010111", -- t[23] = 66225
      "10000010000111011" when "011000", -- t[24] = 66619
      "10000010111001001" when "011001", -- t[25] = 67017
      "10000011101011011" when "011010", -- t[26] = 67419
      "10000100011110010" when "011011", -- t[27] = 67826
      "10000101010001101" when "011100", -- t[28] = 68237
      "10000110000101110" when "011101", -- t[29] = 68654
      "10000110111010011" when "011110", -- t[30] = 69075
      "10000111101111101" when "011111", -- t[31] = 69501
      "10001000100101100" when "100000", -- t[32] = 69932
      "10001001011100000" when "100001", -- t[33] = 70368
      "10001010010011010" when "100010", -- t[34] = 70810
      "10001011001011001" when "100011", -- t[35] = 71257
      "10001100000011101" when "100100", -- t[36] = 71709
      "10001100111100111" when "100101", -- t[37] = 72167
      "10001101110110111" when "100110", -- t[38] = 72631
      "10001110110001101" when "100111", -- t[39] = 73101
      "10001111101101001" when "101000", -- t[40] = 73577
      "10010000101001010" when "101001", -- t[41] = 74058
      "10010001100110010" when "101010", -- t[42] = 74546
      "10010010100100001" when "101011", -- t[43] = 75041
      "10010011100010110" when "101100", -- t[44] = 75542
      "10010100100010010" when "101101", -- t[45] = 76050
      "10010101100010101" when "101110", -- t[46] = 76565
      "10010110100011111" when "101111", -- t[47] = 77087
      "10010111100110000" when "110000", -- t[48] = 77616
      "10011000101001000" when "110001", -- t[49] = 78152
      "10011001101101001" when "110010", -- t[50] = 78697
      "10011010110010001" when "110011", -- t[51] = 79249
      "10011011111000001" when "110100", -- t[52] = 79809
      "10011100111111001" when "110101", -- t[53] = 80377
      "10011110000111010" when "110110", -- t[54] = 80954
      "10011111010000100" when "110111", -- t[55] = 81540
      "10100000011010110" when "111000", -- t[56] = 82134
      "10100001100110010" when "111001", -- t[57] = 82738
      "10100010110010111" when "111010", -- t[58] = 83351
      "10100100000000110" when "111011", -- t[59] = 83974
      "10100101001111111" when "111100", -- t[60] = 84607
      "10100110100000011" when "111101", -- t[61] = 85251
      "10100111110010001" when "111110", -- t[62] = 85905
      "10101001000101010" when "111111", -- t[63] = 86570
      "-----------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_13_to1 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13_to1 is
begin
  with x select
    r <=
      "00100110" when "000000", -- t[0] = 38
      "01110100" when "000001", -- t[1] = 116
      "00100111" when "000010", -- t[2] = 39
      "01110111" when "000011", -- t[3] = 119
      "00101000" when "000100", -- t[4] = 40
      "01111001" when "000101", -- t[5] = 121
      "00101001" when "000110", -- t[6] = 41
      "01111011" when "000111", -- t[7] = 123
      "00101010" when "001000", -- t[8] = 42
      "01111110" when "001001", -- t[9] = 126
      "00101010" when "001010", -- t[10] = 42
      "10000000" when "001011", -- t[11] = 128
      "00101011" when "001100", -- t[12] = 43
      "10000011" when "001101", -- t[13] = 131
      "00101100" when "001110", -- t[14] = 44
      "10000101" when "001111", -- t[15] = 133
      "00101101" when "010000", -- t[16] = 45
      "10001000" when "010001", -- t[17] = 136
      "00101110" when "010010", -- t[18] = 46
      "10001011" when "010011", -- t[19] = 139
      "00101111" when "010100", -- t[20] = 47
      "10001110" when "010101", -- t[21] = 142
      "00110000" when "010110", -- t[22] = 48
      "10010001" when "010111", -- t[23] = 145
      "00110001" when "011000", -- t[24] = 49
      "10010101" when "011001", -- t[25] = 149
      "00110010" when "011010", -- t[26] = 50
      "10011000" when "011011", -- t[27] = 152
      "00110011" when "011100", -- t[28] = 51
      "10011011" when "011101", -- t[29] = 155
      "00110101" when "011110", -- t[30] = 53
      "10011111" when "011111", -- t[31] = 159
      "00110110" when "100000", -- t[32] = 54
      "10100011" when "100001", -- t[33] = 163
      "00110111" when "100010", -- t[34] = 55
      "10100111" when "100011", -- t[35] = 167
      "00111001" when "100100", -- t[36] = 57
      "10101011" when "100101", -- t[37] = 171
      "00111010" when "100110", -- t[38] = 58
      "10101111" when "100111", -- t[39] = 175
      "00111100" when "101000", -- t[40] = 60
      "10110100" when "101001", -- t[41] = 180
      "00111101" when "101010", -- t[42] = 61
      "10111001" when "101011", -- t[43] = 185
      "00111111" when "101100", -- t[44] = 63
      "10111110" when "101101", -- t[45] = 190
      "01000001" when "101110", -- t[46] = 65
      "11000011" when "101111", -- t[47] = 195
      "01000010" when "110000", -- t[48] = 66
      "11001000" when "110001", -- t[49] = 200
      "01000100" when "110010", -- t[50] = 68
      "11001110" when "110011", -- t[51] = 206
      "01000110" when "110100", -- t[52] = 70
      "11010100" when "110101", -- t[53] = 212
      "01001001" when "110110", -- t[54] = 73
      "11011011" when "110111", -- t[55] = 219
      "01001011" when "111000", -- t[56] = 75
      "11100010" when "111001", -- t[57] = 226
      "01001101" when "111010", -- t[58] = 77
      "11101001" when "111011", -- t[59] = 233
      "01010000" when "111100", -- t[60] = 80
      "11110000" when "111101", -- t[61] = 240
      "01010010" when "111110", -- t[62] = 82
      "11111000" when "111111", -- t[63] = 248
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_13_to0 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13_to0 is
begin
  with x select
    r <=
      "0000100" when "000000", -- t[0] = 4
      "0001110" when "000001", -- t[1] = 14
      "0011000" when "000010", -- t[2] = 24
      "0100010" when "000011", -- t[3] = 34
      "0000101" when "000100", -- t[4] = 5
      "0001111" when "000101", -- t[5] = 15
      "0011001" when "000110", -- t[6] = 25
      "0100011" when "000111", -- t[7] = 35
      "0000101" when "001000", -- t[8] = 5
      "0001111" when "001001", -- t[9] = 15
      "0011010" when "001010", -- t[10] = 26
      "0100101" when "001011", -- t[11] = 37
      "0000101" when "001100", -- t[12] = 5
      "0010000" when "001101", -- t[13] = 16
      "0011011" when "001110", -- t[14] = 27
      "0100110" when "001111", -- t[15] = 38
      "0000101" when "010000", -- t[16] = 5
      "0010001" when "010001", -- t[17] = 17
      "0011100" when "010010", -- t[18] = 28
      "0101000" when "010011", -- t[19] = 40
      "0000110" when "010100", -- t[20] = 6
      "0010010" when "010101", -- t[21] = 18
      "0011110" when "010110", -- t[22] = 30
      "0101010" when "010111", -- t[23] = 42
      "0000110" when "011000", -- t[24] = 6
      "0010010" when "011001", -- t[25] = 18
      "0011111" when "011010", -- t[26] = 31
      "0101100" when "011011", -- t[27] = 44
      "0000110" when "011100", -- t[28] = 6
      "0010011" when "011101", -- t[29] = 19
      "0100000" when "011110", -- t[30] = 32
      "0101110" when "011111", -- t[31] = 46
      "0000110" when "100000", -- t[32] = 6
      "0010100" when "100001", -- t[33] = 20
      "0100010" when "100010", -- t[34] = 34
      "0110000" when "100011", -- t[35] = 48
      "0000111" when "100100", -- t[36] = 7
      "0010101" when "100101", -- t[37] = 21
      "0100100" when "100110", -- t[38] = 36
      "0110010" when "100111", -- t[39] = 50
      "0000111" when "101000", -- t[40] = 7
      "0010110" when "101001", -- t[41] = 22
      "0100110" when "101010", -- t[42] = 38
      "0110101" when "101011", -- t[43] = 53
      "0001000" when "101100", -- t[44] = 8
      "0011000" when "101101", -- t[45] = 24
      "0101000" when "101110", -- t[46] = 40
      "0111000" when "101111", -- t[47] = 56
      "0001000" when "110000", -- t[48] = 8
      "0011001" when "110001", -- t[49] = 25
      "0101010" when "110010", -- t[50] = 42
      "0111011" when "110011", -- t[51] = 59
      "0001001" when "110100", -- t[52] = 9
      "0011011" when "110101", -- t[53] = 27
      "0101101" when "110110", -- t[54] = 45
      "0111111" when "110111", -- t[55] = 63
      "0001001" when "111000", -- t[56] = 9
      "0011100" when "111001", -- t[57] = 28
      "0101111" when "111010", -- t[58] = 47
      "1000011" when "111011", -- t[59] = 67
      "0001010" when "111100", -- t[60] = 10
      "0011110" when "111101", -- t[61] = 30
      "0110011" when "111110", -- t[62] = 51
      "1000111" when "111111", -- t[63] = 71
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_13.all;

entity LNSSub_MPT_T5_13_to1_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(7 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T5_13_to1
    port map( x => in_t,
              r => out_t );

  r(16 downto 8) <= (16 downto 8 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_13.all;

entity LNSSub_MPT_T5_13_to0_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(6 downto 0);
begin
  sign <= not b(2);
  in_t(5 downto 2) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T5_13_to0
    port map( x => in_t,
              r => out_t );

  r(16 downto 7) <= (16 downto 7 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_13.all;

entity LNSSub_MPT_T5_13 is
  port( x : in  std_logic_vector(10 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_13 is
  signal in_tiv  : std_logic_vector(5 downto 0);
  signal out_tiv : std_logic_vector(16 downto 0);
  signal a1      : std_logic_vector(4 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(16 downto 0);
  signal a0      : std_logic_vector(3 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(16 downto 0);
  signal sum     : std_logic_vector(16 downto 0);
begin
  in_tiv <= x(10 downto 5);
  inst_tiv : LNSSub_MPT_T5_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(10 downto 6);
  b1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T5_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(10 downto 7);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T5_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(16 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T5_13_Clk is
  port( x   : in  std_logic_vector(10 downto 0);
        r   : out std_logic_vector(11 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T5_13_Clk is
  signal in_tiv_1  : std_logic_vector(5 downto 0);
  signal out_tiv_1 : std_logic_vector(16 downto 0);
  signal out_tiv_2 : std_logic_vector(16 downto 0);
  signal a1_1      : std_logic_vector(4 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(16 downto 0);
  signal out1_2    : std_logic_vector(16 downto 0);
  signal a0_1      : std_logic_vector(3 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(16 downto 0);
  signal out0_2    : std_logic_vector(16 downto 0);
  signal psum1_2     : std_logic_vector(16 downto 0);
  signal psum1_3     : std_logic_vector(16 downto 0);
  signal psum2_2     : std_logic_vector(16 downto 0);
  signal psum2_3     : std_logic_vector(16 downto 0);
  signal sum_3     : std_logic_vector(16 downto 0);
begin
  in_tiv_1 <= x(10 downto 5);
  inst_tiv : LNSSub_MPT_T5_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(10 downto 6);
  b1_1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T5_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(10 downto 7);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T5_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(16 downto 5);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.25 -0.12500000000000003[ -> [0.0 4.0[
-- wI = 10 bits
-- wO = 11 bits
-- Decomposition: 5, 5 / 4, 3 / 2, 3
-- Guard bits: 6
-- Size: 1088 = 17.2^5 + 9.2^5 + 8.2^5

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T6_13 is
  component LNSSub_MPT_T6_13_tiv is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T6_13_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T6_13_to0 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T6_13_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;

  component LNSSub_MPT_T6_13_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(16 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_13_tiv is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13_tiv is
begin
  with x select
    r <=
      "10101010011011110" when "00000", -- t[0] = 87262
      "10101011110001110" when "00001", -- t[1] = 87950
      "10101101001001011" when "00010", -- t[2] = 88651
      "10101110100010011" when "00011", -- t[3] = 89363
      "10101111111101001" when "00100", -- t[4] = 90089
      "10110001011001100" when "00101", -- t[5] = 90828
      "10110010110111100" when "00110", -- t[6] = 91580
      "10110100010111011" when "00111", -- t[7] = 92347
      "10110101111001001" when "01000", -- t[8] = 93129
      "10110111011100110" when "01001", -- t[9] = 93926
      "10111001000010011" when "01010", -- t[10] = 94739
      "10111010101010000" when "01011", -- t[11] = 95568
      "10111100010011110" when "01100", -- t[12] = 96414
      "10111101111111111" when "01101", -- t[13] = 97279
      "10111111101110001" when "01110", -- t[14] = 98161
      "11000001011110111" when "01111", -- t[15] = 99063
      "11000011010010001" when "10000", -- t[16] = 99985
      "11000101001000000" when "10001", -- t[17] = 100928
      "11000111000000101" when "10010", -- t[18] = 101893
      "11001000111100001" when "10011", -- t[19] = 102881
      "11001010111010100" when "10100", -- t[20] = 103892
      "11001100111100001" when "10101", -- t[21] = 104929
      "11001111000000111" when "10110", -- t[22] = 105991
      "11010001001001001" when "10111", -- t[23] = 107081
      "11010011010101000" when "11000", -- t[24] = 108200
      "11010101100100101" when "11001", -- t[25] = 109349
      "11010111111000010" when "11010", -- t[26] = 110530
      "11011010010000001" when "11011", -- t[27] = 111745
      "11011100101100011" when "11100", -- t[28] = 112995
      "11011111001101010" when "11101", -- t[29] = 114282
      "11100001110011001" when "11110", -- t[30] = 115609
      "11100100011110010" when "11111", -- t[31] = 116978
      "-----------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_13_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13_to1 is
begin
  with x select
    r <=
      "001010101" when "00000", -- t[0] = 85
      "100000001" when "00001", -- t[1] = 257
      "001011000" when "00010", -- t[2] = 88
      "100001010" when "00011", -- t[3] = 266
      "001011100" when "00100", -- t[4] = 92
      "100010100" when "00101", -- t[5] = 276
      "001011111" when "00110", -- t[6] = 95
      "100011110" when "00111", -- t[7] = 286
      "001100011" when "01000", -- t[8] = 99
      "100101010" when "01001", -- t[9] = 298
      "001100111" when "01010", -- t[10] = 103
      "100110110" when "01011", -- t[11] = 310
      "001101011" when "01100", -- t[12] = 107
      "101000011" when "01101", -- t[13] = 323
      "001110000" when "01110", -- t[14] = 112
      "101010001" when "01111", -- t[15] = 337
      "001110101" when "10000", -- t[16] = 117
      "101100000" when "10001", -- t[17] = 352
      "001111011" when "10010", -- t[18] = 123
      "101110001" when "10011", -- t[19] = 369
      "010000001" when "10100", -- t[20] = 129
      "110000011" when "10101", -- t[21] = 387
      "010000111" when "10110", -- t[22] = 135
      "110010111" when "10111", -- t[23] = 407
      "010001111" when "11000", -- t[24] = 143
      "110101101" when "11001", -- t[25] = 429
      "010010111" when "11010", -- t[26] = 151
      "111000101" when "11011", -- t[27] = 453
      "010100000" when "11100", -- t[28] = 160
      "111100001" when "11101", -- t[29] = 481
      "010101010" when "11110", -- t[30] = 170
      "111111111" when "11111", -- t[31] = 511
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_13_to0 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13_to0 is
begin
  with x select
    r <=
      "00001010" when "00000", -- t[0] = 10
      "00100000" when "00001", -- t[1] = 32
      "00110110" when "00010", -- t[2] = 54
      "01001100" when "00011", -- t[3] = 76
      "00001011" when "00100", -- t[4] = 11
      "00100011" when "00101", -- t[5] = 35
      "00111010" when "00110", -- t[6] = 58
      "01010010" when "00111", -- t[7] = 82
      "00001100" when "01000", -- t[8] = 12
      "00100110" when "01001", -- t[9] = 38
      "00111111" when "01010", -- t[10] = 63
      "01011000" when "01011", -- t[11] = 88
      "00001101" when "01100", -- t[12] = 13
      "00101001" when "01101", -- t[13] = 41
      "01000100" when "01110", -- t[14] = 68
      "01100000" when "01111", -- t[15] = 96
      "00001111" when "10000", -- t[16] = 15
      "00101101" when "10001", -- t[17] = 45
      "01001011" when "10010", -- t[18] = 75
      "01101001" when "10011", -- t[19] = 105
      "00010000" when "10100", -- t[20] = 16
      "00110001" when "10101", -- t[21] = 49
      "01010010" when "10110", -- t[22] = 82
      "01110100" when "10111", -- t[23] = 116
      "00010010" when "11000", -- t[24] = 18
      "00110111" when "11001", -- t[25] = 55
      "01011100" when "11010", -- t[26] = 92
      "10000001" when "11011", -- t[27] = 129
      "00010100" when "11100", -- t[28] = 20
      "00111110" when "11101", -- t[29] = 62
      "01100111" when "11110", -- t[30] = 103
      "10010001" when "11111", -- t[31] = 145
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_13.all;

entity LNSSub_MPT_T6_13_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(8 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T6_13_to1
    port map( x => in_t,
              r => out_t );

  r(16 downto 9) <= (16 downto 9 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
  r(8) <= out_t(8) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_13.all;

entity LNSSub_MPT_T6_13_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(7 downto 0);
begin
  sign <= not b(2);
  in_t(4 downto 2) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T6_13_to0
    port map( x => in_t,
              r => out_t );

  r(16 downto 8) <= (16 downto 8 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_13.all;

entity LNSSub_MPT_T6_13 is
  port( x : in  std_logic_vector(9 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_13 is
  signal in_tiv  : std_logic_vector(4 downto 0);
  signal out_tiv : std_logic_vector(16 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(16 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(16 downto 0);
  signal sum     : std_logic_vector(16 downto 0);
begin
  in_tiv <= x(9 downto 5);
  inst_tiv : LNSSub_MPT_T6_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(9 downto 6);
  b1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T6_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(9 downto 7);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T6_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(16 downto 6);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T6_13_Clk is
  port( x   : in  std_logic_vector(9 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T6_13_Clk is
  signal in_tiv_1  : std_logic_vector(4 downto 0);
  signal out_tiv_1 : std_logic_vector(16 downto 0);
  signal out_tiv_2 : std_logic_vector(16 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(16 downto 0);
  signal out1_2    : std_logic_vector(16 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(16 downto 0);
  signal out0_2    : std_logic_vector(16 downto 0);
  signal psum1_2     : std_logic_vector(16 downto 0);
  signal psum1_3     : std_logic_vector(16 downto 0);
  signal psum2_2     : std_logic_vector(16 downto 0);
  signal psum2_3     : std_logic_vector(16 downto 0);
  signal sum_3     : std_logic_vector(16 downto 0);
begin
  in_tiv_1 <= x(9 downto 5);
  inst_tiv : LNSSub_MPT_T6_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(9 downto 6);
  b1_1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T6_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(9 downto 7);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T6_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(16 downto 6);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.12500000000000003 -0.0625[ -> [0.0 7.999999999999998[
-- wI = 9 bits
-- wO = 11 bits
-- Decomposition: 4, 5 / 3, 2 / 3, 2
-- Guard bits: 4
-- Size: 528 = 15.2^4 + 8.2^5 + 4.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T7_13 is
  component LNSSub_MPT_T7_13_tiv is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T7_13_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T7_13_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T7_13_to1_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T7_13_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T7_13_tiv is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13_tiv is
begin
  with x select
    r <=
      "011100111010011" when "0000", -- t[0] = 14803
      "011101010001010" when "0001", -- t[1] = 14986
      "011101101000111" when "0010", -- t[2] = 15175
      "011110000001011" when "0011", -- t[3] = 15371
      "011110011010110" when "0100", -- t[4] = 15574
      "011110110101001" when "0101", -- t[5] = 15785
      "011111010000100" when "0110", -- t[6] = 16004
      "011111101101001" when "0111", -- t[7] = 16233
      "100000001010111" when "1000", -- t[8] = 16471
      "100000101010000" when "1001", -- t[9] = 16720
      "100001001010101" when "1010", -- t[10] = 16981
      "100001101100110" when "1011", -- t[11] = 17254
      "100010010000110" when "1100", -- t[12] = 17542
      "100010110110101" when "1101", -- t[13] = 17845
      "100011011110101" when "1110", -- t[14] = 18165
      "100100001001001" when "1111", -- t[15] = 18505
      "---------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T7_13_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13_to1 is
begin
  with x select
    r <=
      "00001011" when "00000", -- t[0] = 11
      "00100010" when "00001", -- t[1] = 34
      "00111000" when "00010", -- t[2] = 56
      "01001111" when "00011", -- t[3] = 79
      "00001100" when "00100", -- t[4] = 12
      "00100100" when "00101", -- t[5] = 36
      "00111101" when "00110", -- t[6] = 61
      "01010101" when "00111", -- t[7] = 85
      "00001101" when "01000", -- t[8] = 13
      "00100111" when "01001", -- t[9] = 39
      "01000001" when "01010", -- t[10] = 65
      "01011100" when "01011", -- t[11] = 92
      "00001110" when "01100", -- t[12] = 14
      "00101010" when "01101", -- t[13] = 42
      "01000111" when "01110", -- t[14] = 71
      "01100011" when "01111", -- t[15] = 99
      "00001111" when "10000", -- t[16] = 15
      "00101110" when "10001", -- t[17] = 46
      "01001101" when "10010", -- t[18] = 77
      "01101100" when "10011", -- t[19] = 108
      "00010001" when "10100", -- t[20] = 17
      "00110011" when "10101", -- t[21] = 51
      "01010101" when "10110", -- t[22] = 85
      "01110111" when "10111", -- t[23] = 119
      "00010010" when "11000", -- t[24] = 18
      "00111000" when "11001", -- t[25] = 56
      "01011110" when "11010", -- t[26] = 94
      "10000100" when "11011", -- t[27] = 132
      "00010101" when "11100", -- t[28] = 21
      "00111111" when "11101", -- t[29] = 63
      "01101001" when "11110", -- t[30] = 105
      "10010100" when "11111", -- t[31] = 148
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T7_13_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13_to0 is
begin
  with x select
    r <=
      "0010" when "000", -- t[0] = 2
      "1000" when "001", -- t[1] = 8
      "0011" when "010", -- t[2] = 3
      "1010" when "011", -- t[3] = 10
      "0100" when "100", -- t[4] = 4
      "1100" when "101", -- t[5] = 12
      "0101" when "110", -- t[6] = 5
      "1111" when "111", -- t[7] = 15
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_13.all;

entity LNSSub_MPT_T7_13_to1_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(7 downto 0);
begin
  sign <= not b(2);
  in_t(4 downto 2) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to1 : LNSSub_MPT_T7_13_to1
    port map( x => in_t,
              r => out_t );

  r(14 downto 8) <= (14 downto 8 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_13.all;

entity LNSSub_MPT_T7_13_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T7_13_to0
    port map( x => in_t,
              r => out_t );

  r(14 downto 4) <= (14 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_13.all;

entity LNSSub_MPT_T7_13 is
  port( x : in  std_logic_vector(8 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_13 is
  signal in_tiv  : std_logic_vector(3 downto 0);
  signal out_tiv : std_logic_vector(14 downto 0);
  signal a1      : std_logic_vector(2 downto 0);
  signal b1      : std_logic_vector(2 downto 0);
  signal out1    : std_logic_vector(14 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(14 downto 0);
  signal sum     : std_logic_vector(14 downto 0);
begin
  in_tiv <= x(8 downto 5);
  inst_tiv : LNSSub_MPT_T7_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(8 downto 6);
  b1 <= x(4 downto 2);
  inst_to1_xor : LNSSub_MPT_T7_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(8 downto 7);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T7_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(14 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T7_13_Clk is
  port( x   : in  std_logic_vector(8 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T7_13_Clk is
  signal in_tiv_1  : std_logic_vector(3 downto 0);
  signal out_tiv_1 : std_logic_vector(14 downto 0);
  signal out_tiv_2 : std_logic_vector(14 downto 0);
  signal a1_1      : std_logic_vector(2 downto 0);
  signal b1_1      : std_logic_vector(2 downto 0);
  signal out1_1    : std_logic_vector(14 downto 0);
  signal out1_2    : std_logic_vector(14 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(14 downto 0);
  signal out0_2    : std_logic_vector(14 downto 0);
  signal psum1_2     : std_logic_vector(14 downto 0);
  signal psum1_3     : std_logic_vector(14 downto 0);
  signal psum2_2     : std_logic_vector(14 downto 0);
  signal psum2_3     : std_logic_vector(14 downto 0);
  signal sum_3     : std_logic_vector(14 downto 0);
begin
  in_tiv_1 <= x(8 downto 5);
  inst_tiv : LNSSub_MPT_T7_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(8 downto 6);
  b1_1 <= x(4 downto 2);
  inst_to1_xor : LNSSub_MPT_T7_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(8 downto 7);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T7_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(14 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.0625 -0.03125[ -> [0.0 7.999999999999998[
-- wI = 8 bits
-- wO = 10 bits
-- Decomposition: 4, 4 / 3, 1 / 2, 2
-- Guard bits: 3
-- Size: 300 = 13.2^4 + 5.2^4 + 3.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T8_13 is
  component LNSSub_MPT_T8_13_tiv is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T8_13_to1 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T8_13_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T8_13_to1_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T8_13_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_13_tiv is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13_tiv is
begin
  with x select
    r <=
      "1001001010111" when "0000", -- t[0] = 4695
      "1001010000110" when "0001", -- t[1] = 4742
      "1001010110110" when "0010", -- t[2] = 4790
      "1001011101000" when "0011", -- t[3] = 4840
      "1001100011100" when "0100", -- t[4] = 4892
      "1001101010010" when "0101", -- t[5] = 4946
      "1001110001001" when "0110", -- t[6] = 5001
      "1001111000011" when "0111", -- t[7] = 5059
      "1010000000000" when "1000", -- t[8] = 5120
      "1010000111111" when "1001", -- t[9] = 5183
      "1010010000001" when "1010", -- t[10] = 5249
      "1010011000110" when "1011", -- t[11] = 5318
      "1010100001111" when "1100", -- t[12] = 5391
      "1010101011100" when "1101", -- t[13] = 5468
      "1010110101101" when "1110", -- t[14] = 5549
      "1011000000011" when "1111", -- t[15] = 5635
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_13_to1 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13_to1 is
begin
  with x select
    r <=
      "00101" when "0000", -- t[0] = 5
      "10001" when "0001", -- t[1] = 17
      "00110" when "0010", -- t[2] = 6
      "10010" when "0011", -- t[3] = 18
      "00110" when "0100", -- t[4] = 6
      "10100" when "0101", -- t[5] = 20
      "00111" when "0110", -- t[6] = 7
      "10101" when "0111", -- t[7] = 21
      "00111" when "1000", -- t[8] = 7
      "10111" when "1001", -- t[9] = 23
      "01000" when "1010", -- t[10] = 8
      "11001" when "1011", -- t[11] = 25
      "01001" when "1100", -- t[12] = 9
      "11100" when "1101", -- t[13] = 28
      "01010" when "1110", -- t[14] = 10
      "11111" when "1111", -- t[15] = 31
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_13_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13_to0 is
begin
  with x select
    r <=
      "001" when "00", -- t[0] = 1
      "100" when "01", -- t[1] = 4
      "010" when "10", -- t[2] = 2
      "110" when "11", -- t[3] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_13.all;

entity LNSSub_MPT_T8_13_to1_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T8_13_to1
    port map( x => in_t,
              r => out_t );

  r(12 downto 5) <= (12 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_13.all;

entity LNSSub_MPT_T8_13_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T8_13_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 3) <= (12 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_13.all;

entity LNSSub_MPT_T8_13 is
  port( x : in  std_logic_vector(7 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_13 is
  signal in_tiv  : std_logic_vector(3 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a1      : std_logic_vector(2 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(7 downto 4);
  inst_tiv : LNSSub_MPT_T8_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(7 downto 5);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T8_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(7 downto 7);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T8_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(12 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T8_13_Clk is
  port( x   : in  std_logic_vector(7 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T8_13_Clk is
  signal in_tiv_1  : std_logic_vector(3 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a1_1      : std_logic_vector(2 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(12 downto 0);
  signal out1_2    : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(7 downto 4);
  inst_tiv : LNSSub_MPT_T8_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(7 downto 5);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T8_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(7 downto 7);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T8_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.03125 -0.015625000000000007[ -> [0.0 7.999999999999998[
-- wI = 7 bits
-- wO = 9 bits
-- Decomposition: 3, 4 / 2, 1 / 2, 2
-- Guard bits: 4
-- Size: 168 = 13.2^3 + 6.2^3 + 4.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T9_13 is
  component LNSSub_MPT_T9_13_tiv is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T9_13_to1 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T9_13_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T9_13_to1_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T9_13_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_13_tiv is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13_tiv is
begin
  with x select
    r <=
      "1011001100010" when "000", -- t[0] = 5730
      "1011011000011" when "001", -- t[1] = 5827
      "1011100101100" when "010", -- t[2] = 5932
      "1011110011101" when "011", -- t[3] = 6045
      "1100000010111" when "100", -- t[4] = 6167
      "1100010011100" when "101", -- t[5] = 6300
      "1100100101111" when "110", -- t[6] = 6447
      "1100111010010" when "111", -- t[7] = 6610
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_13_to1 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13_to1 is
begin
  with x select
    r <=
      "001100" when "000", -- t[0] = 12
      "100100" when "001", -- t[1] = 36
      "001101" when "010", -- t[2] = 13
      "101001" when "011", -- t[3] = 41
      "010000" when "100", -- t[4] = 16
      "110001" when "101", -- t[5] = 49
      "010100" when "110", -- t[6] = 20
      "111100" when "111", -- t[7] = 60
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_13_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13_to0 is
begin
  with x select
    r <=
      "0011" when "00", -- t[0] = 3
      "1001" when "01", -- t[1] = 9
      "0100" when "10", -- t[2] = 4
      "1101" when "11", -- t[3] = 13
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_13.all;

entity LNSSub_MPT_T9_13_to1_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(5 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T9_13_to1
    port map( x => in_t,
              r => out_t );

  r(12 downto 6) <= (12 downto 6 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_13.all;

entity LNSSub_MPT_T9_13_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T9_13_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 4) <= (12 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_13.all;

entity LNSSub_MPT_T9_13 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_13 is
  signal in_tiv  : std_logic_vector(2 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a1      : std_logic_vector(1 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(6 downto 4);
  inst_tiv : LNSSub_MPT_T9_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(6 downto 5);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T9_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(6 downto 6);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T9_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(12 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T9_13_Clk is
  port( x   : in  std_logic_vector(6 downto 0);
        r   : out std_logic_vector(8 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T9_13_Clk is
  signal in_tiv_1  : std_logic_vector(2 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a1_1      : std_logic_vector(1 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(12 downto 0);
  signal out1_2    : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(6 downto 4);
  inst_tiv : LNSSub_MPT_T9_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(6 downto 5);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T9_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(6 downto 6);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T9_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.015625000000000007 -0.007812500000000002[ -> [0.0 7.999999999999998[
-- wI = 6 bits
-- wO = 8 bits
-- Decomposition: 2, 4 / 2, 1 / 2, 2
-- Guard bits: 3
-- Size: 96 = 11.2^2 + 5.2^3 + 3.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T10_13 is
  component LNSSub_MPT_T10_13_tiv is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T10_13_to1 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T10_13_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T10_13_to1_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T10_13_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T10_13_tiv is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13_tiv is
begin
  with x select
    r <=
      "11010100101" when "00", -- t[0] = 1701
      "11011011001" when "01", -- t[1] = 1753
      "11100010111" when "10", -- t[2] = 1815
      "11101100001" when "11", -- t[3] = 1889
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T10_13_to1 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13_to1 is
begin
  with x select
    r <=
      "00110" when "000", -- t[0] = 6
      "10010" when "001", -- t[1] = 18
      "00110" when "010", -- t[2] = 6
      "10100" when "011", -- t[3] = 20
      "01000" when "100", -- t[4] = 8
      "11000" when "101", -- t[5] = 24
      "01001" when "110", -- t[6] = 9
      "11101" when "111", -- t[7] = 29
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T10_13_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13_to0 is
begin
  with x select
    r <=
      "001" when "00", -- t[0] = 1
      "100" when "01", -- t[1] = 4
      "010" when "10", -- t[2] = 2
      "110" when "11", -- t[3] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_13.all;

entity LNSSub_MPT_T10_13_to1_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T10_13_to1
    port map( x => in_t,
              r => out_t );

  r(10 downto 5) <= (10 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_13.all;

entity LNSSub_MPT_T10_13_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T10_13_to0
    port map( x => in_t,
              r => out_t );

  r(10 downto 3) <= (10 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_13.all;

entity LNSSub_MPT_T10_13 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_13 is
  signal in_tiv  : std_logic_vector(1 downto 0);
  signal out_tiv : std_logic_vector(10 downto 0);
  signal a1      : std_logic_vector(1 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(10 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(10 downto 0);
  signal sum     : std_logic_vector(10 downto 0);
begin
  in_tiv <= x(5 downto 4);
  inst_tiv : LNSSub_MPT_T10_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(5 downto 4);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T10_13_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(5 downto 5);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T10_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(10 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T10_13_Clk is
  port( x   : in  std_logic_vector(5 downto 0);
        r   : out std_logic_vector(7 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T10_13_Clk is
  signal in_tiv_1  : std_logic_vector(1 downto 0);
  signal out_tiv_1 : std_logic_vector(10 downto 0);
  signal out_tiv_2 : std_logic_vector(10 downto 0);
  signal a1_1      : std_logic_vector(1 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(10 downto 0);
  signal out1_2    : std_logic_vector(10 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(10 downto 0);
  signal out0_2    : std_logic_vector(10 downto 0);
  signal psum1_2     : std_logic_vector(10 downto 0);
  signal psum1_3     : std_logic_vector(10 downto 0);
  signal psum2_2     : std_logic_vector(10 downto 0);
  signal psum2_3     : std_logic_vector(10 downto 0);
  signal sum_3     : std_logic_vector(10 downto 0);
begin
  in_tiv_1 <= x(5 downto 4);
  inst_tiv : LNSSub_MPT_T10_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(5 downto 4);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T10_13_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(5 downto 5);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T10_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(10 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.007812500000000002 -0.003906250000000001[ -> [0.0 15.999999999999998[
-- wI = 5 bits
-- wO = 8 bits
-- Decomposition: 3, 2 / 1 / 2
-- Guard bits: 3
-- Size: 100 = 11.2^3 + 3.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T11_13 is
  component LNSSub_MPT_T11_13_tiv is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T11_13_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T11_13_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T11_13_tiv is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_13_tiv is
begin
  with x select
    r <=
      "01111001101" when "000", -- t[0] = 973
      "01111011001" when "001", -- t[1] = 985
      "01111100110" when "010", -- t[2] = 998
      "01111110100" when "011", -- t[3] = 1012
      "10000000011" when "100", -- t[4] = 1027
      "10000010100" when "101", -- t[5] = 1044
      "10000100110" when "110", -- t[6] = 1062
      "10000111010" when "111", -- t[7] = 1082
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T11_13_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_13_to0 is
begin
  with x select
    r <=
      "001" when "00", -- t[0] = 1
      "100" when "01", -- t[1] = 4
      "010" when "10", -- t[2] = 2
      "110" when "11", -- t[3] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_13.all;

entity LNSSub_MPT_T11_13_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T11_13_to0
    port map( x => in_t,
              r => out_t );

  r(10 downto 3) <= (10 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_13.all;

entity LNSSub_MPT_T11_13 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_13 is
  signal in_tiv  : std_logic_vector(2 downto 0);
  signal out_tiv : std_logic_vector(10 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(10 downto 0);
  signal sum     : std_logic_vector(10 downto 0);
begin
  in_tiv <= x(4 downto 2);
  inst_tiv : LNSSub_MPT_T11_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a0 <= x(4 downto 4);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T11_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(10 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T11_13_Clk is
  port( x   : in  std_logic_vector(4 downto 0);
        r   : out std_logic_vector(7 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T11_13_Clk is
  signal in_tiv_1  : std_logic_vector(2 downto 0);
  signal out_tiv_1 : std_logic_vector(10 downto 0);
  signal out_tiv_2 : std_logic_vector(10 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(10 downto 0);
  signal out0_2    : std_logic_vector(10 downto 0);
  signal psum1_2     : std_logic_vector(10 downto 0);
  signal psum1_3     : std_logic_vector(10 downto 0);
  signal psum2_2     : std_logic_vector(10 downto 0);
  signal psum2_3     : std_logic_vector(10 downto 0);
  signal sum_3     : std_logic_vector(10 downto 0);
begin
  in_tiv_1 <= x(4 downto 2);
  inst_tiv : LNSSub_MPT_T11_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a0_1 <= x(4 downto 4);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T11_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(10 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.003906250000000001 -0.001953125[ -> [0.0 15.999999999999998[
-- wI = 4 bits
-- wO = 7 bits
-- Decomposition: 1, 3 / 0 / 3
-- Guard bits: 4
-- Size: 42 = 11.2^1 + 5.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T12_13 is
  component LNSSub_MPT_T12_13_tiv is
    port( x : in  std_logic_vector(0 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T12_13_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T12_13_to0_xor is
    port( b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T12_13_tiv is
  port( x : in  std_logic_vector(0 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_13_tiv is
begin
  with x select
    r <=
      "10001100011" when "0", -- t[0] = 1123
      "10010100001" when "1", -- t[1] = 1185
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T12_13_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_13_to0 is
begin
  with x select
    r <=
      "00011" when "00", -- t[0] = 3
      "01011" when "01", -- t[1] = 11
      "10010" when "10", -- t[2] = 18
      "11010" when "11", -- t[3] = 26
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_13.all;

entity LNSSub_MPT_T12_13_to0_xor is
  port( b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(2);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T12_13_to0
    port map( x => in_t,
              r => out_t );

  r(10 downto 5) <= (10 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_13.all;

entity LNSSub_MPT_T12_13 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_13 is
  signal in_tiv  : std_logic_vector(0 downto 0);
  signal out_tiv : std_logic_vector(10 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(10 downto 0);
  signal sum     : std_logic_vector(10 downto 0);
begin
  in_tiv <= x(3 downto 3);
  inst_tiv : LNSSub_MPT_T12_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T12_13_to0_xor
    port map( b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(10 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T12_13_Clk is
  port( x   : in  std_logic_vector(3 downto 0);
        r   : out std_logic_vector(6 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T12_13_Clk is
  signal in_tiv_1  : std_logic_vector(0 downto 0);
  signal out_tiv_1 : std_logic_vector(10 downto 0);
  signal out_tiv_2 : std_logic_vector(10 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(10 downto 0);
  signal out0_2    : std_logic_vector(10 downto 0);
  signal psum1_2     : std_logic_vector(10 downto 0);
  signal psum1_3     : std_logic_vector(10 downto 0);
  signal psum2_2     : std_logic_vector(10 downto 0);
  signal psum2_3     : std_logic_vector(10 downto 0);
  signal sum_3     : std_logic_vector(10 downto 0);
begin
  in_tiv_1 <= x(3 downto 3);
  inst_tiv : LNSSub_MPT_T12_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T12_13_to0_xor
    port map( b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(10 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.001953125 0.0[ -> [0.0 15.999999999999998[
-- wI = 4 bits
-- wO = 7 bits
-- Decomposition: 2, 2 / 2 / 2
-- Guard bits: 0
-- Size: 52 = 7.2^2 + 3.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T13_13 is
  component LNSSub_MPT_T13_13_tiv is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T13_13_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T13_13_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T13_13_tiv is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T13_13_tiv is
begin
  with x select
    r <=
      "1001110" when "00", -- t[0] = 78
      "1010010" when "01", -- t[1] = 82
      "1010111" when "10", -- t[2] = 87
      "1100101" when "11", -- t[3] = 101
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T13_13_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T13_13_to0 is
begin
  with x select
    r <=
      "000" when "000", -- t[0] = 0
      "001" when "001", -- t[1] = 1
      "000" when "010", -- t[2] = 0
      "001" when "011", -- t[3] = 1
      "000" when "100", -- t[4] = 0
      "010" when "101", -- t[5] = 2
      "010" when "110", -- t[6] = 2
      "111" when "111", -- t[7] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T13_13.all;

entity LNSSub_MPT_T13_13_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T13_13_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T13_13_to0
    port map( x => in_t,
              r => out_t );

  r(6 downto 3) <= (6 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T13_13.all;

entity LNSSub_MPT_T13_13 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T13_13 is
  signal in_tiv  : std_logic_vector(1 downto 0);
  signal out_tiv : std_logic_vector(6 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(6 downto 0);
  signal sum     : std_logic_vector(6 downto 0);
begin
  in_tiv <= x(3 downto 2);
  inst_tiv : LNSSub_MPT_T13_13_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a0 <= x(3 downto 2);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T13_13_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(6 downto 0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T13_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T13_13_Clk is
  port( x   : in  std_logic_vector(3 downto 0);
        r   : out std_logic_vector(6 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T13_13_Clk is
  signal in_tiv_1  : std_logic_vector(1 downto 0);
  signal out_tiv_1 : std_logic_vector(6 downto 0);
  signal out_tiv_2 : std_logic_vector(6 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(6 downto 0);
  signal out0_2    : std_logic_vector(6 downto 0);
  signal psum1_2     : std_logic_vector(6 downto 0);
  signal psum1_3     : std_logic_vector(6 downto 0);
  signal psum2_2     : std_logic_vector(6 downto 0);
  signal psum2_3     : std_logic_vector(6 downto 0);
  signal sum_3     : std_logic_vector(6 downto 0);
begin
  in_tiv_1 <= x(3 downto 2);
  inst_tiv : LNSSub_MPT_T13_13_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a0_1 <= x(3 downto 2);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T13_13_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(6 downto 0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnssub_mpt_13.all;

entity LNSSub_MPT_13 is
  port( x : in  std_logic_vector(16 downto 0);
        r : out std_logic_vector(16 downto 0) );
end entity;

architecture arch of LNSSub_MPT_13 is

  signal out_t0 : std_logic_vector(6 downto 0);
  signal out_t1 : std_logic_vector(9 downto 0);
  signal out_t2 : std_logic_vector(11 downto 0);
  signal out_t3 : std_logic_vector(11 downto 0);
  signal out_t4 : std_logic_vector(11 downto 0);
  signal out_t5 : std_logic_vector(11 downto 0);
  signal out_t6 : std_logic_vector(10 downto 0);
  signal out_t7 : std_logic_vector(10 downto 0);
  signal out_t8 : std_logic_vector(9 downto 0);
  signal out_t9 : std_logic_vector(8 downto 0);
  signal out_t10 : std_logic_vector(7 downto 0);
  signal out_t11 : std_logic_vector(7 downto 0);
  signal out_t12 : std_logic_vector(6 downto 0);
  signal out_t13 : std_logic_vector(6 downto 0);
begin
  inst_t0 : LNSSub_MPT_T0_13
    port map( x => x,
              r => out_t0 );

  inst_t1 : LNSSub_MPT_T1_13
    port map( x => x(14 downto 0),
              r => out_t1 );

  inst_t2 : LNSSub_MPT_T2_13
    port map( x => x(13 downto 0),
              r => out_t2 );

  inst_t3 : LNSSub_MPT_T3_13
    port map( x => x(12 downto 0),
              r => out_t3 );

  inst_t4 : LNSSub_MPT_T4_13
    port map( x => x(11 downto 0),
              r => out_t4 );

  inst_t5 : LNSSub_MPT_T5_13
    port map( x => x(10 downto 0),
              r => out_t5 );

  inst_t6 : LNSSub_MPT_T6_13
    port map( x => x(9 downto 0),
              r => out_t6 );

  inst_t7 : LNSSub_MPT_T7_13
    port map( x => x(8 downto 0),
              r => out_t7 );

  inst_t8 : LNSSub_MPT_T8_13
    port map( x => x(7 downto 0),
              r => out_t8 );

  inst_t9 : LNSSub_MPT_T9_13
    port map( x => x(6 downto 0),
              r => out_t9 );

  inst_t10 : LNSSub_MPT_T10_13
    port map( x => x(5 downto 0),
              r => out_t10 );

  inst_t11 : LNSSub_MPT_T11_13
    port map( x => x(4 downto 0),
              r => out_t11 );

  inst_t12 : LNSSub_MPT_T12_13
    port map( x => x(3 downto 0),
              r => out_t12 );

  inst_t13 : LNSSub_MPT_T13_13
    port map( x => x(3 downto 0),
              r => out_t13 );

  r <= (16 downto 7 => '0') & out_t0
         when x(16 downto 16) /= (16 downto 16 => '1') else
       (16 downto 10 => '0') & out_t1
         when x(15) /= '1' else
       (16 downto 12 => '0') & out_t2
         when x(14) /= '1' else
       (16 downto 13 => '0') & out_t3 & (0 downto 0 => '0')
         when x(13) /= '1' else
       (16 downto 14 => '0') & out_t4 & (1 downto 0 => '0')
         when x(12) /= '1' else
       (16 downto 15 => '0') & out_t5 & (2 downto 0 => '0')
         when x(11) /= '1' else
       (16 downto 15 => '0') & out_t6 & (3 downto 0 => '0')
         when x(10) /= '1' else
       (16 downto 16 => '0') & out_t7 & (4 downto 0 => '0')
         when x(9) /= '1' else
       (16 downto 16 => '0') & out_t8 & (5 downto 0 => '0')
         when x(8) /= '1' else
       (16 downto 16 => '0') & out_t9 & (6 downto 0 => '0')
         when x(7) /= '1' else
       (16 downto 16 => '0') & out_t10 & (7 downto 0 => '0')
         when x(6) /= '1' else
       out_t11 & (8 downto 0 => '0')
         when x(5) /= '1' else
       out_t12 & (9 downto 0 => '0')
         when x(4) /= '1' else
       out_t13 & (9 downto 0 => '0');
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnssub_mpt_13.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_13_Clk is
  port( x   : in  std_logic_vector(16 downto 0);
        r   : out std_logic_vector(16 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_13_Clk is
  signal x_1  : std_logic_vector(16 downto 0);
  signal x_10 : std_logic_vector(16 downto 0);

  signal out_t0_1  : std_logic_vector(6 downto 0);
  signal out_t0_10 : std_logic_vector(6 downto 0);
  signal out_t1_10 : std_logic_vector(9 downto 0);
  signal out_t2_10 : std_logic_vector(11 downto 0);
  signal out_t3_10 : std_logic_vector(11 downto 0);
  signal out_t4_10 : std_logic_vector(11 downto 0);
  signal out_t5_10 : std_logic_vector(11 downto 0);
  signal out_t6_10 : std_logic_vector(10 downto 0);
  signal out_t7_10 : std_logic_vector(10 downto 0);
  signal out_t8_10 : std_logic_vector(9 downto 0);
  signal out_t9_10 : std_logic_vector(8 downto 0);
  signal out_t10_10 : std_logic_vector(7 downto 0);
  signal out_t11_10 : std_logic_vector(7 downto 0);
  signal out_t12_10 : std_logic_vector(6 downto 0);
  signal out_t13_10 : std_logic_vector(6 downto 0);
begin
  x_1 <= x;

  inst_t0 : LNSSub_MPT_T0_13
    port map( x   => x_1,
              r   => out_t0_1 );

  out_t0_delay : Delay
    generic map ( w => 7,
                  n => 1 )
    port map ( input  => out_t0_1,
               output => out_t0_10,
               clk    => clk );

  inst_t1 : LNSSub_MPT_T1_13_Clk
    port map( x   => x_1(14 downto 0),
              r   => out_t1_10,
              clk => clk );

  inst_t2 : LNSSub_MPT_T2_13_Clk
    port map( x   => x_1(13 downto 0),
              r   => out_t2_10,
              clk => clk );

  inst_t3 : LNSSub_MPT_T3_13_Clk
    port map( x   => x_1(12 downto 0),
              r   => out_t3_10,
              clk => clk );

  inst_t4 : LNSSub_MPT_T4_13_Clk
    port map( x   => x_1(11 downto 0),
              r   => out_t4_10,
              clk => clk );

  inst_t5 : LNSSub_MPT_T5_13_Clk
    port map( x   => x_1(10 downto 0),
              r   => out_t5_10,
              clk => clk );

  inst_t6 : LNSSub_MPT_T6_13_Clk
    port map( x   => x_1(9 downto 0),
              r   => out_t6_10,
              clk => clk );

  inst_t7 : LNSSub_MPT_T7_13_Clk
    port map( x   => x_1(8 downto 0),
              r   => out_t7_10,
              clk => clk );

  inst_t8 : LNSSub_MPT_T8_13_Clk
    port map( x   => x_1(7 downto 0),
              r   => out_t8_10,
              clk => clk );

  inst_t9 : LNSSub_MPT_T9_13_Clk
    port map( x   => x_1(6 downto 0),
              r   => out_t9_10,
              clk => clk );

  inst_t10 : LNSSub_MPT_T10_13_Clk
    port map( x   => x_1(5 downto 0),
              r   => out_t10_10,
              clk => clk );

  inst_t11 : LNSSub_MPT_T11_13_Clk
    port map( x   => x_1(4 downto 0),
              r   => out_t11_10,
              clk => clk );

  inst_t12 : LNSSub_MPT_T12_13_Clk
    port map( x   => x_1(3 downto 0),
              r   => out_t12_10,
              clk => clk );

  inst_t13 : LNSSub_MPT_T13_13_Clk
    port map( x   => x_1(3 downto 0),
              r   => out_t13_10,
              clk => clk );

  x_delay : Delay
    generic map ( w => 17,
                  n => 1 )
    port map ( input  => x_1,
               output => x_10,
               clk    => clk );

  r <= (16 downto 7 => '0') & out_t0_10
         when x_10(16 downto 16) /= (16 downto 16 => '1') else
       (16 downto 10 => '0') & out_t1_10
         when x_10(15) /= '1' else
       (16 downto 12 => '0') & out_t2_10
         when x_10(14) /= '1' else
       (16 downto 13 => '0') & out_t3_10 & (0 downto 0 => '0')
         when x_10(13) /= '1' else
       (16 downto 14 => '0') & out_t4_10 & (1 downto 0 => '0')
         when x_10(12) /= '1' else
       (16 downto 15 => '0') & out_t5_10 & (2 downto 0 => '0')
         when x_10(11) /= '1' else
       (16 downto 15 => '0') & out_t6_10 & (3 downto 0 => '0')
         when x_10(10) /= '1' else
       (16 downto 16 => '0') & out_t7_10 & (4 downto 0 => '0')
         when x_10(9) /= '1' else
       (16 downto 16 => '0') & out_t8_10 & (5 downto 0 => '0')
         when x_10(8) /= '1' else
       (16 downto 16 => '0') & out_t9_10 & (6 downto 0 => '0')
         when x_10(7) /= '1' else
       (16 downto 16 => '0') & out_t10_10 & (7 downto 0 => '0')
         when x_10(6) /= '1' else
       out_t11_10 & (8 downto 0 => '0')
         when x_10(5) /= '1' else
       out_t12_10 & (9 downto 0 => '0')
         when x_10(4) /= '1' else
       out_t13_10 & (9 downto 0 => '0');
end architecture;
