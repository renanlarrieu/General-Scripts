library verilog;
use verilog.vl_types.all;
entity my_and_vlg_vec_tst is
end my_and_vlg_vec_tst;
