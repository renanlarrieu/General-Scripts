-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of LNS sub function with 8-bit integer part and 11-bit fractional part
-- wI = 15 bits
-- wO = 15 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnssub_mnmx_11 is
  component LNSSub_MNMX_T0_11 is
    port ( x : in  std_logic_vector(14 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11 is
    port ( x : in  std_logic_vector(12 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11 is
    port ( x : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11 is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11 is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11 is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11 is
    port ( x : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11 is
    port ( x : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11 is
    port ( x : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T10_11 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
end package;


-- Simple table: LNS subtraction function [ -16.000000, 0.000000 [ -> [ 0.000000, 0.015625 [
-- (restricted to [ -16.000000, -8.000000 [ )
-- Input:  wE =   4, wF =  11, w =  15
-- Output: wE =  -6, wF =  11, w =   5

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T0_11 is
  port ( x : in  std_logic_vector(14 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T0_11 is
begin
  with x select
    r <=
      "00000" when "000000000000000", -- t[0] = 0
      "00000" when "000000000000001", -- t[1] = 0
      "00000" when "000000000000010", -- t[2] = 0
      "00000" when "000000000000011", -- t[3] = 0
      "00000" when "000000000000100", -- t[4] = 0
      "00000" when "000000000000101", -- t[5] = 0
      "00000" when "000000000000110", -- t[6] = 0
      "00000" when "000000000000111", -- t[7] = 0
      "00000" when "000000000001000", -- t[8] = 0
      "00000" when "000000000001001", -- t[9] = 0
      "00000" when "000000000001010", -- t[10] = 0
      "00000" when "000000000001011", -- t[11] = 0
      "00000" when "000000000001100", -- t[12] = 0
      "00000" when "000000000001101", -- t[13] = 0
      "00000" when "000000000001110", -- t[14] = 0
      "00000" when "000000000001111", -- t[15] = 0
      "00000" when "000000000010000", -- t[16] = 0
      "00000" when "000000000010001", -- t[17] = 0
      "00000" when "000000000010010", -- t[18] = 0
      "00000" when "000000000010011", -- t[19] = 0
      "00000" when "000000000010100", -- t[20] = 0
      "00000" when "000000000010101", -- t[21] = 0
      "00000" when "000000000010110", -- t[22] = 0
      "00000" when "000000000010111", -- t[23] = 0
      "00000" when "000000000011000", -- t[24] = 0
      "00000" when "000000000011001", -- t[25] = 0
      "00000" when "000000000011010", -- t[26] = 0
      "00000" when "000000000011011", -- t[27] = 0
      "00000" when "000000000011100", -- t[28] = 0
      "00000" when "000000000011101", -- t[29] = 0
      "00000" when "000000000011110", -- t[30] = 0
      "00000" when "000000000011111", -- t[31] = 0
      "00000" when "000000000100000", -- t[32] = 0
      "00000" when "000000000100001", -- t[33] = 0
      "00000" when "000000000100010", -- t[34] = 0
      "00000" when "000000000100011", -- t[35] = 0
      "00000" when "000000000100100", -- t[36] = 0
      "00000" when "000000000100101", -- t[37] = 0
      "00000" when "000000000100110", -- t[38] = 0
      "00000" when "000000000100111", -- t[39] = 0
      "00000" when "000000000101000", -- t[40] = 0
      "00000" when "000000000101001", -- t[41] = 0
      "00000" when "000000000101010", -- t[42] = 0
      "00000" when "000000000101011", -- t[43] = 0
      "00000" when "000000000101100", -- t[44] = 0
      "00000" when "000000000101101", -- t[45] = 0
      "00000" when "000000000101110", -- t[46] = 0
      "00000" when "000000000101111", -- t[47] = 0
      "00000" when "000000000110000", -- t[48] = 0
      "00000" when "000000000110001", -- t[49] = 0
      "00000" when "000000000110010", -- t[50] = 0
      "00000" when "000000000110011", -- t[51] = 0
      "00000" when "000000000110100", -- t[52] = 0
      "00000" when "000000000110101", -- t[53] = 0
      "00000" when "000000000110110", -- t[54] = 0
      "00000" when "000000000110111", -- t[55] = 0
      "00000" when "000000000111000", -- t[56] = 0
      "00000" when "000000000111001", -- t[57] = 0
      "00000" when "000000000111010", -- t[58] = 0
      "00000" when "000000000111011", -- t[59] = 0
      "00000" when "000000000111100", -- t[60] = 0
      "00000" when "000000000111101", -- t[61] = 0
      "00000" when "000000000111110", -- t[62] = 0
      "00000" when "000000000111111", -- t[63] = 0
      "00000" when "000000001000000", -- t[64] = 0
      "00000" when "000000001000001", -- t[65] = 0
      "00000" when "000000001000010", -- t[66] = 0
      "00000" when "000000001000011", -- t[67] = 0
      "00000" when "000000001000100", -- t[68] = 0
      "00000" when "000000001000101", -- t[69] = 0
      "00000" when "000000001000110", -- t[70] = 0
      "00000" when "000000001000111", -- t[71] = 0
      "00000" when "000000001001000", -- t[72] = 0
      "00000" when "000000001001001", -- t[73] = 0
      "00000" when "000000001001010", -- t[74] = 0
      "00000" when "000000001001011", -- t[75] = 0
      "00000" when "000000001001100", -- t[76] = 0
      "00000" when "000000001001101", -- t[77] = 0
      "00000" when "000000001001110", -- t[78] = 0
      "00000" when "000000001001111", -- t[79] = 0
      "00000" when "000000001010000", -- t[80] = 0
      "00000" when "000000001010001", -- t[81] = 0
      "00000" when "000000001010010", -- t[82] = 0
      "00000" when "000000001010011", -- t[83] = 0
      "00000" when "000000001010100", -- t[84] = 0
      "00000" when "000000001010101", -- t[85] = 0
      "00000" when "000000001010110", -- t[86] = 0
      "00000" when "000000001010111", -- t[87] = 0
      "00000" when "000000001011000", -- t[88] = 0
      "00000" when "000000001011001", -- t[89] = 0
      "00000" when "000000001011010", -- t[90] = 0
      "00000" when "000000001011011", -- t[91] = 0
      "00000" when "000000001011100", -- t[92] = 0
      "00000" when "000000001011101", -- t[93] = 0
      "00000" when "000000001011110", -- t[94] = 0
      "00000" when "000000001011111", -- t[95] = 0
      "00000" when "000000001100000", -- t[96] = 0
      "00000" when "000000001100001", -- t[97] = 0
      "00000" when "000000001100010", -- t[98] = 0
      "00000" when "000000001100011", -- t[99] = 0
      "00000" when "000000001100100", -- t[100] = 0
      "00000" when "000000001100101", -- t[101] = 0
      "00000" when "000000001100110", -- t[102] = 0
      "00000" when "000000001100111", -- t[103] = 0
      "00000" when "000000001101000", -- t[104] = 0
      "00000" when "000000001101001", -- t[105] = 0
      "00000" when "000000001101010", -- t[106] = 0
      "00000" when "000000001101011", -- t[107] = 0
      "00000" when "000000001101100", -- t[108] = 0
      "00000" when "000000001101101", -- t[109] = 0
      "00000" when "000000001101110", -- t[110] = 0
      "00000" when "000000001101111", -- t[111] = 0
      "00000" when "000000001110000", -- t[112] = 0
      "00000" when "000000001110001", -- t[113] = 0
      "00000" when "000000001110010", -- t[114] = 0
      "00000" when "000000001110011", -- t[115] = 0
      "00000" when "000000001110100", -- t[116] = 0
      "00000" when "000000001110101", -- t[117] = 0
      "00000" when "000000001110110", -- t[118] = 0
      "00000" when "000000001110111", -- t[119] = 0
      "00000" when "000000001111000", -- t[120] = 0
      "00000" when "000000001111001", -- t[121] = 0
      "00000" when "000000001111010", -- t[122] = 0
      "00000" when "000000001111011", -- t[123] = 0
      "00000" when "000000001111100", -- t[124] = 0
      "00000" when "000000001111101", -- t[125] = 0
      "00000" when "000000001111110", -- t[126] = 0
      "00000" when "000000001111111", -- t[127] = 0
      "00000" when "000000010000000", -- t[128] = 0
      "00000" when "000000010000001", -- t[129] = 0
      "00000" when "000000010000010", -- t[130] = 0
      "00000" when "000000010000011", -- t[131] = 0
      "00000" when "000000010000100", -- t[132] = 0
      "00000" when "000000010000101", -- t[133] = 0
      "00000" when "000000010000110", -- t[134] = 0
      "00000" when "000000010000111", -- t[135] = 0
      "00000" when "000000010001000", -- t[136] = 0
      "00000" when "000000010001001", -- t[137] = 0
      "00000" when "000000010001010", -- t[138] = 0
      "00000" when "000000010001011", -- t[139] = 0
      "00000" when "000000010001100", -- t[140] = 0
      "00000" when "000000010001101", -- t[141] = 0
      "00000" when "000000010001110", -- t[142] = 0
      "00000" when "000000010001111", -- t[143] = 0
      "00000" when "000000010010000", -- t[144] = 0
      "00000" when "000000010010001", -- t[145] = 0
      "00000" when "000000010010010", -- t[146] = 0
      "00000" when "000000010010011", -- t[147] = 0
      "00000" when "000000010010100", -- t[148] = 0
      "00000" when "000000010010101", -- t[149] = 0
      "00000" when "000000010010110", -- t[150] = 0
      "00000" when "000000010010111", -- t[151] = 0
      "00000" when "000000010011000", -- t[152] = 0
      "00000" when "000000010011001", -- t[153] = 0
      "00000" when "000000010011010", -- t[154] = 0
      "00000" when "000000010011011", -- t[155] = 0
      "00000" when "000000010011100", -- t[156] = 0
      "00000" when "000000010011101", -- t[157] = 0
      "00000" when "000000010011110", -- t[158] = 0
      "00000" when "000000010011111", -- t[159] = 0
      "00000" when "000000010100000", -- t[160] = 0
      "00000" when "000000010100001", -- t[161] = 0
      "00000" when "000000010100010", -- t[162] = 0
      "00000" when "000000010100011", -- t[163] = 0
      "00000" when "000000010100100", -- t[164] = 0
      "00000" when "000000010100101", -- t[165] = 0
      "00000" when "000000010100110", -- t[166] = 0
      "00000" when "000000010100111", -- t[167] = 0
      "00000" when "000000010101000", -- t[168] = 0
      "00000" when "000000010101001", -- t[169] = 0
      "00000" when "000000010101010", -- t[170] = 0
      "00000" when "000000010101011", -- t[171] = 0
      "00000" when "000000010101100", -- t[172] = 0
      "00000" when "000000010101101", -- t[173] = 0
      "00000" when "000000010101110", -- t[174] = 0
      "00000" when "000000010101111", -- t[175] = 0
      "00000" when "000000010110000", -- t[176] = 0
      "00000" when "000000010110001", -- t[177] = 0
      "00000" when "000000010110010", -- t[178] = 0
      "00000" when "000000010110011", -- t[179] = 0
      "00000" when "000000010110100", -- t[180] = 0
      "00000" when "000000010110101", -- t[181] = 0
      "00000" when "000000010110110", -- t[182] = 0
      "00000" when "000000010110111", -- t[183] = 0
      "00000" when "000000010111000", -- t[184] = 0
      "00000" when "000000010111001", -- t[185] = 0
      "00000" when "000000010111010", -- t[186] = 0
      "00000" when "000000010111011", -- t[187] = 0
      "00000" when "000000010111100", -- t[188] = 0
      "00000" when "000000010111101", -- t[189] = 0
      "00000" when "000000010111110", -- t[190] = 0
      "00000" when "000000010111111", -- t[191] = 0
      "00000" when "000000011000000", -- t[192] = 0
      "00000" when "000000011000001", -- t[193] = 0
      "00000" when "000000011000010", -- t[194] = 0
      "00000" when "000000011000011", -- t[195] = 0
      "00000" when "000000011000100", -- t[196] = 0
      "00000" when "000000011000101", -- t[197] = 0
      "00000" when "000000011000110", -- t[198] = 0
      "00000" when "000000011000111", -- t[199] = 0
      "00000" when "000000011001000", -- t[200] = 0
      "00000" when "000000011001001", -- t[201] = 0
      "00000" when "000000011001010", -- t[202] = 0
      "00000" when "000000011001011", -- t[203] = 0
      "00000" when "000000011001100", -- t[204] = 0
      "00000" when "000000011001101", -- t[205] = 0
      "00000" when "000000011001110", -- t[206] = 0
      "00000" when "000000011001111", -- t[207] = 0
      "00000" when "000000011010000", -- t[208] = 0
      "00000" when "000000011010001", -- t[209] = 0
      "00000" when "000000011010010", -- t[210] = 0
      "00000" when "000000011010011", -- t[211] = 0
      "00000" when "000000011010100", -- t[212] = 0
      "00000" when "000000011010101", -- t[213] = 0
      "00000" when "000000011010110", -- t[214] = 0
      "00000" when "000000011010111", -- t[215] = 0
      "00000" when "000000011011000", -- t[216] = 0
      "00000" when "000000011011001", -- t[217] = 0
      "00000" when "000000011011010", -- t[218] = 0
      "00000" when "000000011011011", -- t[219] = 0
      "00000" when "000000011011100", -- t[220] = 0
      "00000" when "000000011011101", -- t[221] = 0
      "00000" when "000000011011110", -- t[222] = 0
      "00000" when "000000011011111", -- t[223] = 0
      "00000" when "000000011100000", -- t[224] = 0
      "00000" when "000000011100001", -- t[225] = 0
      "00000" when "000000011100010", -- t[226] = 0
      "00000" when "000000011100011", -- t[227] = 0
      "00000" when "000000011100100", -- t[228] = 0
      "00000" when "000000011100101", -- t[229] = 0
      "00000" when "000000011100110", -- t[230] = 0
      "00000" when "000000011100111", -- t[231] = 0
      "00000" when "000000011101000", -- t[232] = 0
      "00000" when "000000011101001", -- t[233] = 0
      "00000" when "000000011101010", -- t[234] = 0
      "00000" when "000000011101011", -- t[235] = 0
      "00000" when "000000011101100", -- t[236] = 0
      "00000" when "000000011101101", -- t[237] = 0
      "00000" when "000000011101110", -- t[238] = 0
      "00000" when "000000011101111", -- t[239] = 0
      "00000" when "000000011110000", -- t[240] = 0
      "00000" when "000000011110001", -- t[241] = 0
      "00000" when "000000011110010", -- t[242] = 0
      "00000" when "000000011110011", -- t[243] = 0
      "00000" when "000000011110100", -- t[244] = 0
      "00000" when "000000011110101", -- t[245] = 0
      "00000" when "000000011110110", -- t[246] = 0
      "00000" when "000000011110111", -- t[247] = 0
      "00000" when "000000011111000", -- t[248] = 0
      "00000" when "000000011111001", -- t[249] = 0
      "00000" when "000000011111010", -- t[250] = 0
      "00000" when "000000011111011", -- t[251] = 0
      "00000" when "000000011111100", -- t[252] = 0
      "00000" when "000000011111101", -- t[253] = 0
      "00000" when "000000011111110", -- t[254] = 0
      "00000" when "000000011111111", -- t[255] = 0
      "00000" when "000000100000000", -- t[256] = 0
      "00000" when "000000100000001", -- t[257] = 0
      "00000" when "000000100000010", -- t[258] = 0
      "00000" when "000000100000011", -- t[259] = 0
      "00000" when "000000100000100", -- t[260] = 0
      "00000" when "000000100000101", -- t[261] = 0
      "00000" when "000000100000110", -- t[262] = 0
      "00000" when "000000100000111", -- t[263] = 0
      "00000" when "000000100001000", -- t[264] = 0
      "00000" when "000000100001001", -- t[265] = 0
      "00000" when "000000100001010", -- t[266] = 0
      "00000" when "000000100001011", -- t[267] = 0
      "00000" when "000000100001100", -- t[268] = 0
      "00000" when "000000100001101", -- t[269] = 0
      "00000" when "000000100001110", -- t[270] = 0
      "00000" when "000000100001111", -- t[271] = 0
      "00000" when "000000100010000", -- t[272] = 0
      "00000" when "000000100010001", -- t[273] = 0
      "00000" when "000000100010010", -- t[274] = 0
      "00000" when "000000100010011", -- t[275] = 0
      "00000" when "000000100010100", -- t[276] = 0
      "00000" when "000000100010101", -- t[277] = 0
      "00000" when "000000100010110", -- t[278] = 0
      "00000" when "000000100010111", -- t[279] = 0
      "00000" when "000000100011000", -- t[280] = 0
      "00000" when "000000100011001", -- t[281] = 0
      "00000" when "000000100011010", -- t[282] = 0
      "00000" when "000000100011011", -- t[283] = 0
      "00000" when "000000100011100", -- t[284] = 0
      "00000" when "000000100011101", -- t[285] = 0
      "00000" when "000000100011110", -- t[286] = 0
      "00000" when "000000100011111", -- t[287] = 0
      "00000" when "000000100100000", -- t[288] = 0
      "00000" when "000000100100001", -- t[289] = 0
      "00000" when "000000100100010", -- t[290] = 0
      "00000" when "000000100100011", -- t[291] = 0
      "00000" when "000000100100100", -- t[292] = 0
      "00000" when "000000100100101", -- t[293] = 0
      "00000" when "000000100100110", -- t[294] = 0
      "00000" when "000000100100111", -- t[295] = 0
      "00000" when "000000100101000", -- t[296] = 0
      "00000" when "000000100101001", -- t[297] = 0
      "00000" when "000000100101010", -- t[298] = 0
      "00000" when "000000100101011", -- t[299] = 0
      "00000" when "000000100101100", -- t[300] = 0
      "00000" when "000000100101101", -- t[301] = 0
      "00000" when "000000100101110", -- t[302] = 0
      "00000" when "000000100101111", -- t[303] = 0
      "00000" when "000000100110000", -- t[304] = 0
      "00000" when "000000100110001", -- t[305] = 0
      "00000" when "000000100110010", -- t[306] = 0
      "00000" when "000000100110011", -- t[307] = 0
      "00000" when "000000100110100", -- t[308] = 0
      "00000" when "000000100110101", -- t[309] = 0
      "00000" when "000000100110110", -- t[310] = 0
      "00000" when "000000100110111", -- t[311] = 0
      "00000" when "000000100111000", -- t[312] = 0
      "00000" when "000000100111001", -- t[313] = 0
      "00000" when "000000100111010", -- t[314] = 0
      "00000" when "000000100111011", -- t[315] = 0
      "00000" when "000000100111100", -- t[316] = 0
      "00000" when "000000100111101", -- t[317] = 0
      "00000" when "000000100111110", -- t[318] = 0
      "00000" when "000000100111111", -- t[319] = 0
      "00000" when "000000101000000", -- t[320] = 0
      "00000" when "000000101000001", -- t[321] = 0
      "00000" when "000000101000010", -- t[322] = 0
      "00000" when "000000101000011", -- t[323] = 0
      "00000" when "000000101000100", -- t[324] = 0
      "00000" when "000000101000101", -- t[325] = 0
      "00000" when "000000101000110", -- t[326] = 0
      "00000" when "000000101000111", -- t[327] = 0
      "00000" when "000000101001000", -- t[328] = 0
      "00000" when "000000101001001", -- t[329] = 0
      "00000" when "000000101001010", -- t[330] = 0
      "00000" when "000000101001011", -- t[331] = 0
      "00000" when "000000101001100", -- t[332] = 0
      "00000" when "000000101001101", -- t[333] = 0
      "00000" when "000000101001110", -- t[334] = 0
      "00000" when "000000101001111", -- t[335] = 0
      "00000" when "000000101010000", -- t[336] = 0
      "00000" when "000000101010001", -- t[337] = 0
      "00000" when "000000101010010", -- t[338] = 0
      "00000" when "000000101010011", -- t[339] = 0
      "00000" when "000000101010100", -- t[340] = 0
      "00000" when "000000101010101", -- t[341] = 0
      "00000" when "000000101010110", -- t[342] = 0
      "00000" when "000000101010111", -- t[343] = 0
      "00000" when "000000101011000", -- t[344] = 0
      "00000" when "000000101011001", -- t[345] = 0
      "00000" when "000000101011010", -- t[346] = 0
      "00000" when "000000101011011", -- t[347] = 0
      "00000" when "000000101011100", -- t[348] = 0
      "00000" when "000000101011101", -- t[349] = 0
      "00000" when "000000101011110", -- t[350] = 0
      "00000" when "000000101011111", -- t[351] = 0
      "00000" when "000000101100000", -- t[352] = 0
      "00000" when "000000101100001", -- t[353] = 0
      "00000" when "000000101100010", -- t[354] = 0
      "00000" when "000000101100011", -- t[355] = 0
      "00000" when "000000101100100", -- t[356] = 0
      "00000" when "000000101100101", -- t[357] = 0
      "00000" when "000000101100110", -- t[358] = 0
      "00000" when "000000101100111", -- t[359] = 0
      "00000" when "000000101101000", -- t[360] = 0
      "00000" when "000000101101001", -- t[361] = 0
      "00000" when "000000101101010", -- t[362] = 0
      "00000" when "000000101101011", -- t[363] = 0
      "00000" when "000000101101100", -- t[364] = 0
      "00000" when "000000101101101", -- t[365] = 0
      "00000" when "000000101101110", -- t[366] = 0
      "00000" when "000000101101111", -- t[367] = 0
      "00000" when "000000101110000", -- t[368] = 0
      "00000" when "000000101110001", -- t[369] = 0
      "00000" when "000000101110010", -- t[370] = 0
      "00000" when "000000101110011", -- t[371] = 0
      "00000" when "000000101110100", -- t[372] = 0
      "00000" when "000000101110101", -- t[373] = 0
      "00000" when "000000101110110", -- t[374] = 0
      "00000" when "000000101110111", -- t[375] = 0
      "00000" when "000000101111000", -- t[376] = 0
      "00000" when "000000101111001", -- t[377] = 0
      "00000" when "000000101111010", -- t[378] = 0
      "00000" when "000000101111011", -- t[379] = 0
      "00000" when "000000101111100", -- t[380] = 0
      "00000" when "000000101111101", -- t[381] = 0
      "00000" when "000000101111110", -- t[382] = 0
      "00000" when "000000101111111", -- t[383] = 0
      "00000" when "000000110000000", -- t[384] = 0
      "00000" when "000000110000001", -- t[385] = 0
      "00000" when "000000110000010", -- t[386] = 0
      "00000" when "000000110000011", -- t[387] = 0
      "00000" when "000000110000100", -- t[388] = 0
      "00000" when "000000110000101", -- t[389] = 0
      "00000" when "000000110000110", -- t[390] = 0
      "00000" when "000000110000111", -- t[391] = 0
      "00000" when "000000110001000", -- t[392] = 0
      "00000" when "000000110001001", -- t[393] = 0
      "00000" when "000000110001010", -- t[394] = 0
      "00000" when "000000110001011", -- t[395] = 0
      "00000" when "000000110001100", -- t[396] = 0
      "00000" when "000000110001101", -- t[397] = 0
      "00000" when "000000110001110", -- t[398] = 0
      "00000" when "000000110001111", -- t[399] = 0
      "00000" when "000000110010000", -- t[400] = 0
      "00000" when "000000110010001", -- t[401] = 0
      "00000" when "000000110010010", -- t[402] = 0
      "00000" when "000000110010011", -- t[403] = 0
      "00000" when "000000110010100", -- t[404] = 0
      "00000" when "000000110010101", -- t[405] = 0
      "00000" when "000000110010110", -- t[406] = 0
      "00000" when "000000110010111", -- t[407] = 0
      "00000" when "000000110011000", -- t[408] = 0
      "00000" when "000000110011001", -- t[409] = 0
      "00000" when "000000110011010", -- t[410] = 0
      "00000" when "000000110011011", -- t[411] = 0
      "00000" when "000000110011100", -- t[412] = 0
      "00000" when "000000110011101", -- t[413] = 0
      "00000" when "000000110011110", -- t[414] = 0
      "00000" when "000000110011111", -- t[415] = 0
      "00000" when "000000110100000", -- t[416] = 0
      "00000" when "000000110100001", -- t[417] = 0
      "00000" when "000000110100010", -- t[418] = 0
      "00000" when "000000110100011", -- t[419] = 0
      "00000" when "000000110100100", -- t[420] = 0
      "00000" when "000000110100101", -- t[421] = 0
      "00000" when "000000110100110", -- t[422] = 0
      "00000" when "000000110100111", -- t[423] = 0
      "00000" when "000000110101000", -- t[424] = 0
      "00000" when "000000110101001", -- t[425] = 0
      "00000" when "000000110101010", -- t[426] = 0
      "00000" when "000000110101011", -- t[427] = 0
      "00000" when "000000110101100", -- t[428] = 0
      "00000" when "000000110101101", -- t[429] = 0
      "00000" when "000000110101110", -- t[430] = 0
      "00000" when "000000110101111", -- t[431] = 0
      "00000" when "000000110110000", -- t[432] = 0
      "00000" when "000000110110001", -- t[433] = 0
      "00000" when "000000110110010", -- t[434] = 0
      "00000" when "000000110110011", -- t[435] = 0
      "00000" when "000000110110100", -- t[436] = 0
      "00000" when "000000110110101", -- t[437] = 0
      "00000" when "000000110110110", -- t[438] = 0
      "00000" when "000000110110111", -- t[439] = 0
      "00000" when "000000110111000", -- t[440] = 0
      "00000" when "000000110111001", -- t[441] = 0
      "00000" when "000000110111010", -- t[442] = 0
      "00000" when "000000110111011", -- t[443] = 0
      "00000" when "000000110111100", -- t[444] = 0
      "00000" when "000000110111101", -- t[445] = 0
      "00000" when "000000110111110", -- t[446] = 0
      "00000" when "000000110111111", -- t[447] = 0
      "00000" when "000000111000000", -- t[448] = 0
      "00000" when "000000111000001", -- t[449] = 0
      "00000" when "000000111000010", -- t[450] = 0
      "00000" when "000000111000011", -- t[451] = 0
      "00000" when "000000111000100", -- t[452] = 0
      "00000" when "000000111000101", -- t[453] = 0
      "00000" when "000000111000110", -- t[454] = 0
      "00000" when "000000111000111", -- t[455] = 0
      "00000" when "000000111001000", -- t[456] = 0
      "00000" when "000000111001001", -- t[457] = 0
      "00000" when "000000111001010", -- t[458] = 0
      "00000" when "000000111001011", -- t[459] = 0
      "00000" when "000000111001100", -- t[460] = 0
      "00000" when "000000111001101", -- t[461] = 0
      "00000" when "000000111001110", -- t[462] = 0
      "00000" when "000000111001111", -- t[463] = 0
      "00000" when "000000111010000", -- t[464] = 0
      "00000" when "000000111010001", -- t[465] = 0
      "00000" when "000000111010010", -- t[466] = 0
      "00000" when "000000111010011", -- t[467] = 0
      "00000" when "000000111010100", -- t[468] = 0
      "00000" when "000000111010101", -- t[469] = 0
      "00000" when "000000111010110", -- t[470] = 0
      "00000" when "000000111010111", -- t[471] = 0
      "00000" when "000000111011000", -- t[472] = 0
      "00000" when "000000111011001", -- t[473] = 0
      "00000" when "000000111011010", -- t[474] = 0
      "00000" when "000000111011011", -- t[475] = 0
      "00000" when "000000111011100", -- t[476] = 0
      "00000" when "000000111011101", -- t[477] = 0
      "00000" when "000000111011110", -- t[478] = 0
      "00000" when "000000111011111", -- t[479] = 0
      "00000" when "000000111100000", -- t[480] = 0
      "00000" when "000000111100001", -- t[481] = 0
      "00000" when "000000111100010", -- t[482] = 0
      "00000" when "000000111100011", -- t[483] = 0
      "00000" when "000000111100100", -- t[484] = 0
      "00000" when "000000111100101", -- t[485] = 0
      "00000" when "000000111100110", -- t[486] = 0
      "00000" when "000000111100111", -- t[487] = 0
      "00000" when "000000111101000", -- t[488] = 0
      "00000" when "000000111101001", -- t[489] = 0
      "00000" when "000000111101010", -- t[490] = 0
      "00000" when "000000111101011", -- t[491] = 0
      "00000" when "000000111101100", -- t[492] = 0
      "00000" when "000000111101101", -- t[493] = 0
      "00000" when "000000111101110", -- t[494] = 0
      "00000" when "000000111101111", -- t[495] = 0
      "00000" when "000000111110000", -- t[496] = 0
      "00000" when "000000111110001", -- t[497] = 0
      "00000" when "000000111110010", -- t[498] = 0
      "00000" when "000000111110011", -- t[499] = 0
      "00000" when "000000111110100", -- t[500] = 0
      "00000" when "000000111110101", -- t[501] = 0
      "00000" when "000000111110110", -- t[502] = 0
      "00000" when "000000111110111", -- t[503] = 0
      "00000" when "000000111111000", -- t[504] = 0
      "00000" when "000000111111001", -- t[505] = 0
      "00000" when "000000111111010", -- t[506] = 0
      "00000" when "000000111111011", -- t[507] = 0
      "00000" when "000000111111100", -- t[508] = 0
      "00000" when "000000111111101", -- t[509] = 0
      "00000" when "000000111111110", -- t[510] = 0
      "00000" when "000000111111111", -- t[511] = 0
      "00000" when "000001000000000", -- t[512] = 0
      "00000" when "000001000000001", -- t[513] = 0
      "00000" when "000001000000010", -- t[514] = 0
      "00000" when "000001000000011", -- t[515] = 0
      "00000" when "000001000000100", -- t[516] = 0
      "00000" when "000001000000101", -- t[517] = 0
      "00000" when "000001000000110", -- t[518] = 0
      "00000" when "000001000000111", -- t[519] = 0
      "00000" when "000001000001000", -- t[520] = 0
      "00000" when "000001000001001", -- t[521] = 0
      "00000" when "000001000001010", -- t[522] = 0
      "00000" when "000001000001011", -- t[523] = 0
      "00000" when "000001000001100", -- t[524] = 0
      "00000" when "000001000001101", -- t[525] = 0
      "00000" when "000001000001110", -- t[526] = 0
      "00000" when "000001000001111", -- t[527] = 0
      "00000" when "000001000010000", -- t[528] = 0
      "00000" when "000001000010001", -- t[529] = 0
      "00000" when "000001000010010", -- t[530] = 0
      "00000" when "000001000010011", -- t[531] = 0
      "00000" when "000001000010100", -- t[532] = 0
      "00000" when "000001000010101", -- t[533] = 0
      "00000" when "000001000010110", -- t[534] = 0
      "00000" when "000001000010111", -- t[535] = 0
      "00000" when "000001000011000", -- t[536] = 0
      "00000" when "000001000011001", -- t[537] = 0
      "00000" when "000001000011010", -- t[538] = 0
      "00000" when "000001000011011", -- t[539] = 0
      "00000" when "000001000011100", -- t[540] = 0
      "00000" when "000001000011101", -- t[541] = 0
      "00000" when "000001000011110", -- t[542] = 0
      "00000" when "000001000011111", -- t[543] = 0
      "00000" when "000001000100000", -- t[544] = 0
      "00000" when "000001000100001", -- t[545] = 0
      "00000" when "000001000100010", -- t[546] = 0
      "00000" when "000001000100011", -- t[547] = 0
      "00000" when "000001000100100", -- t[548] = 0
      "00000" when "000001000100101", -- t[549] = 0
      "00000" when "000001000100110", -- t[550] = 0
      "00000" when "000001000100111", -- t[551] = 0
      "00000" when "000001000101000", -- t[552] = 0
      "00000" when "000001000101001", -- t[553] = 0
      "00000" when "000001000101010", -- t[554] = 0
      "00000" when "000001000101011", -- t[555] = 0
      "00000" when "000001000101100", -- t[556] = 0
      "00000" when "000001000101101", -- t[557] = 0
      "00000" when "000001000101110", -- t[558] = 0
      "00000" when "000001000101111", -- t[559] = 0
      "00000" when "000001000110000", -- t[560] = 0
      "00000" when "000001000110001", -- t[561] = 0
      "00000" when "000001000110010", -- t[562] = 0
      "00000" when "000001000110011", -- t[563] = 0
      "00000" when "000001000110100", -- t[564] = 0
      "00000" when "000001000110101", -- t[565] = 0
      "00000" when "000001000110110", -- t[566] = 0
      "00000" when "000001000110111", -- t[567] = 0
      "00000" when "000001000111000", -- t[568] = 0
      "00000" when "000001000111001", -- t[569] = 0
      "00000" when "000001000111010", -- t[570] = 0
      "00000" when "000001000111011", -- t[571] = 0
      "00000" when "000001000111100", -- t[572] = 0
      "00000" when "000001000111101", -- t[573] = 0
      "00000" when "000001000111110", -- t[574] = 0
      "00000" when "000001000111111", -- t[575] = 0
      "00000" when "000001001000000", -- t[576] = 0
      "00000" when "000001001000001", -- t[577] = 0
      "00000" when "000001001000010", -- t[578] = 0
      "00000" when "000001001000011", -- t[579] = 0
      "00000" when "000001001000100", -- t[580] = 0
      "00000" when "000001001000101", -- t[581] = 0
      "00000" when "000001001000110", -- t[582] = 0
      "00000" when "000001001000111", -- t[583] = 0
      "00000" when "000001001001000", -- t[584] = 0
      "00000" when "000001001001001", -- t[585] = 0
      "00000" when "000001001001010", -- t[586] = 0
      "00000" when "000001001001011", -- t[587] = 0
      "00000" when "000001001001100", -- t[588] = 0
      "00000" when "000001001001101", -- t[589] = 0
      "00000" when "000001001001110", -- t[590] = 0
      "00000" when "000001001001111", -- t[591] = 0
      "00000" when "000001001010000", -- t[592] = 0
      "00000" when "000001001010001", -- t[593] = 0
      "00000" when "000001001010010", -- t[594] = 0
      "00000" when "000001001010011", -- t[595] = 0
      "00000" when "000001001010100", -- t[596] = 0
      "00000" when "000001001010101", -- t[597] = 0
      "00000" when "000001001010110", -- t[598] = 0
      "00000" when "000001001010111", -- t[599] = 0
      "00000" when "000001001011000", -- t[600] = 0
      "00000" when "000001001011001", -- t[601] = 0
      "00000" when "000001001011010", -- t[602] = 0
      "00000" when "000001001011011", -- t[603] = 0
      "00000" when "000001001011100", -- t[604] = 0
      "00000" when "000001001011101", -- t[605] = 0
      "00000" when "000001001011110", -- t[606] = 0
      "00000" when "000001001011111", -- t[607] = 0
      "00000" when "000001001100000", -- t[608] = 0
      "00000" when "000001001100001", -- t[609] = 0
      "00000" when "000001001100010", -- t[610] = 0
      "00000" when "000001001100011", -- t[611] = 0
      "00000" when "000001001100100", -- t[612] = 0
      "00000" when "000001001100101", -- t[613] = 0
      "00000" when "000001001100110", -- t[614] = 0
      "00000" when "000001001100111", -- t[615] = 0
      "00000" when "000001001101000", -- t[616] = 0
      "00000" when "000001001101001", -- t[617] = 0
      "00000" when "000001001101010", -- t[618] = 0
      "00000" when "000001001101011", -- t[619] = 0
      "00000" when "000001001101100", -- t[620] = 0
      "00000" when "000001001101101", -- t[621] = 0
      "00000" when "000001001101110", -- t[622] = 0
      "00000" when "000001001101111", -- t[623] = 0
      "00000" when "000001001110000", -- t[624] = 0
      "00000" when "000001001110001", -- t[625] = 0
      "00000" when "000001001110010", -- t[626] = 0
      "00000" when "000001001110011", -- t[627] = 0
      "00000" when "000001001110100", -- t[628] = 0
      "00000" when "000001001110101", -- t[629] = 0
      "00000" when "000001001110110", -- t[630] = 0
      "00000" when "000001001110111", -- t[631] = 0
      "00000" when "000001001111000", -- t[632] = 0
      "00000" when "000001001111001", -- t[633] = 0
      "00000" when "000001001111010", -- t[634] = 0
      "00000" when "000001001111011", -- t[635] = 0
      "00000" when "000001001111100", -- t[636] = 0
      "00000" when "000001001111101", -- t[637] = 0
      "00000" when "000001001111110", -- t[638] = 0
      "00000" when "000001001111111", -- t[639] = 0
      "00000" when "000001010000000", -- t[640] = 0
      "00000" when "000001010000001", -- t[641] = 0
      "00000" when "000001010000010", -- t[642] = 0
      "00000" when "000001010000011", -- t[643] = 0
      "00000" when "000001010000100", -- t[644] = 0
      "00000" when "000001010000101", -- t[645] = 0
      "00000" when "000001010000110", -- t[646] = 0
      "00000" when "000001010000111", -- t[647] = 0
      "00000" when "000001010001000", -- t[648] = 0
      "00000" when "000001010001001", -- t[649] = 0
      "00000" when "000001010001010", -- t[650] = 0
      "00000" when "000001010001011", -- t[651] = 0
      "00000" when "000001010001100", -- t[652] = 0
      "00000" when "000001010001101", -- t[653] = 0
      "00000" when "000001010001110", -- t[654] = 0
      "00000" when "000001010001111", -- t[655] = 0
      "00000" when "000001010010000", -- t[656] = 0
      "00000" when "000001010010001", -- t[657] = 0
      "00000" when "000001010010010", -- t[658] = 0
      "00000" when "000001010010011", -- t[659] = 0
      "00000" when "000001010010100", -- t[660] = 0
      "00000" when "000001010010101", -- t[661] = 0
      "00000" when "000001010010110", -- t[662] = 0
      "00000" when "000001010010111", -- t[663] = 0
      "00000" when "000001010011000", -- t[664] = 0
      "00000" when "000001010011001", -- t[665] = 0
      "00000" when "000001010011010", -- t[666] = 0
      "00000" when "000001010011011", -- t[667] = 0
      "00000" when "000001010011100", -- t[668] = 0
      "00000" when "000001010011101", -- t[669] = 0
      "00000" when "000001010011110", -- t[670] = 0
      "00000" when "000001010011111", -- t[671] = 0
      "00000" when "000001010100000", -- t[672] = 0
      "00000" when "000001010100001", -- t[673] = 0
      "00000" when "000001010100010", -- t[674] = 0
      "00000" when "000001010100011", -- t[675] = 0
      "00000" when "000001010100100", -- t[676] = 0
      "00000" when "000001010100101", -- t[677] = 0
      "00000" when "000001010100110", -- t[678] = 0
      "00000" when "000001010100111", -- t[679] = 0
      "00000" when "000001010101000", -- t[680] = 0
      "00000" when "000001010101001", -- t[681] = 0
      "00000" when "000001010101010", -- t[682] = 0
      "00000" when "000001010101011", -- t[683] = 0
      "00000" when "000001010101100", -- t[684] = 0
      "00000" when "000001010101101", -- t[685] = 0
      "00000" when "000001010101110", -- t[686] = 0
      "00000" when "000001010101111", -- t[687] = 0
      "00000" when "000001010110000", -- t[688] = 0
      "00000" when "000001010110001", -- t[689] = 0
      "00000" when "000001010110010", -- t[690] = 0
      "00000" when "000001010110011", -- t[691] = 0
      "00000" when "000001010110100", -- t[692] = 0
      "00000" when "000001010110101", -- t[693] = 0
      "00000" when "000001010110110", -- t[694] = 0
      "00000" when "000001010110111", -- t[695] = 0
      "00000" when "000001010111000", -- t[696] = 0
      "00000" when "000001010111001", -- t[697] = 0
      "00000" when "000001010111010", -- t[698] = 0
      "00000" when "000001010111011", -- t[699] = 0
      "00000" when "000001010111100", -- t[700] = 0
      "00000" when "000001010111101", -- t[701] = 0
      "00000" when "000001010111110", -- t[702] = 0
      "00000" when "000001010111111", -- t[703] = 0
      "00000" when "000001011000000", -- t[704] = 0
      "00000" when "000001011000001", -- t[705] = 0
      "00000" when "000001011000010", -- t[706] = 0
      "00000" when "000001011000011", -- t[707] = 0
      "00000" when "000001011000100", -- t[708] = 0
      "00000" when "000001011000101", -- t[709] = 0
      "00000" when "000001011000110", -- t[710] = 0
      "00000" when "000001011000111", -- t[711] = 0
      "00000" when "000001011001000", -- t[712] = 0
      "00000" when "000001011001001", -- t[713] = 0
      "00000" when "000001011001010", -- t[714] = 0
      "00000" when "000001011001011", -- t[715] = 0
      "00000" when "000001011001100", -- t[716] = 0
      "00000" when "000001011001101", -- t[717] = 0
      "00000" when "000001011001110", -- t[718] = 0
      "00000" when "000001011001111", -- t[719] = 0
      "00000" when "000001011010000", -- t[720] = 0
      "00000" when "000001011010001", -- t[721] = 0
      "00000" when "000001011010010", -- t[722] = 0
      "00000" when "000001011010011", -- t[723] = 0
      "00000" when "000001011010100", -- t[724] = 0
      "00000" when "000001011010101", -- t[725] = 0
      "00000" when "000001011010110", -- t[726] = 0
      "00000" when "000001011010111", -- t[727] = 0
      "00000" when "000001011011000", -- t[728] = 0
      "00000" when "000001011011001", -- t[729] = 0
      "00000" when "000001011011010", -- t[730] = 0
      "00000" when "000001011011011", -- t[731] = 0
      "00000" when "000001011011100", -- t[732] = 0
      "00000" when "000001011011101", -- t[733] = 0
      "00000" when "000001011011110", -- t[734] = 0
      "00000" when "000001011011111", -- t[735] = 0
      "00000" when "000001011100000", -- t[736] = 0
      "00000" when "000001011100001", -- t[737] = 0
      "00000" when "000001011100010", -- t[738] = 0
      "00000" when "000001011100011", -- t[739] = 0
      "00000" when "000001011100100", -- t[740] = 0
      "00000" when "000001011100101", -- t[741] = 0
      "00000" when "000001011100110", -- t[742] = 0
      "00000" when "000001011100111", -- t[743] = 0
      "00000" when "000001011101000", -- t[744] = 0
      "00000" when "000001011101001", -- t[745] = 0
      "00000" when "000001011101010", -- t[746] = 0
      "00000" when "000001011101011", -- t[747] = 0
      "00000" when "000001011101100", -- t[748] = 0
      "00000" when "000001011101101", -- t[749] = 0
      "00000" when "000001011101110", -- t[750] = 0
      "00000" when "000001011101111", -- t[751] = 0
      "00000" when "000001011110000", -- t[752] = 0
      "00000" when "000001011110001", -- t[753] = 0
      "00000" when "000001011110010", -- t[754] = 0
      "00000" when "000001011110011", -- t[755] = 0
      "00000" when "000001011110100", -- t[756] = 0
      "00000" when "000001011110101", -- t[757] = 0
      "00000" when "000001011110110", -- t[758] = 0
      "00000" when "000001011110111", -- t[759] = 0
      "00000" when "000001011111000", -- t[760] = 0
      "00000" when "000001011111001", -- t[761] = 0
      "00000" when "000001011111010", -- t[762] = 0
      "00000" when "000001011111011", -- t[763] = 0
      "00000" when "000001011111100", -- t[764] = 0
      "00000" when "000001011111101", -- t[765] = 0
      "00000" when "000001011111110", -- t[766] = 0
      "00000" when "000001011111111", -- t[767] = 0
      "00000" when "000001100000000", -- t[768] = 0
      "00000" when "000001100000001", -- t[769] = 0
      "00000" when "000001100000010", -- t[770] = 0
      "00000" when "000001100000011", -- t[771] = 0
      "00000" when "000001100000100", -- t[772] = 0
      "00000" when "000001100000101", -- t[773] = 0
      "00000" when "000001100000110", -- t[774] = 0
      "00000" when "000001100000111", -- t[775] = 0
      "00000" when "000001100001000", -- t[776] = 0
      "00000" when "000001100001001", -- t[777] = 0
      "00000" when "000001100001010", -- t[778] = 0
      "00000" when "000001100001011", -- t[779] = 0
      "00000" when "000001100001100", -- t[780] = 0
      "00000" when "000001100001101", -- t[781] = 0
      "00000" when "000001100001110", -- t[782] = 0
      "00000" when "000001100001111", -- t[783] = 0
      "00000" when "000001100010000", -- t[784] = 0
      "00000" when "000001100010001", -- t[785] = 0
      "00000" when "000001100010010", -- t[786] = 0
      "00000" when "000001100010011", -- t[787] = 0
      "00000" when "000001100010100", -- t[788] = 0
      "00000" when "000001100010101", -- t[789] = 0
      "00000" when "000001100010110", -- t[790] = 0
      "00000" when "000001100010111", -- t[791] = 0
      "00000" when "000001100011000", -- t[792] = 0
      "00000" when "000001100011001", -- t[793] = 0
      "00000" when "000001100011010", -- t[794] = 0
      "00000" when "000001100011011", -- t[795] = 0
      "00000" when "000001100011100", -- t[796] = 0
      "00000" when "000001100011101", -- t[797] = 0
      "00000" when "000001100011110", -- t[798] = 0
      "00000" when "000001100011111", -- t[799] = 0
      "00000" when "000001100100000", -- t[800] = 0
      "00000" when "000001100100001", -- t[801] = 0
      "00000" when "000001100100010", -- t[802] = 0
      "00000" when "000001100100011", -- t[803] = 0
      "00000" when "000001100100100", -- t[804] = 0
      "00000" when "000001100100101", -- t[805] = 0
      "00000" when "000001100100110", -- t[806] = 0
      "00000" when "000001100100111", -- t[807] = 0
      "00000" when "000001100101000", -- t[808] = 0
      "00000" when "000001100101001", -- t[809] = 0
      "00000" when "000001100101010", -- t[810] = 0
      "00000" when "000001100101011", -- t[811] = 0
      "00000" when "000001100101100", -- t[812] = 0
      "00000" when "000001100101101", -- t[813] = 0
      "00000" when "000001100101110", -- t[814] = 0
      "00000" when "000001100101111", -- t[815] = 0
      "00000" when "000001100110000", -- t[816] = 0
      "00000" when "000001100110001", -- t[817] = 0
      "00000" when "000001100110010", -- t[818] = 0
      "00000" when "000001100110011", -- t[819] = 0
      "00000" when "000001100110100", -- t[820] = 0
      "00000" when "000001100110101", -- t[821] = 0
      "00000" when "000001100110110", -- t[822] = 0
      "00000" when "000001100110111", -- t[823] = 0
      "00000" when "000001100111000", -- t[824] = 0
      "00000" when "000001100111001", -- t[825] = 0
      "00000" when "000001100111010", -- t[826] = 0
      "00000" when "000001100111011", -- t[827] = 0
      "00000" when "000001100111100", -- t[828] = 0
      "00000" when "000001100111101", -- t[829] = 0
      "00000" when "000001100111110", -- t[830] = 0
      "00000" when "000001100111111", -- t[831] = 0
      "00000" when "000001101000000", -- t[832] = 0
      "00000" when "000001101000001", -- t[833] = 0
      "00000" when "000001101000010", -- t[834] = 0
      "00000" when "000001101000011", -- t[835] = 0
      "00000" when "000001101000100", -- t[836] = 0
      "00000" when "000001101000101", -- t[837] = 0
      "00000" when "000001101000110", -- t[838] = 0
      "00000" when "000001101000111", -- t[839] = 0
      "00000" when "000001101001000", -- t[840] = 0
      "00000" when "000001101001001", -- t[841] = 0
      "00000" when "000001101001010", -- t[842] = 0
      "00000" when "000001101001011", -- t[843] = 0
      "00000" when "000001101001100", -- t[844] = 0
      "00000" when "000001101001101", -- t[845] = 0
      "00000" when "000001101001110", -- t[846] = 0
      "00000" when "000001101001111", -- t[847] = 0
      "00000" when "000001101010000", -- t[848] = 0
      "00000" when "000001101010001", -- t[849] = 0
      "00000" when "000001101010010", -- t[850] = 0
      "00000" when "000001101010011", -- t[851] = 0
      "00000" when "000001101010100", -- t[852] = 0
      "00000" when "000001101010101", -- t[853] = 0
      "00000" when "000001101010110", -- t[854] = 0
      "00000" when "000001101010111", -- t[855] = 0
      "00000" when "000001101011000", -- t[856] = 0
      "00000" when "000001101011001", -- t[857] = 0
      "00000" when "000001101011010", -- t[858] = 0
      "00000" when "000001101011011", -- t[859] = 0
      "00000" when "000001101011100", -- t[860] = 0
      "00000" when "000001101011101", -- t[861] = 0
      "00000" when "000001101011110", -- t[862] = 0
      "00000" when "000001101011111", -- t[863] = 0
      "00000" when "000001101100000", -- t[864] = 0
      "00000" when "000001101100001", -- t[865] = 0
      "00000" when "000001101100010", -- t[866] = 0
      "00000" when "000001101100011", -- t[867] = 0
      "00000" when "000001101100100", -- t[868] = 0
      "00000" when "000001101100101", -- t[869] = 0
      "00000" when "000001101100110", -- t[870] = 0
      "00000" when "000001101100111", -- t[871] = 0
      "00000" when "000001101101000", -- t[872] = 0
      "00000" when "000001101101001", -- t[873] = 0
      "00000" when "000001101101010", -- t[874] = 0
      "00000" when "000001101101011", -- t[875] = 0
      "00000" when "000001101101100", -- t[876] = 0
      "00000" when "000001101101101", -- t[877] = 0
      "00000" when "000001101101110", -- t[878] = 0
      "00000" when "000001101101111", -- t[879] = 0
      "00000" when "000001101110000", -- t[880] = 0
      "00000" when "000001101110001", -- t[881] = 0
      "00000" when "000001101110010", -- t[882] = 0
      "00000" when "000001101110011", -- t[883] = 0
      "00000" when "000001101110100", -- t[884] = 0
      "00000" when "000001101110101", -- t[885] = 0
      "00000" when "000001101110110", -- t[886] = 0
      "00000" when "000001101110111", -- t[887] = 0
      "00000" when "000001101111000", -- t[888] = 0
      "00000" when "000001101111001", -- t[889] = 0
      "00000" when "000001101111010", -- t[890] = 0
      "00000" when "000001101111011", -- t[891] = 0
      "00000" when "000001101111100", -- t[892] = 0
      "00000" when "000001101111101", -- t[893] = 0
      "00000" when "000001101111110", -- t[894] = 0
      "00000" when "000001101111111", -- t[895] = 0
      "00000" when "000001110000000", -- t[896] = 0
      "00000" when "000001110000001", -- t[897] = 0
      "00000" when "000001110000010", -- t[898] = 0
      "00000" when "000001110000011", -- t[899] = 0
      "00000" when "000001110000100", -- t[900] = 0
      "00000" when "000001110000101", -- t[901] = 0
      "00000" when "000001110000110", -- t[902] = 0
      "00000" when "000001110000111", -- t[903] = 0
      "00000" when "000001110001000", -- t[904] = 0
      "00000" when "000001110001001", -- t[905] = 0
      "00000" when "000001110001010", -- t[906] = 0
      "00000" when "000001110001011", -- t[907] = 0
      "00000" when "000001110001100", -- t[908] = 0
      "00000" when "000001110001101", -- t[909] = 0
      "00000" when "000001110001110", -- t[910] = 0
      "00000" when "000001110001111", -- t[911] = 0
      "00000" when "000001110010000", -- t[912] = 0
      "00000" when "000001110010001", -- t[913] = 0
      "00000" when "000001110010010", -- t[914] = 0
      "00000" when "000001110010011", -- t[915] = 0
      "00000" when "000001110010100", -- t[916] = 0
      "00000" when "000001110010101", -- t[917] = 0
      "00000" when "000001110010110", -- t[918] = 0
      "00000" when "000001110010111", -- t[919] = 0
      "00000" when "000001110011000", -- t[920] = 0
      "00000" when "000001110011001", -- t[921] = 0
      "00000" when "000001110011010", -- t[922] = 0
      "00000" when "000001110011011", -- t[923] = 0
      "00000" when "000001110011100", -- t[924] = 0
      "00000" when "000001110011101", -- t[925] = 0
      "00000" when "000001110011110", -- t[926] = 0
      "00000" when "000001110011111", -- t[927] = 0
      "00000" when "000001110100000", -- t[928] = 0
      "00000" when "000001110100001", -- t[929] = 0
      "00000" when "000001110100010", -- t[930] = 0
      "00000" when "000001110100011", -- t[931] = 0
      "00000" when "000001110100100", -- t[932] = 0
      "00000" when "000001110100101", -- t[933] = 0
      "00000" when "000001110100110", -- t[934] = 0
      "00000" when "000001110100111", -- t[935] = 0
      "00000" when "000001110101000", -- t[936] = 0
      "00000" when "000001110101001", -- t[937] = 0
      "00000" when "000001110101010", -- t[938] = 0
      "00000" when "000001110101011", -- t[939] = 0
      "00000" when "000001110101100", -- t[940] = 0
      "00000" when "000001110101101", -- t[941] = 0
      "00000" when "000001110101110", -- t[942] = 0
      "00000" when "000001110101111", -- t[943] = 0
      "00000" when "000001110110000", -- t[944] = 0
      "00000" when "000001110110001", -- t[945] = 0
      "00000" when "000001110110010", -- t[946] = 0
      "00000" when "000001110110011", -- t[947] = 0
      "00000" when "000001110110100", -- t[948] = 0
      "00000" when "000001110110101", -- t[949] = 0
      "00000" when "000001110110110", -- t[950] = 0
      "00000" when "000001110110111", -- t[951] = 0
      "00000" when "000001110111000", -- t[952] = 0
      "00000" when "000001110111001", -- t[953] = 0
      "00000" when "000001110111010", -- t[954] = 0
      "00000" when "000001110111011", -- t[955] = 0
      "00000" when "000001110111100", -- t[956] = 0
      "00000" when "000001110111101", -- t[957] = 0
      "00000" when "000001110111110", -- t[958] = 0
      "00000" when "000001110111111", -- t[959] = 0
      "00000" when "000001111000000", -- t[960] = 0
      "00000" when "000001111000001", -- t[961] = 0
      "00000" when "000001111000010", -- t[962] = 0
      "00000" when "000001111000011", -- t[963] = 0
      "00000" when "000001111000100", -- t[964] = 0
      "00000" when "000001111000101", -- t[965] = 0
      "00000" when "000001111000110", -- t[966] = 0
      "00000" when "000001111000111", -- t[967] = 0
      "00000" when "000001111001000", -- t[968] = 0
      "00000" when "000001111001001", -- t[969] = 0
      "00000" when "000001111001010", -- t[970] = 0
      "00000" when "000001111001011", -- t[971] = 0
      "00000" when "000001111001100", -- t[972] = 0
      "00000" when "000001111001101", -- t[973] = 0
      "00000" when "000001111001110", -- t[974] = 0
      "00000" when "000001111001111", -- t[975] = 0
      "00000" when "000001111010000", -- t[976] = 0
      "00000" when "000001111010001", -- t[977] = 0
      "00000" when "000001111010010", -- t[978] = 0
      "00000" when "000001111010011", -- t[979] = 0
      "00000" when "000001111010100", -- t[980] = 0
      "00000" when "000001111010101", -- t[981] = 0
      "00000" when "000001111010110", -- t[982] = 0
      "00000" when "000001111010111", -- t[983] = 0
      "00000" when "000001111011000", -- t[984] = 0
      "00000" when "000001111011001", -- t[985] = 0
      "00000" when "000001111011010", -- t[986] = 0
      "00000" when "000001111011011", -- t[987] = 0
      "00000" when "000001111011100", -- t[988] = 0
      "00000" when "000001111011101", -- t[989] = 0
      "00000" when "000001111011110", -- t[990] = 0
      "00000" when "000001111011111", -- t[991] = 0
      "00000" when "000001111100000", -- t[992] = 0
      "00000" when "000001111100001", -- t[993] = 0
      "00000" when "000001111100010", -- t[994] = 0
      "00000" when "000001111100011", -- t[995] = 0
      "00000" when "000001111100100", -- t[996] = 0
      "00000" when "000001111100101", -- t[997] = 0
      "00000" when "000001111100110", -- t[998] = 0
      "00000" when "000001111100111", -- t[999] = 0
      "00000" when "000001111101000", -- t[1000] = 0
      "00000" when "000001111101001", -- t[1001] = 0
      "00000" when "000001111101010", -- t[1002] = 0
      "00000" when "000001111101011", -- t[1003] = 0
      "00000" when "000001111101100", -- t[1004] = 0
      "00000" when "000001111101101", -- t[1005] = 0
      "00000" when "000001111101110", -- t[1006] = 0
      "00000" when "000001111101111", -- t[1007] = 0
      "00000" when "000001111110000", -- t[1008] = 0
      "00000" when "000001111110001", -- t[1009] = 0
      "00000" when "000001111110010", -- t[1010] = 0
      "00000" when "000001111110011", -- t[1011] = 0
      "00000" when "000001111110100", -- t[1012] = 0
      "00000" when "000001111110101", -- t[1013] = 0
      "00000" when "000001111110110", -- t[1014] = 0
      "00000" when "000001111110111", -- t[1015] = 0
      "00000" when "000001111111000", -- t[1016] = 0
      "00000" when "000001111111001", -- t[1017] = 0
      "00000" when "000001111111010", -- t[1018] = 0
      "00000" when "000001111111011", -- t[1019] = 0
      "00000" when "000001111111100", -- t[1020] = 0
      "00000" when "000001111111101", -- t[1021] = 0
      "00000" when "000001111111110", -- t[1022] = 0
      "00000" when "000001111111111", -- t[1023] = 0
      "00000" when "000010000000000", -- t[1024] = 0
      "00000" when "000010000000001", -- t[1025] = 0
      "00000" when "000010000000010", -- t[1026] = 0
      "00000" when "000010000000011", -- t[1027] = 0
      "00000" when "000010000000100", -- t[1028] = 0
      "00000" when "000010000000101", -- t[1029] = 0
      "00000" when "000010000000110", -- t[1030] = 0
      "00000" when "000010000000111", -- t[1031] = 0
      "00000" when "000010000001000", -- t[1032] = 0
      "00000" when "000010000001001", -- t[1033] = 0
      "00000" when "000010000001010", -- t[1034] = 0
      "00000" when "000010000001011", -- t[1035] = 0
      "00000" when "000010000001100", -- t[1036] = 0
      "00000" when "000010000001101", -- t[1037] = 0
      "00000" when "000010000001110", -- t[1038] = 0
      "00000" when "000010000001111", -- t[1039] = 0
      "00000" when "000010000010000", -- t[1040] = 0
      "00000" when "000010000010001", -- t[1041] = 0
      "00000" when "000010000010010", -- t[1042] = 0
      "00000" when "000010000010011", -- t[1043] = 0
      "00000" when "000010000010100", -- t[1044] = 0
      "00000" when "000010000010101", -- t[1045] = 0
      "00000" when "000010000010110", -- t[1046] = 0
      "00000" when "000010000010111", -- t[1047] = 0
      "00000" when "000010000011000", -- t[1048] = 0
      "00000" when "000010000011001", -- t[1049] = 0
      "00000" when "000010000011010", -- t[1050] = 0
      "00000" when "000010000011011", -- t[1051] = 0
      "00000" when "000010000011100", -- t[1052] = 0
      "00000" when "000010000011101", -- t[1053] = 0
      "00000" when "000010000011110", -- t[1054] = 0
      "00000" when "000010000011111", -- t[1055] = 0
      "00000" when "000010000100000", -- t[1056] = 0
      "00000" when "000010000100001", -- t[1057] = 0
      "00000" when "000010000100010", -- t[1058] = 0
      "00000" when "000010000100011", -- t[1059] = 0
      "00000" when "000010000100100", -- t[1060] = 0
      "00000" when "000010000100101", -- t[1061] = 0
      "00000" when "000010000100110", -- t[1062] = 0
      "00000" when "000010000100111", -- t[1063] = 0
      "00000" when "000010000101000", -- t[1064] = 0
      "00000" when "000010000101001", -- t[1065] = 0
      "00000" when "000010000101010", -- t[1066] = 0
      "00000" when "000010000101011", -- t[1067] = 0
      "00000" when "000010000101100", -- t[1068] = 0
      "00000" when "000010000101101", -- t[1069] = 0
      "00000" when "000010000101110", -- t[1070] = 0
      "00000" when "000010000101111", -- t[1071] = 0
      "00000" when "000010000110000", -- t[1072] = 0
      "00000" when "000010000110001", -- t[1073] = 0
      "00000" when "000010000110010", -- t[1074] = 0
      "00000" when "000010000110011", -- t[1075] = 0
      "00000" when "000010000110100", -- t[1076] = 0
      "00000" when "000010000110101", -- t[1077] = 0
      "00000" when "000010000110110", -- t[1078] = 0
      "00000" when "000010000110111", -- t[1079] = 0
      "00000" when "000010000111000", -- t[1080] = 0
      "00000" when "000010000111001", -- t[1081] = 0
      "00000" when "000010000111010", -- t[1082] = 0
      "00000" when "000010000111011", -- t[1083] = 0
      "00000" when "000010000111100", -- t[1084] = 0
      "00000" when "000010000111101", -- t[1085] = 0
      "00000" when "000010000111110", -- t[1086] = 0
      "00000" when "000010000111111", -- t[1087] = 0
      "00000" when "000010001000000", -- t[1088] = 0
      "00000" when "000010001000001", -- t[1089] = 0
      "00000" when "000010001000010", -- t[1090] = 0
      "00000" when "000010001000011", -- t[1091] = 0
      "00000" when "000010001000100", -- t[1092] = 0
      "00000" when "000010001000101", -- t[1093] = 0
      "00000" when "000010001000110", -- t[1094] = 0
      "00000" when "000010001000111", -- t[1095] = 0
      "00000" when "000010001001000", -- t[1096] = 0
      "00000" when "000010001001001", -- t[1097] = 0
      "00000" when "000010001001010", -- t[1098] = 0
      "00000" when "000010001001011", -- t[1099] = 0
      "00000" when "000010001001100", -- t[1100] = 0
      "00000" when "000010001001101", -- t[1101] = 0
      "00000" when "000010001001110", -- t[1102] = 0
      "00000" when "000010001001111", -- t[1103] = 0
      "00000" when "000010001010000", -- t[1104] = 0
      "00000" when "000010001010001", -- t[1105] = 0
      "00000" when "000010001010010", -- t[1106] = 0
      "00000" when "000010001010011", -- t[1107] = 0
      "00000" when "000010001010100", -- t[1108] = 0
      "00000" when "000010001010101", -- t[1109] = 0
      "00000" when "000010001010110", -- t[1110] = 0
      "00000" when "000010001010111", -- t[1111] = 0
      "00000" when "000010001011000", -- t[1112] = 0
      "00000" when "000010001011001", -- t[1113] = 0
      "00000" when "000010001011010", -- t[1114] = 0
      "00000" when "000010001011011", -- t[1115] = 0
      "00000" when "000010001011100", -- t[1116] = 0
      "00000" when "000010001011101", -- t[1117] = 0
      "00000" when "000010001011110", -- t[1118] = 0
      "00000" when "000010001011111", -- t[1119] = 0
      "00000" when "000010001100000", -- t[1120] = 0
      "00000" when "000010001100001", -- t[1121] = 0
      "00000" when "000010001100010", -- t[1122] = 0
      "00000" when "000010001100011", -- t[1123] = 0
      "00000" when "000010001100100", -- t[1124] = 0
      "00000" when "000010001100101", -- t[1125] = 0
      "00000" when "000010001100110", -- t[1126] = 0
      "00000" when "000010001100111", -- t[1127] = 0
      "00000" when "000010001101000", -- t[1128] = 0
      "00000" when "000010001101001", -- t[1129] = 0
      "00000" when "000010001101010", -- t[1130] = 0
      "00000" when "000010001101011", -- t[1131] = 0
      "00000" when "000010001101100", -- t[1132] = 0
      "00000" when "000010001101101", -- t[1133] = 0
      "00000" when "000010001101110", -- t[1134] = 0
      "00000" when "000010001101111", -- t[1135] = 0
      "00000" when "000010001110000", -- t[1136] = 0
      "00000" when "000010001110001", -- t[1137] = 0
      "00000" when "000010001110010", -- t[1138] = 0
      "00000" when "000010001110011", -- t[1139] = 0
      "00000" when "000010001110100", -- t[1140] = 0
      "00000" when "000010001110101", -- t[1141] = 0
      "00000" when "000010001110110", -- t[1142] = 0
      "00000" when "000010001110111", -- t[1143] = 0
      "00000" when "000010001111000", -- t[1144] = 0
      "00000" when "000010001111001", -- t[1145] = 0
      "00000" when "000010001111010", -- t[1146] = 0
      "00000" when "000010001111011", -- t[1147] = 0
      "00000" when "000010001111100", -- t[1148] = 0
      "00000" when "000010001111101", -- t[1149] = 0
      "00000" when "000010001111110", -- t[1150] = 0
      "00000" when "000010001111111", -- t[1151] = 0
      "00000" when "000010010000000", -- t[1152] = 0
      "00000" when "000010010000001", -- t[1153] = 0
      "00000" when "000010010000010", -- t[1154] = 0
      "00000" when "000010010000011", -- t[1155] = 0
      "00000" when "000010010000100", -- t[1156] = 0
      "00000" when "000010010000101", -- t[1157] = 0
      "00000" when "000010010000110", -- t[1158] = 0
      "00000" when "000010010000111", -- t[1159] = 0
      "00000" when "000010010001000", -- t[1160] = 0
      "00000" when "000010010001001", -- t[1161] = 0
      "00000" when "000010010001010", -- t[1162] = 0
      "00000" when "000010010001011", -- t[1163] = 0
      "00000" when "000010010001100", -- t[1164] = 0
      "00000" when "000010010001101", -- t[1165] = 0
      "00000" when "000010010001110", -- t[1166] = 0
      "00000" when "000010010001111", -- t[1167] = 0
      "00000" when "000010010010000", -- t[1168] = 0
      "00000" when "000010010010001", -- t[1169] = 0
      "00000" when "000010010010010", -- t[1170] = 0
      "00000" when "000010010010011", -- t[1171] = 0
      "00000" when "000010010010100", -- t[1172] = 0
      "00000" when "000010010010101", -- t[1173] = 0
      "00000" when "000010010010110", -- t[1174] = 0
      "00000" when "000010010010111", -- t[1175] = 0
      "00000" when "000010010011000", -- t[1176] = 0
      "00000" when "000010010011001", -- t[1177] = 0
      "00000" when "000010010011010", -- t[1178] = 0
      "00000" when "000010010011011", -- t[1179] = 0
      "00000" when "000010010011100", -- t[1180] = 0
      "00000" when "000010010011101", -- t[1181] = 0
      "00000" when "000010010011110", -- t[1182] = 0
      "00000" when "000010010011111", -- t[1183] = 0
      "00000" when "000010010100000", -- t[1184] = 0
      "00000" when "000010010100001", -- t[1185] = 0
      "00000" when "000010010100010", -- t[1186] = 0
      "00000" when "000010010100011", -- t[1187] = 0
      "00000" when "000010010100100", -- t[1188] = 0
      "00000" when "000010010100101", -- t[1189] = 0
      "00000" when "000010010100110", -- t[1190] = 0
      "00000" when "000010010100111", -- t[1191] = 0
      "00000" when "000010010101000", -- t[1192] = 0
      "00000" when "000010010101001", -- t[1193] = 0
      "00000" when "000010010101010", -- t[1194] = 0
      "00000" when "000010010101011", -- t[1195] = 0
      "00000" when "000010010101100", -- t[1196] = 0
      "00000" when "000010010101101", -- t[1197] = 0
      "00000" when "000010010101110", -- t[1198] = 0
      "00000" when "000010010101111", -- t[1199] = 0
      "00000" when "000010010110000", -- t[1200] = 0
      "00000" when "000010010110001", -- t[1201] = 0
      "00000" when "000010010110010", -- t[1202] = 0
      "00000" when "000010010110011", -- t[1203] = 0
      "00000" when "000010010110100", -- t[1204] = 0
      "00000" when "000010010110101", -- t[1205] = 0
      "00000" when "000010010110110", -- t[1206] = 0
      "00000" when "000010010110111", -- t[1207] = 0
      "00000" when "000010010111000", -- t[1208] = 0
      "00000" when "000010010111001", -- t[1209] = 0
      "00000" when "000010010111010", -- t[1210] = 0
      "00000" when "000010010111011", -- t[1211] = 0
      "00000" when "000010010111100", -- t[1212] = 0
      "00000" when "000010010111101", -- t[1213] = 0
      "00000" when "000010010111110", -- t[1214] = 0
      "00000" when "000010010111111", -- t[1215] = 0
      "00000" when "000010011000000", -- t[1216] = 0
      "00000" when "000010011000001", -- t[1217] = 0
      "00000" when "000010011000010", -- t[1218] = 0
      "00000" when "000010011000011", -- t[1219] = 0
      "00000" when "000010011000100", -- t[1220] = 0
      "00000" when "000010011000101", -- t[1221] = 0
      "00000" when "000010011000110", -- t[1222] = 0
      "00000" when "000010011000111", -- t[1223] = 0
      "00000" when "000010011001000", -- t[1224] = 0
      "00000" when "000010011001001", -- t[1225] = 0
      "00000" when "000010011001010", -- t[1226] = 0
      "00000" when "000010011001011", -- t[1227] = 0
      "00000" when "000010011001100", -- t[1228] = 0
      "00000" when "000010011001101", -- t[1229] = 0
      "00000" when "000010011001110", -- t[1230] = 0
      "00000" when "000010011001111", -- t[1231] = 0
      "00000" when "000010011010000", -- t[1232] = 0
      "00000" when "000010011010001", -- t[1233] = 0
      "00000" when "000010011010010", -- t[1234] = 0
      "00000" when "000010011010011", -- t[1235] = 0
      "00000" when "000010011010100", -- t[1236] = 0
      "00000" when "000010011010101", -- t[1237] = 0
      "00000" when "000010011010110", -- t[1238] = 0
      "00000" when "000010011010111", -- t[1239] = 0
      "00000" when "000010011011000", -- t[1240] = 0
      "00000" when "000010011011001", -- t[1241] = 0
      "00000" when "000010011011010", -- t[1242] = 0
      "00000" when "000010011011011", -- t[1243] = 0
      "00000" when "000010011011100", -- t[1244] = 0
      "00000" when "000010011011101", -- t[1245] = 0
      "00000" when "000010011011110", -- t[1246] = 0
      "00000" when "000010011011111", -- t[1247] = 0
      "00000" when "000010011100000", -- t[1248] = 0
      "00000" when "000010011100001", -- t[1249] = 0
      "00000" when "000010011100010", -- t[1250] = 0
      "00000" when "000010011100011", -- t[1251] = 0
      "00000" when "000010011100100", -- t[1252] = 0
      "00000" when "000010011100101", -- t[1253] = 0
      "00000" when "000010011100110", -- t[1254] = 0
      "00000" when "000010011100111", -- t[1255] = 0
      "00000" when "000010011101000", -- t[1256] = 0
      "00000" when "000010011101001", -- t[1257] = 0
      "00000" when "000010011101010", -- t[1258] = 0
      "00000" when "000010011101011", -- t[1259] = 0
      "00000" when "000010011101100", -- t[1260] = 0
      "00000" when "000010011101101", -- t[1261] = 0
      "00000" when "000010011101110", -- t[1262] = 0
      "00000" when "000010011101111", -- t[1263] = 0
      "00000" when "000010011110000", -- t[1264] = 0
      "00000" when "000010011110001", -- t[1265] = 0
      "00000" when "000010011110010", -- t[1266] = 0
      "00000" when "000010011110011", -- t[1267] = 0
      "00000" when "000010011110100", -- t[1268] = 0
      "00000" when "000010011110101", -- t[1269] = 0
      "00000" when "000010011110110", -- t[1270] = 0
      "00000" when "000010011110111", -- t[1271] = 0
      "00000" when "000010011111000", -- t[1272] = 0
      "00000" when "000010011111001", -- t[1273] = 0
      "00000" when "000010011111010", -- t[1274] = 0
      "00000" when "000010011111011", -- t[1275] = 0
      "00000" when "000010011111100", -- t[1276] = 0
      "00000" when "000010011111101", -- t[1277] = 0
      "00000" when "000010011111110", -- t[1278] = 0
      "00000" when "000010011111111", -- t[1279] = 0
      "00000" when "000010100000000", -- t[1280] = 0
      "00000" when "000010100000001", -- t[1281] = 0
      "00000" when "000010100000010", -- t[1282] = 0
      "00000" when "000010100000011", -- t[1283] = 0
      "00000" when "000010100000100", -- t[1284] = 0
      "00000" when "000010100000101", -- t[1285] = 0
      "00000" when "000010100000110", -- t[1286] = 0
      "00000" when "000010100000111", -- t[1287] = 0
      "00000" when "000010100001000", -- t[1288] = 0
      "00000" when "000010100001001", -- t[1289] = 0
      "00000" when "000010100001010", -- t[1290] = 0
      "00000" when "000010100001011", -- t[1291] = 0
      "00000" when "000010100001100", -- t[1292] = 0
      "00000" when "000010100001101", -- t[1293] = 0
      "00000" when "000010100001110", -- t[1294] = 0
      "00000" when "000010100001111", -- t[1295] = 0
      "00000" when "000010100010000", -- t[1296] = 0
      "00000" when "000010100010001", -- t[1297] = 0
      "00000" when "000010100010010", -- t[1298] = 0
      "00000" when "000010100010011", -- t[1299] = 0
      "00000" when "000010100010100", -- t[1300] = 0
      "00000" when "000010100010101", -- t[1301] = 0
      "00000" when "000010100010110", -- t[1302] = 0
      "00000" when "000010100010111", -- t[1303] = 0
      "00000" when "000010100011000", -- t[1304] = 0
      "00000" when "000010100011001", -- t[1305] = 0
      "00000" when "000010100011010", -- t[1306] = 0
      "00000" when "000010100011011", -- t[1307] = 0
      "00000" when "000010100011100", -- t[1308] = 0
      "00000" when "000010100011101", -- t[1309] = 0
      "00000" when "000010100011110", -- t[1310] = 0
      "00000" when "000010100011111", -- t[1311] = 0
      "00000" when "000010100100000", -- t[1312] = 0
      "00000" when "000010100100001", -- t[1313] = 0
      "00000" when "000010100100010", -- t[1314] = 0
      "00000" when "000010100100011", -- t[1315] = 0
      "00000" when "000010100100100", -- t[1316] = 0
      "00000" when "000010100100101", -- t[1317] = 0
      "00000" when "000010100100110", -- t[1318] = 0
      "00000" when "000010100100111", -- t[1319] = 0
      "00000" when "000010100101000", -- t[1320] = 0
      "00000" when "000010100101001", -- t[1321] = 0
      "00000" when "000010100101010", -- t[1322] = 0
      "00000" when "000010100101011", -- t[1323] = 0
      "00000" when "000010100101100", -- t[1324] = 0
      "00000" when "000010100101101", -- t[1325] = 0
      "00000" when "000010100101110", -- t[1326] = 0
      "00000" when "000010100101111", -- t[1327] = 0
      "00000" when "000010100110000", -- t[1328] = 0
      "00000" when "000010100110001", -- t[1329] = 0
      "00000" when "000010100110010", -- t[1330] = 0
      "00000" when "000010100110011", -- t[1331] = 0
      "00000" when "000010100110100", -- t[1332] = 0
      "00000" when "000010100110101", -- t[1333] = 0
      "00000" when "000010100110110", -- t[1334] = 0
      "00000" when "000010100110111", -- t[1335] = 0
      "00000" when "000010100111000", -- t[1336] = 0
      "00000" when "000010100111001", -- t[1337] = 0
      "00000" when "000010100111010", -- t[1338] = 0
      "00000" when "000010100111011", -- t[1339] = 0
      "00000" when "000010100111100", -- t[1340] = 0
      "00000" when "000010100111101", -- t[1341] = 0
      "00000" when "000010100111110", -- t[1342] = 0
      "00000" when "000010100111111", -- t[1343] = 0
      "00000" when "000010101000000", -- t[1344] = 0
      "00000" when "000010101000001", -- t[1345] = 0
      "00000" when "000010101000010", -- t[1346] = 0
      "00000" when "000010101000011", -- t[1347] = 0
      "00000" when "000010101000100", -- t[1348] = 0
      "00000" when "000010101000101", -- t[1349] = 0
      "00000" when "000010101000110", -- t[1350] = 0
      "00000" when "000010101000111", -- t[1351] = 0
      "00000" when "000010101001000", -- t[1352] = 0
      "00000" when "000010101001001", -- t[1353] = 0
      "00000" when "000010101001010", -- t[1354] = 0
      "00000" when "000010101001011", -- t[1355] = 0
      "00000" when "000010101001100", -- t[1356] = 0
      "00000" when "000010101001101", -- t[1357] = 0
      "00000" when "000010101001110", -- t[1358] = 0
      "00000" when "000010101001111", -- t[1359] = 0
      "00000" when "000010101010000", -- t[1360] = 0
      "00000" when "000010101010001", -- t[1361] = 0
      "00000" when "000010101010010", -- t[1362] = 0
      "00000" when "000010101010011", -- t[1363] = 0
      "00000" when "000010101010100", -- t[1364] = 0
      "00000" when "000010101010101", -- t[1365] = 0
      "00000" when "000010101010110", -- t[1366] = 0
      "00000" when "000010101010111", -- t[1367] = 0
      "00000" when "000010101011000", -- t[1368] = 0
      "00000" when "000010101011001", -- t[1369] = 0
      "00000" when "000010101011010", -- t[1370] = 0
      "00000" when "000010101011011", -- t[1371] = 0
      "00000" when "000010101011100", -- t[1372] = 0
      "00000" when "000010101011101", -- t[1373] = 0
      "00000" when "000010101011110", -- t[1374] = 0
      "00000" when "000010101011111", -- t[1375] = 0
      "00000" when "000010101100000", -- t[1376] = 0
      "00000" when "000010101100001", -- t[1377] = 0
      "00000" when "000010101100010", -- t[1378] = 0
      "00000" when "000010101100011", -- t[1379] = 0
      "00000" when "000010101100100", -- t[1380] = 0
      "00000" when "000010101100101", -- t[1381] = 0
      "00000" when "000010101100110", -- t[1382] = 0
      "00000" when "000010101100111", -- t[1383] = 0
      "00000" when "000010101101000", -- t[1384] = 0
      "00000" when "000010101101001", -- t[1385] = 0
      "00000" when "000010101101010", -- t[1386] = 0
      "00000" when "000010101101011", -- t[1387] = 0
      "00000" when "000010101101100", -- t[1388] = 0
      "00000" when "000010101101101", -- t[1389] = 0
      "00000" when "000010101101110", -- t[1390] = 0
      "00000" when "000010101101111", -- t[1391] = 0
      "00000" when "000010101110000", -- t[1392] = 0
      "00000" when "000010101110001", -- t[1393] = 0
      "00000" when "000010101110010", -- t[1394] = 0
      "00000" when "000010101110011", -- t[1395] = 0
      "00000" when "000010101110100", -- t[1396] = 0
      "00000" when "000010101110101", -- t[1397] = 0
      "00000" when "000010101110110", -- t[1398] = 0
      "00000" when "000010101110111", -- t[1399] = 0
      "00000" when "000010101111000", -- t[1400] = 0
      "00000" when "000010101111001", -- t[1401] = 0
      "00000" when "000010101111010", -- t[1402] = 0
      "00000" when "000010101111011", -- t[1403] = 0
      "00000" when "000010101111100", -- t[1404] = 0
      "00000" when "000010101111101", -- t[1405] = 0
      "00000" when "000010101111110", -- t[1406] = 0
      "00000" when "000010101111111", -- t[1407] = 0
      "00000" when "000010110000000", -- t[1408] = 0
      "00000" when "000010110000001", -- t[1409] = 0
      "00000" when "000010110000010", -- t[1410] = 0
      "00000" when "000010110000011", -- t[1411] = 0
      "00000" when "000010110000100", -- t[1412] = 0
      "00000" when "000010110000101", -- t[1413] = 0
      "00000" when "000010110000110", -- t[1414] = 0
      "00000" when "000010110000111", -- t[1415] = 0
      "00000" when "000010110001000", -- t[1416] = 0
      "00000" when "000010110001001", -- t[1417] = 0
      "00000" when "000010110001010", -- t[1418] = 0
      "00000" when "000010110001011", -- t[1419] = 0
      "00000" when "000010110001100", -- t[1420] = 0
      "00000" when "000010110001101", -- t[1421] = 0
      "00000" when "000010110001110", -- t[1422] = 0
      "00000" when "000010110001111", -- t[1423] = 0
      "00000" when "000010110010000", -- t[1424] = 0
      "00000" when "000010110010001", -- t[1425] = 0
      "00000" when "000010110010010", -- t[1426] = 0
      "00000" when "000010110010011", -- t[1427] = 0
      "00000" when "000010110010100", -- t[1428] = 0
      "00000" when "000010110010101", -- t[1429] = 0
      "00000" when "000010110010110", -- t[1430] = 0
      "00000" when "000010110010111", -- t[1431] = 0
      "00000" when "000010110011000", -- t[1432] = 0
      "00000" when "000010110011001", -- t[1433] = 0
      "00000" when "000010110011010", -- t[1434] = 0
      "00000" when "000010110011011", -- t[1435] = 0
      "00000" when "000010110011100", -- t[1436] = 0
      "00000" when "000010110011101", -- t[1437] = 0
      "00000" when "000010110011110", -- t[1438] = 0
      "00000" when "000010110011111", -- t[1439] = 0
      "00000" when "000010110100000", -- t[1440] = 0
      "00000" when "000010110100001", -- t[1441] = 0
      "00000" when "000010110100010", -- t[1442] = 0
      "00000" when "000010110100011", -- t[1443] = 0
      "00000" when "000010110100100", -- t[1444] = 0
      "00000" when "000010110100101", -- t[1445] = 0
      "00000" when "000010110100110", -- t[1446] = 0
      "00000" when "000010110100111", -- t[1447] = 0
      "00000" when "000010110101000", -- t[1448] = 0
      "00000" when "000010110101001", -- t[1449] = 0
      "00000" when "000010110101010", -- t[1450] = 0
      "00000" when "000010110101011", -- t[1451] = 0
      "00000" when "000010110101100", -- t[1452] = 0
      "00000" when "000010110101101", -- t[1453] = 0
      "00000" when "000010110101110", -- t[1454] = 0
      "00000" when "000010110101111", -- t[1455] = 0
      "00000" when "000010110110000", -- t[1456] = 0
      "00000" when "000010110110001", -- t[1457] = 0
      "00000" when "000010110110010", -- t[1458] = 0
      "00000" when "000010110110011", -- t[1459] = 0
      "00000" when "000010110110100", -- t[1460] = 0
      "00000" when "000010110110101", -- t[1461] = 0
      "00000" when "000010110110110", -- t[1462] = 0
      "00000" when "000010110110111", -- t[1463] = 0
      "00000" when "000010110111000", -- t[1464] = 0
      "00000" when "000010110111001", -- t[1465] = 0
      "00000" when "000010110111010", -- t[1466] = 0
      "00000" when "000010110111011", -- t[1467] = 0
      "00000" when "000010110111100", -- t[1468] = 0
      "00000" when "000010110111101", -- t[1469] = 0
      "00000" when "000010110111110", -- t[1470] = 0
      "00000" when "000010110111111", -- t[1471] = 0
      "00000" when "000010111000000", -- t[1472] = 0
      "00000" when "000010111000001", -- t[1473] = 0
      "00000" when "000010111000010", -- t[1474] = 0
      "00000" when "000010111000011", -- t[1475] = 0
      "00000" when "000010111000100", -- t[1476] = 0
      "00000" when "000010111000101", -- t[1477] = 0
      "00000" when "000010111000110", -- t[1478] = 0
      "00000" when "000010111000111", -- t[1479] = 0
      "00000" when "000010111001000", -- t[1480] = 0
      "00000" when "000010111001001", -- t[1481] = 0
      "00000" when "000010111001010", -- t[1482] = 0
      "00000" when "000010111001011", -- t[1483] = 0
      "00000" when "000010111001100", -- t[1484] = 0
      "00000" when "000010111001101", -- t[1485] = 0
      "00000" when "000010111001110", -- t[1486] = 0
      "00000" when "000010111001111", -- t[1487] = 0
      "00000" when "000010111010000", -- t[1488] = 0
      "00000" when "000010111010001", -- t[1489] = 0
      "00000" when "000010111010010", -- t[1490] = 0
      "00000" when "000010111010011", -- t[1491] = 0
      "00000" when "000010111010100", -- t[1492] = 0
      "00000" when "000010111010101", -- t[1493] = 0
      "00000" when "000010111010110", -- t[1494] = 0
      "00000" when "000010111010111", -- t[1495] = 0
      "00000" when "000010111011000", -- t[1496] = 0
      "00000" when "000010111011001", -- t[1497] = 0
      "00000" when "000010111011010", -- t[1498] = 0
      "00000" when "000010111011011", -- t[1499] = 0
      "00000" when "000010111011100", -- t[1500] = 0
      "00000" when "000010111011101", -- t[1501] = 0
      "00000" when "000010111011110", -- t[1502] = 0
      "00000" when "000010111011111", -- t[1503] = 0
      "00000" when "000010111100000", -- t[1504] = 0
      "00000" when "000010111100001", -- t[1505] = 0
      "00000" when "000010111100010", -- t[1506] = 0
      "00000" when "000010111100011", -- t[1507] = 0
      "00000" when "000010111100100", -- t[1508] = 0
      "00000" when "000010111100101", -- t[1509] = 0
      "00000" when "000010111100110", -- t[1510] = 0
      "00000" when "000010111100111", -- t[1511] = 0
      "00000" when "000010111101000", -- t[1512] = 0
      "00000" when "000010111101001", -- t[1513] = 0
      "00000" when "000010111101010", -- t[1514] = 0
      "00000" when "000010111101011", -- t[1515] = 0
      "00000" when "000010111101100", -- t[1516] = 0
      "00000" when "000010111101101", -- t[1517] = 0
      "00000" when "000010111101110", -- t[1518] = 0
      "00000" when "000010111101111", -- t[1519] = 0
      "00000" when "000010111110000", -- t[1520] = 0
      "00000" when "000010111110001", -- t[1521] = 0
      "00000" when "000010111110010", -- t[1522] = 0
      "00000" when "000010111110011", -- t[1523] = 0
      "00000" when "000010111110100", -- t[1524] = 0
      "00000" when "000010111110101", -- t[1525] = 0
      "00000" when "000010111110110", -- t[1526] = 0
      "00000" when "000010111110111", -- t[1527] = 0
      "00000" when "000010111111000", -- t[1528] = 0
      "00000" when "000010111111001", -- t[1529] = 0
      "00000" when "000010111111010", -- t[1530] = 0
      "00000" when "000010111111011", -- t[1531] = 0
      "00000" when "000010111111100", -- t[1532] = 0
      "00000" when "000010111111101", -- t[1533] = 0
      "00000" when "000010111111110", -- t[1534] = 0
      "00000" when "000010111111111", -- t[1535] = 0
      "00000" when "000011000000000", -- t[1536] = 0
      "00000" when "000011000000001", -- t[1537] = 0
      "00000" when "000011000000010", -- t[1538] = 0
      "00000" when "000011000000011", -- t[1539] = 0
      "00000" when "000011000000100", -- t[1540] = 0
      "00000" when "000011000000101", -- t[1541] = 0
      "00000" when "000011000000110", -- t[1542] = 0
      "00000" when "000011000000111", -- t[1543] = 0
      "00000" when "000011000001000", -- t[1544] = 0
      "00000" when "000011000001001", -- t[1545] = 0
      "00000" when "000011000001010", -- t[1546] = 0
      "00000" when "000011000001011", -- t[1547] = 0
      "00000" when "000011000001100", -- t[1548] = 0
      "00000" when "000011000001101", -- t[1549] = 0
      "00000" when "000011000001110", -- t[1550] = 0
      "00000" when "000011000001111", -- t[1551] = 0
      "00000" when "000011000010000", -- t[1552] = 0
      "00000" when "000011000010001", -- t[1553] = 0
      "00000" when "000011000010010", -- t[1554] = 0
      "00000" when "000011000010011", -- t[1555] = 0
      "00000" when "000011000010100", -- t[1556] = 0
      "00000" when "000011000010101", -- t[1557] = 0
      "00000" when "000011000010110", -- t[1558] = 0
      "00000" when "000011000010111", -- t[1559] = 0
      "00000" when "000011000011000", -- t[1560] = 0
      "00000" when "000011000011001", -- t[1561] = 0
      "00000" when "000011000011010", -- t[1562] = 0
      "00000" when "000011000011011", -- t[1563] = 0
      "00000" when "000011000011100", -- t[1564] = 0
      "00000" when "000011000011101", -- t[1565] = 0
      "00000" when "000011000011110", -- t[1566] = 0
      "00000" when "000011000011111", -- t[1567] = 0
      "00000" when "000011000100000", -- t[1568] = 0
      "00000" when "000011000100001", -- t[1569] = 0
      "00000" when "000011000100010", -- t[1570] = 0
      "00000" when "000011000100011", -- t[1571] = 0
      "00000" when "000011000100100", -- t[1572] = 0
      "00000" when "000011000100101", -- t[1573] = 0
      "00000" when "000011000100110", -- t[1574] = 0
      "00000" when "000011000100111", -- t[1575] = 0
      "00000" when "000011000101000", -- t[1576] = 0
      "00000" when "000011000101001", -- t[1577] = 0
      "00000" when "000011000101010", -- t[1578] = 0
      "00000" when "000011000101011", -- t[1579] = 0
      "00000" when "000011000101100", -- t[1580] = 0
      "00000" when "000011000101101", -- t[1581] = 0
      "00000" when "000011000101110", -- t[1582] = 0
      "00000" when "000011000101111", -- t[1583] = 0
      "00000" when "000011000110000", -- t[1584] = 0
      "00000" when "000011000110001", -- t[1585] = 0
      "00000" when "000011000110010", -- t[1586] = 0
      "00000" when "000011000110011", -- t[1587] = 0
      "00000" when "000011000110100", -- t[1588] = 0
      "00000" when "000011000110101", -- t[1589] = 0
      "00000" when "000011000110110", -- t[1590] = 0
      "00000" when "000011000110111", -- t[1591] = 0
      "00000" when "000011000111000", -- t[1592] = 0
      "00000" when "000011000111001", -- t[1593] = 0
      "00000" when "000011000111010", -- t[1594] = 0
      "00000" when "000011000111011", -- t[1595] = 0
      "00000" when "000011000111100", -- t[1596] = 0
      "00000" when "000011000111101", -- t[1597] = 0
      "00000" when "000011000111110", -- t[1598] = 0
      "00000" when "000011000111111", -- t[1599] = 0
      "00000" when "000011001000000", -- t[1600] = 0
      "00000" when "000011001000001", -- t[1601] = 0
      "00000" when "000011001000010", -- t[1602] = 0
      "00000" when "000011001000011", -- t[1603] = 0
      "00000" when "000011001000100", -- t[1604] = 0
      "00000" when "000011001000101", -- t[1605] = 0
      "00000" when "000011001000110", -- t[1606] = 0
      "00000" when "000011001000111", -- t[1607] = 0
      "00000" when "000011001001000", -- t[1608] = 0
      "00000" when "000011001001001", -- t[1609] = 0
      "00000" when "000011001001010", -- t[1610] = 0
      "00000" when "000011001001011", -- t[1611] = 0
      "00000" when "000011001001100", -- t[1612] = 0
      "00000" when "000011001001101", -- t[1613] = 0
      "00000" when "000011001001110", -- t[1614] = 0
      "00000" when "000011001001111", -- t[1615] = 0
      "00000" when "000011001010000", -- t[1616] = 0
      "00000" when "000011001010001", -- t[1617] = 0
      "00000" when "000011001010010", -- t[1618] = 0
      "00000" when "000011001010011", -- t[1619] = 0
      "00000" when "000011001010100", -- t[1620] = 0
      "00000" when "000011001010101", -- t[1621] = 0
      "00000" when "000011001010110", -- t[1622] = 0
      "00000" when "000011001010111", -- t[1623] = 0
      "00000" when "000011001011000", -- t[1624] = 0
      "00000" when "000011001011001", -- t[1625] = 0
      "00000" when "000011001011010", -- t[1626] = 0
      "00000" when "000011001011011", -- t[1627] = 0
      "00000" when "000011001011100", -- t[1628] = 0
      "00000" when "000011001011101", -- t[1629] = 0
      "00000" when "000011001011110", -- t[1630] = 0
      "00000" when "000011001011111", -- t[1631] = 0
      "00000" when "000011001100000", -- t[1632] = 0
      "00000" when "000011001100001", -- t[1633] = 0
      "00000" when "000011001100010", -- t[1634] = 0
      "00000" when "000011001100011", -- t[1635] = 0
      "00000" when "000011001100100", -- t[1636] = 0
      "00000" when "000011001100101", -- t[1637] = 0
      "00000" when "000011001100110", -- t[1638] = 0
      "00000" when "000011001100111", -- t[1639] = 0
      "00000" when "000011001101000", -- t[1640] = 0
      "00000" when "000011001101001", -- t[1641] = 0
      "00000" when "000011001101010", -- t[1642] = 0
      "00000" when "000011001101011", -- t[1643] = 0
      "00000" when "000011001101100", -- t[1644] = 0
      "00000" when "000011001101101", -- t[1645] = 0
      "00000" when "000011001101110", -- t[1646] = 0
      "00000" when "000011001101111", -- t[1647] = 0
      "00000" when "000011001110000", -- t[1648] = 0
      "00000" when "000011001110001", -- t[1649] = 0
      "00000" when "000011001110010", -- t[1650] = 0
      "00000" when "000011001110011", -- t[1651] = 0
      "00000" when "000011001110100", -- t[1652] = 0
      "00000" when "000011001110101", -- t[1653] = 0
      "00000" when "000011001110110", -- t[1654] = 0
      "00000" when "000011001110111", -- t[1655] = 0
      "00000" when "000011001111000", -- t[1656] = 0
      "00000" when "000011001111001", -- t[1657] = 0
      "00000" when "000011001111010", -- t[1658] = 0
      "00000" when "000011001111011", -- t[1659] = 0
      "00000" when "000011001111100", -- t[1660] = 0
      "00000" when "000011001111101", -- t[1661] = 0
      "00000" when "000011001111110", -- t[1662] = 0
      "00000" when "000011001111111", -- t[1663] = 0
      "00000" when "000011010000000", -- t[1664] = 0
      "00000" when "000011010000001", -- t[1665] = 0
      "00000" when "000011010000010", -- t[1666] = 0
      "00000" when "000011010000011", -- t[1667] = 0
      "00000" when "000011010000100", -- t[1668] = 0
      "00000" when "000011010000101", -- t[1669] = 0
      "00000" when "000011010000110", -- t[1670] = 0
      "00000" when "000011010000111", -- t[1671] = 0
      "00000" when "000011010001000", -- t[1672] = 0
      "00000" when "000011010001001", -- t[1673] = 0
      "00000" when "000011010001010", -- t[1674] = 0
      "00000" when "000011010001011", -- t[1675] = 0
      "00000" when "000011010001100", -- t[1676] = 0
      "00000" when "000011010001101", -- t[1677] = 0
      "00000" when "000011010001110", -- t[1678] = 0
      "00000" when "000011010001111", -- t[1679] = 0
      "00000" when "000011010010000", -- t[1680] = 0
      "00000" when "000011010010001", -- t[1681] = 0
      "00000" when "000011010010010", -- t[1682] = 0
      "00000" when "000011010010011", -- t[1683] = 0
      "00000" when "000011010010100", -- t[1684] = 0
      "00000" when "000011010010101", -- t[1685] = 0
      "00000" when "000011010010110", -- t[1686] = 0
      "00000" when "000011010010111", -- t[1687] = 0
      "00000" when "000011010011000", -- t[1688] = 0
      "00000" when "000011010011001", -- t[1689] = 0
      "00000" when "000011010011010", -- t[1690] = 0
      "00000" when "000011010011011", -- t[1691] = 0
      "00000" when "000011010011100", -- t[1692] = 0
      "00000" when "000011010011101", -- t[1693] = 0
      "00000" when "000011010011110", -- t[1694] = 0
      "00000" when "000011010011111", -- t[1695] = 0
      "00000" when "000011010100000", -- t[1696] = 0
      "00000" when "000011010100001", -- t[1697] = 0
      "00000" when "000011010100010", -- t[1698] = 0
      "00000" when "000011010100011", -- t[1699] = 0
      "00000" when "000011010100100", -- t[1700] = 0
      "00000" when "000011010100101", -- t[1701] = 0
      "00000" when "000011010100110", -- t[1702] = 0
      "00000" when "000011010100111", -- t[1703] = 0
      "00000" when "000011010101000", -- t[1704] = 0
      "00000" when "000011010101001", -- t[1705] = 0
      "00000" when "000011010101010", -- t[1706] = 0
      "00000" when "000011010101011", -- t[1707] = 0
      "00000" when "000011010101100", -- t[1708] = 0
      "00000" when "000011010101101", -- t[1709] = 0
      "00000" when "000011010101110", -- t[1710] = 0
      "00000" when "000011010101111", -- t[1711] = 0
      "00000" when "000011010110000", -- t[1712] = 0
      "00000" when "000011010110001", -- t[1713] = 0
      "00000" when "000011010110010", -- t[1714] = 0
      "00000" when "000011010110011", -- t[1715] = 0
      "00000" when "000011010110100", -- t[1716] = 0
      "00000" when "000011010110101", -- t[1717] = 0
      "00000" when "000011010110110", -- t[1718] = 0
      "00000" when "000011010110111", -- t[1719] = 0
      "00000" when "000011010111000", -- t[1720] = 0
      "00000" when "000011010111001", -- t[1721] = 0
      "00000" when "000011010111010", -- t[1722] = 0
      "00000" when "000011010111011", -- t[1723] = 0
      "00000" when "000011010111100", -- t[1724] = 0
      "00000" when "000011010111101", -- t[1725] = 0
      "00000" when "000011010111110", -- t[1726] = 0
      "00000" when "000011010111111", -- t[1727] = 0
      "00000" when "000011011000000", -- t[1728] = 0
      "00000" when "000011011000001", -- t[1729] = 0
      "00000" when "000011011000010", -- t[1730] = 0
      "00000" when "000011011000011", -- t[1731] = 0
      "00000" when "000011011000100", -- t[1732] = 0
      "00000" when "000011011000101", -- t[1733] = 0
      "00000" when "000011011000110", -- t[1734] = 0
      "00000" when "000011011000111", -- t[1735] = 0
      "00000" when "000011011001000", -- t[1736] = 0
      "00000" when "000011011001001", -- t[1737] = 0
      "00000" when "000011011001010", -- t[1738] = 0
      "00000" when "000011011001011", -- t[1739] = 0
      "00000" when "000011011001100", -- t[1740] = 0
      "00000" when "000011011001101", -- t[1741] = 0
      "00000" when "000011011001110", -- t[1742] = 0
      "00000" when "000011011001111", -- t[1743] = 0
      "00000" when "000011011010000", -- t[1744] = 0
      "00000" when "000011011010001", -- t[1745] = 0
      "00000" when "000011011010010", -- t[1746] = 0
      "00000" when "000011011010011", -- t[1747] = 0
      "00000" when "000011011010100", -- t[1748] = 0
      "00000" when "000011011010101", -- t[1749] = 0
      "00000" when "000011011010110", -- t[1750] = 0
      "00000" when "000011011010111", -- t[1751] = 0
      "00000" when "000011011011000", -- t[1752] = 0
      "00000" when "000011011011001", -- t[1753] = 0
      "00000" when "000011011011010", -- t[1754] = 0
      "00000" when "000011011011011", -- t[1755] = 0
      "00000" when "000011011011100", -- t[1756] = 0
      "00000" when "000011011011101", -- t[1757] = 0
      "00000" when "000011011011110", -- t[1758] = 0
      "00000" when "000011011011111", -- t[1759] = 0
      "00000" when "000011011100000", -- t[1760] = 0
      "00000" when "000011011100001", -- t[1761] = 0
      "00000" when "000011011100010", -- t[1762] = 0
      "00000" when "000011011100011", -- t[1763] = 0
      "00000" when "000011011100100", -- t[1764] = 0
      "00000" when "000011011100101", -- t[1765] = 0
      "00000" when "000011011100110", -- t[1766] = 0
      "00000" when "000011011100111", -- t[1767] = 0
      "00000" when "000011011101000", -- t[1768] = 0
      "00000" when "000011011101001", -- t[1769] = 0
      "00000" when "000011011101010", -- t[1770] = 0
      "00000" when "000011011101011", -- t[1771] = 0
      "00000" when "000011011101100", -- t[1772] = 0
      "00000" when "000011011101101", -- t[1773] = 0
      "00000" when "000011011101110", -- t[1774] = 0
      "00000" when "000011011101111", -- t[1775] = 0
      "00000" when "000011011110000", -- t[1776] = 0
      "00000" when "000011011110001", -- t[1777] = 0
      "00000" when "000011011110010", -- t[1778] = 0
      "00000" when "000011011110011", -- t[1779] = 0
      "00000" when "000011011110100", -- t[1780] = 0
      "00000" when "000011011110101", -- t[1781] = 0
      "00000" when "000011011110110", -- t[1782] = 0
      "00000" when "000011011110111", -- t[1783] = 0
      "00000" when "000011011111000", -- t[1784] = 0
      "00000" when "000011011111001", -- t[1785] = 0
      "00000" when "000011011111010", -- t[1786] = 0
      "00000" when "000011011111011", -- t[1787] = 0
      "00000" when "000011011111100", -- t[1788] = 0
      "00000" when "000011011111101", -- t[1789] = 0
      "00000" when "000011011111110", -- t[1790] = 0
      "00000" when "000011011111111", -- t[1791] = 0
      "00000" when "000011100000000", -- t[1792] = 0
      "00000" when "000011100000001", -- t[1793] = 0
      "00000" when "000011100000010", -- t[1794] = 0
      "00000" when "000011100000011", -- t[1795] = 0
      "00000" when "000011100000100", -- t[1796] = 0
      "00000" when "000011100000101", -- t[1797] = 0
      "00000" when "000011100000110", -- t[1798] = 0
      "00000" when "000011100000111", -- t[1799] = 0
      "00000" when "000011100001000", -- t[1800] = 0
      "00000" when "000011100001001", -- t[1801] = 0
      "00000" when "000011100001010", -- t[1802] = 0
      "00000" when "000011100001011", -- t[1803] = 0
      "00000" when "000011100001100", -- t[1804] = 0
      "00000" when "000011100001101", -- t[1805] = 0
      "00000" when "000011100001110", -- t[1806] = 0
      "00000" when "000011100001111", -- t[1807] = 0
      "00000" when "000011100010000", -- t[1808] = 0
      "00000" when "000011100010001", -- t[1809] = 0
      "00000" when "000011100010010", -- t[1810] = 0
      "00000" when "000011100010011", -- t[1811] = 0
      "00000" when "000011100010100", -- t[1812] = 0
      "00000" when "000011100010101", -- t[1813] = 0
      "00000" when "000011100010110", -- t[1814] = 0
      "00000" when "000011100010111", -- t[1815] = 0
      "00000" when "000011100011000", -- t[1816] = 0
      "00000" when "000011100011001", -- t[1817] = 0
      "00000" when "000011100011010", -- t[1818] = 0
      "00000" when "000011100011011", -- t[1819] = 0
      "00000" when "000011100011100", -- t[1820] = 0
      "00000" when "000011100011101", -- t[1821] = 0
      "00000" when "000011100011110", -- t[1822] = 0
      "00000" when "000011100011111", -- t[1823] = 0
      "00000" when "000011100100000", -- t[1824] = 0
      "00000" when "000011100100001", -- t[1825] = 0
      "00000" when "000011100100010", -- t[1826] = 0
      "00000" when "000011100100011", -- t[1827] = 0
      "00000" when "000011100100100", -- t[1828] = 0
      "00000" when "000011100100101", -- t[1829] = 0
      "00000" when "000011100100110", -- t[1830] = 0
      "00000" when "000011100100111", -- t[1831] = 0
      "00000" when "000011100101000", -- t[1832] = 0
      "00000" when "000011100101001", -- t[1833] = 0
      "00000" when "000011100101010", -- t[1834] = 0
      "00000" when "000011100101011", -- t[1835] = 0
      "00000" when "000011100101100", -- t[1836] = 0
      "00000" when "000011100101101", -- t[1837] = 0
      "00000" when "000011100101110", -- t[1838] = 0
      "00000" when "000011100101111", -- t[1839] = 0
      "00000" when "000011100110000", -- t[1840] = 0
      "00000" when "000011100110001", -- t[1841] = 0
      "00000" when "000011100110010", -- t[1842] = 0
      "00000" when "000011100110011", -- t[1843] = 0
      "00000" when "000011100110100", -- t[1844] = 0
      "00000" when "000011100110101", -- t[1845] = 0
      "00000" when "000011100110110", -- t[1846] = 0
      "00000" when "000011100110111", -- t[1847] = 0
      "00000" when "000011100111000", -- t[1848] = 0
      "00000" when "000011100111001", -- t[1849] = 0
      "00000" when "000011100111010", -- t[1850] = 0
      "00000" when "000011100111011", -- t[1851] = 0
      "00000" when "000011100111100", -- t[1852] = 0
      "00000" when "000011100111101", -- t[1853] = 0
      "00000" when "000011100111110", -- t[1854] = 0
      "00000" when "000011100111111", -- t[1855] = 0
      "00000" when "000011101000000", -- t[1856] = 0
      "00000" when "000011101000001", -- t[1857] = 0
      "00000" when "000011101000010", -- t[1858] = 0
      "00000" when "000011101000011", -- t[1859] = 0
      "00000" when "000011101000100", -- t[1860] = 0
      "00000" when "000011101000101", -- t[1861] = 0
      "00000" when "000011101000110", -- t[1862] = 0
      "00000" when "000011101000111", -- t[1863] = 0
      "00000" when "000011101001000", -- t[1864] = 0
      "00000" when "000011101001001", -- t[1865] = 0
      "00000" when "000011101001010", -- t[1866] = 0
      "00000" when "000011101001011", -- t[1867] = 0
      "00000" when "000011101001100", -- t[1868] = 0
      "00000" when "000011101001101", -- t[1869] = 0
      "00000" when "000011101001110", -- t[1870] = 0
      "00000" when "000011101001111", -- t[1871] = 0
      "00000" when "000011101010000", -- t[1872] = 0
      "00000" when "000011101010001", -- t[1873] = 0
      "00000" when "000011101010010", -- t[1874] = 0
      "00000" when "000011101010011", -- t[1875] = 0
      "00000" when "000011101010100", -- t[1876] = 0
      "00000" when "000011101010101", -- t[1877] = 0
      "00000" when "000011101010110", -- t[1878] = 0
      "00000" when "000011101010111", -- t[1879] = 0
      "00000" when "000011101011000", -- t[1880] = 0
      "00000" when "000011101011001", -- t[1881] = 0
      "00000" when "000011101011010", -- t[1882] = 0
      "00000" when "000011101011011", -- t[1883] = 0
      "00000" when "000011101011100", -- t[1884] = 0
      "00000" when "000011101011101", -- t[1885] = 0
      "00000" when "000011101011110", -- t[1886] = 0
      "00000" when "000011101011111", -- t[1887] = 0
      "00000" when "000011101100000", -- t[1888] = 0
      "00000" when "000011101100001", -- t[1889] = 0
      "00000" when "000011101100010", -- t[1890] = 0
      "00000" when "000011101100011", -- t[1891] = 0
      "00000" when "000011101100100", -- t[1892] = 0
      "00000" when "000011101100101", -- t[1893] = 0
      "00000" when "000011101100110", -- t[1894] = 0
      "00000" when "000011101100111", -- t[1895] = 0
      "00000" when "000011101101000", -- t[1896] = 0
      "00000" when "000011101101001", -- t[1897] = 0
      "00000" when "000011101101010", -- t[1898] = 0
      "00000" when "000011101101011", -- t[1899] = 0
      "00000" when "000011101101100", -- t[1900] = 0
      "00000" when "000011101101101", -- t[1901] = 0
      "00000" when "000011101101110", -- t[1902] = 0
      "00000" when "000011101101111", -- t[1903] = 0
      "00000" when "000011101110000", -- t[1904] = 0
      "00000" when "000011101110001", -- t[1905] = 0
      "00000" when "000011101110010", -- t[1906] = 0
      "00000" when "000011101110011", -- t[1907] = 0
      "00000" when "000011101110100", -- t[1908] = 0
      "00000" when "000011101110101", -- t[1909] = 0
      "00000" when "000011101110110", -- t[1910] = 0
      "00000" when "000011101110111", -- t[1911] = 0
      "00000" when "000011101111000", -- t[1912] = 0
      "00000" when "000011101111001", -- t[1913] = 0
      "00000" when "000011101111010", -- t[1914] = 0
      "00000" when "000011101111011", -- t[1915] = 0
      "00000" when "000011101111100", -- t[1916] = 0
      "00000" when "000011101111101", -- t[1917] = 0
      "00000" when "000011101111110", -- t[1918] = 0
      "00000" when "000011101111111", -- t[1919] = 0
      "00000" when "000011110000000", -- t[1920] = 0
      "00000" when "000011110000001", -- t[1921] = 0
      "00000" when "000011110000010", -- t[1922] = 0
      "00000" when "000011110000011", -- t[1923] = 0
      "00000" when "000011110000100", -- t[1924] = 0
      "00000" when "000011110000101", -- t[1925] = 0
      "00000" when "000011110000110", -- t[1926] = 0
      "00000" when "000011110000111", -- t[1927] = 0
      "00000" when "000011110001000", -- t[1928] = 0
      "00000" when "000011110001001", -- t[1929] = 0
      "00000" when "000011110001010", -- t[1930] = 0
      "00000" when "000011110001011", -- t[1931] = 0
      "00000" when "000011110001100", -- t[1932] = 0
      "00000" when "000011110001101", -- t[1933] = 0
      "00000" when "000011110001110", -- t[1934] = 0
      "00000" when "000011110001111", -- t[1935] = 0
      "00000" when "000011110010000", -- t[1936] = 0
      "00000" when "000011110010001", -- t[1937] = 0
      "00000" when "000011110010010", -- t[1938] = 0
      "00000" when "000011110010011", -- t[1939] = 0
      "00000" when "000011110010100", -- t[1940] = 0
      "00000" when "000011110010101", -- t[1941] = 0
      "00000" when "000011110010110", -- t[1942] = 0
      "00000" when "000011110010111", -- t[1943] = 0
      "00000" when "000011110011000", -- t[1944] = 0
      "00000" when "000011110011001", -- t[1945] = 0
      "00000" when "000011110011010", -- t[1946] = 0
      "00000" when "000011110011011", -- t[1947] = 0
      "00000" when "000011110011100", -- t[1948] = 0
      "00000" when "000011110011101", -- t[1949] = 0
      "00000" when "000011110011110", -- t[1950] = 0
      "00000" when "000011110011111", -- t[1951] = 0
      "00000" when "000011110100000", -- t[1952] = 0
      "00000" when "000011110100001", -- t[1953] = 0
      "00000" when "000011110100010", -- t[1954] = 0
      "00000" when "000011110100011", -- t[1955] = 0
      "00000" when "000011110100100", -- t[1956] = 0
      "00000" when "000011110100101", -- t[1957] = 0
      "00000" when "000011110100110", -- t[1958] = 0
      "00000" when "000011110100111", -- t[1959] = 0
      "00000" when "000011110101000", -- t[1960] = 0
      "00000" when "000011110101001", -- t[1961] = 0
      "00000" when "000011110101010", -- t[1962] = 0
      "00000" when "000011110101011", -- t[1963] = 0
      "00000" when "000011110101100", -- t[1964] = 0
      "00000" when "000011110101101", -- t[1965] = 0
      "00000" when "000011110101110", -- t[1966] = 0
      "00000" when "000011110101111", -- t[1967] = 0
      "00000" when "000011110110000", -- t[1968] = 0
      "00000" when "000011110110001", -- t[1969] = 0
      "00000" when "000011110110010", -- t[1970] = 0
      "00000" when "000011110110011", -- t[1971] = 0
      "00000" when "000011110110100", -- t[1972] = 0
      "00000" when "000011110110101", -- t[1973] = 0
      "00000" when "000011110110110", -- t[1974] = 0
      "00000" when "000011110110111", -- t[1975] = 0
      "00000" when "000011110111000", -- t[1976] = 0
      "00000" when "000011110111001", -- t[1977] = 0
      "00000" when "000011110111010", -- t[1978] = 0
      "00000" when "000011110111011", -- t[1979] = 0
      "00000" when "000011110111100", -- t[1980] = 0
      "00000" when "000011110111101", -- t[1981] = 0
      "00000" when "000011110111110", -- t[1982] = 0
      "00000" when "000011110111111", -- t[1983] = 0
      "00000" when "000011111000000", -- t[1984] = 0
      "00000" when "000011111000001", -- t[1985] = 0
      "00000" when "000011111000010", -- t[1986] = 0
      "00000" when "000011111000011", -- t[1987] = 0
      "00000" when "000011111000100", -- t[1988] = 0
      "00000" when "000011111000101", -- t[1989] = 0
      "00000" when "000011111000110", -- t[1990] = 0
      "00000" when "000011111000111", -- t[1991] = 0
      "00000" when "000011111001000", -- t[1992] = 0
      "00000" when "000011111001001", -- t[1993] = 0
      "00000" when "000011111001010", -- t[1994] = 0
      "00000" when "000011111001011", -- t[1995] = 0
      "00000" when "000011111001100", -- t[1996] = 0
      "00000" when "000011111001101", -- t[1997] = 0
      "00000" when "000011111001110", -- t[1998] = 0
      "00000" when "000011111001111", -- t[1999] = 0
      "00000" when "000011111010000", -- t[2000] = 0
      "00000" when "000011111010001", -- t[2001] = 0
      "00000" when "000011111010010", -- t[2002] = 0
      "00000" when "000011111010011", -- t[2003] = 0
      "00000" when "000011111010100", -- t[2004] = 0
      "00000" when "000011111010101", -- t[2005] = 0
      "00000" when "000011111010110", -- t[2006] = 0
      "00000" when "000011111010111", -- t[2007] = 0
      "00000" when "000011111011000", -- t[2008] = 0
      "00000" when "000011111011001", -- t[2009] = 0
      "00000" when "000011111011010", -- t[2010] = 0
      "00000" when "000011111011011", -- t[2011] = 0
      "00000" when "000011111011100", -- t[2012] = 0
      "00000" when "000011111011101", -- t[2013] = 0
      "00000" when "000011111011110", -- t[2014] = 0
      "00000" when "000011111011111", -- t[2015] = 0
      "00000" when "000011111100000", -- t[2016] = 0
      "00000" when "000011111100001", -- t[2017] = 0
      "00000" when "000011111100010", -- t[2018] = 0
      "00000" when "000011111100011", -- t[2019] = 0
      "00000" when "000011111100100", -- t[2020] = 0
      "00000" when "000011111100101", -- t[2021] = 0
      "00000" when "000011111100110", -- t[2022] = 0
      "00000" when "000011111100111", -- t[2023] = 0
      "00000" when "000011111101000", -- t[2024] = 0
      "00000" when "000011111101001", -- t[2025] = 0
      "00000" when "000011111101010", -- t[2026] = 0
      "00000" when "000011111101011", -- t[2027] = 0
      "00000" when "000011111101100", -- t[2028] = 0
      "00000" when "000011111101101", -- t[2029] = 0
      "00000" when "000011111101110", -- t[2030] = 0
      "00000" when "000011111101111", -- t[2031] = 0
      "00000" when "000011111110000", -- t[2032] = 0
      "00000" when "000011111110001", -- t[2033] = 0
      "00000" when "000011111110010", -- t[2034] = 0
      "00000" when "000011111110011", -- t[2035] = 0
      "00000" when "000011111110100", -- t[2036] = 0
      "00000" when "000011111110101", -- t[2037] = 0
      "00000" when "000011111110110", -- t[2038] = 0
      "00000" when "000011111110111", -- t[2039] = 0
      "00000" when "000011111111000", -- t[2040] = 0
      "00000" when "000011111111001", -- t[2041] = 0
      "00000" when "000011111111010", -- t[2042] = 0
      "00000" when "000011111111011", -- t[2043] = 0
      "00000" when "000011111111100", -- t[2044] = 0
      "00000" when "000011111111101", -- t[2045] = 0
      "00000" when "000011111111110", -- t[2046] = 0
      "00000" when "000011111111111", -- t[2047] = 0
      "00000" when "000100000000000", -- t[2048] = 0
      "00000" when "000100000000001", -- t[2049] = 0
      "00000" when "000100000000010", -- t[2050] = 0
      "00000" when "000100000000011", -- t[2051] = 0
      "00000" when "000100000000100", -- t[2052] = 0
      "00000" when "000100000000101", -- t[2053] = 0
      "00000" when "000100000000110", -- t[2054] = 0
      "00000" when "000100000000111", -- t[2055] = 0
      "00000" when "000100000001000", -- t[2056] = 0
      "00000" when "000100000001001", -- t[2057] = 0
      "00000" when "000100000001010", -- t[2058] = 0
      "00000" when "000100000001011", -- t[2059] = 0
      "00000" when "000100000001100", -- t[2060] = 0
      "00000" when "000100000001101", -- t[2061] = 0
      "00000" when "000100000001110", -- t[2062] = 0
      "00000" when "000100000001111", -- t[2063] = 0
      "00000" when "000100000010000", -- t[2064] = 0
      "00000" when "000100000010001", -- t[2065] = 0
      "00000" when "000100000010010", -- t[2066] = 0
      "00000" when "000100000010011", -- t[2067] = 0
      "00000" when "000100000010100", -- t[2068] = 0
      "00000" when "000100000010101", -- t[2069] = 0
      "00000" when "000100000010110", -- t[2070] = 0
      "00000" when "000100000010111", -- t[2071] = 0
      "00000" when "000100000011000", -- t[2072] = 0
      "00000" when "000100000011001", -- t[2073] = 0
      "00000" when "000100000011010", -- t[2074] = 0
      "00000" when "000100000011011", -- t[2075] = 0
      "00000" when "000100000011100", -- t[2076] = 0
      "00000" when "000100000011101", -- t[2077] = 0
      "00000" when "000100000011110", -- t[2078] = 0
      "00000" when "000100000011111", -- t[2079] = 0
      "00000" when "000100000100000", -- t[2080] = 0
      "00000" when "000100000100001", -- t[2081] = 0
      "00000" when "000100000100010", -- t[2082] = 0
      "00000" when "000100000100011", -- t[2083] = 0
      "00000" when "000100000100100", -- t[2084] = 0
      "00000" when "000100000100101", -- t[2085] = 0
      "00000" when "000100000100110", -- t[2086] = 0
      "00000" when "000100000100111", -- t[2087] = 0
      "00000" when "000100000101000", -- t[2088] = 0
      "00000" when "000100000101001", -- t[2089] = 0
      "00000" when "000100000101010", -- t[2090] = 0
      "00000" when "000100000101011", -- t[2091] = 0
      "00000" when "000100000101100", -- t[2092] = 0
      "00000" when "000100000101101", -- t[2093] = 0
      "00000" when "000100000101110", -- t[2094] = 0
      "00000" when "000100000101111", -- t[2095] = 0
      "00000" when "000100000110000", -- t[2096] = 0
      "00000" when "000100000110001", -- t[2097] = 0
      "00000" when "000100000110010", -- t[2098] = 0
      "00000" when "000100000110011", -- t[2099] = 0
      "00000" when "000100000110100", -- t[2100] = 0
      "00000" when "000100000110101", -- t[2101] = 0
      "00000" when "000100000110110", -- t[2102] = 0
      "00000" when "000100000110111", -- t[2103] = 0
      "00000" when "000100000111000", -- t[2104] = 0
      "00000" when "000100000111001", -- t[2105] = 0
      "00000" when "000100000111010", -- t[2106] = 0
      "00000" when "000100000111011", -- t[2107] = 0
      "00000" when "000100000111100", -- t[2108] = 0
      "00000" when "000100000111101", -- t[2109] = 0
      "00000" when "000100000111110", -- t[2110] = 0
      "00000" when "000100000111111", -- t[2111] = 0
      "00000" when "000100001000000", -- t[2112] = 0
      "00000" when "000100001000001", -- t[2113] = 0
      "00000" when "000100001000010", -- t[2114] = 0
      "00000" when "000100001000011", -- t[2115] = 0
      "00000" when "000100001000100", -- t[2116] = 0
      "00000" when "000100001000101", -- t[2117] = 0
      "00000" when "000100001000110", -- t[2118] = 0
      "00000" when "000100001000111", -- t[2119] = 0
      "00000" when "000100001001000", -- t[2120] = 0
      "00000" when "000100001001001", -- t[2121] = 0
      "00000" when "000100001001010", -- t[2122] = 0
      "00000" when "000100001001011", -- t[2123] = 0
      "00000" when "000100001001100", -- t[2124] = 0
      "00000" when "000100001001101", -- t[2125] = 0
      "00000" when "000100001001110", -- t[2126] = 0
      "00000" when "000100001001111", -- t[2127] = 0
      "00000" when "000100001010000", -- t[2128] = 0
      "00000" when "000100001010001", -- t[2129] = 0
      "00000" when "000100001010010", -- t[2130] = 0
      "00000" when "000100001010011", -- t[2131] = 0
      "00000" when "000100001010100", -- t[2132] = 0
      "00000" when "000100001010101", -- t[2133] = 0
      "00000" when "000100001010110", -- t[2134] = 0
      "00000" when "000100001010111", -- t[2135] = 0
      "00000" when "000100001011000", -- t[2136] = 0
      "00000" when "000100001011001", -- t[2137] = 0
      "00000" when "000100001011010", -- t[2138] = 0
      "00000" when "000100001011011", -- t[2139] = 0
      "00000" when "000100001011100", -- t[2140] = 0
      "00000" when "000100001011101", -- t[2141] = 0
      "00000" when "000100001011110", -- t[2142] = 0
      "00000" when "000100001011111", -- t[2143] = 0
      "00000" when "000100001100000", -- t[2144] = 0
      "00000" when "000100001100001", -- t[2145] = 0
      "00000" when "000100001100010", -- t[2146] = 0
      "00000" when "000100001100011", -- t[2147] = 0
      "00000" when "000100001100100", -- t[2148] = 0
      "00000" when "000100001100101", -- t[2149] = 0
      "00000" when "000100001100110", -- t[2150] = 0
      "00000" when "000100001100111", -- t[2151] = 0
      "00000" when "000100001101000", -- t[2152] = 0
      "00000" when "000100001101001", -- t[2153] = 0
      "00000" when "000100001101010", -- t[2154] = 0
      "00000" when "000100001101011", -- t[2155] = 0
      "00000" when "000100001101100", -- t[2156] = 0
      "00000" when "000100001101101", -- t[2157] = 0
      "00000" when "000100001101110", -- t[2158] = 0
      "00000" when "000100001101111", -- t[2159] = 0
      "00000" when "000100001110000", -- t[2160] = 0
      "00000" when "000100001110001", -- t[2161] = 0
      "00000" when "000100001110010", -- t[2162] = 0
      "00000" when "000100001110011", -- t[2163] = 0
      "00000" when "000100001110100", -- t[2164] = 0
      "00000" when "000100001110101", -- t[2165] = 0
      "00000" when "000100001110110", -- t[2166] = 0
      "00000" when "000100001110111", -- t[2167] = 0
      "00000" when "000100001111000", -- t[2168] = 0
      "00000" when "000100001111001", -- t[2169] = 0
      "00000" when "000100001111010", -- t[2170] = 0
      "00000" when "000100001111011", -- t[2171] = 0
      "00000" when "000100001111100", -- t[2172] = 0
      "00000" when "000100001111101", -- t[2173] = 0
      "00000" when "000100001111110", -- t[2174] = 0
      "00000" when "000100001111111", -- t[2175] = 0
      "00000" when "000100010000000", -- t[2176] = 0
      "00000" when "000100010000001", -- t[2177] = 0
      "00000" when "000100010000010", -- t[2178] = 0
      "00000" when "000100010000011", -- t[2179] = 0
      "00000" when "000100010000100", -- t[2180] = 0
      "00000" when "000100010000101", -- t[2181] = 0
      "00000" when "000100010000110", -- t[2182] = 0
      "00000" when "000100010000111", -- t[2183] = 0
      "00000" when "000100010001000", -- t[2184] = 0
      "00000" when "000100010001001", -- t[2185] = 0
      "00000" when "000100010001010", -- t[2186] = 0
      "00000" when "000100010001011", -- t[2187] = 0
      "00000" when "000100010001100", -- t[2188] = 0
      "00000" when "000100010001101", -- t[2189] = 0
      "00000" when "000100010001110", -- t[2190] = 0
      "00000" when "000100010001111", -- t[2191] = 0
      "00000" when "000100010010000", -- t[2192] = 0
      "00000" when "000100010010001", -- t[2193] = 0
      "00000" when "000100010010010", -- t[2194] = 0
      "00000" when "000100010010011", -- t[2195] = 0
      "00000" when "000100010010100", -- t[2196] = 0
      "00000" when "000100010010101", -- t[2197] = 0
      "00000" when "000100010010110", -- t[2198] = 0
      "00000" when "000100010010111", -- t[2199] = 0
      "00000" when "000100010011000", -- t[2200] = 0
      "00000" when "000100010011001", -- t[2201] = 0
      "00000" when "000100010011010", -- t[2202] = 0
      "00000" when "000100010011011", -- t[2203] = 0
      "00000" when "000100010011100", -- t[2204] = 0
      "00000" when "000100010011101", -- t[2205] = 0
      "00000" when "000100010011110", -- t[2206] = 0
      "00000" when "000100010011111", -- t[2207] = 0
      "00000" when "000100010100000", -- t[2208] = 0
      "00000" when "000100010100001", -- t[2209] = 0
      "00000" when "000100010100010", -- t[2210] = 0
      "00000" when "000100010100011", -- t[2211] = 0
      "00000" when "000100010100100", -- t[2212] = 0
      "00000" when "000100010100101", -- t[2213] = 0
      "00000" when "000100010100110", -- t[2214] = 0
      "00000" when "000100010100111", -- t[2215] = 0
      "00000" when "000100010101000", -- t[2216] = 0
      "00000" when "000100010101001", -- t[2217] = 0
      "00000" when "000100010101010", -- t[2218] = 0
      "00000" when "000100010101011", -- t[2219] = 0
      "00000" when "000100010101100", -- t[2220] = 0
      "00000" when "000100010101101", -- t[2221] = 0
      "00000" when "000100010101110", -- t[2222] = 0
      "00000" when "000100010101111", -- t[2223] = 0
      "00000" when "000100010110000", -- t[2224] = 0
      "00000" when "000100010110001", -- t[2225] = 0
      "00000" when "000100010110010", -- t[2226] = 0
      "00000" when "000100010110011", -- t[2227] = 0
      "00000" when "000100010110100", -- t[2228] = 0
      "00000" when "000100010110101", -- t[2229] = 0
      "00000" when "000100010110110", -- t[2230] = 0
      "00000" when "000100010110111", -- t[2231] = 0
      "00000" when "000100010111000", -- t[2232] = 0
      "00000" when "000100010111001", -- t[2233] = 0
      "00000" when "000100010111010", -- t[2234] = 0
      "00000" when "000100010111011", -- t[2235] = 0
      "00000" when "000100010111100", -- t[2236] = 0
      "00000" when "000100010111101", -- t[2237] = 0
      "00000" when "000100010111110", -- t[2238] = 0
      "00000" when "000100010111111", -- t[2239] = 0
      "00000" when "000100011000000", -- t[2240] = 0
      "00000" when "000100011000001", -- t[2241] = 0
      "00000" when "000100011000010", -- t[2242] = 0
      "00000" when "000100011000011", -- t[2243] = 0
      "00000" when "000100011000100", -- t[2244] = 0
      "00000" when "000100011000101", -- t[2245] = 0
      "00000" when "000100011000110", -- t[2246] = 0
      "00000" when "000100011000111", -- t[2247] = 0
      "00000" when "000100011001000", -- t[2248] = 0
      "00000" when "000100011001001", -- t[2249] = 0
      "00000" when "000100011001010", -- t[2250] = 0
      "00000" when "000100011001011", -- t[2251] = 0
      "00000" when "000100011001100", -- t[2252] = 0
      "00000" when "000100011001101", -- t[2253] = 0
      "00000" when "000100011001110", -- t[2254] = 0
      "00000" when "000100011001111", -- t[2255] = 0
      "00000" when "000100011010000", -- t[2256] = 0
      "00000" when "000100011010001", -- t[2257] = 0
      "00000" when "000100011010010", -- t[2258] = 0
      "00000" when "000100011010011", -- t[2259] = 0
      "00000" when "000100011010100", -- t[2260] = 0
      "00000" when "000100011010101", -- t[2261] = 0
      "00000" when "000100011010110", -- t[2262] = 0
      "00000" when "000100011010111", -- t[2263] = 0
      "00000" when "000100011011000", -- t[2264] = 0
      "00000" when "000100011011001", -- t[2265] = 0
      "00000" when "000100011011010", -- t[2266] = 0
      "00000" when "000100011011011", -- t[2267] = 0
      "00000" when "000100011011100", -- t[2268] = 0
      "00000" when "000100011011101", -- t[2269] = 0
      "00000" when "000100011011110", -- t[2270] = 0
      "00000" when "000100011011111", -- t[2271] = 0
      "00000" when "000100011100000", -- t[2272] = 0
      "00000" when "000100011100001", -- t[2273] = 0
      "00000" when "000100011100010", -- t[2274] = 0
      "00000" when "000100011100011", -- t[2275] = 0
      "00000" when "000100011100100", -- t[2276] = 0
      "00000" when "000100011100101", -- t[2277] = 0
      "00000" when "000100011100110", -- t[2278] = 0
      "00000" when "000100011100111", -- t[2279] = 0
      "00000" when "000100011101000", -- t[2280] = 0
      "00000" when "000100011101001", -- t[2281] = 0
      "00000" when "000100011101010", -- t[2282] = 0
      "00000" when "000100011101011", -- t[2283] = 0
      "00000" when "000100011101100", -- t[2284] = 0
      "00000" when "000100011101101", -- t[2285] = 0
      "00000" when "000100011101110", -- t[2286] = 0
      "00000" when "000100011101111", -- t[2287] = 0
      "00000" when "000100011110000", -- t[2288] = 0
      "00000" when "000100011110001", -- t[2289] = 0
      "00000" when "000100011110010", -- t[2290] = 0
      "00000" when "000100011110011", -- t[2291] = 0
      "00000" when "000100011110100", -- t[2292] = 0
      "00000" when "000100011110101", -- t[2293] = 0
      "00000" when "000100011110110", -- t[2294] = 0
      "00000" when "000100011110111", -- t[2295] = 0
      "00000" when "000100011111000", -- t[2296] = 0
      "00000" when "000100011111001", -- t[2297] = 0
      "00000" when "000100011111010", -- t[2298] = 0
      "00000" when "000100011111011", -- t[2299] = 0
      "00000" when "000100011111100", -- t[2300] = 0
      "00000" when "000100011111101", -- t[2301] = 0
      "00000" when "000100011111110", -- t[2302] = 0
      "00000" when "000100011111111", -- t[2303] = 0
      "00000" when "000100100000000", -- t[2304] = 0
      "00000" when "000100100000001", -- t[2305] = 0
      "00000" when "000100100000010", -- t[2306] = 0
      "00000" when "000100100000011", -- t[2307] = 0
      "00000" when "000100100000100", -- t[2308] = 0
      "00000" when "000100100000101", -- t[2309] = 0
      "00000" when "000100100000110", -- t[2310] = 0
      "00000" when "000100100000111", -- t[2311] = 0
      "00000" when "000100100001000", -- t[2312] = 0
      "00000" when "000100100001001", -- t[2313] = 0
      "00000" when "000100100001010", -- t[2314] = 0
      "00000" when "000100100001011", -- t[2315] = 0
      "00000" when "000100100001100", -- t[2316] = 0
      "00000" when "000100100001101", -- t[2317] = 0
      "00000" when "000100100001110", -- t[2318] = 0
      "00000" when "000100100001111", -- t[2319] = 0
      "00000" when "000100100010000", -- t[2320] = 0
      "00000" when "000100100010001", -- t[2321] = 0
      "00000" when "000100100010010", -- t[2322] = 0
      "00000" when "000100100010011", -- t[2323] = 0
      "00000" when "000100100010100", -- t[2324] = 0
      "00000" when "000100100010101", -- t[2325] = 0
      "00000" when "000100100010110", -- t[2326] = 0
      "00000" when "000100100010111", -- t[2327] = 0
      "00000" when "000100100011000", -- t[2328] = 0
      "00000" when "000100100011001", -- t[2329] = 0
      "00000" when "000100100011010", -- t[2330] = 0
      "00000" when "000100100011011", -- t[2331] = 0
      "00000" when "000100100011100", -- t[2332] = 0
      "00000" when "000100100011101", -- t[2333] = 0
      "00000" when "000100100011110", -- t[2334] = 0
      "00000" when "000100100011111", -- t[2335] = 0
      "00000" when "000100100100000", -- t[2336] = 0
      "00000" when "000100100100001", -- t[2337] = 0
      "00000" when "000100100100010", -- t[2338] = 0
      "00000" when "000100100100011", -- t[2339] = 0
      "00000" when "000100100100100", -- t[2340] = 0
      "00000" when "000100100100101", -- t[2341] = 0
      "00000" when "000100100100110", -- t[2342] = 0
      "00000" when "000100100100111", -- t[2343] = 0
      "00000" when "000100100101000", -- t[2344] = 0
      "00000" when "000100100101001", -- t[2345] = 0
      "00000" when "000100100101010", -- t[2346] = 0
      "00000" when "000100100101011", -- t[2347] = 0
      "00000" when "000100100101100", -- t[2348] = 0
      "00000" when "000100100101101", -- t[2349] = 0
      "00000" when "000100100101110", -- t[2350] = 0
      "00000" when "000100100101111", -- t[2351] = 0
      "00000" when "000100100110000", -- t[2352] = 0
      "00000" when "000100100110001", -- t[2353] = 0
      "00000" when "000100100110010", -- t[2354] = 0
      "00000" when "000100100110011", -- t[2355] = 0
      "00000" when "000100100110100", -- t[2356] = 0
      "00000" when "000100100110101", -- t[2357] = 0
      "00000" when "000100100110110", -- t[2358] = 0
      "00000" when "000100100110111", -- t[2359] = 0
      "00000" when "000100100111000", -- t[2360] = 0
      "00000" when "000100100111001", -- t[2361] = 0
      "00000" when "000100100111010", -- t[2362] = 0
      "00000" when "000100100111011", -- t[2363] = 0
      "00000" when "000100100111100", -- t[2364] = 0
      "00000" when "000100100111101", -- t[2365] = 0
      "00000" when "000100100111110", -- t[2366] = 0
      "00000" when "000100100111111", -- t[2367] = 0
      "00000" when "000100101000000", -- t[2368] = 0
      "00000" when "000100101000001", -- t[2369] = 0
      "00000" when "000100101000010", -- t[2370] = 0
      "00000" when "000100101000011", -- t[2371] = 0
      "00000" when "000100101000100", -- t[2372] = 0
      "00000" when "000100101000101", -- t[2373] = 0
      "00000" when "000100101000110", -- t[2374] = 0
      "00000" when "000100101000111", -- t[2375] = 0
      "00000" when "000100101001000", -- t[2376] = 0
      "00000" when "000100101001001", -- t[2377] = 0
      "00000" when "000100101001010", -- t[2378] = 0
      "00000" when "000100101001011", -- t[2379] = 0
      "00000" when "000100101001100", -- t[2380] = 0
      "00000" when "000100101001101", -- t[2381] = 0
      "00000" when "000100101001110", -- t[2382] = 0
      "00000" when "000100101001111", -- t[2383] = 0
      "00000" when "000100101010000", -- t[2384] = 0
      "00000" when "000100101010001", -- t[2385] = 0
      "00000" when "000100101010010", -- t[2386] = 0
      "00000" when "000100101010011", -- t[2387] = 0
      "00000" when "000100101010100", -- t[2388] = 0
      "00000" when "000100101010101", -- t[2389] = 0
      "00000" when "000100101010110", -- t[2390] = 0
      "00000" when "000100101010111", -- t[2391] = 0
      "00000" when "000100101011000", -- t[2392] = 0
      "00000" when "000100101011001", -- t[2393] = 0
      "00000" when "000100101011010", -- t[2394] = 0
      "00000" when "000100101011011", -- t[2395] = 0
      "00000" when "000100101011100", -- t[2396] = 0
      "00000" when "000100101011101", -- t[2397] = 0
      "00000" when "000100101011110", -- t[2398] = 0
      "00000" when "000100101011111", -- t[2399] = 0
      "00000" when "000100101100000", -- t[2400] = 0
      "00000" when "000100101100001", -- t[2401] = 0
      "00000" when "000100101100010", -- t[2402] = 0
      "00000" when "000100101100011", -- t[2403] = 0
      "00000" when "000100101100100", -- t[2404] = 0
      "00000" when "000100101100101", -- t[2405] = 0
      "00000" when "000100101100110", -- t[2406] = 0
      "00000" when "000100101100111", -- t[2407] = 0
      "00000" when "000100101101000", -- t[2408] = 0
      "00000" when "000100101101001", -- t[2409] = 0
      "00000" when "000100101101010", -- t[2410] = 0
      "00000" when "000100101101011", -- t[2411] = 0
      "00000" when "000100101101100", -- t[2412] = 0
      "00000" when "000100101101101", -- t[2413] = 0
      "00000" when "000100101101110", -- t[2414] = 0
      "00000" when "000100101101111", -- t[2415] = 0
      "00000" when "000100101110000", -- t[2416] = 0
      "00000" when "000100101110001", -- t[2417] = 0
      "00000" when "000100101110010", -- t[2418] = 0
      "00000" when "000100101110011", -- t[2419] = 0
      "00000" when "000100101110100", -- t[2420] = 0
      "00000" when "000100101110101", -- t[2421] = 0
      "00000" when "000100101110110", -- t[2422] = 0
      "00000" when "000100101110111", -- t[2423] = 0
      "00000" when "000100101111000", -- t[2424] = 0
      "00000" when "000100101111001", -- t[2425] = 0
      "00000" when "000100101111010", -- t[2426] = 0
      "00000" when "000100101111011", -- t[2427] = 0
      "00000" when "000100101111100", -- t[2428] = 0
      "00000" when "000100101111101", -- t[2429] = 0
      "00000" when "000100101111110", -- t[2430] = 0
      "00000" when "000100101111111", -- t[2431] = 0
      "00000" when "000100110000000", -- t[2432] = 0
      "00000" when "000100110000001", -- t[2433] = 0
      "00000" when "000100110000010", -- t[2434] = 0
      "00000" when "000100110000011", -- t[2435] = 0
      "00000" when "000100110000100", -- t[2436] = 0
      "00000" when "000100110000101", -- t[2437] = 0
      "00000" when "000100110000110", -- t[2438] = 0
      "00000" when "000100110000111", -- t[2439] = 0
      "00000" when "000100110001000", -- t[2440] = 0
      "00000" when "000100110001001", -- t[2441] = 0
      "00000" when "000100110001010", -- t[2442] = 0
      "00000" when "000100110001011", -- t[2443] = 0
      "00000" when "000100110001100", -- t[2444] = 0
      "00000" when "000100110001101", -- t[2445] = 0
      "00000" when "000100110001110", -- t[2446] = 0
      "00000" when "000100110001111", -- t[2447] = 0
      "00000" when "000100110010000", -- t[2448] = 0
      "00000" when "000100110010001", -- t[2449] = 0
      "00000" when "000100110010010", -- t[2450] = 0
      "00000" when "000100110010011", -- t[2451] = 0
      "00000" when "000100110010100", -- t[2452] = 0
      "00000" when "000100110010101", -- t[2453] = 0
      "00000" when "000100110010110", -- t[2454] = 0
      "00000" when "000100110010111", -- t[2455] = 0
      "00000" when "000100110011000", -- t[2456] = 0
      "00000" when "000100110011001", -- t[2457] = 0
      "00000" when "000100110011010", -- t[2458] = 0
      "00000" when "000100110011011", -- t[2459] = 0
      "00000" when "000100110011100", -- t[2460] = 0
      "00000" when "000100110011101", -- t[2461] = 0
      "00000" when "000100110011110", -- t[2462] = 0
      "00000" when "000100110011111", -- t[2463] = 0
      "00000" when "000100110100000", -- t[2464] = 0
      "00000" when "000100110100001", -- t[2465] = 0
      "00000" when "000100110100010", -- t[2466] = 0
      "00000" when "000100110100011", -- t[2467] = 0
      "00000" when "000100110100100", -- t[2468] = 0
      "00000" when "000100110100101", -- t[2469] = 0
      "00000" when "000100110100110", -- t[2470] = 0
      "00000" when "000100110100111", -- t[2471] = 0
      "00000" when "000100110101000", -- t[2472] = 0
      "00000" when "000100110101001", -- t[2473] = 0
      "00000" when "000100110101010", -- t[2474] = 0
      "00000" when "000100110101011", -- t[2475] = 0
      "00000" when "000100110101100", -- t[2476] = 0
      "00000" when "000100110101101", -- t[2477] = 0
      "00000" when "000100110101110", -- t[2478] = 0
      "00000" when "000100110101111", -- t[2479] = 0
      "00000" when "000100110110000", -- t[2480] = 0
      "00000" when "000100110110001", -- t[2481] = 0
      "00000" when "000100110110010", -- t[2482] = 0
      "00000" when "000100110110011", -- t[2483] = 0
      "00000" when "000100110110100", -- t[2484] = 0
      "00000" when "000100110110101", -- t[2485] = 0
      "00000" when "000100110110110", -- t[2486] = 0
      "00000" when "000100110110111", -- t[2487] = 0
      "00000" when "000100110111000", -- t[2488] = 0
      "00000" when "000100110111001", -- t[2489] = 0
      "00000" when "000100110111010", -- t[2490] = 0
      "00000" when "000100110111011", -- t[2491] = 0
      "00000" when "000100110111100", -- t[2492] = 0
      "00000" when "000100110111101", -- t[2493] = 0
      "00000" when "000100110111110", -- t[2494] = 0
      "00000" when "000100110111111", -- t[2495] = 0
      "00000" when "000100111000000", -- t[2496] = 0
      "00000" when "000100111000001", -- t[2497] = 0
      "00000" when "000100111000010", -- t[2498] = 0
      "00000" when "000100111000011", -- t[2499] = 0
      "00000" when "000100111000100", -- t[2500] = 0
      "00000" when "000100111000101", -- t[2501] = 0
      "00000" when "000100111000110", -- t[2502] = 0
      "00000" when "000100111000111", -- t[2503] = 0
      "00000" when "000100111001000", -- t[2504] = 0
      "00000" when "000100111001001", -- t[2505] = 0
      "00000" when "000100111001010", -- t[2506] = 0
      "00000" when "000100111001011", -- t[2507] = 0
      "00000" when "000100111001100", -- t[2508] = 0
      "00000" when "000100111001101", -- t[2509] = 0
      "00000" when "000100111001110", -- t[2510] = 0
      "00000" when "000100111001111", -- t[2511] = 0
      "00000" when "000100111010000", -- t[2512] = 0
      "00000" when "000100111010001", -- t[2513] = 0
      "00000" when "000100111010010", -- t[2514] = 0
      "00000" when "000100111010011", -- t[2515] = 0
      "00000" when "000100111010100", -- t[2516] = 0
      "00000" when "000100111010101", -- t[2517] = 0
      "00000" when "000100111010110", -- t[2518] = 0
      "00000" when "000100111010111", -- t[2519] = 0
      "00000" when "000100111011000", -- t[2520] = 0
      "00000" when "000100111011001", -- t[2521] = 0
      "00000" when "000100111011010", -- t[2522] = 0
      "00000" when "000100111011011", -- t[2523] = 0
      "00000" when "000100111011100", -- t[2524] = 0
      "00000" when "000100111011101", -- t[2525] = 0
      "00000" when "000100111011110", -- t[2526] = 0
      "00000" when "000100111011111", -- t[2527] = 0
      "00000" when "000100111100000", -- t[2528] = 0
      "00000" when "000100111100001", -- t[2529] = 0
      "00000" when "000100111100010", -- t[2530] = 0
      "00000" when "000100111100011", -- t[2531] = 0
      "00000" when "000100111100100", -- t[2532] = 0
      "00000" when "000100111100101", -- t[2533] = 0
      "00000" when "000100111100110", -- t[2534] = 0
      "00000" when "000100111100111", -- t[2535] = 0
      "00000" when "000100111101000", -- t[2536] = 0
      "00000" when "000100111101001", -- t[2537] = 0
      "00000" when "000100111101010", -- t[2538] = 0
      "00000" when "000100111101011", -- t[2539] = 0
      "00000" when "000100111101100", -- t[2540] = 0
      "00000" when "000100111101101", -- t[2541] = 0
      "00000" when "000100111101110", -- t[2542] = 0
      "00000" when "000100111101111", -- t[2543] = 0
      "00000" when "000100111110000", -- t[2544] = 0
      "00000" when "000100111110001", -- t[2545] = 0
      "00000" when "000100111110010", -- t[2546] = 0
      "00000" when "000100111110011", -- t[2547] = 0
      "00000" when "000100111110100", -- t[2548] = 0
      "00000" when "000100111110101", -- t[2549] = 0
      "00000" when "000100111110110", -- t[2550] = 0
      "00000" when "000100111110111", -- t[2551] = 0
      "00000" when "000100111111000", -- t[2552] = 0
      "00000" when "000100111111001", -- t[2553] = 0
      "00000" when "000100111111010", -- t[2554] = 0
      "00000" when "000100111111011", -- t[2555] = 0
      "00000" when "000100111111100", -- t[2556] = 0
      "00000" when "000100111111101", -- t[2557] = 0
      "00000" when "000100111111110", -- t[2558] = 0
      "00000" when "000100111111111", -- t[2559] = 0
      "00000" when "000101000000000", -- t[2560] = 0
      "00000" when "000101000000001", -- t[2561] = 0
      "00000" when "000101000000010", -- t[2562] = 0
      "00000" when "000101000000011", -- t[2563] = 0
      "00000" when "000101000000100", -- t[2564] = 0
      "00000" when "000101000000101", -- t[2565] = 0
      "00000" when "000101000000110", -- t[2566] = 0
      "00000" when "000101000000111", -- t[2567] = 0
      "00000" when "000101000001000", -- t[2568] = 0
      "00000" when "000101000001001", -- t[2569] = 0
      "00000" when "000101000001010", -- t[2570] = 0
      "00000" when "000101000001011", -- t[2571] = 0
      "00000" when "000101000001100", -- t[2572] = 0
      "00000" when "000101000001101", -- t[2573] = 0
      "00000" when "000101000001110", -- t[2574] = 0
      "00000" when "000101000001111", -- t[2575] = 0
      "00000" when "000101000010000", -- t[2576] = 0
      "00000" when "000101000010001", -- t[2577] = 0
      "00000" when "000101000010010", -- t[2578] = 0
      "00000" when "000101000010011", -- t[2579] = 0
      "00000" when "000101000010100", -- t[2580] = 0
      "00000" when "000101000010101", -- t[2581] = 0
      "00000" when "000101000010110", -- t[2582] = 0
      "00000" when "000101000010111", -- t[2583] = 0
      "00000" when "000101000011000", -- t[2584] = 0
      "00000" when "000101000011001", -- t[2585] = 0
      "00000" when "000101000011010", -- t[2586] = 0
      "00000" when "000101000011011", -- t[2587] = 0
      "00000" when "000101000011100", -- t[2588] = 0
      "00000" when "000101000011101", -- t[2589] = 0
      "00000" when "000101000011110", -- t[2590] = 0
      "00000" when "000101000011111", -- t[2591] = 0
      "00000" when "000101000100000", -- t[2592] = 0
      "00000" when "000101000100001", -- t[2593] = 0
      "00000" when "000101000100010", -- t[2594] = 0
      "00000" when "000101000100011", -- t[2595] = 0
      "00000" when "000101000100100", -- t[2596] = 0
      "00000" when "000101000100101", -- t[2597] = 0
      "00000" when "000101000100110", -- t[2598] = 0
      "00000" when "000101000100111", -- t[2599] = 0
      "00000" when "000101000101000", -- t[2600] = 0
      "00000" when "000101000101001", -- t[2601] = 0
      "00000" when "000101000101010", -- t[2602] = 0
      "00000" when "000101000101011", -- t[2603] = 0
      "00000" when "000101000101100", -- t[2604] = 0
      "00000" when "000101000101101", -- t[2605] = 0
      "00000" when "000101000101110", -- t[2606] = 0
      "00000" when "000101000101111", -- t[2607] = 0
      "00000" when "000101000110000", -- t[2608] = 0
      "00000" when "000101000110001", -- t[2609] = 0
      "00000" when "000101000110010", -- t[2610] = 0
      "00000" when "000101000110011", -- t[2611] = 0
      "00000" when "000101000110100", -- t[2612] = 0
      "00000" when "000101000110101", -- t[2613] = 0
      "00000" when "000101000110110", -- t[2614] = 0
      "00000" when "000101000110111", -- t[2615] = 0
      "00000" when "000101000111000", -- t[2616] = 0
      "00000" when "000101000111001", -- t[2617] = 0
      "00000" when "000101000111010", -- t[2618] = 0
      "00000" when "000101000111011", -- t[2619] = 0
      "00000" when "000101000111100", -- t[2620] = 0
      "00000" when "000101000111101", -- t[2621] = 0
      "00000" when "000101000111110", -- t[2622] = 0
      "00000" when "000101000111111", -- t[2623] = 0
      "00000" when "000101001000000", -- t[2624] = 0
      "00000" when "000101001000001", -- t[2625] = 0
      "00000" when "000101001000010", -- t[2626] = 0
      "00000" when "000101001000011", -- t[2627] = 0
      "00000" when "000101001000100", -- t[2628] = 0
      "00000" when "000101001000101", -- t[2629] = 0
      "00000" when "000101001000110", -- t[2630] = 0
      "00000" when "000101001000111", -- t[2631] = 0
      "00000" when "000101001001000", -- t[2632] = 0
      "00000" when "000101001001001", -- t[2633] = 0
      "00000" when "000101001001010", -- t[2634] = 0
      "00000" when "000101001001011", -- t[2635] = 0
      "00000" when "000101001001100", -- t[2636] = 0
      "00000" when "000101001001101", -- t[2637] = 0
      "00000" when "000101001001110", -- t[2638] = 0
      "00000" when "000101001001111", -- t[2639] = 0
      "00000" when "000101001010000", -- t[2640] = 0
      "00000" when "000101001010001", -- t[2641] = 0
      "00000" when "000101001010010", -- t[2642] = 0
      "00000" when "000101001010011", -- t[2643] = 0
      "00000" when "000101001010100", -- t[2644] = 0
      "00000" when "000101001010101", -- t[2645] = 0
      "00000" when "000101001010110", -- t[2646] = 0
      "00000" when "000101001010111", -- t[2647] = 0
      "00000" when "000101001011000", -- t[2648] = 0
      "00000" when "000101001011001", -- t[2649] = 0
      "00000" when "000101001011010", -- t[2650] = 0
      "00000" when "000101001011011", -- t[2651] = 0
      "00000" when "000101001011100", -- t[2652] = 0
      "00000" when "000101001011101", -- t[2653] = 0
      "00000" when "000101001011110", -- t[2654] = 0
      "00000" when "000101001011111", -- t[2655] = 0
      "00000" when "000101001100000", -- t[2656] = 0
      "00000" when "000101001100001", -- t[2657] = 0
      "00000" when "000101001100010", -- t[2658] = 0
      "00000" when "000101001100011", -- t[2659] = 0
      "00000" when "000101001100100", -- t[2660] = 0
      "00000" when "000101001100101", -- t[2661] = 0
      "00000" when "000101001100110", -- t[2662] = 0
      "00000" when "000101001100111", -- t[2663] = 0
      "00000" when "000101001101000", -- t[2664] = 0
      "00000" when "000101001101001", -- t[2665] = 0
      "00000" when "000101001101010", -- t[2666] = 0
      "00000" when "000101001101011", -- t[2667] = 0
      "00000" when "000101001101100", -- t[2668] = 0
      "00000" when "000101001101101", -- t[2669] = 0
      "00000" when "000101001101110", -- t[2670] = 0
      "00000" when "000101001101111", -- t[2671] = 0
      "00000" when "000101001110000", -- t[2672] = 0
      "00000" when "000101001110001", -- t[2673] = 0
      "00000" when "000101001110010", -- t[2674] = 0
      "00000" when "000101001110011", -- t[2675] = 0
      "00000" when "000101001110100", -- t[2676] = 0
      "00000" when "000101001110101", -- t[2677] = 0
      "00000" when "000101001110110", -- t[2678] = 0
      "00000" when "000101001110111", -- t[2679] = 0
      "00000" when "000101001111000", -- t[2680] = 0
      "00000" when "000101001111001", -- t[2681] = 0
      "00000" when "000101001111010", -- t[2682] = 0
      "00000" when "000101001111011", -- t[2683] = 0
      "00000" when "000101001111100", -- t[2684] = 0
      "00000" when "000101001111101", -- t[2685] = 0
      "00000" when "000101001111110", -- t[2686] = 0
      "00000" when "000101001111111", -- t[2687] = 0
      "00000" when "000101010000000", -- t[2688] = 0
      "00000" when "000101010000001", -- t[2689] = 0
      "00000" when "000101010000010", -- t[2690] = 0
      "00000" when "000101010000011", -- t[2691] = 0
      "00000" when "000101010000100", -- t[2692] = 0
      "00000" when "000101010000101", -- t[2693] = 0
      "00000" when "000101010000110", -- t[2694] = 0
      "00000" when "000101010000111", -- t[2695] = 0
      "00000" when "000101010001000", -- t[2696] = 0
      "00000" when "000101010001001", -- t[2697] = 0
      "00000" when "000101010001010", -- t[2698] = 0
      "00000" when "000101010001011", -- t[2699] = 0
      "00000" when "000101010001100", -- t[2700] = 0
      "00000" when "000101010001101", -- t[2701] = 0
      "00000" when "000101010001110", -- t[2702] = 0
      "00000" when "000101010001111", -- t[2703] = 0
      "00000" when "000101010010000", -- t[2704] = 0
      "00000" when "000101010010001", -- t[2705] = 0
      "00000" when "000101010010010", -- t[2706] = 0
      "00000" when "000101010010011", -- t[2707] = 0
      "00000" when "000101010010100", -- t[2708] = 0
      "00000" when "000101010010101", -- t[2709] = 0
      "00000" when "000101010010110", -- t[2710] = 0
      "00000" when "000101010010111", -- t[2711] = 0
      "00000" when "000101010011000", -- t[2712] = 0
      "00000" when "000101010011001", -- t[2713] = 0
      "00000" when "000101010011010", -- t[2714] = 0
      "00000" when "000101010011011", -- t[2715] = 0
      "00000" when "000101010011100", -- t[2716] = 0
      "00000" when "000101010011101", -- t[2717] = 0
      "00000" when "000101010011110", -- t[2718] = 0
      "00000" when "000101010011111", -- t[2719] = 0
      "00000" when "000101010100000", -- t[2720] = 0
      "00000" when "000101010100001", -- t[2721] = 0
      "00000" when "000101010100010", -- t[2722] = 0
      "00000" when "000101010100011", -- t[2723] = 0
      "00000" when "000101010100100", -- t[2724] = 0
      "00000" when "000101010100101", -- t[2725] = 0
      "00000" when "000101010100110", -- t[2726] = 0
      "00000" when "000101010100111", -- t[2727] = 0
      "00000" when "000101010101000", -- t[2728] = 0
      "00000" when "000101010101001", -- t[2729] = 0
      "00000" when "000101010101010", -- t[2730] = 0
      "00000" when "000101010101011", -- t[2731] = 0
      "00000" when "000101010101100", -- t[2732] = 0
      "00000" when "000101010101101", -- t[2733] = 0
      "00000" when "000101010101110", -- t[2734] = 0
      "00000" when "000101010101111", -- t[2735] = 0
      "00000" when "000101010110000", -- t[2736] = 0
      "00000" when "000101010110001", -- t[2737] = 0
      "00000" when "000101010110010", -- t[2738] = 0
      "00000" when "000101010110011", -- t[2739] = 0
      "00000" when "000101010110100", -- t[2740] = 0
      "00000" when "000101010110101", -- t[2741] = 0
      "00000" when "000101010110110", -- t[2742] = 0
      "00000" when "000101010110111", -- t[2743] = 0
      "00000" when "000101010111000", -- t[2744] = 0
      "00000" when "000101010111001", -- t[2745] = 0
      "00000" when "000101010111010", -- t[2746] = 0
      "00000" when "000101010111011", -- t[2747] = 0
      "00000" when "000101010111100", -- t[2748] = 0
      "00000" when "000101010111101", -- t[2749] = 0
      "00000" when "000101010111110", -- t[2750] = 0
      "00000" when "000101010111111", -- t[2751] = 0
      "00000" when "000101011000000", -- t[2752] = 0
      "00000" when "000101011000001", -- t[2753] = 0
      "00000" when "000101011000010", -- t[2754] = 0
      "00000" when "000101011000011", -- t[2755] = 0
      "00000" when "000101011000100", -- t[2756] = 0
      "00000" when "000101011000101", -- t[2757] = 0
      "00000" when "000101011000110", -- t[2758] = 0
      "00000" when "000101011000111", -- t[2759] = 0
      "00000" when "000101011001000", -- t[2760] = 0
      "00000" when "000101011001001", -- t[2761] = 0
      "00000" when "000101011001010", -- t[2762] = 0
      "00000" when "000101011001011", -- t[2763] = 0
      "00000" when "000101011001100", -- t[2764] = 0
      "00000" when "000101011001101", -- t[2765] = 0
      "00000" when "000101011001110", -- t[2766] = 0
      "00000" when "000101011001111", -- t[2767] = 0
      "00000" when "000101011010000", -- t[2768] = 0
      "00000" when "000101011010001", -- t[2769] = 0
      "00000" when "000101011010010", -- t[2770] = 0
      "00000" when "000101011010011", -- t[2771] = 0
      "00000" when "000101011010100", -- t[2772] = 0
      "00000" when "000101011010101", -- t[2773] = 0
      "00000" when "000101011010110", -- t[2774] = 0
      "00000" when "000101011010111", -- t[2775] = 0
      "00000" when "000101011011000", -- t[2776] = 0
      "00000" when "000101011011001", -- t[2777] = 0
      "00000" when "000101011011010", -- t[2778] = 0
      "00000" when "000101011011011", -- t[2779] = 0
      "00000" when "000101011011100", -- t[2780] = 0
      "00000" when "000101011011101", -- t[2781] = 0
      "00000" when "000101011011110", -- t[2782] = 0
      "00000" when "000101011011111", -- t[2783] = 0
      "00000" when "000101011100000", -- t[2784] = 0
      "00000" when "000101011100001", -- t[2785] = 0
      "00000" when "000101011100010", -- t[2786] = 0
      "00000" when "000101011100011", -- t[2787] = 0
      "00000" when "000101011100100", -- t[2788] = 0
      "00000" when "000101011100101", -- t[2789] = 0
      "00000" when "000101011100110", -- t[2790] = 0
      "00000" when "000101011100111", -- t[2791] = 0
      "00000" when "000101011101000", -- t[2792] = 0
      "00000" when "000101011101001", -- t[2793] = 0
      "00000" when "000101011101010", -- t[2794] = 0
      "00000" when "000101011101011", -- t[2795] = 0
      "00000" when "000101011101100", -- t[2796] = 0
      "00000" when "000101011101101", -- t[2797] = 0
      "00000" when "000101011101110", -- t[2798] = 0
      "00000" when "000101011101111", -- t[2799] = 0
      "00000" when "000101011110000", -- t[2800] = 0
      "00000" when "000101011110001", -- t[2801] = 0
      "00000" when "000101011110010", -- t[2802] = 0
      "00000" when "000101011110011", -- t[2803] = 0
      "00000" when "000101011110100", -- t[2804] = 0
      "00000" when "000101011110101", -- t[2805] = 0
      "00000" when "000101011110110", -- t[2806] = 0
      "00000" when "000101011110111", -- t[2807] = 0
      "00000" when "000101011111000", -- t[2808] = 0
      "00000" when "000101011111001", -- t[2809] = 0
      "00000" when "000101011111010", -- t[2810] = 0
      "00000" when "000101011111011", -- t[2811] = 0
      "00000" when "000101011111100", -- t[2812] = 0
      "00000" when "000101011111101", -- t[2813] = 0
      "00000" when "000101011111110", -- t[2814] = 0
      "00000" when "000101011111111", -- t[2815] = 0
      "00000" when "000101100000000", -- t[2816] = 0
      "00000" when "000101100000001", -- t[2817] = 0
      "00000" when "000101100000010", -- t[2818] = 0
      "00000" when "000101100000011", -- t[2819] = 0
      "00000" when "000101100000100", -- t[2820] = 0
      "00000" when "000101100000101", -- t[2821] = 0
      "00000" when "000101100000110", -- t[2822] = 0
      "00000" when "000101100000111", -- t[2823] = 0
      "00000" when "000101100001000", -- t[2824] = 0
      "00000" when "000101100001001", -- t[2825] = 0
      "00000" when "000101100001010", -- t[2826] = 0
      "00000" when "000101100001011", -- t[2827] = 0
      "00000" when "000101100001100", -- t[2828] = 0
      "00000" when "000101100001101", -- t[2829] = 0
      "00000" when "000101100001110", -- t[2830] = 0
      "00000" when "000101100001111", -- t[2831] = 0
      "00000" when "000101100010000", -- t[2832] = 0
      "00000" when "000101100010001", -- t[2833] = 0
      "00000" when "000101100010010", -- t[2834] = 0
      "00000" when "000101100010011", -- t[2835] = 0
      "00000" when "000101100010100", -- t[2836] = 0
      "00000" when "000101100010101", -- t[2837] = 0
      "00000" when "000101100010110", -- t[2838] = 0
      "00000" when "000101100010111", -- t[2839] = 0
      "00000" when "000101100011000", -- t[2840] = 0
      "00000" when "000101100011001", -- t[2841] = 0
      "00000" when "000101100011010", -- t[2842] = 0
      "00000" when "000101100011011", -- t[2843] = 0
      "00000" when "000101100011100", -- t[2844] = 0
      "00000" when "000101100011101", -- t[2845] = 0
      "00000" when "000101100011110", -- t[2846] = 0
      "00000" when "000101100011111", -- t[2847] = 0
      "00000" when "000101100100000", -- t[2848] = 0
      "00000" when "000101100100001", -- t[2849] = 0
      "00000" when "000101100100010", -- t[2850] = 0
      "00000" when "000101100100011", -- t[2851] = 0
      "00000" when "000101100100100", -- t[2852] = 0
      "00000" when "000101100100101", -- t[2853] = 0
      "00000" when "000101100100110", -- t[2854] = 0
      "00000" when "000101100100111", -- t[2855] = 0
      "00000" when "000101100101000", -- t[2856] = 0
      "00000" when "000101100101001", -- t[2857] = 0
      "00000" when "000101100101010", -- t[2858] = 0
      "00000" when "000101100101011", -- t[2859] = 0
      "00000" when "000101100101100", -- t[2860] = 0
      "00000" when "000101100101101", -- t[2861] = 0
      "00000" when "000101100101110", -- t[2862] = 0
      "00000" when "000101100101111", -- t[2863] = 0
      "00000" when "000101100110000", -- t[2864] = 0
      "00000" when "000101100110001", -- t[2865] = 0
      "00000" when "000101100110010", -- t[2866] = 0
      "00000" when "000101100110011", -- t[2867] = 0
      "00000" when "000101100110100", -- t[2868] = 0
      "00000" when "000101100110101", -- t[2869] = 0
      "00000" when "000101100110110", -- t[2870] = 0
      "00000" when "000101100110111", -- t[2871] = 0
      "00000" when "000101100111000", -- t[2872] = 0
      "00000" when "000101100111001", -- t[2873] = 0
      "00000" when "000101100111010", -- t[2874] = 0
      "00000" when "000101100111011", -- t[2875] = 0
      "00000" when "000101100111100", -- t[2876] = 0
      "00000" when "000101100111101", -- t[2877] = 0
      "00000" when "000101100111110", -- t[2878] = 0
      "00000" when "000101100111111", -- t[2879] = 0
      "00000" when "000101101000000", -- t[2880] = 0
      "00000" when "000101101000001", -- t[2881] = 0
      "00000" when "000101101000010", -- t[2882] = 0
      "00000" when "000101101000011", -- t[2883] = 0
      "00000" when "000101101000100", -- t[2884] = 0
      "00000" when "000101101000101", -- t[2885] = 0
      "00000" when "000101101000110", -- t[2886] = 0
      "00000" when "000101101000111", -- t[2887] = 0
      "00000" when "000101101001000", -- t[2888] = 0
      "00000" when "000101101001001", -- t[2889] = 0
      "00000" when "000101101001010", -- t[2890] = 0
      "00000" when "000101101001011", -- t[2891] = 0
      "00000" when "000101101001100", -- t[2892] = 0
      "00000" when "000101101001101", -- t[2893] = 0
      "00000" when "000101101001110", -- t[2894] = 0
      "00000" when "000101101001111", -- t[2895] = 0
      "00000" when "000101101010000", -- t[2896] = 0
      "00000" when "000101101010001", -- t[2897] = 0
      "00000" when "000101101010010", -- t[2898] = 0
      "00000" when "000101101010011", -- t[2899] = 0
      "00000" when "000101101010100", -- t[2900] = 0
      "00000" when "000101101010101", -- t[2901] = 0
      "00000" when "000101101010110", -- t[2902] = 0
      "00000" when "000101101010111", -- t[2903] = 0
      "00000" when "000101101011000", -- t[2904] = 0
      "00000" when "000101101011001", -- t[2905] = 0
      "00000" when "000101101011010", -- t[2906] = 0
      "00000" when "000101101011011", -- t[2907] = 0
      "00000" when "000101101011100", -- t[2908] = 0
      "00000" when "000101101011101", -- t[2909] = 0
      "00000" when "000101101011110", -- t[2910] = 0
      "00000" when "000101101011111", -- t[2911] = 0
      "00000" when "000101101100000", -- t[2912] = 0
      "00000" when "000101101100001", -- t[2913] = 0
      "00000" when "000101101100010", -- t[2914] = 0
      "00000" when "000101101100011", -- t[2915] = 0
      "00000" when "000101101100100", -- t[2916] = 0
      "00000" when "000101101100101", -- t[2917] = 0
      "00000" when "000101101100110", -- t[2918] = 0
      "00000" when "000101101100111", -- t[2919] = 0
      "00000" when "000101101101000", -- t[2920] = 0
      "00000" when "000101101101001", -- t[2921] = 0
      "00000" when "000101101101010", -- t[2922] = 0
      "00000" when "000101101101011", -- t[2923] = 0
      "00000" when "000101101101100", -- t[2924] = 0
      "00000" when "000101101101101", -- t[2925] = 0
      "00000" when "000101101101110", -- t[2926] = 0
      "00000" when "000101101101111", -- t[2927] = 0
      "00000" when "000101101110000", -- t[2928] = 0
      "00000" when "000101101110001", -- t[2929] = 0
      "00000" when "000101101110010", -- t[2930] = 0
      "00000" when "000101101110011", -- t[2931] = 0
      "00000" when "000101101110100", -- t[2932] = 0
      "00000" when "000101101110101", -- t[2933] = 0
      "00000" when "000101101110110", -- t[2934] = 0
      "00000" when "000101101110111", -- t[2935] = 0
      "00000" when "000101101111000", -- t[2936] = 0
      "00000" when "000101101111001", -- t[2937] = 0
      "00000" when "000101101111010", -- t[2938] = 0
      "00000" when "000101101111011", -- t[2939] = 0
      "00000" when "000101101111100", -- t[2940] = 0
      "00000" when "000101101111101", -- t[2941] = 0
      "00000" when "000101101111110", -- t[2942] = 0
      "00000" when "000101101111111", -- t[2943] = 0
      "00000" when "000101110000000", -- t[2944] = 0
      "00000" when "000101110000001", -- t[2945] = 0
      "00000" when "000101110000010", -- t[2946] = 0
      "00000" when "000101110000011", -- t[2947] = 0
      "00000" when "000101110000100", -- t[2948] = 0
      "00000" when "000101110000101", -- t[2949] = 0
      "00000" when "000101110000110", -- t[2950] = 0
      "00000" when "000101110000111", -- t[2951] = 0
      "00000" when "000101110001000", -- t[2952] = 0
      "00000" when "000101110001001", -- t[2953] = 0
      "00000" when "000101110001010", -- t[2954] = 0
      "00000" when "000101110001011", -- t[2955] = 0
      "00000" when "000101110001100", -- t[2956] = 0
      "00000" when "000101110001101", -- t[2957] = 0
      "00000" when "000101110001110", -- t[2958] = 0
      "00000" when "000101110001111", -- t[2959] = 0
      "00000" when "000101110010000", -- t[2960] = 0
      "00000" when "000101110010001", -- t[2961] = 0
      "00000" when "000101110010010", -- t[2962] = 0
      "00000" when "000101110010011", -- t[2963] = 0
      "00000" when "000101110010100", -- t[2964] = 0
      "00000" when "000101110010101", -- t[2965] = 0
      "00000" when "000101110010110", -- t[2966] = 0
      "00000" when "000101110010111", -- t[2967] = 0
      "00000" when "000101110011000", -- t[2968] = 0
      "00000" when "000101110011001", -- t[2969] = 0
      "00000" when "000101110011010", -- t[2970] = 0
      "00000" when "000101110011011", -- t[2971] = 0
      "00000" when "000101110011100", -- t[2972] = 0
      "00000" when "000101110011101", -- t[2973] = 0
      "00000" when "000101110011110", -- t[2974] = 0
      "00000" when "000101110011111", -- t[2975] = 0
      "00000" when "000101110100000", -- t[2976] = 0
      "00000" when "000101110100001", -- t[2977] = 0
      "00000" when "000101110100010", -- t[2978] = 0
      "00000" when "000101110100011", -- t[2979] = 0
      "00000" when "000101110100100", -- t[2980] = 0
      "00000" when "000101110100101", -- t[2981] = 0
      "00000" when "000101110100110", -- t[2982] = 0
      "00000" when "000101110100111", -- t[2983] = 0
      "00000" when "000101110101000", -- t[2984] = 0
      "00000" when "000101110101001", -- t[2985] = 0
      "00000" when "000101110101010", -- t[2986] = 0
      "00000" when "000101110101011", -- t[2987] = 0
      "00000" when "000101110101100", -- t[2988] = 0
      "00000" when "000101110101101", -- t[2989] = 0
      "00000" when "000101110101110", -- t[2990] = 0
      "00000" when "000101110101111", -- t[2991] = 0
      "00000" when "000101110110000", -- t[2992] = 0
      "00000" when "000101110110001", -- t[2993] = 0
      "00000" when "000101110110010", -- t[2994] = 0
      "00000" when "000101110110011", -- t[2995] = 0
      "00000" when "000101110110100", -- t[2996] = 0
      "00000" when "000101110110101", -- t[2997] = 0
      "00000" when "000101110110110", -- t[2998] = 0
      "00000" when "000101110110111", -- t[2999] = 0
      "00000" when "000101110111000", -- t[3000] = 0
      "00000" when "000101110111001", -- t[3001] = 0
      "00000" when "000101110111010", -- t[3002] = 0
      "00000" when "000101110111011", -- t[3003] = 0
      "00000" when "000101110111100", -- t[3004] = 0
      "00000" when "000101110111101", -- t[3005] = 0
      "00000" when "000101110111110", -- t[3006] = 0
      "00000" when "000101110111111", -- t[3007] = 0
      "00000" when "000101111000000", -- t[3008] = 0
      "00000" when "000101111000001", -- t[3009] = 0
      "00000" when "000101111000010", -- t[3010] = 0
      "00000" when "000101111000011", -- t[3011] = 0
      "00000" when "000101111000100", -- t[3012] = 0
      "00000" when "000101111000101", -- t[3013] = 0
      "00000" when "000101111000110", -- t[3014] = 0
      "00000" when "000101111000111", -- t[3015] = 0
      "00000" when "000101111001000", -- t[3016] = 0
      "00000" when "000101111001001", -- t[3017] = 0
      "00000" when "000101111001010", -- t[3018] = 0
      "00000" when "000101111001011", -- t[3019] = 0
      "00000" when "000101111001100", -- t[3020] = 0
      "00000" when "000101111001101", -- t[3021] = 0
      "00000" when "000101111001110", -- t[3022] = 0
      "00000" when "000101111001111", -- t[3023] = 0
      "00000" when "000101111010000", -- t[3024] = 0
      "00000" when "000101111010001", -- t[3025] = 0
      "00000" when "000101111010010", -- t[3026] = 0
      "00000" when "000101111010011", -- t[3027] = 0
      "00000" when "000101111010100", -- t[3028] = 0
      "00000" when "000101111010101", -- t[3029] = 0
      "00000" when "000101111010110", -- t[3030] = 0
      "00000" when "000101111010111", -- t[3031] = 0
      "00000" when "000101111011000", -- t[3032] = 0
      "00000" when "000101111011001", -- t[3033] = 0
      "00000" when "000101111011010", -- t[3034] = 0
      "00000" when "000101111011011", -- t[3035] = 0
      "00000" when "000101111011100", -- t[3036] = 0
      "00000" when "000101111011101", -- t[3037] = 0
      "00000" when "000101111011110", -- t[3038] = 0
      "00000" when "000101111011111", -- t[3039] = 0
      "00000" when "000101111100000", -- t[3040] = 0
      "00000" when "000101111100001", -- t[3041] = 0
      "00000" when "000101111100010", -- t[3042] = 0
      "00000" when "000101111100011", -- t[3043] = 0
      "00000" when "000101111100100", -- t[3044] = 0
      "00000" when "000101111100101", -- t[3045] = 0
      "00000" when "000101111100110", -- t[3046] = 0
      "00000" when "000101111100111", -- t[3047] = 0
      "00000" when "000101111101000", -- t[3048] = 0
      "00000" when "000101111101001", -- t[3049] = 0
      "00000" when "000101111101010", -- t[3050] = 0
      "00000" when "000101111101011", -- t[3051] = 0
      "00000" when "000101111101100", -- t[3052] = 0
      "00000" when "000101111101101", -- t[3053] = 0
      "00000" when "000101111101110", -- t[3054] = 0
      "00000" when "000101111101111", -- t[3055] = 0
      "00000" when "000101111110000", -- t[3056] = 0
      "00000" when "000101111110001", -- t[3057] = 0
      "00000" when "000101111110010", -- t[3058] = 0
      "00000" when "000101111110011", -- t[3059] = 0
      "00000" when "000101111110100", -- t[3060] = 0
      "00000" when "000101111110101", -- t[3061] = 0
      "00000" when "000101111110110", -- t[3062] = 0
      "00000" when "000101111110111", -- t[3063] = 0
      "00000" when "000101111111000", -- t[3064] = 0
      "00000" when "000101111111001", -- t[3065] = 0
      "00000" when "000101111111010", -- t[3066] = 0
      "00000" when "000101111111011", -- t[3067] = 0
      "00000" when "000101111111100", -- t[3068] = 0
      "00000" when "000101111111101", -- t[3069] = 0
      "00000" when "000101111111110", -- t[3070] = 0
      "00000" when "000101111111111", -- t[3071] = 0
      "00000" when "000110000000000", -- t[3072] = 0
      "00000" when "000110000000001", -- t[3073] = 0
      "00000" when "000110000000010", -- t[3074] = 0
      "00000" when "000110000000011", -- t[3075] = 0
      "00000" when "000110000000100", -- t[3076] = 0
      "00000" when "000110000000101", -- t[3077] = 0
      "00000" when "000110000000110", -- t[3078] = 0
      "00000" when "000110000000111", -- t[3079] = 0
      "00000" when "000110000001000", -- t[3080] = 0
      "00000" when "000110000001001", -- t[3081] = 0
      "00000" when "000110000001010", -- t[3082] = 0
      "00000" when "000110000001011", -- t[3083] = 0
      "00000" when "000110000001100", -- t[3084] = 0
      "00000" when "000110000001101", -- t[3085] = 0
      "00000" when "000110000001110", -- t[3086] = 0
      "00000" when "000110000001111", -- t[3087] = 0
      "00000" when "000110000010000", -- t[3088] = 0
      "00000" when "000110000010001", -- t[3089] = 0
      "00000" when "000110000010010", -- t[3090] = 0
      "00000" when "000110000010011", -- t[3091] = 0
      "00000" when "000110000010100", -- t[3092] = 0
      "00000" when "000110000010101", -- t[3093] = 0
      "00000" when "000110000010110", -- t[3094] = 0
      "00000" when "000110000010111", -- t[3095] = 0
      "00000" when "000110000011000", -- t[3096] = 0
      "00000" when "000110000011001", -- t[3097] = 0
      "00000" when "000110000011010", -- t[3098] = 0
      "00000" when "000110000011011", -- t[3099] = 0
      "00000" when "000110000011100", -- t[3100] = 0
      "00000" when "000110000011101", -- t[3101] = 0
      "00000" when "000110000011110", -- t[3102] = 0
      "00000" when "000110000011111", -- t[3103] = 0
      "00000" when "000110000100000", -- t[3104] = 0
      "00000" when "000110000100001", -- t[3105] = 0
      "00000" when "000110000100010", -- t[3106] = 0
      "00000" when "000110000100011", -- t[3107] = 0
      "00000" when "000110000100100", -- t[3108] = 0
      "00000" when "000110000100101", -- t[3109] = 0
      "00000" when "000110000100110", -- t[3110] = 0
      "00000" when "000110000100111", -- t[3111] = 0
      "00000" when "000110000101000", -- t[3112] = 0
      "00000" when "000110000101001", -- t[3113] = 0
      "00000" when "000110000101010", -- t[3114] = 0
      "00000" when "000110000101011", -- t[3115] = 0
      "00000" when "000110000101100", -- t[3116] = 0
      "00000" when "000110000101101", -- t[3117] = 0
      "00000" when "000110000101110", -- t[3118] = 0
      "00000" when "000110000101111", -- t[3119] = 0
      "00000" when "000110000110000", -- t[3120] = 0
      "00000" when "000110000110001", -- t[3121] = 0
      "00000" when "000110000110010", -- t[3122] = 0
      "00000" when "000110000110011", -- t[3123] = 0
      "00000" when "000110000110100", -- t[3124] = 0
      "00000" when "000110000110101", -- t[3125] = 0
      "00000" when "000110000110110", -- t[3126] = 0
      "00000" when "000110000110111", -- t[3127] = 0
      "00000" when "000110000111000", -- t[3128] = 0
      "00000" when "000110000111001", -- t[3129] = 0
      "00000" when "000110000111010", -- t[3130] = 0
      "00000" when "000110000111011", -- t[3131] = 0
      "00000" when "000110000111100", -- t[3132] = 0
      "00000" when "000110000111101", -- t[3133] = 0
      "00000" when "000110000111110", -- t[3134] = 0
      "00000" when "000110000111111", -- t[3135] = 0
      "00000" when "000110001000000", -- t[3136] = 0
      "00000" when "000110001000001", -- t[3137] = 0
      "00000" when "000110001000010", -- t[3138] = 0
      "00000" when "000110001000011", -- t[3139] = 0
      "00000" when "000110001000100", -- t[3140] = 0
      "00000" when "000110001000101", -- t[3141] = 0
      "00000" when "000110001000110", -- t[3142] = 0
      "00000" when "000110001000111", -- t[3143] = 0
      "00000" when "000110001001000", -- t[3144] = 0
      "00000" when "000110001001001", -- t[3145] = 0
      "00000" when "000110001001010", -- t[3146] = 0
      "00000" when "000110001001011", -- t[3147] = 0
      "00000" when "000110001001100", -- t[3148] = 0
      "00000" when "000110001001101", -- t[3149] = 0
      "00000" when "000110001001110", -- t[3150] = 0
      "00000" when "000110001001111", -- t[3151] = 0
      "00000" when "000110001010000", -- t[3152] = 0
      "00000" when "000110001010001", -- t[3153] = 0
      "00000" when "000110001010010", -- t[3154] = 0
      "00000" when "000110001010011", -- t[3155] = 0
      "00000" when "000110001010100", -- t[3156] = 0
      "00000" when "000110001010101", -- t[3157] = 0
      "00000" when "000110001010110", -- t[3158] = 0
      "00000" when "000110001010111", -- t[3159] = 0
      "00000" when "000110001011000", -- t[3160] = 0
      "00000" when "000110001011001", -- t[3161] = 0
      "00000" when "000110001011010", -- t[3162] = 0
      "00000" when "000110001011011", -- t[3163] = 0
      "00000" when "000110001011100", -- t[3164] = 0
      "00000" when "000110001011101", -- t[3165] = 0
      "00000" when "000110001011110", -- t[3166] = 0
      "00000" when "000110001011111", -- t[3167] = 0
      "00000" when "000110001100000", -- t[3168] = 0
      "00000" when "000110001100001", -- t[3169] = 0
      "00000" when "000110001100010", -- t[3170] = 0
      "00000" when "000110001100011", -- t[3171] = 0
      "00000" when "000110001100100", -- t[3172] = 0
      "00000" when "000110001100101", -- t[3173] = 0
      "00000" when "000110001100110", -- t[3174] = 0
      "00000" when "000110001100111", -- t[3175] = 0
      "00000" when "000110001101000", -- t[3176] = 0
      "00000" when "000110001101001", -- t[3177] = 0
      "00000" when "000110001101010", -- t[3178] = 0
      "00000" when "000110001101011", -- t[3179] = 0
      "00000" when "000110001101100", -- t[3180] = 0
      "00000" when "000110001101101", -- t[3181] = 0
      "00000" when "000110001101110", -- t[3182] = 0
      "00000" when "000110001101111", -- t[3183] = 0
      "00000" when "000110001110000", -- t[3184] = 0
      "00000" when "000110001110001", -- t[3185] = 0
      "00000" when "000110001110010", -- t[3186] = 0
      "00000" when "000110001110011", -- t[3187] = 0
      "00000" when "000110001110100", -- t[3188] = 0
      "00000" when "000110001110101", -- t[3189] = 0
      "00000" when "000110001110110", -- t[3190] = 0
      "00000" when "000110001110111", -- t[3191] = 0
      "00000" when "000110001111000", -- t[3192] = 0
      "00000" when "000110001111001", -- t[3193] = 0
      "00000" when "000110001111010", -- t[3194] = 0
      "00000" when "000110001111011", -- t[3195] = 0
      "00000" when "000110001111100", -- t[3196] = 0
      "00000" when "000110001111101", -- t[3197] = 0
      "00000" when "000110001111110", -- t[3198] = 0
      "00000" when "000110001111111", -- t[3199] = 0
      "00000" when "000110010000000", -- t[3200] = 0
      "00000" when "000110010000001", -- t[3201] = 0
      "00000" when "000110010000010", -- t[3202] = 0
      "00000" when "000110010000011", -- t[3203] = 0
      "00000" when "000110010000100", -- t[3204] = 0
      "00000" when "000110010000101", -- t[3205] = 0
      "00000" when "000110010000110", -- t[3206] = 0
      "00000" when "000110010000111", -- t[3207] = 0
      "00000" when "000110010001000", -- t[3208] = 0
      "00000" when "000110010001001", -- t[3209] = 0
      "00000" when "000110010001010", -- t[3210] = 0
      "00000" when "000110010001011", -- t[3211] = 0
      "00000" when "000110010001100", -- t[3212] = 0
      "00000" when "000110010001101", -- t[3213] = 0
      "00000" when "000110010001110", -- t[3214] = 0
      "00000" when "000110010001111", -- t[3215] = 0
      "00000" when "000110010010000", -- t[3216] = 0
      "00000" when "000110010010001", -- t[3217] = 0
      "00000" when "000110010010010", -- t[3218] = 0
      "00000" when "000110010010011", -- t[3219] = 0
      "00000" when "000110010010100", -- t[3220] = 0
      "00000" when "000110010010101", -- t[3221] = 0
      "00000" when "000110010010110", -- t[3222] = 0
      "00000" when "000110010010111", -- t[3223] = 0
      "00000" when "000110010011000", -- t[3224] = 0
      "00000" when "000110010011001", -- t[3225] = 0
      "00000" when "000110010011010", -- t[3226] = 0
      "00000" when "000110010011011", -- t[3227] = 0
      "00000" when "000110010011100", -- t[3228] = 0
      "00000" when "000110010011101", -- t[3229] = 0
      "00000" when "000110010011110", -- t[3230] = 0
      "00000" when "000110010011111", -- t[3231] = 0
      "00000" when "000110010100000", -- t[3232] = 0
      "00000" when "000110010100001", -- t[3233] = 0
      "00000" when "000110010100010", -- t[3234] = 0
      "00000" when "000110010100011", -- t[3235] = 0
      "00000" when "000110010100100", -- t[3236] = 0
      "00000" when "000110010100101", -- t[3237] = 0
      "00000" when "000110010100110", -- t[3238] = 0
      "00000" when "000110010100111", -- t[3239] = 0
      "00000" when "000110010101000", -- t[3240] = 0
      "00000" when "000110010101001", -- t[3241] = 0
      "00000" when "000110010101010", -- t[3242] = 0
      "00000" when "000110010101011", -- t[3243] = 0
      "00000" when "000110010101100", -- t[3244] = 0
      "00000" when "000110010101101", -- t[3245] = 0
      "00000" when "000110010101110", -- t[3246] = 0
      "00000" when "000110010101111", -- t[3247] = 0
      "00000" when "000110010110000", -- t[3248] = 0
      "00000" when "000110010110001", -- t[3249] = 0
      "00000" when "000110010110010", -- t[3250] = 0
      "00000" when "000110010110011", -- t[3251] = 0
      "00000" when "000110010110100", -- t[3252] = 0
      "00000" when "000110010110101", -- t[3253] = 0
      "00000" when "000110010110110", -- t[3254] = 0
      "00000" when "000110010110111", -- t[3255] = 0
      "00000" when "000110010111000", -- t[3256] = 0
      "00000" when "000110010111001", -- t[3257] = 0
      "00000" when "000110010111010", -- t[3258] = 0
      "00000" when "000110010111011", -- t[3259] = 0
      "00000" when "000110010111100", -- t[3260] = 0
      "00000" when "000110010111101", -- t[3261] = 0
      "00000" when "000110010111110", -- t[3262] = 0
      "00000" when "000110010111111", -- t[3263] = 0
      "00000" when "000110011000000", -- t[3264] = 0
      "00000" when "000110011000001", -- t[3265] = 0
      "00000" when "000110011000010", -- t[3266] = 0
      "00000" when "000110011000011", -- t[3267] = 0
      "00000" when "000110011000100", -- t[3268] = 0
      "00000" when "000110011000101", -- t[3269] = 0
      "00000" when "000110011000110", -- t[3270] = 0
      "00000" when "000110011000111", -- t[3271] = 0
      "00000" when "000110011001000", -- t[3272] = 0
      "00000" when "000110011001001", -- t[3273] = 0
      "00000" when "000110011001010", -- t[3274] = 0
      "00000" when "000110011001011", -- t[3275] = 0
      "00000" when "000110011001100", -- t[3276] = 0
      "00000" when "000110011001101", -- t[3277] = 0
      "00000" when "000110011001110", -- t[3278] = 0
      "00000" when "000110011001111", -- t[3279] = 0
      "00000" when "000110011010000", -- t[3280] = 0
      "00000" when "000110011010001", -- t[3281] = 0
      "00000" when "000110011010010", -- t[3282] = 0
      "00000" when "000110011010011", -- t[3283] = 0
      "00000" when "000110011010100", -- t[3284] = 0
      "00000" when "000110011010101", -- t[3285] = 0
      "00000" when "000110011010110", -- t[3286] = 0
      "00000" when "000110011010111", -- t[3287] = 0
      "00000" when "000110011011000", -- t[3288] = 0
      "00000" when "000110011011001", -- t[3289] = 0
      "00000" when "000110011011010", -- t[3290] = 0
      "00000" when "000110011011011", -- t[3291] = 0
      "00000" when "000110011011100", -- t[3292] = 0
      "00000" when "000110011011101", -- t[3293] = 0
      "00000" when "000110011011110", -- t[3294] = 0
      "00000" when "000110011011111", -- t[3295] = 0
      "00000" when "000110011100000", -- t[3296] = 0
      "00000" when "000110011100001", -- t[3297] = 0
      "00000" when "000110011100010", -- t[3298] = 0
      "00000" when "000110011100011", -- t[3299] = 0
      "00000" when "000110011100100", -- t[3300] = 0
      "00000" when "000110011100101", -- t[3301] = 0
      "00000" when "000110011100110", -- t[3302] = 0
      "00000" when "000110011100111", -- t[3303] = 0
      "00000" when "000110011101000", -- t[3304] = 0
      "00000" when "000110011101001", -- t[3305] = 0
      "00000" when "000110011101010", -- t[3306] = 0
      "00000" when "000110011101011", -- t[3307] = 0
      "00000" when "000110011101100", -- t[3308] = 0
      "00000" when "000110011101101", -- t[3309] = 0
      "00000" when "000110011101110", -- t[3310] = 0
      "00000" when "000110011101111", -- t[3311] = 0
      "00000" when "000110011110000", -- t[3312] = 0
      "00000" when "000110011110001", -- t[3313] = 0
      "00000" when "000110011110010", -- t[3314] = 0
      "00000" when "000110011110011", -- t[3315] = 0
      "00000" when "000110011110100", -- t[3316] = 0
      "00000" when "000110011110101", -- t[3317] = 0
      "00000" when "000110011110110", -- t[3318] = 0
      "00000" when "000110011110111", -- t[3319] = 0
      "00000" when "000110011111000", -- t[3320] = 0
      "00000" when "000110011111001", -- t[3321] = 0
      "00000" when "000110011111010", -- t[3322] = 0
      "00000" when "000110011111011", -- t[3323] = 0
      "00000" when "000110011111100", -- t[3324] = 0
      "00000" when "000110011111101", -- t[3325] = 0
      "00000" when "000110011111110", -- t[3326] = 0
      "00000" when "000110011111111", -- t[3327] = 0
      "00000" when "000110100000000", -- t[3328] = 0
      "00000" when "000110100000001", -- t[3329] = 0
      "00000" when "000110100000010", -- t[3330] = 0
      "00000" when "000110100000011", -- t[3331] = 0
      "00000" when "000110100000100", -- t[3332] = 0
      "00000" when "000110100000101", -- t[3333] = 0
      "00000" when "000110100000110", -- t[3334] = 0
      "00000" when "000110100000111", -- t[3335] = 0
      "00000" when "000110100001000", -- t[3336] = 0
      "00000" when "000110100001001", -- t[3337] = 0
      "00000" when "000110100001010", -- t[3338] = 0
      "00000" when "000110100001011", -- t[3339] = 0
      "00000" when "000110100001100", -- t[3340] = 0
      "00000" when "000110100001101", -- t[3341] = 0
      "00000" when "000110100001110", -- t[3342] = 0
      "00000" when "000110100001111", -- t[3343] = 0
      "00000" when "000110100010000", -- t[3344] = 0
      "00000" when "000110100010001", -- t[3345] = 0
      "00000" when "000110100010010", -- t[3346] = 0
      "00000" when "000110100010011", -- t[3347] = 0
      "00000" when "000110100010100", -- t[3348] = 0
      "00000" when "000110100010101", -- t[3349] = 0
      "00000" when "000110100010110", -- t[3350] = 0
      "00000" when "000110100010111", -- t[3351] = 0
      "00000" when "000110100011000", -- t[3352] = 0
      "00000" when "000110100011001", -- t[3353] = 0
      "00000" when "000110100011010", -- t[3354] = 0
      "00000" when "000110100011011", -- t[3355] = 0
      "00000" when "000110100011100", -- t[3356] = 0
      "00000" when "000110100011101", -- t[3357] = 0
      "00000" when "000110100011110", -- t[3358] = 0
      "00000" when "000110100011111", -- t[3359] = 0
      "00000" when "000110100100000", -- t[3360] = 0
      "00000" when "000110100100001", -- t[3361] = 0
      "00000" when "000110100100010", -- t[3362] = 0
      "00000" when "000110100100011", -- t[3363] = 0
      "00000" when "000110100100100", -- t[3364] = 0
      "00000" when "000110100100101", -- t[3365] = 0
      "00000" when "000110100100110", -- t[3366] = 0
      "00000" when "000110100100111", -- t[3367] = 0
      "00000" when "000110100101000", -- t[3368] = 0
      "00000" when "000110100101001", -- t[3369] = 0
      "00000" when "000110100101010", -- t[3370] = 0
      "00000" when "000110100101011", -- t[3371] = 0
      "00000" when "000110100101100", -- t[3372] = 0
      "00000" when "000110100101101", -- t[3373] = 0
      "00000" when "000110100101110", -- t[3374] = 0
      "00000" when "000110100101111", -- t[3375] = 0
      "00000" when "000110100110000", -- t[3376] = 0
      "00000" when "000110100110001", -- t[3377] = 0
      "00000" when "000110100110010", -- t[3378] = 0
      "00000" when "000110100110011", -- t[3379] = 0
      "00000" when "000110100110100", -- t[3380] = 0
      "00000" when "000110100110101", -- t[3381] = 0
      "00000" when "000110100110110", -- t[3382] = 0
      "00000" when "000110100110111", -- t[3383] = 0
      "00000" when "000110100111000", -- t[3384] = 0
      "00000" when "000110100111001", -- t[3385] = 0
      "00000" when "000110100111010", -- t[3386] = 0
      "00000" when "000110100111011", -- t[3387] = 0
      "00000" when "000110100111100", -- t[3388] = 0
      "00000" when "000110100111101", -- t[3389] = 0
      "00000" when "000110100111110", -- t[3390] = 0
      "00000" when "000110100111111", -- t[3391] = 0
      "00000" when "000110101000000", -- t[3392] = 0
      "00000" when "000110101000001", -- t[3393] = 0
      "00000" when "000110101000010", -- t[3394] = 0
      "00000" when "000110101000011", -- t[3395] = 0
      "00000" when "000110101000100", -- t[3396] = 0
      "00000" when "000110101000101", -- t[3397] = 0
      "00000" when "000110101000110", -- t[3398] = 0
      "00000" when "000110101000111", -- t[3399] = 0
      "00000" when "000110101001000", -- t[3400] = 0
      "00000" when "000110101001001", -- t[3401] = 0
      "00000" when "000110101001010", -- t[3402] = 0
      "00000" when "000110101001011", -- t[3403] = 0
      "00000" when "000110101001100", -- t[3404] = 0
      "00000" when "000110101001101", -- t[3405] = 0
      "00000" when "000110101001110", -- t[3406] = 0
      "00000" when "000110101001111", -- t[3407] = 0
      "00000" when "000110101010000", -- t[3408] = 0
      "00000" when "000110101010001", -- t[3409] = 0
      "00000" when "000110101010010", -- t[3410] = 0
      "00000" when "000110101010011", -- t[3411] = 0
      "00000" when "000110101010100", -- t[3412] = 0
      "00000" when "000110101010101", -- t[3413] = 0
      "00000" when "000110101010110", -- t[3414] = 0
      "00000" when "000110101010111", -- t[3415] = 0
      "00000" when "000110101011000", -- t[3416] = 0
      "00000" when "000110101011001", -- t[3417] = 0
      "00000" when "000110101011010", -- t[3418] = 0
      "00000" when "000110101011011", -- t[3419] = 0
      "00000" when "000110101011100", -- t[3420] = 0
      "00000" when "000110101011101", -- t[3421] = 0
      "00000" when "000110101011110", -- t[3422] = 0
      "00000" when "000110101011111", -- t[3423] = 0
      "00000" when "000110101100000", -- t[3424] = 0
      "00000" when "000110101100001", -- t[3425] = 0
      "00000" when "000110101100010", -- t[3426] = 0
      "00000" when "000110101100011", -- t[3427] = 0
      "00000" when "000110101100100", -- t[3428] = 0
      "00000" when "000110101100101", -- t[3429] = 0
      "00000" when "000110101100110", -- t[3430] = 0
      "00000" when "000110101100111", -- t[3431] = 0
      "00000" when "000110101101000", -- t[3432] = 0
      "00000" when "000110101101001", -- t[3433] = 0
      "00000" when "000110101101010", -- t[3434] = 0
      "00000" when "000110101101011", -- t[3435] = 0
      "00000" when "000110101101100", -- t[3436] = 0
      "00000" when "000110101101101", -- t[3437] = 0
      "00000" when "000110101101110", -- t[3438] = 0
      "00000" when "000110101101111", -- t[3439] = 0
      "00000" when "000110101110000", -- t[3440] = 0
      "00000" when "000110101110001", -- t[3441] = 0
      "00000" when "000110101110010", -- t[3442] = 0
      "00000" when "000110101110011", -- t[3443] = 0
      "00000" when "000110101110100", -- t[3444] = 0
      "00000" when "000110101110101", -- t[3445] = 0
      "00000" when "000110101110110", -- t[3446] = 0
      "00000" when "000110101110111", -- t[3447] = 0
      "00000" when "000110101111000", -- t[3448] = 0
      "00000" when "000110101111001", -- t[3449] = 0
      "00000" when "000110101111010", -- t[3450] = 0
      "00000" when "000110101111011", -- t[3451] = 0
      "00000" when "000110101111100", -- t[3452] = 0
      "00000" when "000110101111101", -- t[3453] = 0
      "00000" when "000110101111110", -- t[3454] = 0
      "00000" when "000110101111111", -- t[3455] = 0
      "00000" when "000110110000000", -- t[3456] = 0
      "00000" when "000110110000001", -- t[3457] = 0
      "00000" when "000110110000010", -- t[3458] = 0
      "00000" when "000110110000011", -- t[3459] = 0
      "00000" when "000110110000100", -- t[3460] = 0
      "00000" when "000110110000101", -- t[3461] = 0
      "00000" when "000110110000110", -- t[3462] = 0
      "00000" when "000110110000111", -- t[3463] = 0
      "00000" when "000110110001000", -- t[3464] = 0
      "00000" when "000110110001001", -- t[3465] = 0
      "00000" when "000110110001010", -- t[3466] = 0
      "00000" when "000110110001011", -- t[3467] = 0
      "00000" when "000110110001100", -- t[3468] = 0
      "00000" when "000110110001101", -- t[3469] = 0
      "00000" when "000110110001110", -- t[3470] = 0
      "00000" when "000110110001111", -- t[3471] = 0
      "00000" when "000110110010000", -- t[3472] = 0
      "00000" when "000110110010001", -- t[3473] = 0
      "00000" when "000110110010010", -- t[3474] = 0
      "00000" when "000110110010011", -- t[3475] = 0
      "00000" when "000110110010100", -- t[3476] = 0
      "00000" when "000110110010101", -- t[3477] = 0
      "00000" when "000110110010110", -- t[3478] = 0
      "00000" when "000110110010111", -- t[3479] = 0
      "00000" when "000110110011000", -- t[3480] = 0
      "00000" when "000110110011001", -- t[3481] = 0
      "00000" when "000110110011010", -- t[3482] = 0
      "00000" when "000110110011011", -- t[3483] = 0
      "00000" when "000110110011100", -- t[3484] = 0
      "00000" when "000110110011101", -- t[3485] = 0
      "00000" when "000110110011110", -- t[3486] = 0
      "00000" when "000110110011111", -- t[3487] = 0
      "00000" when "000110110100000", -- t[3488] = 0
      "00000" when "000110110100001", -- t[3489] = 0
      "00000" when "000110110100010", -- t[3490] = 0
      "00000" when "000110110100011", -- t[3491] = 0
      "00000" when "000110110100100", -- t[3492] = 0
      "00000" when "000110110100101", -- t[3493] = 0
      "00000" when "000110110100110", -- t[3494] = 0
      "00000" when "000110110100111", -- t[3495] = 0
      "00000" when "000110110101000", -- t[3496] = 0
      "00000" when "000110110101001", -- t[3497] = 0
      "00000" when "000110110101010", -- t[3498] = 0
      "00000" when "000110110101011", -- t[3499] = 0
      "00000" when "000110110101100", -- t[3500] = 0
      "00000" when "000110110101101", -- t[3501] = 0
      "00000" when "000110110101110", -- t[3502] = 0
      "00000" when "000110110101111", -- t[3503] = 0
      "00000" when "000110110110000", -- t[3504] = 0
      "00000" when "000110110110001", -- t[3505] = 0
      "00000" when "000110110110010", -- t[3506] = 0
      "00000" when "000110110110011", -- t[3507] = 0
      "00000" when "000110110110100", -- t[3508] = 0
      "00000" when "000110110110101", -- t[3509] = 0
      "00000" when "000110110110110", -- t[3510] = 0
      "00000" when "000110110110111", -- t[3511] = 0
      "00000" when "000110110111000", -- t[3512] = 0
      "00000" when "000110110111001", -- t[3513] = 0
      "00000" when "000110110111010", -- t[3514] = 0
      "00000" when "000110110111011", -- t[3515] = 0
      "00000" when "000110110111100", -- t[3516] = 0
      "00000" when "000110110111101", -- t[3517] = 0
      "00000" when "000110110111110", -- t[3518] = 0
      "00000" when "000110110111111", -- t[3519] = 0
      "00000" when "000110111000000", -- t[3520] = 0
      "00000" when "000110111000001", -- t[3521] = 0
      "00000" when "000110111000010", -- t[3522] = 0
      "00000" when "000110111000011", -- t[3523] = 0
      "00000" when "000110111000100", -- t[3524] = 0
      "00000" when "000110111000101", -- t[3525] = 0
      "00000" when "000110111000110", -- t[3526] = 0
      "00000" when "000110111000111", -- t[3527] = 0
      "00000" when "000110111001000", -- t[3528] = 0
      "00000" when "000110111001001", -- t[3529] = 0
      "00000" when "000110111001010", -- t[3530] = 0
      "00000" when "000110111001011", -- t[3531] = 0
      "00000" when "000110111001100", -- t[3532] = 0
      "00000" when "000110111001101", -- t[3533] = 0
      "00000" when "000110111001110", -- t[3534] = 0
      "00000" when "000110111001111", -- t[3535] = 0
      "00000" when "000110111010000", -- t[3536] = 0
      "00000" when "000110111010001", -- t[3537] = 0
      "00000" when "000110111010010", -- t[3538] = 0
      "00000" when "000110111010011", -- t[3539] = 0
      "00000" when "000110111010100", -- t[3540] = 0
      "00000" when "000110111010101", -- t[3541] = 0
      "00000" when "000110111010110", -- t[3542] = 0
      "00000" when "000110111010111", -- t[3543] = 0
      "00000" when "000110111011000", -- t[3544] = 0
      "00000" when "000110111011001", -- t[3545] = 0
      "00000" when "000110111011010", -- t[3546] = 0
      "00000" when "000110111011011", -- t[3547] = 0
      "00000" when "000110111011100", -- t[3548] = 0
      "00000" when "000110111011101", -- t[3549] = 0
      "00000" when "000110111011110", -- t[3550] = 0
      "00000" when "000110111011111", -- t[3551] = 0
      "00000" when "000110111100000", -- t[3552] = 0
      "00000" when "000110111100001", -- t[3553] = 0
      "00000" when "000110111100010", -- t[3554] = 0
      "00000" when "000110111100011", -- t[3555] = 0
      "00000" when "000110111100100", -- t[3556] = 0
      "00000" when "000110111100101", -- t[3557] = 0
      "00000" when "000110111100110", -- t[3558] = 0
      "00000" when "000110111100111", -- t[3559] = 0
      "00000" when "000110111101000", -- t[3560] = 0
      "00000" when "000110111101001", -- t[3561] = 0
      "00000" when "000110111101010", -- t[3562] = 0
      "00000" when "000110111101011", -- t[3563] = 0
      "00000" when "000110111101100", -- t[3564] = 0
      "00000" when "000110111101101", -- t[3565] = 0
      "00000" when "000110111101110", -- t[3566] = 0
      "00000" when "000110111101111", -- t[3567] = 0
      "00000" when "000110111110000", -- t[3568] = 0
      "00000" when "000110111110001", -- t[3569] = 0
      "00000" when "000110111110010", -- t[3570] = 0
      "00000" when "000110111110011", -- t[3571] = 0
      "00000" when "000110111110100", -- t[3572] = 0
      "00000" when "000110111110101", -- t[3573] = 0
      "00000" when "000110111110110", -- t[3574] = 0
      "00000" when "000110111110111", -- t[3575] = 0
      "00000" when "000110111111000", -- t[3576] = 0
      "00000" when "000110111111001", -- t[3577] = 0
      "00000" when "000110111111010", -- t[3578] = 0
      "00000" when "000110111111011", -- t[3579] = 0
      "00000" when "000110111111100", -- t[3580] = 0
      "00000" when "000110111111101", -- t[3581] = 0
      "00000" when "000110111111110", -- t[3582] = 0
      "00000" when "000110111111111", -- t[3583] = 0
      "00000" when "000111000000000", -- t[3584] = 0
      "00000" when "000111000000001", -- t[3585] = 0
      "00000" when "000111000000010", -- t[3586] = 0
      "00000" when "000111000000011", -- t[3587] = 0
      "00000" when "000111000000100", -- t[3588] = 0
      "00000" when "000111000000101", -- t[3589] = 0
      "00000" when "000111000000110", -- t[3590] = 0
      "00000" when "000111000000111", -- t[3591] = 0
      "00000" when "000111000001000", -- t[3592] = 0
      "00000" when "000111000001001", -- t[3593] = 0
      "00000" when "000111000001010", -- t[3594] = 0
      "00000" when "000111000001011", -- t[3595] = 0
      "00000" when "000111000001100", -- t[3596] = 0
      "00000" when "000111000001101", -- t[3597] = 0
      "00000" when "000111000001110", -- t[3598] = 0
      "00000" when "000111000001111", -- t[3599] = 0
      "00000" when "000111000010000", -- t[3600] = 0
      "00000" when "000111000010001", -- t[3601] = 0
      "00000" when "000111000010010", -- t[3602] = 0
      "00000" when "000111000010011", -- t[3603] = 0
      "00000" when "000111000010100", -- t[3604] = 0
      "00000" when "000111000010101", -- t[3605] = 0
      "00000" when "000111000010110", -- t[3606] = 0
      "00000" when "000111000010111", -- t[3607] = 0
      "00000" when "000111000011000", -- t[3608] = 0
      "00000" when "000111000011001", -- t[3609] = 0
      "00000" when "000111000011010", -- t[3610] = 0
      "00000" when "000111000011011", -- t[3611] = 0
      "00000" when "000111000011100", -- t[3612] = 0
      "00000" when "000111000011101", -- t[3613] = 0
      "00000" when "000111000011110", -- t[3614] = 0
      "00000" when "000111000011111", -- t[3615] = 0
      "00000" when "000111000100000", -- t[3616] = 0
      "00000" when "000111000100001", -- t[3617] = 0
      "00000" when "000111000100010", -- t[3618] = 0
      "00000" when "000111000100011", -- t[3619] = 0
      "00000" when "000111000100100", -- t[3620] = 0
      "00000" when "000111000100101", -- t[3621] = 0
      "00000" when "000111000100110", -- t[3622] = 0
      "00000" when "000111000100111", -- t[3623] = 0
      "00000" when "000111000101000", -- t[3624] = 0
      "00000" when "000111000101001", -- t[3625] = 0
      "00000" when "000111000101010", -- t[3626] = 0
      "00000" when "000111000101011", -- t[3627] = 0
      "00000" when "000111000101100", -- t[3628] = 0
      "00000" when "000111000101101", -- t[3629] = 0
      "00000" when "000111000101110", -- t[3630] = 0
      "00000" when "000111000101111", -- t[3631] = 0
      "00000" when "000111000110000", -- t[3632] = 0
      "00000" when "000111000110001", -- t[3633] = 0
      "00000" when "000111000110010", -- t[3634] = 0
      "00000" when "000111000110011", -- t[3635] = 0
      "00000" when "000111000110100", -- t[3636] = 0
      "00000" when "000111000110101", -- t[3637] = 0
      "00000" when "000111000110110", -- t[3638] = 0
      "00000" when "000111000110111", -- t[3639] = 0
      "00000" when "000111000111000", -- t[3640] = 0
      "00000" when "000111000111001", -- t[3641] = 0
      "00000" when "000111000111010", -- t[3642] = 0
      "00000" when "000111000111011", -- t[3643] = 0
      "00000" when "000111000111100", -- t[3644] = 0
      "00000" when "000111000111101", -- t[3645] = 0
      "00000" when "000111000111110", -- t[3646] = 0
      "00000" when "000111000111111", -- t[3647] = 0
      "00000" when "000111001000000", -- t[3648] = 0
      "00000" when "000111001000001", -- t[3649] = 0
      "00000" when "000111001000010", -- t[3650] = 0
      "00000" when "000111001000011", -- t[3651] = 0
      "00000" when "000111001000100", -- t[3652] = 0
      "00000" when "000111001000101", -- t[3653] = 0
      "00000" when "000111001000110", -- t[3654] = 0
      "00000" when "000111001000111", -- t[3655] = 0
      "00000" when "000111001001000", -- t[3656] = 0
      "00000" when "000111001001001", -- t[3657] = 0
      "00000" when "000111001001010", -- t[3658] = 0
      "00000" when "000111001001011", -- t[3659] = 0
      "00000" when "000111001001100", -- t[3660] = 0
      "00000" when "000111001001101", -- t[3661] = 0
      "00000" when "000111001001110", -- t[3662] = 0
      "00000" when "000111001001111", -- t[3663] = 0
      "00000" when "000111001010000", -- t[3664] = 0
      "00000" when "000111001010001", -- t[3665] = 0
      "00000" when "000111001010010", -- t[3666] = 0
      "00000" when "000111001010011", -- t[3667] = 0
      "00000" when "000111001010100", -- t[3668] = 0
      "00000" when "000111001010101", -- t[3669] = 0
      "00000" when "000111001010110", -- t[3670] = 0
      "00000" when "000111001010111", -- t[3671] = 0
      "00000" when "000111001011000", -- t[3672] = 0
      "00000" when "000111001011001", -- t[3673] = 0
      "00000" when "000111001011010", -- t[3674] = 0
      "00000" when "000111001011011", -- t[3675] = 0
      "00000" when "000111001011100", -- t[3676] = 0
      "00000" when "000111001011101", -- t[3677] = 0
      "00000" when "000111001011110", -- t[3678] = 0
      "00000" when "000111001011111", -- t[3679] = 0
      "00000" when "000111001100000", -- t[3680] = 0
      "00000" when "000111001100001", -- t[3681] = 0
      "00000" when "000111001100010", -- t[3682] = 0
      "00000" when "000111001100011", -- t[3683] = 0
      "00000" when "000111001100100", -- t[3684] = 0
      "00000" when "000111001100101", -- t[3685] = 0
      "00000" when "000111001100110", -- t[3686] = 0
      "00000" when "000111001100111", -- t[3687] = 0
      "00000" when "000111001101000", -- t[3688] = 0
      "00000" when "000111001101001", -- t[3689] = 0
      "00000" when "000111001101010", -- t[3690] = 0
      "00000" when "000111001101011", -- t[3691] = 0
      "00000" when "000111001101100", -- t[3692] = 0
      "00000" when "000111001101101", -- t[3693] = 0
      "00000" when "000111001101110", -- t[3694] = 0
      "00000" when "000111001101111", -- t[3695] = 0
      "00000" when "000111001110000", -- t[3696] = 0
      "00000" when "000111001110001", -- t[3697] = 0
      "00000" when "000111001110010", -- t[3698] = 0
      "00000" when "000111001110011", -- t[3699] = 0
      "00000" when "000111001110100", -- t[3700] = 0
      "00000" when "000111001110101", -- t[3701] = 0
      "00000" when "000111001110110", -- t[3702] = 0
      "00000" when "000111001110111", -- t[3703] = 0
      "00000" when "000111001111000", -- t[3704] = 0
      "00000" when "000111001111001", -- t[3705] = 0
      "00000" when "000111001111010", -- t[3706] = 0
      "00000" when "000111001111011", -- t[3707] = 0
      "00000" when "000111001111100", -- t[3708] = 0
      "00000" when "000111001111101", -- t[3709] = 0
      "00000" when "000111001111110", -- t[3710] = 0
      "00000" when "000111001111111", -- t[3711] = 0
      "00000" when "000111010000000", -- t[3712] = 0
      "00000" when "000111010000001", -- t[3713] = 0
      "00000" when "000111010000010", -- t[3714] = 0
      "00000" when "000111010000011", -- t[3715] = 0
      "00000" when "000111010000100", -- t[3716] = 0
      "00000" when "000111010000101", -- t[3717] = 0
      "00000" when "000111010000110", -- t[3718] = 0
      "00000" when "000111010000111", -- t[3719] = 0
      "00000" when "000111010001000", -- t[3720] = 0
      "00000" when "000111010001001", -- t[3721] = 0
      "00000" when "000111010001010", -- t[3722] = 0
      "00000" when "000111010001011", -- t[3723] = 0
      "00000" when "000111010001100", -- t[3724] = 0
      "00000" when "000111010001101", -- t[3725] = 0
      "00000" when "000111010001110", -- t[3726] = 0
      "00000" when "000111010001111", -- t[3727] = 0
      "00000" when "000111010010000", -- t[3728] = 0
      "00000" when "000111010010001", -- t[3729] = 0
      "00000" when "000111010010010", -- t[3730] = 0
      "00000" when "000111010010011", -- t[3731] = 0
      "00000" when "000111010010100", -- t[3732] = 0
      "00000" when "000111010010101", -- t[3733] = 0
      "00000" when "000111010010110", -- t[3734] = 0
      "00000" when "000111010010111", -- t[3735] = 0
      "00000" when "000111010011000", -- t[3736] = 0
      "00000" when "000111010011001", -- t[3737] = 0
      "00000" when "000111010011010", -- t[3738] = 0
      "00000" when "000111010011011", -- t[3739] = 0
      "00000" when "000111010011100", -- t[3740] = 0
      "00000" when "000111010011101", -- t[3741] = 0
      "00000" when "000111010011110", -- t[3742] = 0
      "00000" when "000111010011111", -- t[3743] = 0
      "00000" when "000111010100000", -- t[3744] = 0
      "00000" when "000111010100001", -- t[3745] = 0
      "00000" when "000111010100010", -- t[3746] = 0
      "00000" when "000111010100011", -- t[3747] = 0
      "00000" when "000111010100100", -- t[3748] = 0
      "00000" when "000111010100101", -- t[3749] = 0
      "00000" when "000111010100110", -- t[3750] = 0
      "00000" when "000111010100111", -- t[3751] = 0
      "00000" when "000111010101000", -- t[3752] = 0
      "00000" when "000111010101001", -- t[3753] = 0
      "00000" when "000111010101010", -- t[3754] = 0
      "00000" when "000111010101011", -- t[3755] = 0
      "00000" when "000111010101100", -- t[3756] = 0
      "00000" when "000111010101101", -- t[3757] = 0
      "00000" when "000111010101110", -- t[3758] = 0
      "00000" when "000111010101111", -- t[3759] = 0
      "00000" when "000111010110000", -- t[3760] = 0
      "00000" when "000111010110001", -- t[3761] = 0
      "00000" when "000111010110010", -- t[3762] = 0
      "00000" when "000111010110011", -- t[3763] = 0
      "00000" when "000111010110100", -- t[3764] = 0
      "00000" when "000111010110101", -- t[3765] = 0
      "00000" when "000111010110110", -- t[3766] = 0
      "00000" when "000111010110111", -- t[3767] = 0
      "00000" when "000111010111000", -- t[3768] = 0
      "00000" when "000111010111001", -- t[3769] = 0
      "00000" when "000111010111010", -- t[3770] = 0
      "00000" when "000111010111011", -- t[3771] = 0
      "00000" when "000111010111100", -- t[3772] = 0
      "00000" when "000111010111101", -- t[3773] = 0
      "00000" when "000111010111110", -- t[3774] = 0
      "00000" when "000111010111111", -- t[3775] = 0
      "00000" when "000111011000000", -- t[3776] = 0
      "00000" when "000111011000001", -- t[3777] = 0
      "00000" when "000111011000010", -- t[3778] = 0
      "00000" when "000111011000011", -- t[3779] = 0
      "00000" when "000111011000100", -- t[3780] = 0
      "00000" when "000111011000101", -- t[3781] = 0
      "00000" when "000111011000110", -- t[3782] = 0
      "00000" when "000111011000111", -- t[3783] = 0
      "00000" when "000111011001000", -- t[3784] = 0
      "00000" when "000111011001001", -- t[3785] = 0
      "00000" when "000111011001010", -- t[3786] = 0
      "00000" when "000111011001011", -- t[3787] = 0
      "00000" when "000111011001100", -- t[3788] = 0
      "00000" when "000111011001101", -- t[3789] = 0
      "00000" when "000111011001110", -- t[3790] = 0
      "00000" when "000111011001111", -- t[3791] = 0
      "00000" when "000111011010000", -- t[3792] = 0
      "00000" when "000111011010001", -- t[3793] = 0
      "00000" when "000111011010010", -- t[3794] = 0
      "00000" when "000111011010011", -- t[3795] = 0
      "00000" when "000111011010100", -- t[3796] = 0
      "00000" when "000111011010101", -- t[3797] = 0
      "00000" when "000111011010110", -- t[3798] = 0
      "00000" when "000111011010111", -- t[3799] = 0
      "00000" when "000111011011000", -- t[3800] = 0
      "00000" when "000111011011001", -- t[3801] = 0
      "00000" when "000111011011010", -- t[3802] = 0
      "00000" when "000111011011011", -- t[3803] = 0
      "00000" when "000111011011100", -- t[3804] = 0
      "00000" when "000111011011101", -- t[3805] = 0
      "00000" when "000111011011110", -- t[3806] = 0
      "00000" when "000111011011111", -- t[3807] = 0
      "00000" when "000111011100000", -- t[3808] = 0
      "00000" when "000111011100001", -- t[3809] = 0
      "00000" when "000111011100010", -- t[3810] = 0
      "00000" when "000111011100011", -- t[3811] = 0
      "00000" when "000111011100100", -- t[3812] = 0
      "00000" when "000111011100101", -- t[3813] = 0
      "00000" when "000111011100110", -- t[3814] = 0
      "00000" when "000111011100111", -- t[3815] = 0
      "00000" when "000111011101000", -- t[3816] = 0
      "00000" when "000111011101001", -- t[3817] = 0
      "00000" when "000111011101010", -- t[3818] = 0
      "00000" when "000111011101011", -- t[3819] = 0
      "00000" when "000111011101100", -- t[3820] = 0
      "00000" when "000111011101101", -- t[3821] = 0
      "00000" when "000111011101110", -- t[3822] = 0
      "00000" when "000111011101111", -- t[3823] = 0
      "00000" when "000111011110000", -- t[3824] = 0
      "00000" when "000111011110001", -- t[3825] = 0
      "00000" when "000111011110010", -- t[3826] = 0
      "00000" when "000111011110011", -- t[3827] = 0
      "00000" when "000111011110100", -- t[3828] = 0
      "00000" when "000111011110101", -- t[3829] = 0
      "00000" when "000111011110110", -- t[3830] = 0
      "00000" when "000111011110111", -- t[3831] = 0
      "00000" when "000111011111000", -- t[3832] = 0
      "00000" when "000111011111001", -- t[3833] = 0
      "00000" when "000111011111010", -- t[3834] = 0
      "00000" when "000111011111011", -- t[3835] = 0
      "00000" when "000111011111100", -- t[3836] = 0
      "00000" when "000111011111101", -- t[3837] = 0
      "00000" when "000111011111110", -- t[3838] = 0
      "00000" when "000111011111111", -- t[3839] = 0
      "00000" when "000111100000000", -- t[3840] = 0
      "00000" when "000111100000001", -- t[3841] = 0
      "00000" when "000111100000010", -- t[3842] = 0
      "00000" when "000111100000011", -- t[3843] = 0
      "00000" when "000111100000100", -- t[3844] = 0
      "00000" when "000111100000101", -- t[3845] = 0
      "00000" when "000111100000110", -- t[3846] = 0
      "00000" when "000111100000111", -- t[3847] = 0
      "00000" when "000111100001000", -- t[3848] = 0
      "00000" when "000111100001001", -- t[3849] = 0
      "00000" when "000111100001010", -- t[3850] = 0
      "00000" when "000111100001011", -- t[3851] = 0
      "00000" when "000111100001100", -- t[3852] = 0
      "00000" when "000111100001101", -- t[3853] = 0
      "00000" when "000111100001110", -- t[3854] = 0
      "00000" when "000111100001111", -- t[3855] = 0
      "00000" when "000111100010000", -- t[3856] = 0
      "00000" when "000111100010001", -- t[3857] = 0
      "00000" when "000111100010010", -- t[3858] = 0
      "00000" when "000111100010011", -- t[3859] = 0
      "00000" when "000111100010100", -- t[3860] = 0
      "00000" when "000111100010101", -- t[3861] = 0
      "00000" when "000111100010110", -- t[3862] = 0
      "00000" when "000111100010111", -- t[3863] = 0
      "00000" when "000111100011000", -- t[3864] = 0
      "00000" when "000111100011001", -- t[3865] = 0
      "00000" when "000111100011010", -- t[3866] = 0
      "00000" when "000111100011011", -- t[3867] = 0
      "00000" when "000111100011100", -- t[3868] = 0
      "00000" when "000111100011101", -- t[3869] = 0
      "00000" when "000111100011110", -- t[3870] = 0
      "00000" when "000111100011111", -- t[3871] = 0
      "00000" when "000111100100000", -- t[3872] = 0
      "00000" when "000111100100001", -- t[3873] = 0
      "00000" when "000111100100010", -- t[3874] = 0
      "00000" when "000111100100011", -- t[3875] = 0
      "00000" when "000111100100100", -- t[3876] = 0
      "00000" when "000111100100101", -- t[3877] = 0
      "00000" when "000111100100110", -- t[3878] = 0
      "00000" when "000111100100111", -- t[3879] = 0
      "00000" when "000111100101000", -- t[3880] = 0
      "00000" when "000111100101001", -- t[3881] = 0
      "00000" when "000111100101010", -- t[3882] = 0
      "00000" when "000111100101011", -- t[3883] = 0
      "00000" when "000111100101100", -- t[3884] = 0
      "00000" when "000111100101101", -- t[3885] = 0
      "00000" when "000111100101110", -- t[3886] = 0
      "00000" when "000111100101111", -- t[3887] = 0
      "00000" when "000111100110000", -- t[3888] = 0
      "00000" when "000111100110001", -- t[3889] = 0
      "00000" when "000111100110010", -- t[3890] = 0
      "00000" when "000111100110011", -- t[3891] = 0
      "00000" when "000111100110100", -- t[3892] = 0
      "00000" when "000111100110101", -- t[3893] = 0
      "00000" when "000111100110110", -- t[3894] = 0
      "00000" when "000111100110111", -- t[3895] = 0
      "00000" when "000111100111000", -- t[3896] = 0
      "00000" when "000111100111001", -- t[3897] = 0
      "00000" when "000111100111010", -- t[3898] = 0
      "00000" when "000111100111011", -- t[3899] = 0
      "00000" when "000111100111100", -- t[3900] = 0
      "00000" when "000111100111101", -- t[3901] = 0
      "00000" when "000111100111110", -- t[3902] = 0
      "00000" when "000111100111111", -- t[3903] = 0
      "00000" when "000111101000000", -- t[3904] = 0
      "00000" when "000111101000001", -- t[3905] = 0
      "00000" when "000111101000010", -- t[3906] = 0
      "00000" when "000111101000011", -- t[3907] = 0
      "00000" when "000111101000100", -- t[3908] = 0
      "00000" when "000111101000101", -- t[3909] = 0
      "00000" when "000111101000110", -- t[3910] = 0
      "00000" when "000111101000111", -- t[3911] = 0
      "00000" when "000111101001000", -- t[3912] = 0
      "00000" when "000111101001001", -- t[3913] = 0
      "00000" when "000111101001010", -- t[3914] = 0
      "00000" when "000111101001011", -- t[3915] = 0
      "00000" when "000111101001100", -- t[3916] = 0
      "00000" when "000111101001101", -- t[3917] = 0
      "00000" when "000111101001110", -- t[3918] = 0
      "00000" when "000111101001111", -- t[3919] = 0
      "00000" when "000111101010000", -- t[3920] = 0
      "00000" when "000111101010001", -- t[3921] = 0
      "00000" when "000111101010010", -- t[3922] = 0
      "00000" when "000111101010011", -- t[3923] = 0
      "00000" when "000111101010100", -- t[3924] = 0
      "00000" when "000111101010101", -- t[3925] = 0
      "00000" when "000111101010110", -- t[3926] = 0
      "00000" when "000111101010111", -- t[3927] = 0
      "00000" when "000111101011000", -- t[3928] = 0
      "00000" when "000111101011001", -- t[3929] = 0
      "00000" when "000111101011010", -- t[3930] = 0
      "00000" when "000111101011011", -- t[3931] = 0
      "00000" when "000111101011100", -- t[3932] = 0
      "00000" when "000111101011101", -- t[3933] = 0
      "00000" when "000111101011110", -- t[3934] = 0
      "00000" when "000111101011111", -- t[3935] = 0
      "00000" when "000111101100000", -- t[3936] = 0
      "00000" when "000111101100001", -- t[3937] = 0
      "00000" when "000111101100010", -- t[3938] = 0
      "00000" when "000111101100011", -- t[3939] = 0
      "00000" when "000111101100100", -- t[3940] = 0
      "00000" when "000111101100101", -- t[3941] = 0
      "00000" when "000111101100110", -- t[3942] = 0
      "00000" when "000111101100111", -- t[3943] = 0
      "00000" when "000111101101000", -- t[3944] = 0
      "00000" when "000111101101001", -- t[3945] = 0
      "00000" when "000111101101010", -- t[3946] = 0
      "00000" when "000111101101011", -- t[3947] = 0
      "00000" when "000111101101100", -- t[3948] = 0
      "00000" when "000111101101101", -- t[3949] = 0
      "00000" when "000111101101110", -- t[3950] = 0
      "00000" when "000111101101111", -- t[3951] = 0
      "00000" when "000111101110000", -- t[3952] = 0
      "00000" when "000111101110001", -- t[3953] = 0
      "00000" when "000111101110010", -- t[3954] = 0
      "00000" when "000111101110011", -- t[3955] = 0
      "00000" when "000111101110100", -- t[3956] = 0
      "00000" when "000111101110101", -- t[3957] = 0
      "00000" when "000111101110110", -- t[3958] = 0
      "00000" when "000111101110111", -- t[3959] = 0
      "00000" when "000111101111000", -- t[3960] = 0
      "00000" when "000111101111001", -- t[3961] = 0
      "00000" when "000111101111010", -- t[3962] = 0
      "00000" when "000111101111011", -- t[3963] = 0
      "00000" when "000111101111100", -- t[3964] = 0
      "00000" when "000111101111101", -- t[3965] = 0
      "00000" when "000111101111110", -- t[3966] = 0
      "00000" when "000111101111111", -- t[3967] = 0
      "00000" when "000111110000000", -- t[3968] = 0
      "00000" when "000111110000001", -- t[3969] = 0
      "00000" when "000111110000010", -- t[3970] = 0
      "00000" when "000111110000011", -- t[3971] = 0
      "00000" when "000111110000100", -- t[3972] = 0
      "00000" when "000111110000101", -- t[3973] = 0
      "00000" when "000111110000110", -- t[3974] = 0
      "00000" when "000111110000111", -- t[3975] = 0
      "00000" when "000111110001000", -- t[3976] = 0
      "00000" when "000111110001001", -- t[3977] = 0
      "00000" when "000111110001010", -- t[3978] = 0
      "00000" when "000111110001011", -- t[3979] = 0
      "00000" when "000111110001100", -- t[3980] = 0
      "00000" when "000111110001101", -- t[3981] = 0
      "00000" when "000111110001110", -- t[3982] = 0
      "00000" when "000111110001111", -- t[3983] = 0
      "00000" when "000111110010000", -- t[3984] = 0
      "00000" when "000111110010001", -- t[3985] = 0
      "00000" when "000111110010010", -- t[3986] = 0
      "00000" when "000111110010011", -- t[3987] = 0
      "00000" when "000111110010100", -- t[3988] = 0
      "00000" when "000111110010101", -- t[3989] = 0
      "00000" when "000111110010110", -- t[3990] = 0
      "00000" when "000111110010111", -- t[3991] = 0
      "00000" when "000111110011000", -- t[3992] = 0
      "00000" when "000111110011001", -- t[3993] = 0
      "00000" when "000111110011010", -- t[3994] = 0
      "00000" when "000111110011011", -- t[3995] = 0
      "00000" when "000111110011100", -- t[3996] = 0
      "00000" when "000111110011101", -- t[3997] = 0
      "00000" when "000111110011110", -- t[3998] = 0
      "00000" when "000111110011111", -- t[3999] = 0
      "00000" when "000111110100000", -- t[4000] = 0
      "00000" when "000111110100001", -- t[4001] = 0
      "00000" when "000111110100010", -- t[4002] = 0
      "00000" when "000111110100011", -- t[4003] = 0
      "00000" when "000111110100100", -- t[4004] = 0
      "00000" when "000111110100101", -- t[4005] = 0
      "00000" when "000111110100110", -- t[4006] = 0
      "00000" when "000111110100111", -- t[4007] = 0
      "00000" when "000111110101000", -- t[4008] = 0
      "00000" when "000111110101001", -- t[4009] = 0
      "00000" when "000111110101010", -- t[4010] = 0
      "00000" when "000111110101011", -- t[4011] = 0
      "00000" when "000111110101100", -- t[4012] = 0
      "00000" when "000111110101101", -- t[4013] = 0
      "00000" when "000111110101110", -- t[4014] = 0
      "00000" when "000111110101111", -- t[4015] = 0
      "00000" when "000111110110000", -- t[4016] = 0
      "00000" when "000111110110001", -- t[4017] = 0
      "00000" when "000111110110010", -- t[4018] = 0
      "00000" when "000111110110011", -- t[4019] = 0
      "00000" when "000111110110100", -- t[4020] = 0
      "00000" when "000111110110101", -- t[4021] = 0
      "00000" when "000111110110110", -- t[4022] = 0
      "00000" when "000111110110111", -- t[4023] = 0
      "00000" when "000111110111000", -- t[4024] = 0
      "00000" when "000111110111001", -- t[4025] = 0
      "00000" when "000111110111010", -- t[4026] = 0
      "00000" when "000111110111011", -- t[4027] = 0
      "00000" when "000111110111100", -- t[4028] = 0
      "00000" when "000111110111101", -- t[4029] = 0
      "00000" when "000111110111110", -- t[4030] = 0
      "00000" when "000111110111111", -- t[4031] = 0
      "00000" when "000111111000000", -- t[4032] = 0
      "00000" when "000111111000001", -- t[4033] = 0
      "00000" when "000111111000010", -- t[4034] = 0
      "00000" when "000111111000011", -- t[4035] = 0
      "00000" when "000111111000100", -- t[4036] = 0
      "00000" when "000111111000101", -- t[4037] = 0
      "00000" when "000111111000110", -- t[4038] = 0
      "00000" when "000111111000111", -- t[4039] = 0
      "00000" when "000111111001000", -- t[4040] = 0
      "00000" when "000111111001001", -- t[4041] = 0
      "00000" when "000111111001010", -- t[4042] = 0
      "00000" when "000111111001011", -- t[4043] = 0
      "00000" when "000111111001100", -- t[4044] = 0
      "00000" when "000111111001101", -- t[4045] = 0
      "00000" when "000111111001110", -- t[4046] = 0
      "00000" when "000111111001111", -- t[4047] = 0
      "00000" when "000111111010000", -- t[4048] = 0
      "00000" when "000111111010001", -- t[4049] = 0
      "00000" when "000111111010010", -- t[4050] = 0
      "00000" when "000111111010011", -- t[4051] = 0
      "00000" when "000111111010100", -- t[4052] = 0
      "00000" when "000111111010101", -- t[4053] = 0
      "00000" when "000111111010110", -- t[4054] = 0
      "00000" when "000111111010111", -- t[4055] = 0
      "00000" when "000111111011000", -- t[4056] = 0
      "00000" when "000111111011001", -- t[4057] = 0
      "00000" when "000111111011010", -- t[4058] = 0
      "00000" when "000111111011011", -- t[4059] = 0
      "00000" when "000111111011100", -- t[4060] = 0
      "00000" when "000111111011101", -- t[4061] = 0
      "00000" when "000111111011110", -- t[4062] = 0
      "00000" when "000111111011111", -- t[4063] = 0
      "00000" when "000111111100000", -- t[4064] = 0
      "00000" when "000111111100001", -- t[4065] = 0
      "00000" when "000111111100010", -- t[4066] = 0
      "00000" when "000111111100011", -- t[4067] = 0
      "00000" when "000111111100100", -- t[4068] = 0
      "00000" when "000111111100101", -- t[4069] = 0
      "00000" when "000111111100110", -- t[4070] = 0
      "00000" when "000111111100111", -- t[4071] = 0
      "00000" when "000111111101000", -- t[4072] = 0
      "00000" when "000111111101001", -- t[4073] = 0
      "00000" when "000111111101010", -- t[4074] = 0
      "00000" when "000111111101011", -- t[4075] = 0
      "00000" when "000111111101100", -- t[4076] = 0
      "00000" when "000111111101101", -- t[4077] = 0
      "00000" when "000111111101110", -- t[4078] = 0
      "00000" when "000111111101111", -- t[4079] = 0
      "00000" when "000111111110000", -- t[4080] = 0
      "00000" when "000111111110001", -- t[4081] = 0
      "00000" when "000111111110010", -- t[4082] = 0
      "00000" when "000111111110011", -- t[4083] = 0
      "00000" when "000111111110100", -- t[4084] = 0
      "00000" when "000111111110101", -- t[4085] = 0
      "00000" when "000111111110110", -- t[4086] = 0
      "00000" when "000111111110111", -- t[4087] = 0
      "00000" when "000111111111000", -- t[4088] = 0
      "00000" when "000111111111001", -- t[4089] = 0
      "00000" when "000111111111010", -- t[4090] = 0
      "00000" when "000111111111011", -- t[4091] = 0
      "00000" when "000111111111100", -- t[4092] = 0
      "00000" when "000111111111101", -- t[4093] = 0
      "00000" when "000111111111110", -- t[4094] = 0
      "00000" when "000111111111111", -- t[4095] = 0
      "00000" when "001000000000000", -- t[4096] = 0
      "00000" when "001000000000001", -- t[4097] = 0
      "00000" when "001000000000010", -- t[4098] = 0
      "00000" when "001000000000011", -- t[4099] = 0
      "00000" when "001000000000100", -- t[4100] = 0
      "00000" when "001000000000101", -- t[4101] = 0
      "00000" when "001000000000110", -- t[4102] = 0
      "00000" when "001000000000111", -- t[4103] = 0
      "00000" when "001000000001000", -- t[4104] = 0
      "00000" when "001000000001001", -- t[4105] = 0
      "00000" when "001000000001010", -- t[4106] = 0
      "00000" when "001000000001011", -- t[4107] = 0
      "00000" when "001000000001100", -- t[4108] = 0
      "00000" when "001000000001101", -- t[4109] = 0
      "00000" when "001000000001110", -- t[4110] = 0
      "00000" when "001000000001111", -- t[4111] = 0
      "00000" when "001000000010000", -- t[4112] = 0
      "00000" when "001000000010001", -- t[4113] = 0
      "00000" when "001000000010010", -- t[4114] = 0
      "00000" when "001000000010011", -- t[4115] = 0
      "00000" when "001000000010100", -- t[4116] = 0
      "00000" when "001000000010101", -- t[4117] = 0
      "00000" when "001000000010110", -- t[4118] = 0
      "00000" when "001000000010111", -- t[4119] = 0
      "00000" when "001000000011000", -- t[4120] = 0
      "00000" when "001000000011001", -- t[4121] = 0
      "00000" when "001000000011010", -- t[4122] = 0
      "00000" when "001000000011011", -- t[4123] = 0
      "00000" when "001000000011100", -- t[4124] = 0
      "00000" when "001000000011101", -- t[4125] = 0
      "00000" when "001000000011110", -- t[4126] = 0
      "00000" when "001000000011111", -- t[4127] = 0
      "00000" when "001000000100000", -- t[4128] = 0
      "00000" when "001000000100001", -- t[4129] = 0
      "00000" when "001000000100010", -- t[4130] = 0
      "00000" when "001000000100011", -- t[4131] = 0
      "00000" when "001000000100100", -- t[4132] = 0
      "00000" when "001000000100101", -- t[4133] = 0
      "00000" when "001000000100110", -- t[4134] = 0
      "00000" when "001000000100111", -- t[4135] = 0
      "00000" when "001000000101000", -- t[4136] = 0
      "00000" when "001000000101001", -- t[4137] = 0
      "00000" when "001000000101010", -- t[4138] = 0
      "00000" when "001000000101011", -- t[4139] = 0
      "00000" when "001000000101100", -- t[4140] = 0
      "00000" when "001000000101101", -- t[4141] = 0
      "00000" when "001000000101110", -- t[4142] = 0
      "00000" when "001000000101111", -- t[4143] = 0
      "00000" when "001000000110000", -- t[4144] = 0
      "00000" when "001000000110001", -- t[4145] = 0
      "00000" when "001000000110010", -- t[4146] = 0
      "00000" when "001000000110011", -- t[4147] = 0
      "00000" when "001000000110100", -- t[4148] = 0
      "00000" when "001000000110101", -- t[4149] = 0
      "00000" when "001000000110110", -- t[4150] = 0
      "00000" when "001000000110111", -- t[4151] = 0
      "00000" when "001000000111000", -- t[4152] = 0
      "00000" when "001000000111001", -- t[4153] = 0
      "00000" when "001000000111010", -- t[4154] = 0
      "00000" when "001000000111011", -- t[4155] = 0
      "00000" when "001000000111100", -- t[4156] = 0
      "00000" when "001000000111101", -- t[4157] = 0
      "00000" when "001000000111110", -- t[4158] = 0
      "00000" when "001000000111111", -- t[4159] = 0
      "00000" when "001000001000000", -- t[4160] = 0
      "00000" when "001000001000001", -- t[4161] = 0
      "00000" when "001000001000010", -- t[4162] = 0
      "00000" when "001000001000011", -- t[4163] = 0
      "00000" when "001000001000100", -- t[4164] = 0
      "00000" when "001000001000101", -- t[4165] = 0
      "00000" when "001000001000110", -- t[4166] = 0
      "00000" when "001000001000111", -- t[4167] = 0
      "00000" when "001000001001000", -- t[4168] = 0
      "00000" when "001000001001001", -- t[4169] = 0
      "00000" when "001000001001010", -- t[4170] = 0
      "00000" when "001000001001011", -- t[4171] = 0
      "00000" when "001000001001100", -- t[4172] = 0
      "00000" when "001000001001101", -- t[4173] = 0
      "00000" when "001000001001110", -- t[4174] = 0
      "00000" when "001000001001111", -- t[4175] = 0
      "00000" when "001000001010000", -- t[4176] = 0
      "00000" when "001000001010001", -- t[4177] = 0
      "00000" when "001000001010010", -- t[4178] = 0
      "00000" when "001000001010011", -- t[4179] = 0
      "00000" when "001000001010100", -- t[4180] = 0
      "00000" when "001000001010101", -- t[4181] = 0
      "00000" when "001000001010110", -- t[4182] = 0
      "00000" when "001000001010111", -- t[4183] = 0
      "00000" when "001000001011000", -- t[4184] = 0
      "00000" when "001000001011001", -- t[4185] = 0
      "00000" when "001000001011010", -- t[4186] = 0
      "00000" when "001000001011011", -- t[4187] = 0
      "00000" when "001000001011100", -- t[4188] = 0
      "00000" when "001000001011101", -- t[4189] = 0
      "00000" when "001000001011110", -- t[4190] = 0
      "00000" when "001000001011111", -- t[4191] = 0
      "00000" when "001000001100000", -- t[4192] = 0
      "00000" when "001000001100001", -- t[4193] = 0
      "00000" when "001000001100010", -- t[4194] = 0
      "00000" when "001000001100011", -- t[4195] = 0
      "00000" when "001000001100100", -- t[4196] = 0
      "00000" when "001000001100101", -- t[4197] = 0
      "00000" when "001000001100110", -- t[4198] = 0
      "00000" when "001000001100111", -- t[4199] = 0
      "00000" when "001000001101000", -- t[4200] = 0
      "00000" when "001000001101001", -- t[4201] = 0
      "00000" when "001000001101010", -- t[4202] = 0
      "00000" when "001000001101011", -- t[4203] = 0
      "00000" when "001000001101100", -- t[4204] = 0
      "00000" when "001000001101101", -- t[4205] = 0
      "00000" when "001000001101110", -- t[4206] = 0
      "00000" when "001000001101111", -- t[4207] = 0
      "00000" when "001000001110000", -- t[4208] = 0
      "00000" when "001000001110001", -- t[4209] = 0
      "00000" when "001000001110010", -- t[4210] = 0
      "00000" when "001000001110011", -- t[4211] = 0
      "00000" when "001000001110100", -- t[4212] = 0
      "00000" when "001000001110101", -- t[4213] = 0
      "00000" when "001000001110110", -- t[4214] = 0
      "00000" when "001000001110111", -- t[4215] = 0
      "00000" when "001000001111000", -- t[4216] = 0
      "00000" when "001000001111001", -- t[4217] = 0
      "00000" when "001000001111010", -- t[4218] = 0
      "00000" when "001000001111011", -- t[4219] = 0
      "00000" when "001000001111100", -- t[4220] = 0
      "00000" when "001000001111101", -- t[4221] = 0
      "00000" when "001000001111110", -- t[4222] = 0
      "00000" when "001000001111111", -- t[4223] = 0
      "00000" when "001000010000000", -- t[4224] = 0
      "00000" when "001000010000001", -- t[4225] = 0
      "00000" when "001000010000010", -- t[4226] = 0
      "00000" when "001000010000011", -- t[4227] = 0
      "00000" when "001000010000100", -- t[4228] = 0
      "00000" when "001000010000101", -- t[4229] = 0
      "00000" when "001000010000110", -- t[4230] = 0
      "00000" when "001000010000111", -- t[4231] = 0
      "00000" when "001000010001000", -- t[4232] = 0
      "00000" when "001000010001001", -- t[4233] = 0
      "00000" when "001000010001010", -- t[4234] = 0
      "00000" when "001000010001011", -- t[4235] = 0
      "00000" when "001000010001100", -- t[4236] = 0
      "00000" when "001000010001101", -- t[4237] = 0
      "00000" when "001000010001110", -- t[4238] = 0
      "00000" when "001000010001111", -- t[4239] = 0
      "00000" when "001000010010000", -- t[4240] = 0
      "00000" when "001000010010001", -- t[4241] = 0
      "00000" when "001000010010010", -- t[4242] = 0
      "00000" when "001000010010011", -- t[4243] = 0
      "00000" when "001000010010100", -- t[4244] = 0
      "00000" when "001000010010101", -- t[4245] = 0
      "00000" when "001000010010110", -- t[4246] = 0
      "00000" when "001000010010111", -- t[4247] = 0
      "00000" when "001000010011000", -- t[4248] = 0
      "00000" when "001000010011001", -- t[4249] = 0
      "00000" when "001000010011010", -- t[4250] = 0
      "00000" when "001000010011011", -- t[4251] = 0
      "00000" when "001000010011100", -- t[4252] = 0
      "00000" when "001000010011101", -- t[4253] = 0
      "00000" when "001000010011110", -- t[4254] = 0
      "00000" when "001000010011111", -- t[4255] = 0
      "00000" when "001000010100000", -- t[4256] = 0
      "00000" when "001000010100001", -- t[4257] = 0
      "00000" when "001000010100010", -- t[4258] = 0
      "00000" when "001000010100011", -- t[4259] = 0
      "00000" when "001000010100100", -- t[4260] = 0
      "00000" when "001000010100101", -- t[4261] = 0
      "00000" when "001000010100110", -- t[4262] = 0
      "00000" when "001000010100111", -- t[4263] = 0
      "00000" when "001000010101000", -- t[4264] = 0
      "00000" when "001000010101001", -- t[4265] = 0
      "00000" when "001000010101010", -- t[4266] = 0
      "00000" when "001000010101011", -- t[4267] = 0
      "00000" when "001000010101100", -- t[4268] = 0
      "00000" when "001000010101101", -- t[4269] = 0
      "00000" when "001000010101110", -- t[4270] = 0
      "00000" when "001000010101111", -- t[4271] = 0
      "00000" when "001000010110000", -- t[4272] = 0
      "00000" when "001000010110001", -- t[4273] = 0
      "00000" when "001000010110010", -- t[4274] = 0
      "00000" when "001000010110011", -- t[4275] = 0
      "00000" when "001000010110100", -- t[4276] = 0
      "00000" when "001000010110101", -- t[4277] = 0
      "00000" when "001000010110110", -- t[4278] = 0
      "00000" when "001000010110111", -- t[4279] = 0
      "00000" when "001000010111000", -- t[4280] = 0
      "00000" when "001000010111001", -- t[4281] = 0
      "00000" when "001000010111010", -- t[4282] = 0
      "00000" when "001000010111011", -- t[4283] = 0
      "00000" when "001000010111100", -- t[4284] = 0
      "00000" when "001000010111101", -- t[4285] = 0
      "00000" when "001000010111110", -- t[4286] = 0
      "00000" when "001000010111111", -- t[4287] = 0
      "00000" when "001000011000000", -- t[4288] = 0
      "00000" when "001000011000001", -- t[4289] = 0
      "00000" when "001000011000010", -- t[4290] = 0
      "00000" when "001000011000011", -- t[4291] = 0
      "00000" when "001000011000100", -- t[4292] = 0
      "00000" when "001000011000101", -- t[4293] = 0
      "00000" when "001000011000110", -- t[4294] = 0
      "00000" when "001000011000111", -- t[4295] = 0
      "00000" when "001000011001000", -- t[4296] = 0
      "00000" when "001000011001001", -- t[4297] = 0
      "00000" when "001000011001010", -- t[4298] = 0
      "00000" when "001000011001011", -- t[4299] = 0
      "00000" when "001000011001100", -- t[4300] = 0
      "00000" when "001000011001101", -- t[4301] = 0
      "00000" when "001000011001110", -- t[4302] = 0
      "00000" when "001000011001111", -- t[4303] = 0
      "00000" when "001000011010000", -- t[4304] = 0
      "00000" when "001000011010001", -- t[4305] = 0
      "00000" when "001000011010010", -- t[4306] = 0
      "00000" when "001000011010011", -- t[4307] = 0
      "00000" when "001000011010100", -- t[4308] = 0
      "00000" when "001000011010101", -- t[4309] = 0
      "00000" when "001000011010110", -- t[4310] = 0
      "00000" when "001000011010111", -- t[4311] = 0
      "00000" when "001000011011000", -- t[4312] = 0
      "00000" when "001000011011001", -- t[4313] = 0
      "00000" when "001000011011010", -- t[4314] = 0
      "00000" when "001000011011011", -- t[4315] = 0
      "00000" when "001000011011100", -- t[4316] = 0
      "00000" when "001000011011101", -- t[4317] = 0
      "00000" when "001000011011110", -- t[4318] = 0
      "00000" when "001000011011111", -- t[4319] = 0
      "00000" when "001000011100000", -- t[4320] = 0
      "00000" when "001000011100001", -- t[4321] = 0
      "00000" when "001000011100010", -- t[4322] = 0
      "00000" when "001000011100011", -- t[4323] = 0
      "00000" when "001000011100100", -- t[4324] = 0
      "00000" when "001000011100101", -- t[4325] = 0
      "00000" when "001000011100110", -- t[4326] = 0
      "00000" when "001000011100111", -- t[4327] = 0
      "00000" when "001000011101000", -- t[4328] = 0
      "00000" when "001000011101001", -- t[4329] = 0
      "00000" when "001000011101010", -- t[4330] = 0
      "00000" when "001000011101011", -- t[4331] = 0
      "00000" when "001000011101100", -- t[4332] = 0
      "00000" when "001000011101101", -- t[4333] = 0
      "00000" when "001000011101110", -- t[4334] = 0
      "00000" when "001000011101111", -- t[4335] = 0
      "00000" when "001000011110000", -- t[4336] = 0
      "00000" when "001000011110001", -- t[4337] = 0
      "00000" when "001000011110010", -- t[4338] = 0
      "00000" when "001000011110011", -- t[4339] = 0
      "00000" when "001000011110100", -- t[4340] = 0
      "00000" when "001000011110101", -- t[4341] = 0
      "00000" when "001000011110110", -- t[4342] = 0
      "00000" when "001000011110111", -- t[4343] = 0
      "00000" when "001000011111000", -- t[4344] = 0
      "00000" when "001000011111001", -- t[4345] = 0
      "00000" when "001000011111010", -- t[4346] = 0
      "00000" when "001000011111011", -- t[4347] = 0
      "00000" when "001000011111100", -- t[4348] = 0
      "00000" when "001000011111101", -- t[4349] = 0
      "00000" when "001000011111110", -- t[4350] = 0
      "00000" when "001000011111111", -- t[4351] = 0
      "00000" when "001000100000000", -- t[4352] = 0
      "00000" when "001000100000001", -- t[4353] = 0
      "00000" when "001000100000010", -- t[4354] = 0
      "00000" when "001000100000011", -- t[4355] = 0
      "00000" when "001000100000100", -- t[4356] = 0
      "00000" when "001000100000101", -- t[4357] = 0
      "00000" when "001000100000110", -- t[4358] = 0
      "00000" when "001000100000111", -- t[4359] = 0
      "00000" when "001000100001000", -- t[4360] = 0
      "00000" when "001000100001001", -- t[4361] = 0
      "00000" when "001000100001010", -- t[4362] = 0
      "00000" when "001000100001011", -- t[4363] = 0
      "00000" when "001000100001100", -- t[4364] = 0
      "00000" when "001000100001101", -- t[4365] = 0
      "00000" when "001000100001110", -- t[4366] = 0
      "00000" when "001000100001111", -- t[4367] = 0
      "00000" when "001000100010000", -- t[4368] = 0
      "00000" when "001000100010001", -- t[4369] = 0
      "00000" when "001000100010010", -- t[4370] = 0
      "00000" when "001000100010011", -- t[4371] = 0
      "00000" when "001000100010100", -- t[4372] = 0
      "00000" when "001000100010101", -- t[4373] = 0
      "00000" when "001000100010110", -- t[4374] = 0
      "00000" when "001000100010111", -- t[4375] = 0
      "00000" when "001000100011000", -- t[4376] = 0
      "00000" when "001000100011001", -- t[4377] = 0
      "00000" when "001000100011010", -- t[4378] = 0
      "00000" when "001000100011011", -- t[4379] = 0
      "00000" when "001000100011100", -- t[4380] = 0
      "00000" when "001000100011101", -- t[4381] = 0
      "00000" when "001000100011110", -- t[4382] = 0
      "00000" when "001000100011111", -- t[4383] = 0
      "00000" when "001000100100000", -- t[4384] = 0
      "00000" when "001000100100001", -- t[4385] = 0
      "00000" when "001000100100010", -- t[4386] = 0
      "00000" when "001000100100011", -- t[4387] = 0
      "00000" when "001000100100100", -- t[4388] = 0
      "00000" when "001000100100101", -- t[4389] = 0
      "00000" when "001000100100110", -- t[4390] = 0
      "00000" when "001000100100111", -- t[4391] = 0
      "00000" when "001000100101000", -- t[4392] = 0
      "00000" when "001000100101001", -- t[4393] = 0
      "00000" when "001000100101010", -- t[4394] = 0
      "00000" when "001000100101011", -- t[4395] = 0
      "00000" when "001000100101100", -- t[4396] = 0
      "00000" when "001000100101101", -- t[4397] = 0
      "00000" when "001000100101110", -- t[4398] = 0
      "00000" when "001000100101111", -- t[4399] = 0
      "00000" when "001000100110000", -- t[4400] = 0
      "00000" when "001000100110001", -- t[4401] = 0
      "00000" when "001000100110010", -- t[4402] = 0
      "00000" when "001000100110011", -- t[4403] = 0
      "00000" when "001000100110100", -- t[4404] = 0
      "00000" when "001000100110101", -- t[4405] = 0
      "00000" when "001000100110110", -- t[4406] = 0
      "00000" when "001000100110111", -- t[4407] = 0
      "00000" when "001000100111000", -- t[4408] = 0
      "00000" when "001000100111001", -- t[4409] = 0
      "00000" when "001000100111010", -- t[4410] = 0
      "00000" when "001000100111011", -- t[4411] = 0
      "00000" when "001000100111100", -- t[4412] = 0
      "00000" when "001000100111101", -- t[4413] = 0
      "00000" when "001000100111110", -- t[4414] = 0
      "00000" when "001000100111111", -- t[4415] = 0
      "00000" when "001000101000000", -- t[4416] = 0
      "00000" when "001000101000001", -- t[4417] = 0
      "00000" when "001000101000010", -- t[4418] = 0
      "00000" when "001000101000011", -- t[4419] = 0
      "00000" when "001000101000100", -- t[4420] = 0
      "00000" when "001000101000101", -- t[4421] = 0
      "00000" when "001000101000110", -- t[4422] = 0
      "00000" when "001000101000111", -- t[4423] = 0
      "00000" when "001000101001000", -- t[4424] = 0
      "00000" when "001000101001001", -- t[4425] = 0
      "00000" when "001000101001010", -- t[4426] = 0
      "00000" when "001000101001011", -- t[4427] = 0
      "00000" when "001000101001100", -- t[4428] = 0
      "00000" when "001000101001101", -- t[4429] = 0
      "00000" when "001000101001110", -- t[4430] = 0
      "00000" when "001000101001111", -- t[4431] = 0
      "00000" when "001000101010000", -- t[4432] = 0
      "00000" when "001000101010001", -- t[4433] = 0
      "00000" when "001000101010010", -- t[4434] = 0
      "00000" when "001000101010011", -- t[4435] = 0
      "00000" when "001000101010100", -- t[4436] = 0
      "00000" when "001000101010101", -- t[4437] = 0
      "00000" when "001000101010110", -- t[4438] = 0
      "00000" when "001000101010111", -- t[4439] = 0
      "00000" when "001000101011000", -- t[4440] = 0
      "00000" when "001000101011001", -- t[4441] = 0
      "00000" when "001000101011010", -- t[4442] = 0
      "00000" when "001000101011011", -- t[4443] = 0
      "00000" when "001000101011100", -- t[4444] = 0
      "00000" when "001000101011101", -- t[4445] = 0
      "00000" when "001000101011110", -- t[4446] = 0
      "00000" when "001000101011111", -- t[4447] = 0
      "00000" when "001000101100000", -- t[4448] = 0
      "00000" when "001000101100001", -- t[4449] = 0
      "00000" when "001000101100010", -- t[4450] = 0
      "00000" when "001000101100011", -- t[4451] = 0
      "00000" when "001000101100100", -- t[4452] = 0
      "00000" when "001000101100101", -- t[4453] = 0
      "00000" when "001000101100110", -- t[4454] = 0
      "00000" when "001000101100111", -- t[4455] = 0
      "00000" when "001000101101000", -- t[4456] = 0
      "00000" when "001000101101001", -- t[4457] = 0
      "00000" when "001000101101010", -- t[4458] = 0
      "00000" when "001000101101011", -- t[4459] = 0
      "00000" when "001000101101100", -- t[4460] = 0
      "00000" when "001000101101101", -- t[4461] = 0
      "00000" when "001000101101110", -- t[4462] = 0
      "00000" when "001000101101111", -- t[4463] = 0
      "00000" when "001000101110000", -- t[4464] = 0
      "00000" when "001000101110001", -- t[4465] = 0
      "00000" when "001000101110010", -- t[4466] = 0
      "00000" when "001000101110011", -- t[4467] = 0
      "00000" when "001000101110100", -- t[4468] = 0
      "00000" when "001000101110101", -- t[4469] = 0
      "00000" when "001000101110110", -- t[4470] = 0
      "00000" when "001000101110111", -- t[4471] = 0
      "00000" when "001000101111000", -- t[4472] = 0
      "00000" when "001000101111001", -- t[4473] = 0
      "00000" when "001000101111010", -- t[4474] = 0
      "00000" when "001000101111011", -- t[4475] = 0
      "00000" when "001000101111100", -- t[4476] = 0
      "00000" when "001000101111101", -- t[4477] = 0
      "00000" when "001000101111110", -- t[4478] = 0
      "00000" when "001000101111111", -- t[4479] = 0
      "00000" when "001000110000000", -- t[4480] = 0
      "00000" when "001000110000001", -- t[4481] = 0
      "00000" when "001000110000010", -- t[4482] = 0
      "00000" when "001000110000011", -- t[4483] = 0
      "00000" when "001000110000100", -- t[4484] = 0
      "00000" when "001000110000101", -- t[4485] = 0
      "00000" when "001000110000110", -- t[4486] = 0
      "00000" when "001000110000111", -- t[4487] = 0
      "00000" when "001000110001000", -- t[4488] = 0
      "00000" when "001000110001001", -- t[4489] = 0
      "00000" when "001000110001010", -- t[4490] = 0
      "00000" when "001000110001011", -- t[4491] = 0
      "00000" when "001000110001100", -- t[4492] = 0
      "00000" when "001000110001101", -- t[4493] = 0
      "00000" when "001000110001110", -- t[4494] = 0
      "00000" when "001000110001111", -- t[4495] = 0
      "00000" when "001000110010000", -- t[4496] = 0
      "00000" when "001000110010001", -- t[4497] = 0
      "00000" when "001000110010010", -- t[4498] = 0
      "00000" when "001000110010011", -- t[4499] = 0
      "00000" when "001000110010100", -- t[4500] = 0
      "00000" when "001000110010101", -- t[4501] = 0
      "00000" when "001000110010110", -- t[4502] = 0
      "00000" when "001000110010111", -- t[4503] = 0
      "00000" when "001000110011000", -- t[4504] = 0
      "00000" when "001000110011001", -- t[4505] = 0
      "00000" when "001000110011010", -- t[4506] = 0
      "00000" when "001000110011011", -- t[4507] = 0
      "00000" when "001000110011100", -- t[4508] = 0
      "00000" when "001000110011101", -- t[4509] = 0
      "00000" when "001000110011110", -- t[4510] = 0
      "00000" when "001000110011111", -- t[4511] = 0
      "00000" when "001000110100000", -- t[4512] = 0
      "00000" when "001000110100001", -- t[4513] = 0
      "00000" when "001000110100010", -- t[4514] = 0
      "00000" when "001000110100011", -- t[4515] = 0
      "00000" when "001000110100100", -- t[4516] = 0
      "00000" when "001000110100101", -- t[4517] = 0
      "00000" when "001000110100110", -- t[4518] = 0
      "00000" when "001000110100111", -- t[4519] = 0
      "00000" when "001000110101000", -- t[4520] = 0
      "00000" when "001000110101001", -- t[4521] = 0
      "00000" when "001000110101010", -- t[4522] = 0
      "00000" when "001000110101011", -- t[4523] = 0
      "00000" when "001000110101100", -- t[4524] = 0
      "00000" when "001000110101101", -- t[4525] = 0
      "00000" when "001000110101110", -- t[4526] = 0
      "00000" when "001000110101111", -- t[4527] = 0
      "00000" when "001000110110000", -- t[4528] = 0
      "00000" when "001000110110001", -- t[4529] = 0
      "00000" when "001000110110010", -- t[4530] = 0
      "00000" when "001000110110011", -- t[4531] = 0
      "00000" when "001000110110100", -- t[4532] = 0
      "00000" when "001000110110101", -- t[4533] = 0
      "00000" when "001000110110110", -- t[4534] = 0
      "00000" when "001000110110111", -- t[4535] = 0
      "00000" when "001000110111000", -- t[4536] = 0
      "00000" when "001000110111001", -- t[4537] = 0
      "00000" when "001000110111010", -- t[4538] = 0
      "00000" when "001000110111011", -- t[4539] = 0
      "00000" when "001000110111100", -- t[4540] = 0
      "00000" when "001000110111101", -- t[4541] = 0
      "00000" when "001000110111110", -- t[4542] = 0
      "00000" when "001000110111111", -- t[4543] = 0
      "00000" when "001000111000000", -- t[4544] = 0
      "00000" when "001000111000001", -- t[4545] = 0
      "00000" when "001000111000010", -- t[4546] = 0
      "00000" when "001000111000011", -- t[4547] = 0
      "00000" when "001000111000100", -- t[4548] = 0
      "00000" when "001000111000101", -- t[4549] = 0
      "00000" when "001000111000110", -- t[4550] = 0
      "00000" when "001000111000111", -- t[4551] = 0
      "00000" when "001000111001000", -- t[4552] = 0
      "00000" when "001000111001001", -- t[4553] = 0
      "00000" when "001000111001010", -- t[4554] = 0
      "00000" when "001000111001011", -- t[4555] = 0
      "00000" when "001000111001100", -- t[4556] = 0
      "00000" when "001000111001101", -- t[4557] = 0
      "00000" when "001000111001110", -- t[4558] = 0
      "00000" when "001000111001111", -- t[4559] = 0
      "00000" when "001000111010000", -- t[4560] = 0
      "00000" when "001000111010001", -- t[4561] = 0
      "00000" when "001000111010010", -- t[4562] = 0
      "00000" when "001000111010011", -- t[4563] = 0
      "00000" when "001000111010100", -- t[4564] = 0
      "00000" when "001000111010101", -- t[4565] = 0
      "00000" when "001000111010110", -- t[4566] = 0
      "00000" when "001000111010111", -- t[4567] = 0
      "00000" when "001000111011000", -- t[4568] = 0
      "00000" when "001000111011001", -- t[4569] = 0
      "00000" when "001000111011010", -- t[4570] = 0
      "00000" when "001000111011011", -- t[4571] = 0
      "00000" when "001000111011100", -- t[4572] = 0
      "00000" when "001000111011101", -- t[4573] = 0
      "00000" when "001000111011110", -- t[4574] = 0
      "00000" when "001000111011111", -- t[4575] = 0
      "00000" when "001000111100000", -- t[4576] = 0
      "00000" when "001000111100001", -- t[4577] = 0
      "00000" when "001000111100010", -- t[4578] = 0
      "00000" when "001000111100011", -- t[4579] = 0
      "00000" when "001000111100100", -- t[4580] = 0
      "00000" when "001000111100101", -- t[4581] = 0
      "00000" when "001000111100110", -- t[4582] = 0
      "00000" when "001000111100111", -- t[4583] = 0
      "00000" when "001000111101000", -- t[4584] = 0
      "00000" when "001000111101001", -- t[4585] = 0
      "00000" when "001000111101010", -- t[4586] = 0
      "00000" when "001000111101011", -- t[4587] = 0
      "00000" when "001000111101100", -- t[4588] = 0
      "00000" when "001000111101101", -- t[4589] = 0
      "00000" when "001000111101110", -- t[4590] = 0
      "00000" when "001000111101111", -- t[4591] = 0
      "00000" when "001000111110000", -- t[4592] = 0
      "00000" when "001000111110001", -- t[4593] = 0
      "00000" when "001000111110010", -- t[4594] = 0
      "00000" when "001000111110011", -- t[4595] = 0
      "00000" when "001000111110100", -- t[4596] = 0
      "00000" when "001000111110101", -- t[4597] = 0
      "00000" when "001000111110110", -- t[4598] = 0
      "00000" when "001000111110111", -- t[4599] = 0
      "00000" when "001000111111000", -- t[4600] = 0
      "00000" when "001000111111001", -- t[4601] = 0
      "00000" when "001000111111010", -- t[4602] = 0
      "00000" when "001000111111011", -- t[4603] = 0
      "00000" when "001000111111100", -- t[4604] = 0
      "00000" when "001000111111101", -- t[4605] = 0
      "00000" when "001000111111110", -- t[4606] = 0
      "00000" when "001000111111111", -- t[4607] = 0
      "00000" when "001001000000000", -- t[4608] = 0
      "00000" when "001001000000001", -- t[4609] = 0
      "00000" when "001001000000010", -- t[4610] = 0
      "00000" when "001001000000011", -- t[4611] = 0
      "00000" when "001001000000100", -- t[4612] = 0
      "00000" when "001001000000101", -- t[4613] = 0
      "00000" when "001001000000110", -- t[4614] = 0
      "00000" when "001001000000111", -- t[4615] = 0
      "00000" when "001001000001000", -- t[4616] = 0
      "00000" when "001001000001001", -- t[4617] = 0
      "00000" when "001001000001010", -- t[4618] = 0
      "00000" when "001001000001011", -- t[4619] = 0
      "00000" when "001001000001100", -- t[4620] = 0
      "00000" when "001001000001101", -- t[4621] = 0
      "00000" when "001001000001110", -- t[4622] = 0
      "00000" when "001001000001111", -- t[4623] = 0
      "00000" when "001001000010000", -- t[4624] = 0
      "00000" when "001001000010001", -- t[4625] = 0
      "00000" when "001001000010010", -- t[4626] = 0
      "00000" when "001001000010011", -- t[4627] = 0
      "00000" when "001001000010100", -- t[4628] = 0
      "00000" when "001001000010101", -- t[4629] = 0
      "00000" when "001001000010110", -- t[4630] = 0
      "00000" when "001001000010111", -- t[4631] = 0
      "00000" when "001001000011000", -- t[4632] = 0
      "00000" when "001001000011001", -- t[4633] = 0
      "00000" when "001001000011010", -- t[4634] = 0
      "00000" when "001001000011011", -- t[4635] = 0
      "00000" when "001001000011100", -- t[4636] = 0
      "00000" when "001001000011101", -- t[4637] = 0
      "00000" when "001001000011110", -- t[4638] = 0
      "00000" when "001001000011111", -- t[4639] = 0
      "00000" when "001001000100000", -- t[4640] = 0
      "00000" when "001001000100001", -- t[4641] = 0
      "00000" when "001001000100010", -- t[4642] = 0
      "00000" when "001001000100011", -- t[4643] = 0
      "00000" when "001001000100100", -- t[4644] = 0
      "00000" when "001001000100101", -- t[4645] = 0
      "00000" when "001001000100110", -- t[4646] = 0
      "00000" when "001001000100111", -- t[4647] = 0
      "00000" when "001001000101000", -- t[4648] = 0
      "00000" when "001001000101001", -- t[4649] = 0
      "00000" when "001001000101010", -- t[4650] = 0
      "00000" when "001001000101011", -- t[4651] = 0
      "00000" when "001001000101100", -- t[4652] = 0
      "00000" when "001001000101101", -- t[4653] = 0
      "00000" when "001001000101110", -- t[4654] = 0
      "00000" when "001001000101111", -- t[4655] = 0
      "00000" when "001001000110000", -- t[4656] = 0
      "00000" when "001001000110001", -- t[4657] = 0
      "00000" when "001001000110010", -- t[4658] = 0
      "00000" when "001001000110011", -- t[4659] = 0
      "00000" when "001001000110100", -- t[4660] = 0
      "00000" when "001001000110101", -- t[4661] = 0
      "00000" when "001001000110110", -- t[4662] = 0
      "00000" when "001001000110111", -- t[4663] = 0
      "00000" when "001001000111000", -- t[4664] = 0
      "00000" when "001001000111001", -- t[4665] = 0
      "00000" when "001001000111010", -- t[4666] = 0
      "00000" when "001001000111011", -- t[4667] = 0
      "00000" when "001001000111100", -- t[4668] = 0
      "00000" when "001001000111101", -- t[4669] = 0
      "00000" when "001001000111110", -- t[4670] = 0
      "00000" when "001001000111111", -- t[4671] = 0
      "00000" when "001001001000000", -- t[4672] = 0
      "00000" when "001001001000001", -- t[4673] = 0
      "00000" when "001001001000010", -- t[4674] = 0
      "00000" when "001001001000011", -- t[4675] = 0
      "00000" when "001001001000100", -- t[4676] = 0
      "00000" when "001001001000101", -- t[4677] = 0
      "00000" when "001001001000110", -- t[4678] = 0
      "00000" when "001001001000111", -- t[4679] = 0
      "00000" when "001001001001000", -- t[4680] = 0
      "00000" when "001001001001001", -- t[4681] = 0
      "00000" when "001001001001010", -- t[4682] = 0
      "00000" when "001001001001011", -- t[4683] = 0
      "00000" when "001001001001100", -- t[4684] = 0
      "00000" when "001001001001101", -- t[4685] = 0
      "00000" when "001001001001110", -- t[4686] = 0
      "00000" when "001001001001111", -- t[4687] = 0
      "00000" when "001001001010000", -- t[4688] = 0
      "00000" when "001001001010001", -- t[4689] = 0
      "00000" when "001001001010010", -- t[4690] = 0
      "00000" when "001001001010011", -- t[4691] = 0
      "00000" when "001001001010100", -- t[4692] = 0
      "00000" when "001001001010101", -- t[4693] = 0
      "00000" when "001001001010110", -- t[4694] = 0
      "00000" when "001001001010111", -- t[4695] = 0
      "00000" when "001001001011000", -- t[4696] = 0
      "00000" when "001001001011001", -- t[4697] = 0
      "00000" when "001001001011010", -- t[4698] = 0
      "00000" when "001001001011011", -- t[4699] = 0
      "00000" when "001001001011100", -- t[4700] = 0
      "00000" when "001001001011101", -- t[4701] = 0
      "00000" when "001001001011110", -- t[4702] = 0
      "00000" when "001001001011111", -- t[4703] = 0
      "00000" when "001001001100000", -- t[4704] = 0
      "00000" when "001001001100001", -- t[4705] = 0
      "00000" when "001001001100010", -- t[4706] = 0
      "00000" when "001001001100011", -- t[4707] = 0
      "00000" when "001001001100100", -- t[4708] = 0
      "00000" when "001001001100101", -- t[4709] = 0
      "00000" when "001001001100110", -- t[4710] = 0
      "00000" when "001001001100111", -- t[4711] = 0
      "00000" when "001001001101000", -- t[4712] = 0
      "00000" when "001001001101001", -- t[4713] = 0
      "00000" when "001001001101010", -- t[4714] = 0
      "00000" when "001001001101011", -- t[4715] = 0
      "00000" when "001001001101100", -- t[4716] = 0
      "00000" when "001001001101101", -- t[4717] = 0
      "00000" when "001001001101110", -- t[4718] = 0
      "00000" when "001001001101111", -- t[4719] = 0
      "00000" when "001001001110000", -- t[4720] = 0
      "00000" when "001001001110001", -- t[4721] = 0
      "00000" when "001001001110010", -- t[4722] = 0
      "00000" when "001001001110011", -- t[4723] = 0
      "00000" when "001001001110100", -- t[4724] = 0
      "00000" when "001001001110101", -- t[4725] = 0
      "00000" when "001001001110110", -- t[4726] = 0
      "00000" when "001001001110111", -- t[4727] = 0
      "00000" when "001001001111000", -- t[4728] = 0
      "00000" when "001001001111001", -- t[4729] = 0
      "00000" when "001001001111010", -- t[4730] = 0
      "00000" when "001001001111011", -- t[4731] = 0
      "00000" when "001001001111100", -- t[4732] = 0
      "00000" when "001001001111101", -- t[4733] = 0
      "00000" when "001001001111110", -- t[4734] = 0
      "00000" when "001001001111111", -- t[4735] = 0
      "00000" when "001001010000000", -- t[4736] = 0
      "00000" when "001001010000001", -- t[4737] = 0
      "00000" when "001001010000010", -- t[4738] = 0
      "00000" when "001001010000011", -- t[4739] = 0
      "00000" when "001001010000100", -- t[4740] = 0
      "00000" when "001001010000101", -- t[4741] = 0
      "00000" when "001001010000110", -- t[4742] = 0
      "00000" when "001001010000111", -- t[4743] = 0
      "00000" when "001001010001000", -- t[4744] = 0
      "00000" when "001001010001001", -- t[4745] = 0
      "00000" when "001001010001010", -- t[4746] = 0
      "00000" when "001001010001011", -- t[4747] = 0
      "00000" when "001001010001100", -- t[4748] = 0
      "00000" when "001001010001101", -- t[4749] = 0
      "00000" when "001001010001110", -- t[4750] = 0
      "00000" when "001001010001111", -- t[4751] = 0
      "00000" when "001001010010000", -- t[4752] = 0
      "00000" when "001001010010001", -- t[4753] = 0
      "00000" when "001001010010010", -- t[4754] = 0
      "00000" when "001001010010011", -- t[4755] = 0
      "00000" when "001001010010100", -- t[4756] = 0
      "00000" when "001001010010101", -- t[4757] = 0
      "00000" when "001001010010110", -- t[4758] = 0
      "00000" when "001001010010111", -- t[4759] = 0
      "00000" when "001001010011000", -- t[4760] = 0
      "00000" when "001001010011001", -- t[4761] = 0
      "00000" when "001001010011010", -- t[4762] = 0
      "00000" when "001001010011011", -- t[4763] = 0
      "00000" when "001001010011100", -- t[4764] = 0
      "00000" when "001001010011101", -- t[4765] = 0
      "00000" when "001001010011110", -- t[4766] = 0
      "00000" when "001001010011111", -- t[4767] = 0
      "00000" when "001001010100000", -- t[4768] = 0
      "00000" when "001001010100001", -- t[4769] = 0
      "00000" when "001001010100010", -- t[4770] = 0
      "00000" when "001001010100011", -- t[4771] = 0
      "00000" when "001001010100100", -- t[4772] = 0
      "00000" when "001001010100101", -- t[4773] = 0
      "00000" when "001001010100110", -- t[4774] = 0
      "00000" when "001001010100111", -- t[4775] = 0
      "00000" when "001001010101000", -- t[4776] = 0
      "00000" when "001001010101001", -- t[4777] = 0
      "00000" when "001001010101010", -- t[4778] = 0
      "00000" when "001001010101011", -- t[4779] = 0
      "00000" when "001001010101100", -- t[4780] = 0
      "00000" when "001001010101101", -- t[4781] = 0
      "00000" when "001001010101110", -- t[4782] = 0
      "00000" when "001001010101111", -- t[4783] = 0
      "00000" when "001001010110000", -- t[4784] = 0
      "00000" when "001001010110001", -- t[4785] = 0
      "00000" when "001001010110010", -- t[4786] = 0
      "00000" when "001001010110011", -- t[4787] = 0
      "00000" when "001001010110100", -- t[4788] = 0
      "00000" when "001001010110101", -- t[4789] = 0
      "00000" when "001001010110110", -- t[4790] = 0
      "00000" when "001001010110111", -- t[4791] = 0
      "00000" when "001001010111000", -- t[4792] = 0
      "00000" when "001001010111001", -- t[4793] = 0
      "00000" when "001001010111010", -- t[4794] = 0
      "00000" when "001001010111011", -- t[4795] = 0
      "00000" when "001001010111100", -- t[4796] = 0
      "00000" when "001001010111101", -- t[4797] = 0
      "00000" when "001001010111110", -- t[4798] = 0
      "00000" when "001001010111111", -- t[4799] = 0
      "00000" when "001001011000000", -- t[4800] = 0
      "00000" when "001001011000001", -- t[4801] = 0
      "00000" when "001001011000010", -- t[4802] = 0
      "00000" when "001001011000011", -- t[4803] = 0
      "00000" when "001001011000100", -- t[4804] = 0
      "00000" when "001001011000101", -- t[4805] = 0
      "00000" when "001001011000110", -- t[4806] = 0
      "00000" when "001001011000111", -- t[4807] = 0
      "00000" when "001001011001000", -- t[4808] = 0
      "00000" when "001001011001001", -- t[4809] = 0
      "00000" when "001001011001010", -- t[4810] = 0
      "00000" when "001001011001011", -- t[4811] = 0
      "00000" when "001001011001100", -- t[4812] = 0
      "00000" when "001001011001101", -- t[4813] = 0
      "00000" when "001001011001110", -- t[4814] = 0
      "00000" when "001001011001111", -- t[4815] = 0
      "00000" when "001001011010000", -- t[4816] = 0
      "00000" when "001001011010001", -- t[4817] = 0
      "00000" when "001001011010010", -- t[4818] = 0
      "00000" when "001001011010011", -- t[4819] = 0
      "00000" when "001001011010100", -- t[4820] = 0
      "00000" when "001001011010101", -- t[4821] = 0
      "00000" when "001001011010110", -- t[4822] = 0
      "00000" when "001001011010111", -- t[4823] = 0
      "00000" when "001001011011000", -- t[4824] = 0
      "00000" when "001001011011001", -- t[4825] = 0
      "00000" when "001001011011010", -- t[4826] = 0
      "00000" when "001001011011011", -- t[4827] = 0
      "00000" when "001001011011100", -- t[4828] = 0
      "00000" when "001001011011101", -- t[4829] = 0
      "00000" when "001001011011110", -- t[4830] = 0
      "00000" when "001001011011111", -- t[4831] = 0
      "00000" when "001001011100000", -- t[4832] = 0
      "00000" when "001001011100001", -- t[4833] = 0
      "00000" when "001001011100010", -- t[4834] = 0
      "00000" when "001001011100011", -- t[4835] = 0
      "00000" when "001001011100100", -- t[4836] = 0
      "00000" when "001001011100101", -- t[4837] = 0
      "00000" when "001001011100110", -- t[4838] = 0
      "00000" when "001001011100111", -- t[4839] = 0
      "00000" when "001001011101000", -- t[4840] = 0
      "00000" when "001001011101001", -- t[4841] = 0
      "00000" when "001001011101010", -- t[4842] = 0
      "00000" when "001001011101011", -- t[4843] = 0
      "00000" when "001001011101100", -- t[4844] = 0
      "00000" when "001001011101101", -- t[4845] = 0
      "00000" when "001001011101110", -- t[4846] = 0
      "00000" when "001001011101111", -- t[4847] = 0
      "00000" when "001001011110000", -- t[4848] = 0
      "00000" when "001001011110001", -- t[4849] = 0
      "00000" when "001001011110010", -- t[4850] = 0
      "00000" when "001001011110011", -- t[4851] = 0
      "00000" when "001001011110100", -- t[4852] = 0
      "00000" when "001001011110101", -- t[4853] = 0
      "00000" when "001001011110110", -- t[4854] = 0
      "00000" when "001001011110111", -- t[4855] = 0
      "00000" when "001001011111000", -- t[4856] = 0
      "00000" when "001001011111001", -- t[4857] = 0
      "00000" when "001001011111010", -- t[4858] = 0
      "00000" when "001001011111011", -- t[4859] = 0
      "00000" when "001001011111100", -- t[4860] = 0
      "00000" when "001001011111101", -- t[4861] = 0
      "00000" when "001001011111110", -- t[4862] = 0
      "00000" when "001001011111111", -- t[4863] = 0
      "00000" when "001001100000000", -- t[4864] = 0
      "00000" when "001001100000001", -- t[4865] = 0
      "00000" when "001001100000010", -- t[4866] = 0
      "00000" when "001001100000011", -- t[4867] = 0
      "00000" when "001001100000100", -- t[4868] = 0
      "00000" when "001001100000101", -- t[4869] = 0
      "00000" when "001001100000110", -- t[4870] = 0
      "00000" when "001001100000111", -- t[4871] = 0
      "00000" when "001001100001000", -- t[4872] = 0
      "00000" when "001001100001001", -- t[4873] = 0
      "00000" when "001001100001010", -- t[4874] = 0
      "00000" when "001001100001011", -- t[4875] = 0
      "00000" when "001001100001100", -- t[4876] = 0
      "00000" when "001001100001101", -- t[4877] = 0
      "00000" when "001001100001110", -- t[4878] = 0
      "00000" when "001001100001111", -- t[4879] = 0
      "00000" when "001001100010000", -- t[4880] = 0
      "00000" when "001001100010001", -- t[4881] = 0
      "00000" when "001001100010010", -- t[4882] = 0
      "00000" when "001001100010011", -- t[4883] = 0
      "00000" when "001001100010100", -- t[4884] = 0
      "00000" when "001001100010101", -- t[4885] = 0
      "00000" when "001001100010110", -- t[4886] = 0
      "00000" when "001001100010111", -- t[4887] = 0
      "00000" when "001001100011000", -- t[4888] = 0
      "00000" when "001001100011001", -- t[4889] = 0
      "00000" when "001001100011010", -- t[4890] = 0
      "00000" when "001001100011011", -- t[4891] = 0
      "00000" when "001001100011100", -- t[4892] = 0
      "00000" when "001001100011101", -- t[4893] = 0
      "00000" when "001001100011110", -- t[4894] = 0
      "00000" when "001001100011111", -- t[4895] = 0
      "00000" when "001001100100000", -- t[4896] = 0
      "00000" when "001001100100001", -- t[4897] = 0
      "00000" when "001001100100010", -- t[4898] = 0
      "00000" when "001001100100011", -- t[4899] = 0
      "00000" when "001001100100100", -- t[4900] = 0
      "00000" when "001001100100101", -- t[4901] = 0
      "00000" when "001001100100110", -- t[4902] = 0
      "00000" when "001001100100111", -- t[4903] = 0
      "00000" when "001001100101000", -- t[4904] = 0
      "00000" when "001001100101001", -- t[4905] = 0
      "00000" when "001001100101010", -- t[4906] = 0
      "00000" when "001001100101011", -- t[4907] = 0
      "00000" when "001001100101100", -- t[4908] = 0
      "00000" when "001001100101101", -- t[4909] = 0
      "00000" when "001001100101110", -- t[4910] = 0
      "00000" when "001001100101111", -- t[4911] = 0
      "00000" when "001001100110000", -- t[4912] = 0
      "00000" when "001001100110001", -- t[4913] = 0
      "00000" when "001001100110010", -- t[4914] = 0
      "00000" when "001001100110011", -- t[4915] = 0
      "00000" when "001001100110100", -- t[4916] = 0
      "00000" when "001001100110101", -- t[4917] = 0
      "00000" when "001001100110110", -- t[4918] = 0
      "00000" when "001001100110111", -- t[4919] = 0
      "00000" when "001001100111000", -- t[4920] = 0
      "00000" when "001001100111001", -- t[4921] = 0
      "00000" when "001001100111010", -- t[4922] = 0
      "00000" when "001001100111011", -- t[4923] = 0
      "00000" when "001001100111100", -- t[4924] = 0
      "00000" when "001001100111101", -- t[4925] = 0
      "00000" when "001001100111110", -- t[4926] = 0
      "00000" when "001001100111111", -- t[4927] = 0
      "00000" when "001001101000000", -- t[4928] = 0
      "00000" when "001001101000001", -- t[4929] = 0
      "00000" when "001001101000010", -- t[4930] = 0
      "00000" when "001001101000011", -- t[4931] = 0
      "00000" when "001001101000100", -- t[4932] = 0
      "00000" when "001001101000101", -- t[4933] = 0
      "00000" when "001001101000110", -- t[4934] = 0
      "00000" when "001001101000111", -- t[4935] = 0
      "00000" when "001001101001000", -- t[4936] = 0
      "00000" when "001001101001001", -- t[4937] = 0
      "00000" when "001001101001010", -- t[4938] = 0
      "00000" when "001001101001011", -- t[4939] = 0
      "00000" when "001001101001100", -- t[4940] = 0
      "00000" when "001001101001101", -- t[4941] = 0
      "00000" when "001001101001110", -- t[4942] = 0
      "00000" when "001001101001111", -- t[4943] = 0
      "00000" when "001001101010000", -- t[4944] = 0
      "00000" when "001001101010001", -- t[4945] = 0
      "00000" when "001001101010010", -- t[4946] = 0
      "00000" when "001001101010011", -- t[4947] = 0
      "00000" when "001001101010100", -- t[4948] = 0
      "00000" when "001001101010101", -- t[4949] = 0
      "00000" when "001001101010110", -- t[4950] = 0
      "00000" when "001001101010111", -- t[4951] = 0
      "00000" when "001001101011000", -- t[4952] = 0
      "00000" when "001001101011001", -- t[4953] = 0
      "00000" when "001001101011010", -- t[4954] = 0
      "00000" when "001001101011011", -- t[4955] = 0
      "00000" when "001001101011100", -- t[4956] = 0
      "00000" when "001001101011101", -- t[4957] = 0
      "00000" when "001001101011110", -- t[4958] = 0
      "00000" when "001001101011111", -- t[4959] = 0
      "00000" when "001001101100000", -- t[4960] = 0
      "00000" when "001001101100001", -- t[4961] = 0
      "00000" when "001001101100010", -- t[4962] = 0
      "00000" when "001001101100011", -- t[4963] = 0
      "00000" when "001001101100100", -- t[4964] = 0
      "00000" when "001001101100101", -- t[4965] = 0
      "00000" when "001001101100110", -- t[4966] = 0
      "00000" when "001001101100111", -- t[4967] = 0
      "00000" when "001001101101000", -- t[4968] = 0
      "00000" when "001001101101001", -- t[4969] = 0
      "00000" when "001001101101010", -- t[4970] = 0
      "00000" when "001001101101011", -- t[4971] = 0
      "00000" when "001001101101100", -- t[4972] = 0
      "00000" when "001001101101101", -- t[4973] = 0
      "00000" when "001001101101110", -- t[4974] = 0
      "00000" when "001001101101111", -- t[4975] = 0
      "00000" when "001001101110000", -- t[4976] = 0
      "00000" when "001001101110001", -- t[4977] = 0
      "00000" when "001001101110010", -- t[4978] = 0
      "00000" when "001001101110011", -- t[4979] = 0
      "00000" when "001001101110100", -- t[4980] = 0
      "00000" when "001001101110101", -- t[4981] = 0
      "00000" when "001001101110110", -- t[4982] = 0
      "00000" when "001001101110111", -- t[4983] = 0
      "00000" when "001001101111000", -- t[4984] = 0
      "00000" when "001001101111001", -- t[4985] = 0
      "00000" when "001001101111010", -- t[4986] = 0
      "00000" when "001001101111011", -- t[4987] = 0
      "00000" when "001001101111100", -- t[4988] = 0
      "00000" when "001001101111101", -- t[4989] = 0
      "00000" when "001001101111110", -- t[4990] = 0
      "00000" when "001001101111111", -- t[4991] = 0
      "00000" when "001001110000000", -- t[4992] = 0
      "00000" when "001001110000001", -- t[4993] = 0
      "00000" when "001001110000010", -- t[4994] = 0
      "00000" when "001001110000011", -- t[4995] = 0
      "00000" when "001001110000100", -- t[4996] = 0
      "00000" when "001001110000101", -- t[4997] = 0
      "00000" when "001001110000110", -- t[4998] = 0
      "00000" when "001001110000111", -- t[4999] = 0
      "00000" when "001001110001000", -- t[5000] = 0
      "00000" when "001001110001001", -- t[5001] = 0
      "00000" when "001001110001010", -- t[5002] = 0
      "00000" when "001001110001011", -- t[5003] = 0
      "00000" when "001001110001100", -- t[5004] = 0
      "00000" when "001001110001101", -- t[5005] = 0
      "00000" when "001001110001110", -- t[5006] = 0
      "00000" when "001001110001111", -- t[5007] = 0
      "00000" when "001001110010000", -- t[5008] = 0
      "00000" when "001001110010001", -- t[5009] = 0
      "00000" when "001001110010010", -- t[5010] = 0
      "00000" when "001001110010011", -- t[5011] = 0
      "00000" when "001001110010100", -- t[5012] = 0
      "00000" when "001001110010101", -- t[5013] = 0
      "00000" when "001001110010110", -- t[5014] = 0
      "00000" when "001001110010111", -- t[5015] = 0
      "00000" when "001001110011000", -- t[5016] = 0
      "00000" when "001001110011001", -- t[5017] = 0
      "00000" when "001001110011010", -- t[5018] = 0
      "00000" when "001001110011011", -- t[5019] = 0
      "00000" when "001001110011100", -- t[5020] = 0
      "00000" when "001001110011101", -- t[5021] = 0
      "00000" when "001001110011110", -- t[5022] = 0
      "00000" when "001001110011111", -- t[5023] = 0
      "00000" when "001001110100000", -- t[5024] = 0
      "00000" when "001001110100001", -- t[5025] = 0
      "00000" when "001001110100010", -- t[5026] = 0
      "00000" when "001001110100011", -- t[5027] = 0
      "00000" when "001001110100100", -- t[5028] = 0
      "00000" when "001001110100101", -- t[5029] = 0
      "00000" when "001001110100110", -- t[5030] = 0
      "00000" when "001001110100111", -- t[5031] = 0
      "00000" when "001001110101000", -- t[5032] = 0
      "00000" when "001001110101001", -- t[5033] = 0
      "00000" when "001001110101010", -- t[5034] = 0
      "00000" when "001001110101011", -- t[5035] = 0
      "00000" when "001001110101100", -- t[5036] = 0
      "00000" when "001001110101101", -- t[5037] = 0
      "00000" when "001001110101110", -- t[5038] = 0
      "00000" when "001001110101111", -- t[5039] = 0
      "00000" when "001001110110000", -- t[5040] = 0
      "00000" when "001001110110001", -- t[5041] = 0
      "00000" when "001001110110010", -- t[5042] = 0
      "00000" when "001001110110011", -- t[5043] = 0
      "00000" when "001001110110100", -- t[5044] = 0
      "00000" when "001001110110101", -- t[5045] = 0
      "00000" when "001001110110110", -- t[5046] = 0
      "00000" when "001001110110111", -- t[5047] = 0
      "00000" when "001001110111000", -- t[5048] = 0
      "00000" when "001001110111001", -- t[5049] = 0
      "00000" when "001001110111010", -- t[5050] = 0
      "00000" when "001001110111011", -- t[5051] = 0
      "00000" when "001001110111100", -- t[5052] = 0
      "00000" when "001001110111101", -- t[5053] = 0
      "00000" when "001001110111110", -- t[5054] = 0
      "00000" when "001001110111111", -- t[5055] = 0
      "00000" when "001001111000000", -- t[5056] = 0
      "00000" when "001001111000001", -- t[5057] = 0
      "00000" when "001001111000010", -- t[5058] = 0
      "00000" when "001001111000011", -- t[5059] = 0
      "00000" when "001001111000100", -- t[5060] = 0
      "00000" when "001001111000101", -- t[5061] = 0
      "00000" when "001001111000110", -- t[5062] = 0
      "00000" when "001001111000111", -- t[5063] = 0
      "00000" when "001001111001000", -- t[5064] = 0
      "00000" when "001001111001001", -- t[5065] = 0
      "00000" when "001001111001010", -- t[5066] = 0
      "00000" when "001001111001011", -- t[5067] = 0
      "00000" when "001001111001100", -- t[5068] = 0
      "00000" when "001001111001101", -- t[5069] = 0
      "00000" when "001001111001110", -- t[5070] = 0
      "00000" when "001001111001111", -- t[5071] = 0
      "00000" when "001001111010000", -- t[5072] = 0
      "00000" when "001001111010001", -- t[5073] = 0
      "00000" when "001001111010010", -- t[5074] = 0
      "00000" when "001001111010011", -- t[5075] = 0
      "00000" when "001001111010100", -- t[5076] = 0
      "00000" when "001001111010101", -- t[5077] = 0
      "00000" when "001001111010110", -- t[5078] = 0
      "00000" when "001001111010111", -- t[5079] = 0
      "00000" when "001001111011000", -- t[5080] = 0
      "00000" when "001001111011001", -- t[5081] = 0
      "00000" when "001001111011010", -- t[5082] = 0
      "00000" when "001001111011011", -- t[5083] = 0
      "00000" when "001001111011100", -- t[5084] = 0
      "00000" when "001001111011101", -- t[5085] = 0
      "00000" when "001001111011110", -- t[5086] = 0
      "00000" when "001001111011111", -- t[5087] = 0
      "00000" when "001001111100000", -- t[5088] = 0
      "00000" when "001001111100001", -- t[5089] = 0
      "00000" when "001001111100010", -- t[5090] = 0
      "00000" when "001001111100011", -- t[5091] = 0
      "00000" when "001001111100100", -- t[5092] = 0
      "00000" when "001001111100101", -- t[5093] = 0
      "00000" when "001001111100110", -- t[5094] = 0
      "00000" when "001001111100111", -- t[5095] = 0
      "00000" when "001001111101000", -- t[5096] = 0
      "00000" when "001001111101001", -- t[5097] = 0
      "00000" when "001001111101010", -- t[5098] = 0
      "00000" when "001001111101011", -- t[5099] = 0
      "00000" when "001001111101100", -- t[5100] = 0
      "00000" when "001001111101101", -- t[5101] = 0
      "00000" when "001001111101110", -- t[5102] = 0
      "00000" when "001001111101111", -- t[5103] = 0
      "00000" when "001001111110000", -- t[5104] = 0
      "00000" when "001001111110001", -- t[5105] = 0
      "00000" when "001001111110010", -- t[5106] = 0
      "00000" when "001001111110011", -- t[5107] = 0
      "00000" when "001001111110100", -- t[5108] = 0
      "00000" when "001001111110101", -- t[5109] = 0
      "00000" when "001001111110110", -- t[5110] = 0
      "00000" when "001001111110111", -- t[5111] = 0
      "00000" when "001001111111000", -- t[5112] = 0
      "00000" when "001001111111001", -- t[5113] = 0
      "00000" when "001001111111010", -- t[5114] = 0
      "00000" when "001001111111011", -- t[5115] = 0
      "00000" when "001001111111100", -- t[5116] = 0
      "00000" when "001001111111101", -- t[5117] = 0
      "00000" when "001001111111110", -- t[5118] = 0
      "00000" when "001001111111111", -- t[5119] = 0
      "00000" when "001010000000000", -- t[5120] = 0
      "00000" when "001010000000001", -- t[5121] = 0
      "00000" when "001010000000010", -- t[5122] = 0
      "00000" when "001010000000011", -- t[5123] = 0
      "00000" when "001010000000100", -- t[5124] = 0
      "00000" when "001010000000101", -- t[5125] = 0
      "00000" when "001010000000110", -- t[5126] = 0
      "00000" when "001010000000111", -- t[5127] = 0
      "00000" when "001010000001000", -- t[5128] = 0
      "00000" when "001010000001001", -- t[5129] = 0
      "00000" when "001010000001010", -- t[5130] = 0
      "00000" when "001010000001011", -- t[5131] = 0
      "00000" when "001010000001100", -- t[5132] = 0
      "00000" when "001010000001101", -- t[5133] = 0
      "00000" when "001010000001110", -- t[5134] = 0
      "00000" when "001010000001111", -- t[5135] = 0
      "00000" when "001010000010000", -- t[5136] = 0
      "00000" when "001010000010001", -- t[5137] = 0
      "00000" when "001010000010010", -- t[5138] = 0
      "00000" when "001010000010011", -- t[5139] = 0
      "00000" when "001010000010100", -- t[5140] = 0
      "00000" when "001010000010101", -- t[5141] = 0
      "00000" when "001010000010110", -- t[5142] = 0
      "00000" when "001010000010111", -- t[5143] = 0
      "00000" when "001010000011000", -- t[5144] = 0
      "00000" when "001010000011001", -- t[5145] = 0
      "00000" when "001010000011010", -- t[5146] = 0
      "00000" when "001010000011011", -- t[5147] = 0
      "00000" when "001010000011100", -- t[5148] = 0
      "00000" when "001010000011101", -- t[5149] = 0
      "00000" when "001010000011110", -- t[5150] = 0
      "00000" when "001010000011111", -- t[5151] = 0
      "00000" when "001010000100000", -- t[5152] = 0
      "00000" when "001010000100001", -- t[5153] = 0
      "00000" when "001010000100010", -- t[5154] = 0
      "00000" when "001010000100011", -- t[5155] = 0
      "00000" when "001010000100100", -- t[5156] = 0
      "00000" when "001010000100101", -- t[5157] = 0
      "00000" when "001010000100110", -- t[5158] = 0
      "00000" when "001010000100111", -- t[5159] = 0
      "00000" when "001010000101000", -- t[5160] = 0
      "00000" when "001010000101001", -- t[5161] = 0
      "00000" when "001010000101010", -- t[5162] = 0
      "00000" when "001010000101011", -- t[5163] = 0
      "00000" when "001010000101100", -- t[5164] = 0
      "00000" when "001010000101101", -- t[5165] = 0
      "00000" when "001010000101110", -- t[5166] = 0
      "00000" when "001010000101111", -- t[5167] = 0
      "00000" when "001010000110000", -- t[5168] = 0
      "00000" when "001010000110001", -- t[5169] = 0
      "00000" when "001010000110010", -- t[5170] = 0
      "00000" when "001010000110011", -- t[5171] = 0
      "00000" when "001010000110100", -- t[5172] = 0
      "00000" when "001010000110101", -- t[5173] = 0
      "00000" when "001010000110110", -- t[5174] = 0
      "00000" when "001010000110111", -- t[5175] = 0
      "00000" when "001010000111000", -- t[5176] = 0
      "00000" when "001010000111001", -- t[5177] = 0
      "00000" when "001010000111010", -- t[5178] = 0
      "00000" when "001010000111011", -- t[5179] = 0
      "00000" when "001010000111100", -- t[5180] = 0
      "00000" when "001010000111101", -- t[5181] = 0
      "00000" when "001010000111110", -- t[5182] = 0
      "00000" when "001010000111111", -- t[5183] = 0
      "00000" when "001010001000000", -- t[5184] = 0
      "00000" when "001010001000001", -- t[5185] = 0
      "00000" when "001010001000010", -- t[5186] = 0
      "00000" when "001010001000011", -- t[5187] = 0
      "00000" when "001010001000100", -- t[5188] = 0
      "00000" when "001010001000101", -- t[5189] = 0
      "00000" when "001010001000110", -- t[5190] = 0
      "00000" when "001010001000111", -- t[5191] = 0
      "00000" when "001010001001000", -- t[5192] = 0
      "00000" when "001010001001001", -- t[5193] = 0
      "00000" when "001010001001010", -- t[5194] = 0
      "00000" when "001010001001011", -- t[5195] = 0
      "00000" when "001010001001100", -- t[5196] = 0
      "00000" when "001010001001101", -- t[5197] = 0
      "00000" when "001010001001110", -- t[5198] = 0
      "00000" when "001010001001111", -- t[5199] = 0
      "00000" when "001010001010000", -- t[5200] = 0
      "00000" when "001010001010001", -- t[5201] = 0
      "00000" when "001010001010010", -- t[5202] = 0
      "00000" when "001010001010011", -- t[5203] = 0
      "00000" when "001010001010100", -- t[5204] = 0
      "00000" when "001010001010101", -- t[5205] = 0
      "00000" when "001010001010110", -- t[5206] = 0
      "00000" when "001010001010111", -- t[5207] = 0
      "00000" when "001010001011000", -- t[5208] = 0
      "00000" when "001010001011001", -- t[5209] = 0
      "00000" when "001010001011010", -- t[5210] = 0
      "00000" when "001010001011011", -- t[5211] = 0
      "00000" when "001010001011100", -- t[5212] = 0
      "00000" when "001010001011101", -- t[5213] = 0
      "00000" when "001010001011110", -- t[5214] = 0
      "00000" when "001010001011111", -- t[5215] = 0
      "00000" when "001010001100000", -- t[5216] = 0
      "00000" when "001010001100001", -- t[5217] = 0
      "00000" when "001010001100010", -- t[5218] = 0
      "00000" when "001010001100011", -- t[5219] = 0
      "00000" when "001010001100100", -- t[5220] = 0
      "00000" when "001010001100101", -- t[5221] = 0
      "00000" when "001010001100110", -- t[5222] = 0
      "00000" when "001010001100111", -- t[5223] = 0
      "00000" when "001010001101000", -- t[5224] = 0
      "00000" when "001010001101001", -- t[5225] = 0
      "00000" when "001010001101010", -- t[5226] = 0
      "00000" when "001010001101011", -- t[5227] = 0
      "00000" when "001010001101100", -- t[5228] = 0
      "00000" when "001010001101101", -- t[5229] = 0
      "00000" when "001010001101110", -- t[5230] = 0
      "00000" when "001010001101111", -- t[5231] = 0
      "00000" when "001010001110000", -- t[5232] = 0
      "00000" when "001010001110001", -- t[5233] = 0
      "00000" when "001010001110010", -- t[5234] = 0
      "00000" when "001010001110011", -- t[5235] = 0
      "00000" when "001010001110100", -- t[5236] = 0
      "00000" when "001010001110101", -- t[5237] = 0
      "00000" when "001010001110110", -- t[5238] = 0
      "00000" when "001010001110111", -- t[5239] = 0
      "00000" when "001010001111000", -- t[5240] = 0
      "00000" when "001010001111001", -- t[5241] = 0
      "00000" when "001010001111010", -- t[5242] = 0
      "00000" when "001010001111011", -- t[5243] = 0
      "00000" when "001010001111100", -- t[5244] = 0
      "00000" when "001010001111101", -- t[5245] = 0
      "00000" when "001010001111110", -- t[5246] = 0
      "00000" when "001010001111111", -- t[5247] = 0
      "00000" when "001010010000000", -- t[5248] = 0
      "00000" when "001010010000001", -- t[5249] = 0
      "00000" when "001010010000010", -- t[5250] = 0
      "00000" when "001010010000011", -- t[5251] = 0
      "00000" when "001010010000100", -- t[5252] = 0
      "00000" when "001010010000101", -- t[5253] = 0
      "00000" when "001010010000110", -- t[5254] = 0
      "00000" when "001010010000111", -- t[5255] = 0
      "00000" when "001010010001000", -- t[5256] = 0
      "00000" when "001010010001001", -- t[5257] = 0
      "00000" when "001010010001010", -- t[5258] = 0
      "00000" when "001010010001011", -- t[5259] = 0
      "00000" when "001010010001100", -- t[5260] = 0
      "00000" when "001010010001101", -- t[5261] = 0
      "00000" when "001010010001110", -- t[5262] = 0
      "00000" when "001010010001111", -- t[5263] = 0
      "00000" when "001010010010000", -- t[5264] = 0
      "00000" when "001010010010001", -- t[5265] = 0
      "00000" when "001010010010010", -- t[5266] = 0
      "00000" when "001010010010011", -- t[5267] = 0
      "00000" when "001010010010100", -- t[5268] = 0
      "00000" when "001010010010101", -- t[5269] = 0
      "00000" when "001010010010110", -- t[5270] = 0
      "00000" when "001010010010111", -- t[5271] = 0
      "00000" when "001010010011000", -- t[5272] = 0
      "00000" when "001010010011001", -- t[5273] = 0
      "00000" when "001010010011010", -- t[5274] = 0
      "00000" when "001010010011011", -- t[5275] = 0
      "00000" when "001010010011100", -- t[5276] = 0
      "00000" when "001010010011101", -- t[5277] = 0
      "00000" when "001010010011110", -- t[5278] = 0
      "00000" when "001010010011111", -- t[5279] = 0
      "00000" when "001010010100000", -- t[5280] = 0
      "00000" when "001010010100001", -- t[5281] = 0
      "00000" when "001010010100010", -- t[5282] = 0
      "00000" when "001010010100011", -- t[5283] = 0
      "00000" when "001010010100100", -- t[5284] = 0
      "00000" when "001010010100101", -- t[5285] = 0
      "00000" when "001010010100110", -- t[5286] = 0
      "00000" when "001010010100111", -- t[5287] = 0
      "00000" when "001010010101000", -- t[5288] = 0
      "00000" when "001010010101001", -- t[5289] = 0
      "00000" when "001010010101010", -- t[5290] = 0
      "00000" when "001010010101011", -- t[5291] = 0
      "00000" when "001010010101100", -- t[5292] = 0
      "00000" when "001010010101101", -- t[5293] = 0
      "00000" when "001010010101110", -- t[5294] = 0
      "00000" when "001010010101111", -- t[5295] = 0
      "00000" when "001010010110000", -- t[5296] = 0
      "00000" when "001010010110001", -- t[5297] = 0
      "00000" when "001010010110010", -- t[5298] = 0
      "00000" when "001010010110011", -- t[5299] = 0
      "00000" when "001010010110100", -- t[5300] = 0
      "00000" when "001010010110101", -- t[5301] = 0
      "00000" when "001010010110110", -- t[5302] = 0
      "00000" when "001010010110111", -- t[5303] = 0
      "00000" when "001010010111000", -- t[5304] = 0
      "00000" when "001010010111001", -- t[5305] = 0
      "00000" when "001010010111010", -- t[5306] = 0
      "00000" when "001010010111011", -- t[5307] = 0
      "00000" when "001010010111100", -- t[5308] = 0
      "00000" when "001010010111101", -- t[5309] = 0
      "00000" when "001010010111110", -- t[5310] = 0
      "00000" when "001010010111111", -- t[5311] = 0
      "00000" when "001010011000000", -- t[5312] = 0
      "00000" when "001010011000001", -- t[5313] = 0
      "00000" when "001010011000010", -- t[5314] = 0
      "00000" when "001010011000011", -- t[5315] = 0
      "00000" when "001010011000100", -- t[5316] = 0
      "00000" when "001010011000101", -- t[5317] = 0
      "00000" when "001010011000110", -- t[5318] = 0
      "00000" when "001010011000111", -- t[5319] = 0
      "00000" when "001010011001000", -- t[5320] = 0
      "00000" when "001010011001001", -- t[5321] = 0
      "00000" when "001010011001010", -- t[5322] = 0
      "00000" when "001010011001011", -- t[5323] = 0
      "00000" when "001010011001100", -- t[5324] = 0
      "00000" when "001010011001101", -- t[5325] = 0
      "00000" when "001010011001110", -- t[5326] = 0
      "00000" when "001010011001111", -- t[5327] = 0
      "00000" when "001010011010000", -- t[5328] = 0
      "00000" when "001010011010001", -- t[5329] = 0
      "00000" when "001010011010010", -- t[5330] = 0
      "00000" when "001010011010011", -- t[5331] = 0
      "00000" when "001010011010100", -- t[5332] = 0
      "00000" when "001010011010101", -- t[5333] = 0
      "00000" when "001010011010110", -- t[5334] = 0
      "00000" when "001010011010111", -- t[5335] = 0
      "00000" when "001010011011000", -- t[5336] = 0
      "00000" when "001010011011001", -- t[5337] = 0
      "00000" when "001010011011010", -- t[5338] = 0
      "00000" when "001010011011011", -- t[5339] = 0
      "00000" when "001010011011100", -- t[5340] = 0
      "00000" when "001010011011101", -- t[5341] = 0
      "00000" when "001010011011110", -- t[5342] = 0
      "00000" when "001010011011111", -- t[5343] = 0
      "00000" when "001010011100000", -- t[5344] = 0
      "00000" when "001010011100001", -- t[5345] = 0
      "00000" when "001010011100010", -- t[5346] = 0
      "00000" when "001010011100011", -- t[5347] = 0
      "00000" when "001010011100100", -- t[5348] = 0
      "00000" when "001010011100101", -- t[5349] = 0
      "00000" when "001010011100110", -- t[5350] = 0
      "00000" when "001010011100111", -- t[5351] = 0
      "00000" when "001010011101000", -- t[5352] = 0
      "00000" when "001010011101001", -- t[5353] = 0
      "00000" when "001010011101010", -- t[5354] = 0
      "00000" when "001010011101011", -- t[5355] = 0
      "00000" when "001010011101100", -- t[5356] = 0
      "00000" when "001010011101101", -- t[5357] = 0
      "00000" when "001010011101110", -- t[5358] = 0
      "00000" when "001010011101111", -- t[5359] = 0
      "00000" when "001010011110000", -- t[5360] = 0
      "00000" when "001010011110001", -- t[5361] = 0
      "00000" when "001010011110010", -- t[5362] = 0
      "00000" when "001010011110011", -- t[5363] = 0
      "00000" when "001010011110100", -- t[5364] = 0
      "00000" when "001010011110101", -- t[5365] = 0
      "00000" when "001010011110110", -- t[5366] = 0
      "00000" when "001010011110111", -- t[5367] = 0
      "00000" when "001010011111000", -- t[5368] = 0
      "00000" when "001010011111001", -- t[5369] = 0
      "00000" when "001010011111010", -- t[5370] = 0
      "00000" when "001010011111011", -- t[5371] = 0
      "00000" when "001010011111100", -- t[5372] = 0
      "00000" when "001010011111101", -- t[5373] = 0
      "00000" when "001010011111110", -- t[5374] = 0
      "00000" when "001010011111111", -- t[5375] = 0
      "00000" when "001010100000000", -- t[5376] = 0
      "00000" when "001010100000001", -- t[5377] = 0
      "00000" when "001010100000010", -- t[5378] = 0
      "00000" when "001010100000011", -- t[5379] = 0
      "00000" when "001010100000100", -- t[5380] = 0
      "00000" when "001010100000101", -- t[5381] = 0
      "00000" when "001010100000110", -- t[5382] = 0
      "00000" when "001010100000111", -- t[5383] = 0
      "00000" when "001010100001000", -- t[5384] = 0
      "00000" when "001010100001001", -- t[5385] = 0
      "00000" when "001010100001010", -- t[5386] = 0
      "00000" when "001010100001011", -- t[5387] = 0
      "00000" when "001010100001100", -- t[5388] = 0
      "00000" when "001010100001101", -- t[5389] = 0
      "00000" when "001010100001110", -- t[5390] = 0
      "00000" when "001010100001111", -- t[5391] = 0
      "00000" when "001010100010000", -- t[5392] = 0
      "00000" when "001010100010001", -- t[5393] = 0
      "00000" when "001010100010010", -- t[5394] = 0
      "00000" when "001010100010011", -- t[5395] = 0
      "00000" when "001010100010100", -- t[5396] = 0
      "00000" when "001010100010101", -- t[5397] = 0
      "00000" when "001010100010110", -- t[5398] = 0
      "00000" when "001010100010111", -- t[5399] = 0
      "00000" when "001010100011000", -- t[5400] = 0
      "00000" when "001010100011001", -- t[5401] = 0
      "00000" when "001010100011010", -- t[5402] = 0
      "00000" when "001010100011011", -- t[5403] = 0
      "00000" when "001010100011100", -- t[5404] = 0
      "00000" when "001010100011101", -- t[5405] = 0
      "00000" when "001010100011110", -- t[5406] = 0
      "00000" when "001010100011111", -- t[5407] = 0
      "00000" when "001010100100000", -- t[5408] = 0
      "00000" when "001010100100001", -- t[5409] = 0
      "00000" when "001010100100010", -- t[5410] = 0
      "00000" when "001010100100011", -- t[5411] = 0
      "00000" when "001010100100100", -- t[5412] = 0
      "00000" when "001010100100101", -- t[5413] = 0
      "00000" when "001010100100110", -- t[5414] = 0
      "00000" when "001010100100111", -- t[5415] = 0
      "00000" when "001010100101000", -- t[5416] = 0
      "00000" when "001010100101001", -- t[5417] = 0
      "00000" when "001010100101010", -- t[5418] = 0
      "00000" when "001010100101011", -- t[5419] = 0
      "00000" when "001010100101100", -- t[5420] = 0
      "00000" when "001010100101101", -- t[5421] = 0
      "00000" when "001010100101110", -- t[5422] = 0
      "00000" when "001010100101111", -- t[5423] = 0
      "00000" when "001010100110000", -- t[5424] = 0
      "00000" when "001010100110001", -- t[5425] = 0
      "00000" when "001010100110010", -- t[5426] = 0
      "00000" when "001010100110011", -- t[5427] = 0
      "00000" when "001010100110100", -- t[5428] = 0
      "00000" when "001010100110101", -- t[5429] = 0
      "00000" when "001010100110110", -- t[5430] = 0
      "00000" when "001010100110111", -- t[5431] = 0
      "00000" when "001010100111000", -- t[5432] = 0
      "00000" when "001010100111001", -- t[5433] = 0
      "00000" when "001010100111010", -- t[5434] = 0
      "00000" when "001010100111011", -- t[5435] = 0
      "00000" when "001010100111100", -- t[5436] = 0
      "00000" when "001010100111101", -- t[5437] = 0
      "00000" when "001010100111110", -- t[5438] = 0
      "00000" when "001010100111111", -- t[5439] = 0
      "00000" when "001010101000000", -- t[5440] = 0
      "00000" when "001010101000001", -- t[5441] = 0
      "00000" when "001010101000010", -- t[5442] = 0
      "00000" when "001010101000011", -- t[5443] = 0
      "00000" when "001010101000100", -- t[5444] = 0
      "00000" when "001010101000101", -- t[5445] = 0
      "00000" when "001010101000110", -- t[5446] = 0
      "00000" when "001010101000111", -- t[5447] = 0
      "00000" when "001010101001000", -- t[5448] = 0
      "00000" when "001010101001001", -- t[5449] = 0
      "00000" when "001010101001010", -- t[5450] = 0
      "00000" when "001010101001011", -- t[5451] = 0
      "00000" when "001010101001100", -- t[5452] = 0
      "00000" when "001010101001101", -- t[5453] = 0
      "00000" when "001010101001110", -- t[5454] = 0
      "00000" when "001010101001111", -- t[5455] = 0
      "00000" when "001010101010000", -- t[5456] = 0
      "00000" when "001010101010001", -- t[5457] = 0
      "00000" when "001010101010010", -- t[5458] = 0
      "00000" when "001010101010011", -- t[5459] = 0
      "00000" when "001010101010100", -- t[5460] = 0
      "00000" when "001010101010101", -- t[5461] = 0
      "00000" when "001010101010110", -- t[5462] = 0
      "00000" when "001010101010111", -- t[5463] = 0
      "00000" when "001010101011000", -- t[5464] = 0
      "00000" when "001010101011001", -- t[5465] = 0
      "00000" when "001010101011010", -- t[5466] = 0
      "00000" when "001010101011011", -- t[5467] = 0
      "00000" when "001010101011100", -- t[5468] = 0
      "00000" when "001010101011101", -- t[5469] = 0
      "00000" when "001010101011110", -- t[5470] = 0
      "00000" when "001010101011111", -- t[5471] = 0
      "00000" when "001010101100000", -- t[5472] = 0
      "00000" when "001010101100001", -- t[5473] = 0
      "00000" when "001010101100010", -- t[5474] = 0
      "00000" when "001010101100011", -- t[5475] = 0
      "00000" when "001010101100100", -- t[5476] = 0
      "00000" when "001010101100101", -- t[5477] = 0
      "00000" when "001010101100110", -- t[5478] = 0
      "00000" when "001010101100111", -- t[5479] = 0
      "00000" when "001010101101000", -- t[5480] = 0
      "00000" when "001010101101001", -- t[5481] = 0
      "00000" when "001010101101010", -- t[5482] = 0
      "00000" when "001010101101011", -- t[5483] = 0
      "00000" when "001010101101100", -- t[5484] = 0
      "00000" when "001010101101101", -- t[5485] = 0
      "00000" when "001010101101110", -- t[5486] = 0
      "00000" when "001010101101111", -- t[5487] = 0
      "00000" when "001010101110000", -- t[5488] = 0
      "00000" when "001010101110001", -- t[5489] = 0
      "00000" when "001010101110010", -- t[5490] = 0
      "00000" when "001010101110011", -- t[5491] = 0
      "00000" when "001010101110100", -- t[5492] = 0
      "00000" when "001010101110101", -- t[5493] = 0
      "00000" when "001010101110110", -- t[5494] = 0
      "00000" when "001010101110111", -- t[5495] = 0
      "00000" when "001010101111000", -- t[5496] = 0
      "00000" when "001010101111001", -- t[5497] = 0
      "00000" when "001010101111010", -- t[5498] = 0
      "00000" when "001010101111011", -- t[5499] = 0
      "00000" when "001010101111100", -- t[5500] = 0
      "00000" when "001010101111101", -- t[5501] = 0
      "00000" when "001010101111110", -- t[5502] = 0
      "00000" when "001010101111111", -- t[5503] = 0
      "00000" when "001010110000000", -- t[5504] = 0
      "00000" when "001010110000001", -- t[5505] = 0
      "00000" when "001010110000010", -- t[5506] = 0
      "00000" when "001010110000011", -- t[5507] = 0
      "00000" when "001010110000100", -- t[5508] = 0
      "00000" when "001010110000101", -- t[5509] = 0
      "00000" when "001010110000110", -- t[5510] = 0
      "00000" when "001010110000111", -- t[5511] = 0
      "00000" when "001010110001000", -- t[5512] = 0
      "00000" when "001010110001001", -- t[5513] = 0
      "00000" when "001010110001010", -- t[5514] = 0
      "00000" when "001010110001011", -- t[5515] = 0
      "00000" when "001010110001100", -- t[5516] = 0
      "00000" when "001010110001101", -- t[5517] = 0
      "00000" when "001010110001110", -- t[5518] = 0
      "00000" when "001010110001111", -- t[5519] = 0
      "00000" when "001010110010000", -- t[5520] = 0
      "00000" when "001010110010001", -- t[5521] = 0
      "00000" when "001010110010010", -- t[5522] = 0
      "00000" when "001010110010011", -- t[5523] = 0
      "00000" when "001010110010100", -- t[5524] = 0
      "00000" when "001010110010101", -- t[5525] = 0
      "00000" when "001010110010110", -- t[5526] = 0
      "00000" when "001010110010111", -- t[5527] = 0
      "00000" when "001010110011000", -- t[5528] = 0
      "00000" when "001010110011001", -- t[5529] = 0
      "00000" when "001010110011010", -- t[5530] = 0
      "00000" when "001010110011011", -- t[5531] = 0
      "00000" when "001010110011100", -- t[5532] = 0
      "00000" when "001010110011101", -- t[5533] = 0
      "00000" when "001010110011110", -- t[5534] = 0
      "00000" when "001010110011111", -- t[5535] = 0
      "00000" when "001010110100000", -- t[5536] = 0
      "00000" when "001010110100001", -- t[5537] = 0
      "00000" when "001010110100010", -- t[5538] = 0
      "00000" when "001010110100011", -- t[5539] = 0
      "00000" when "001010110100100", -- t[5540] = 0
      "00000" when "001010110100101", -- t[5541] = 0
      "00000" when "001010110100110", -- t[5542] = 0
      "00000" when "001010110100111", -- t[5543] = 0
      "00000" when "001010110101000", -- t[5544] = 0
      "00000" when "001010110101001", -- t[5545] = 0
      "00000" when "001010110101010", -- t[5546] = 0
      "00000" when "001010110101011", -- t[5547] = 0
      "00000" when "001010110101100", -- t[5548] = 0
      "00000" when "001010110101101", -- t[5549] = 0
      "00000" when "001010110101110", -- t[5550] = 0
      "00000" when "001010110101111", -- t[5551] = 0
      "00000" when "001010110110000", -- t[5552] = 0
      "00000" when "001010110110001", -- t[5553] = 0
      "00000" when "001010110110010", -- t[5554] = 0
      "00000" when "001010110110011", -- t[5555] = 0
      "00000" when "001010110110100", -- t[5556] = 0
      "00000" when "001010110110101", -- t[5557] = 0
      "00000" when "001010110110110", -- t[5558] = 0
      "00000" when "001010110110111", -- t[5559] = 0
      "00000" when "001010110111000", -- t[5560] = 0
      "00000" when "001010110111001", -- t[5561] = 0
      "00000" when "001010110111010", -- t[5562] = 0
      "00000" when "001010110111011", -- t[5563] = 0
      "00000" when "001010110111100", -- t[5564] = 0
      "00000" when "001010110111101", -- t[5565] = 0
      "00000" when "001010110111110", -- t[5566] = 0
      "00000" when "001010110111111", -- t[5567] = 0
      "00000" when "001010111000000", -- t[5568] = 0
      "00000" when "001010111000001", -- t[5569] = 0
      "00000" when "001010111000010", -- t[5570] = 0
      "00000" when "001010111000011", -- t[5571] = 0
      "00000" when "001010111000100", -- t[5572] = 0
      "00000" when "001010111000101", -- t[5573] = 0
      "00000" when "001010111000110", -- t[5574] = 0
      "00000" when "001010111000111", -- t[5575] = 0
      "00000" when "001010111001000", -- t[5576] = 0
      "00000" when "001010111001001", -- t[5577] = 0
      "00000" when "001010111001010", -- t[5578] = 0
      "00000" when "001010111001011", -- t[5579] = 0
      "00000" when "001010111001100", -- t[5580] = 0
      "00000" when "001010111001101", -- t[5581] = 0
      "00000" when "001010111001110", -- t[5582] = 0
      "00000" when "001010111001111", -- t[5583] = 0
      "00000" when "001010111010000", -- t[5584] = 0
      "00000" when "001010111010001", -- t[5585] = 0
      "00000" when "001010111010010", -- t[5586] = 0
      "00000" when "001010111010011", -- t[5587] = 0
      "00000" when "001010111010100", -- t[5588] = 0
      "00000" when "001010111010101", -- t[5589] = 0
      "00000" when "001010111010110", -- t[5590] = 0
      "00000" when "001010111010111", -- t[5591] = 0
      "00000" when "001010111011000", -- t[5592] = 0
      "00000" when "001010111011001", -- t[5593] = 0
      "00000" when "001010111011010", -- t[5594] = 0
      "00000" when "001010111011011", -- t[5595] = 0
      "00000" when "001010111011100", -- t[5596] = 0
      "00000" when "001010111011101", -- t[5597] = 0
      "00000" when "001010111011110", -- t[5598] = 0
      "00000" when "001010111011111", -- t[5599] = 0
      "00000" when "001010111100000", -- t[5600] = 0
      "00000" when "001010111100001", -- t[5601] = 0
      "00000" when "001010111100010", -- t[5602] = 0
      "00000" when "001010111100011", -- t[5603] = 0
      "00000" when "001010111100100", -- t[5604] = 0
      "00000" when "001010111100101", -- t[5605] = 0
      "00000" when "001010111100110", -- t[5606] = 0
      "00000" when "001010111100111", -- t[5607] = 0
      "00000" when "001010111101000", -- t[5608] = 0
      "00000" when "001010111101001", -- t[5609] = 0
      "00000" when "001010111101010", -- t[5610] = 0
      "00000" when "001010111101011", -- t[5611] = 0
      "00000" when "001010111101100", -- t[5612] = 0
      "00000" when "001010111101101", -- t[5613] = 0
      "00000" when "001010111101110", -- t[5614] = 0
      "00000" when "001010111101111", -- t[5615] = 0
      "00000" when "001010111110000", -- t[5616] = 0
      "00000" when "001010111110001", -- t[5617] = 0
      "00000" when "001010111110010", -- t[5618] = 0
      "00000" when "001010111110011", -- t[5619] = 0
      "00000" when "001010111110100", -- t[5620] = 0
      "00000" when "001010111110101", -- t[5621] = 0
      "00000" when "001010111110110", -- t[5622] = 0
      "00000" when "001010111110111", -- t[5623] = 0
      "00000" when "001010111111000", -- t[5624] = 0
      "00000" when "001010111111001", -- t[5625] = 0
      "00000" when "001010111111010", -- t[5626] = 0
      "00000" when "001010111111011", -- t[5627] = 0
      "00000" when "001010111111100", -- t[5628] = 0
      "00000" when "001010111111101", -- t[5629] = 0
      "00000" when "001010111111110", -- t[5630] = 0
      "00000" when "001010111111111", -- t[5631] = 0
      "00000" when "001011000000000", -- t[5632] = 0
      "00000" when "001011000000001", -- t[5633] = 0
      "00000" when "001011000000010", -- t[5634] = 0
      "00000" when "001011000000011", -- t[5635] = 0
      "00000" when "001011000000100", -- t[5636] = 0
      "00000" when "001011000000101", -- t[5637] = 0
      "00000" when "001011000000110", -- t[5638] = 0
      "00000" when "001011000000111", -- t[5639] = 0
      "00000" when "001011000001000", -- t[5640] = 0
      "00000" when "001011000001001", -- t[5641] = 0
      "00000" when "001011000001010", -- t[5642] = 0
      "00000" when "001011000001011", -- t[5643] = 0
      "00000" when "001011000001100", -- t[5644] = 0
      "00000" when "001011000001101", -- t[5645] = 0
      "00000" when "001011000001110", -- t[5646] = 0
      "00000" when "001011000001111", -- t[5647] = 0
      "00000" when "001011000010000", -- t[5648] = 0
      "00000" when "001011000010001", -- t[5649] = 0
      "00000" when "001011000010010", -- t[5650] = 0
      "00000" when "001011000010011", -- t[5651] = 0
      "00000" when "001011000010100", -- t[5652] = 0
      "00000" when "001011000010101", -- t[5653] = 0
      "00000" when "001011000010110", -- t[5654] = 0
      "00000" when "001011000010111", -- t[5655] = 0
      "00000" when "001011000011000", -- t[5656] = 0
      "00000" when "001011000011001", -- t[5657] = 0
      "00000" when "001011000011010", -- t[5658] = 0
      "00000" when "001011000011011", -- t[5659] = 0
      "00000" when "001011000011100", -- t[5660] = 0
      "00000" when "001011000011101", -- t[5661] = 0
      "00000" when "001011000011110", -- t[5662] = 0
      "00000" when "001011000011111", -- t[5663] = 0
      "00000" when "001011000100000", -- t[5664] = 0
      "00000" when "001011000100001", -- t[5665] = 0
      "00000" when "001011000100010", -- t[5666] = 0
      "00000" when "001011000100011", -- t[5667] = 0
      "00000" when "001011000100100", -- t[5668] = 0
      "00000" when "001011000100101", -- t[5669] = 0
      "00000" when "001011000100110", -- t[5670] = 0
      "00000" when "001011000100111", -- t[5671] = 0
      "00000" when "001011000101000", -- t[5672] = 0
      "00000" when "001011000101001", -- t[5673] = 0
      "00000" when "001011000101010", -- t[5674] = 0
      "00000" when "001011000101011", -- t[5675] = 0
      "00000" when "001011000101100", -- t[5676] = 0
      "00000" when "001011000101101", -- t[5677] = 0
      "00000" when "001011000101110", -- t[5678] = 0
      "00000" when "001011000101111", -- t[5679] = 0
      "00000" when "001011000110000", -- t[5680] = 0
      "00000" when "001011000110001", -- t[5681] = 0
      "00000" when "001011000110010", -- t[5682] = 0
      "00000" when "001011000110011", -- t[5683] = 0
      "00000" when "001011000110100", -- t[5684] = 0
      "00000" when "001011000110101", -- t[5685] = 0
      "00000" when "001011000110110", -- t[5686] = 0
      "00000" when "001011000110111", -- t[5687] = 0
      "00000" when "001011000111000", -- t[5688] = 0
      "00000" when "001011000111001", -- t[5689] = 0
      "00000" when "001011000111010", -- t[5690] = 0
      "00000" when "001011000111011", -- t[5691] = 0
      "00000" when "001011000111100", -- t[5692] = 0
      "00000" when "001011000111101", -- t[5693] = 0
      "00000" when "001011000111110", -- t[5694] = 0
      "00000" when "001011000111111", -- t[5695] = 0
      "00000" when "001011001000000", -- t[5696] = 0
      "00000" when "001011001000001", -- t[5697] = 0
      "00000" when "001011001000010", -- t[5698] = 0
      "00000" when "001011001000011", -- t[5699] = 0
      "00000" when "001011001000100", -- t[5700] = 0
      "00000" when "001011001000101", -- t[5701] = 0
      "00000" when "001011001000110", -- t[5702] = 0
      "00000" when "001011001000111", -- t[5703] = 0
      "00000" when "001011001001000", -- t[5704] = 0
      "00000" when "001011001001001", -- t[5705] = 0
      "00000" when "001011001001010", -- t[5706] = 0
      "00000" when "001011001001011", -- t[5707] = 0
      "00000" when "001011001001100", -- t[5708] = 0
      "00000" when "001011001001101", -- t[5709] = 0
      "00000" when "001011001001110", -- t[5710] = 0
      "00000" when "001011001001111", -- t[5711] = 0
      "00000" when "001011001010000", -- t[5712] = 0
      "00000" when "001011001010001", -- t[5713] = 0
      "00000" when "001011001010010", -- t[5714] = 0
      "00000" when "001011001010011", -- t[5715] = 0
      "00000" when "001011001010100", -- t[5716] = 0
      "00000" when "001011001010101", -- t[5717] = 0
      "00000" when "001011001010110", -- t[5718] = 0
      "00000" when "001011001010111", -- t[5719] = 0
      "00000" when "001011001011000", -- t[5720] = 0
      "00000" when "001011001011001", -- t[5721] = 0
      "00000" when "001011001011010", -- t[5722] = 0
      "00000" when "001011001011011", -- t[5723] = 0
      "00000" when "001011001011100", -- t[5724] = 0
      "00000" when "001011001011101", -- t[5725] = 0
      "00000" when "001011001011110", -- t[5726] = 0
      "00000" when "001011001011111", -- t[5727] = 0
      "00000" when "001011001100000", -- t[5728] = 0
      "00000" when "001011001100001", -- t[5729] = 0
      "00000" when "001011001100010", -- t[5730] = 0
      "00000" when "001011001100011", -- t[5731] = 0
      "00000" when "001011001100100", -- t[5732] = 0
      "00000" when "001011001100101", -- t[5733] = 0
      "00000" when "001011001100110", -- t[5734] = 0
      "00000" when "001011001100111", -- t[5735] = 0
      "00000" when "001011001101000", -- t[5736] = 0
      "00000" when "001011001101001", -- t[5737] = 0
      "00000" when "001011001101010", -- t[5738] = 0
      "00000" when "001011001101011", -- t[5739] = 0
      "00000" when "001011001101100", -- t[5740] = 0
      "00000" when "001011001101101", -- t[5741] = 0
      "00000" when "001011001101110", -- t[5742] = 0
      "00000" when "001011001101111", -- t[5743] = 0
      "00000" when "001011001110000", -- t[5744] = 0
      "00000" when "001011001110001", -- t[5745] = 0
      "00000" when "001011001110010", -- t[5746] = 0
      "00000" when "001011001110011", -- t[5747] = 0
      "00000" when "001011001110100", -- t[5748] = 0
      "00000" when "001011001110101", -- t[5749] = 0
      "00000" when "001011001110110", -- t[5750] = 0
      "00000" when "001011001110111", -- t[5751] = 0
      "00000" when "001011001111000", -- t[5752] = 0
      "00000" when "001011001111001", -- t[5753] = 0
      "00000" when "001011001111010", -- t[5754] = 0
      "00000" when "001011001111011", -- t[5755] = 0
      "00000" when "001011001111100", -- t[5756] = 0
      "00000" when "001011001111101", -- t[5757] = 0
      "00000" when "001011001111110", -- t[5758] = 0
      "00000" when "001011001111111", -- t[5759] = 0
      "00000" when "001011010000000", -- t[5760] = 0
      "00000" when "001011010000001", -- t[5761] = 0
      "00000" when "001011010000010", -- t[5762] = 0
      "00000" when "001011010000011", -- t[5763] = 0
      "00000" when "001011010000100", -- t[5764] = 0
      "00000" when "001011010000101", -- t[5765] = 0
      "00000" when "001011010000110", -- t[5766] = 0
      "00000" when "001011010000111", -- t[5767] = 0
      "00000" when "001011010001000", -- t[5768] = 0
      "00000" when "001011010001001", -- t[5769] = 0
      "00000" when "001011010001010", -- t[5770] = 0
      "00000" when "001011010001011", -- t[5771] = 0
      "00000" when "001011010001100", -- t[5772] = 0
      "00000" when "001011010001101", -- t[5773] = 0
      "00000" when "001011010001110", -- t[5774] = 0
      "00000" when "001011010001111", -- t[5775] = 0
      "00000" when "001011010010000", -- t[5776] = 0
      "00000" when "001011010010001", -- t[5777] = 0
      "00000" when "001011010010010", -- t[5778] = 0
      "00000" when "001011010010011", -- t[5779] = 0
      "00000" when "001011010010100", -- t[5780] = 0
      "00000" when "001011010010101", -- t[5781] = 0
      "00000" when "001011010010110", -- t[5782] = 0
      "00000" when "001011010010111", -- t[5783] = 0
      "00000" when "001011010011000", -- t[5784] = 0
      "00000" when "001011010011001", -- t[5785] = 0
      "00000" when "001011010011010", -- t[5786] = 0
      "00000" when "001011010011011", -- t[5787] = 0
      "00000" when "001011010011100", -- t[5788] = 0
      "00000" when "001011010011101", -- t[5789] = 0
      "00000" when "001011010011110", -- t[5790] = 0
      "00000" when "001011010011111", -- t[5791] = 0
      "00000" when "001011010100000", -- t[5792] = 0
      "00000" when "001011010100001", -- t[5793] = 0
      "00000" when "001011010100010", -- t[5794] = 0
      "00000" when "001011010100011", -- t[5795] = 0
      "00000" when "001011010100100", -- t[5796] = 0
      "00000" when "001011010100101", -- t[5797] = 0
      "00000" when "001011010100110", -- t[5798] = 0
      "00000" when "001011010100111", -- t[5799] = 0
      "00000" when "001011010101000", -- t[5800] = 0
      "00000" when "001011010101001", -- t[5801] = 0
      "00000" when "001011010101010", -- t[5802] = 0
      "00000" when "001011010101011", -- t[5803] = 0
      "00000" when "001011010101100", -- t[5804] = 0
      "00000" when "001011010101101", -- t[5805] = 0
      "00000" when "001011010101110", -- t[5806] = 0
      "00000" when "001011010101111", -- t[5807] = 0
      "00000" when "001011010110000", -- t[5808] = 0
      "00000" when "001011010110001", -- t[5809] = 0
      "00000" when "001011010110010", -- t[5810] = 0
      "00000" when "001011010110011", -- t[5811] = 0
      "00000" when "001011010110100", -- t[5812] = 0
      "00000" when "001011010110101", -- t[5813] = 0
      "00000" when "001011010110110", -- t[5814] = 0
      "00000" when "001011010110111", -- t[5815] = 0
      "00000" when "001011010111000", -- t[5816] = 0
      "00000" when "001011010111001", -- t[5817] = 0
      "00000" when "001011010111010", -- t[5818] = 0
      "00000" when "001011010111011", -- t[5819] = 0
      "00000" when "001011010111100", -- t[5820] = 0
      "00000" when "001011010111101", -- t[5821] = 0
      "00000" when "001011010111110", -- t[5822] = 0
      "00000" when "001011010111111", -- t[5823] = 0
      "00000" when "001011011000000", -- t[5824] = 0
      "00000" when "001011011000001", -- t[5825] = 0
      "00000" when "001011011000010", -- t[5826] = 0
      "00000" when "001011011000011", -- t[5827] = 0
      "00000" when "001011011000100", -- t[5828] = 0
      "00000" when "001011011000101", -- t[5829] = 0
      "00000" when "001011011000110", -- t[5830] = 0
      "00000" when "001011011000111", -- t[5831] = 0
      "00000" when "001011011001000", -- t[5832] = 0
      "00000" when "001011011001001", -- t[5833] = 0
      "00000" when "001011011001010", -- t[5834] = 0
      "00000" when "001011011001011", -- t[5835] = 0
      "00000" when "001011011001100", -- t[5836] = 0
      "00000" when "001011011001101", -- t[5837] = 0
      "00000" when "001011011001110", -- t[5838] = 0
      "00000" when "001011011001111", -- t[5839] = 0
      "00000" when "001011011010000", -- t[5840] = 0
      "00000" when "001011011010001", -- t[5841] = 0
      "00000" when "001011011010010", -- t[5842] = 0
      "00000" when "001011011010011", -- t[5843] = 0
      "00000" when "001011011010100", -- t[5844] = 0
      "00000" when "001011011010101", -- t[5845] = 0
      "00000" when "001011011010110", -- t[5846] = 0
      "00000" when "001011011010111", -- t[5847] = 0
      "00000" when "001011011011000", -- t[5848] = 0
      "00000" when "001011011011001", -- t[5849] = 0
      "00000" when "001011011011010", -- t[5850] = 0
      "00000" when "001011011011011", -- t[5851] = 0
      "00000" when "001011011011100", -- t[5852] = 0
      "00000" when "001011011011101", -- t[5853] = 0
      "00000" when "001011011011110", -- t[5854] = 0
      "00000" when "001011011011111", -- t[5855] = 0
      "00000" when "001011011100000", -- t[5856] = 0
      "00000" when "001011011100001", -- t[5857] = 0
      "00000" when "001011011100010", -- t[5858] = 0
      "00000" when "001011011100011", -- t[5859] = 0
      "00000" when "001011011100100", -- t[5860] = 0
      "00000" when "001011011100101", -- t[5861] = 0
      "00000" when "001011011100110", -- t[5862] = 0
      "00000" when "001011011100111", -- t[5863] = 0
      "00000" when "001011011101000", -- t[5864] = 0
      "00000" when "001011011101001", -- t[5865] = 0
      "00000" when "001011011101010", -- t[5866] = 0
      "00000" when "001011011101011", -- t[5867] = 0
      "00000" when "001011011101100", -- t[5868] = 0
      "00000" when "001011011101101", -- t[5869] = 0
      "00000" when "001011011101110", -- t[5870] = 0
      "00000" when "001011011101111", -- t[5871] = 0
      "00000" when "001011011110000", -- t[5872] = 0
      "00000" when "001011011110001", -- t[5873] = 0
      "00000" when "001011011110010", -- t[5874] = 0
      "00000" when "001011011110011", -- t[5875] = 0
      "00000" when "001011011110100", -- t[5876] = 0
      "00000" when "001011011110101", -- t[5877] = 0
      "00000" when "001011011110110", -- t[5878] = 0
      "00000" when "001011011110111", -- t[5879] = 0
      "00000" when "001011011111000", -- t[5880] = 0
      "00000" when "001011011111001", -- t[5881] = 0
      "00000" when "001011011111010", -- t[5882] = 0
      "00000" when "001011011111011", -- t[5883] = 0
      "00000" when "001011011111100", -- t[5884] = 0
      "00000" when "001011011111101", -- t[5885] = 0
      "00000" when "001011011111110", -- t[5886] = 0
      "00000" when "001011011111111", -- t[5887] = 0
      "00000" when "001011100000000", -- t[5888] = 0
      "00000" when "001011100000001", -- t[5889] = 0
      "00000" when "001011100000010", -- t[5890] = 0
      "00000" when "001011100000011", -- t[5891] = 0
      "00000" when "001011100000100", -- t[5892] = 0
      "00000" when "001011100000101", -- t[5893] = 0
      "00000" when "001011100000110", -- t[5894] = 0
      "00000" when "001011100000111", -- t[5895] = 0
      "00000" when "001011100001000", -- t[5896] = 0
      "00000" when "001011100001001", -- t[5897] = 0
      "00000" when "001011100001010", -- t[5898] = 0
      "00000" when "001011100001011", -- t[5899] = 0
      "00000" when "001011100001100", -- t[5900] = 0
      "00000" when "001011100001101", -- t[5901] = 0
      "00000" when "001011100001110", -- t[5902] = 0
      "00000" when "001011100001111", -- t[5903] = 0
      "00000" when "001011100010000", -- t[5904] = 0
      "00000" when "001011100010001", -- t[5905] = 0
      "00000" when "001011100010010", -- t[5906] = 0
      "00000" when "001011100010011", -- t[5907] = 0
      "00000" when "001011100010100", -- t[5908] = 0
      "00000" when "001011100010101", -- t[5909] = 0
      "00000" when "001011100010110", -- t[5910] = 0
      "00000" when "001011100010111", -- t[5911] = 0
      "00000" when "001011100011000", -- t[5912] = 0
      "00000" when "001011100011001", -- t[5913] = 0
      "00000" when "001011100011010", -- t[5914] = 0
      "00000" when "001011100011011", -- t[5915] = 0
      "00000" when "001011100011100", -- t[5916] = 0
      "00000" when "001011100011101", -- t[5917] = 0
      "00000" when "001011100011110", -- t[5918] = 0
      "00000" when "001011100011111", -- t[5919] = 0
      "00000" when "001011100100000", -- t[5920] = 0
      "00000" when "001011100100001", -- t[5921] = 0
      "00000" when "001011100100010", -- t[5922] = 0
      "00000" when "001011100100011", -- t[5923] = 0
      "00000" when "001011100100100", -- t[5924] = 0
      "00000" when "001011100100101", -- t[5925] = 0
      "00000" when "001011100100110", -- t[5926] = 0
      "00000" when "001011100100111", -- t[5927] = 0
      "00000" when "001011100101000", -- t[5928] = 0
      "00000" when "001011100101001", -- t[5929] = 0
      "00000" when "001011100101010", -- t[5930] = 0
      "00000" when "001011100101011", -- t[5931] = 0
      "00000" when "001011100101100", -- t[5932] = 0
      "00000" when "001011100101101", -- t[5933] = 0
      "00000" when "001011100101110", -- t[5934] = 0
      "00000" when "001011100101111", -- t[5935] = 0
      "00000" when "001011100110000", -- t[5936] = 0
      "00000" when "001011100110001", -- t[5937] = 0
      "00000" when "001011100110010", -- t[5938] = 0
      "00000" when "001011100110011", -- t[5939] = 0
      "00000" when "001011100110100", -- t[5940] = 0
      "00000" when "001011100110101", -- t[5941] = 0
      "00000" when "001011100110110", -- t[5942] = 0
      "00000" when "001011100110111", -- t[5943] = 0
      "00000" when "001011100111000", -- t[5944] = 0
      "00000" when "001011100111001", -- t[5945] = 0
      "00000" when "001011100111010", -- t[5946] = 0
      "00000" when "001011100111011", -- t[5947] = 0
      "00000" when "001011100111100", -- t[5948] = 0
      "00000" when "001011100111101", -- t[5949] = 0
      "00000" when "001011100111110", -- t[5950] = 0
      "00000" when "001011100111111", -- t[5951] = 0
      "00000" when "001011101000000", -- t[5952] = 0
      "00000" when "001011101000001", -- t[5953] = 0
      "00000" when "001011101000010", -- t[5954] = 0
      "00000" when "001011101000011", -- t[5955] = 0
      "00000" when "001011101000100", -- t[5956] = 0
      "00000" when "001011101000101", -- t[5957] = 0
      "00000" when "001011101000110", -- t[5958] = 0
      "00000" when "001011101000111", -- t[5959] = 0
      "00000" when "001011101001000", -- t[5960] = 0
      "00000" when "001011101001001", -- t[5961] = 0
      "00000" when "001011101001010", -- t[5962] = 0
      "00000" when "001011101001011", -- t[5963] = 0
      "00000" when "001011101001100", -- t[5964] = 0
      "00000" when "001011101001101", -- t[5965] = 0
      "00000" when "001011101001110", -- t[5966] = 0
      "00000" when "001011101001111", -- t[5967] = 0
      "00000" when "001011101010000", -- t[5968] = 0
      "00000" when "001011101010001", -- t[5969] = 0
      "00000" when "001011101010010", -- t[5970] = 0
      "00000" when "001011101010011", -- t[5971] = 0
      "00000" when "001011101010100", -- t[5972] = 0
      "00000" when "001011101010101", -- t[5973] = 0
      "00000" when "001011101010110", -- t[5974] = 0
      "00000" when "001011101010111", -- t[5975] = 0
      "00000" when "001011101011000", -- t[5976] = 0
      "00000" when "001011101011001", -- t[5977] = 0
      "00000" when "001011101011010", -- t[5978] = 0
      "00000" when "001011101011011", -- t[5979] = 0
      "00000" when "001011101011100", -- t[5980] = 0
      "00000" when "001011101011101", -- t[5981] = 0
      "00000" when "001011101011110", -- t[5982] = 0
      "00000" when "001011101011111", -- t[5983] = 0
      "00000" when "001011101100000", -- t[5984] = 0
      "00000" when "001011101100001", -- t[5985] = 0
      "00000" when "001011101100010", -- t[5986] = 0
      "00000" when "001011101100011", -- t[5987] = 0
      "00000" when "001011101100100", -- t[5988] = 0
      "00000" when "001011101100101", -- t[5989] = 0
      "00000" when "001011101100110", -- t[5990] = 0
      "00000" when "001011101100111", -- t[5991] = 0
      "00000" when "001011101101000", -- t[5992] = 0
      "00000" when "001011101101001", -- t[5993] = 0
      "00000" when "001011101101010", -- t[5994] = 0
      "00000" when "001011101101011", -- t[5995] = 0
      "00000" when "001011101101100", -- t[5996] = 0
      "00000" when "001011101101101", -- t[5997] = 0
      "00000" when "001011101101110", -- t[5998] = 0
      "00000" when "001011101101111", -- t[5999] = 0
      "00000" when "001011101110000", -- t[6000] = 0
      "00000" when "001011101110001", -- t[6001] = 0
      "00000" when "001011101110010", -- t[6002] = 0
      "00000" when "001011101110011", -- t[6003] = 0
      "00000" when "001011101110100", -- t[6004] = 0
      "00000" when "001011101110101", -- t[6005] = 0
      "00000" when "001011101110110", -- t[6006] = 0
      "00000" when "001011101110111", -- t[6007] = 0
      "00000" when "001011101111000", -- t[6008] = 0
      "00000" when "001011101111001", -- t[6009] = 0
      "00000" when "001011101111010", -- t[6010] = 0
      "00000" when "001011101111011", -- t[6011] = 0
      "00000" when "001011101111100", -- t[6012] = 0
      "00000" when "001011101111101", -- t[6013] = 0
      "00000" when "001011101111110", -- t[6014] = 0
      "00000" when "001011101111111", -- t[6015] = 0
      "00000" when "001011110000000", -- t[6016] = 0
      "00000" when "001011110000001", -- t[6017] = 0
      "00000" when "001011110000010", -- t[6018] = 0
      "00000" when "001011110000011", -- t[6019] = 0
      "00000" when "001011110000100", -- t[6020] = 0
      "00000" when "001011110000101", -- t[6021] = 0
      "00000" when "001011110000110", -- t[6022] = 0
      "00000" when "001011110000111", -- t[6023] = 0
      "00000" when "001011110001000", -- t[6024] = 0
      "00000" when "001011110001001", -- t[6025] = 0
      "00000" when "001011110001010", -- t[6026] = 0
      "00000" when "001011110001011", -- t[6027] = 0
      "00000" when "001011110001100", -- t[6028] = 0
      "00000" when "001011110001101", -- t[6029] = 0
      "00000" when "001011110001110", -- t[6030] = 0
      "00000" when "001011110001111", -- t[6031] = 0
      "00000" when "001011110010000", -- t[6032] = 0
      "00000" when "001011110010001", -- t[6033] = 0
      "00000" when "001011110010010", -- t[6034] = 0
      "00000" when "001011110010011", -- t[6035] = 0
      "00000" when "001011110010100", -- t[6036] = 0
      "00000" when "001011110010101", -- t[6037] = 0
      "00000" when "001011110010110", -- t[6038] = 0
      "00000" when "001011110010111", -- t[6039] = 0
      "00000" when "001011110011000", -- t[6040] = 0
      "00000" when "001011110011001", -- t[6041] = 0
      "00000" when "001011110011010", -- t[6042] = 0
      "00000" when "001011110011011", -- t[6043] = 0
      "00000" when "001011110011100", -- t[6044] = 0
      "00000" when "001011110011101", -- t[6045] = 0
      "00000" when "001011110011110", -- t[6046] = 0
      "00000" when "001011110011111", -- t[6047] = 0
      "00000" when "001011110100000", -- t[6048] = 0
      "00000" when "001011110100001", -- t[6049] = 0
      "00000" when "001011110100010", -- t[6050] = 0
      "00000" when "001011110100011", -- t[6051] = 0
      "00000" when "001011110100100", -- t[6052] = 0
      "00000" when "001011110100101", -- t[6053] = 0
      "00000" when "001011110100110", -- t[6054] = 0
      "00000" when "001011110100111", -- t[6055] = 0
      "00000" when "001011110101000", -- t[6056] = 0
      "00000" when "001011110101001", -- t[6057] = 0
      "00000" when "001011110101010", -- t[6058] = 0
      "00000" when "001011110101011", -- t[6059] = 0
      "00000" when "001011110101100", -- t[6060] = 0
      "00000" when "001011110101101", -- t[6061] = 0
      "00000" when "001011110101110", -- t[6062] = 0
      "00000" when "001011110101111", -- t[6063] = 0
      "00000" when "001011110110000", -- t[6064] = 0
      "00000" when "001011110110001", -- t[6065] = 0
      "00000" when "001011110110010", -- t[6066] = 0
      "00000" when "001011110110011", -- t[6067] = 0
      "00000" when "001011110110100", -- t[6068] = 0
      "00000" when "001011110110101", -- t[6069] = 0
      "00000" when "001011110110110", -- t[6070] = 0
      "00000" when "001011110110111", -- t[6071] = 0
      "00000" when "001011110111000", -- t[6072] = 0
      "00000" when "001011110111001", -- t[6073] = 0
      "00000" when "001011110111010", -- t[6074] = 0
      "00000" when "001011110111011", -- t[6075] = 0
      "00000" when "001011110111100", -- t[6076] = 0
      "00000" when "001011110111101", -- t[6077] = 0
      "00000" when "001011110111110", -- t[6078] = 0
      "00000" when "001011110111111", -- t[6079] = 0
      "00000" when "001011111000000", -- t[6080] = 0
      "00000" when "001011111000001", -- t[6081] = 0
      "00000" when "001011111000010", -- t[6082] = 0
      "00000" when "001011111000011", -- t[6083] = 0
      "00000" when "001011111000100", -- t[6084] = 0
      "00000" when "001011111000101", -- t[6085] = 0
      "00000" when "001011111000110", -- t[6086] = 0
      "00000" when "001011111000111", -- t[6087] = 0
      "00000" when "001011111001000", -- t[6088] = 0
      "00000" when "001011111001001", -- t[6089] = 0
      "00000" when "001011111001010", -- t[6090] = 0
      "00000" when "001011111001011", -- t[6091] = 0
      "00000" when "001011111001100", -- t[6092] = 0
      "00000" when "001011111001101", -- t[6093] = 0
      "00000" when "001011111001110", -- t[6094] = 0
      "00000" when "001011111001111", -- t[6095] = 0
      "00000" when "001011111010000", -- t[6096] = 0
      "00000" when "001011111010001", -- t[6097] = 0
      "00000" when "001011111010010", -- t[6098] = 0
      "00000" when "001011111010011", -- t[6099] = 0
      "00000" when "001011111010100", -- t[6100] = 0
      "00000" when "001011111010101", -- t[6101] = 0
      "00000" when "001011111010110", -- t[6102] = 0
      "00000" when "001011111010111", -- t[6103] = 0
      "00000" when "001011111011000", -- t[6104] = 0
      "00000" when "001011111011001", -- t[6105] = 0
      "00000" when "001011111011010", -- t[6106] = 0
      "00000" when "001011111011011", -- t[6107] = 0
      "00000" when "001011111011100", -- t[6108] = 0
      "00000" when "001011111011101", -- t[6109] = 0
      "00000" when "001011111011110", -- t[6110] = 0
      "00000" when "001011111011111", -- t[6111] = 0
      "00000" when "001011111100000", -- t[6112] = 0
      "00000" when "001011111100001", -- t[6113] = 0
      "00000" when "001011111100010", -- t[6114] = 0
      "00000" when "001011111100011", -- t[6115] = 0
      "00000" when "001011111100100", -- t[6116] = 0
      "00000" when "001011111100101", -- t[6117] = 0
      "00000" when "001011111100110", -- t[6118] = 0
      "00000" when "001011111100111", -- t[6119] = 0
      "00000" when "001011111101000", -- t[6120] = 0
      "00000" when "001011111101001", -- t[6121] = 0
      "00000" when "001011111101010", -- t[6122] = 0
      "00000" when "001011111101011", -- t[6123] = 0
      "00000" when "001011111101100", -- t[6124] = 0
      "00000" when "001011111101101", -- t[6125] = 0
      "00000" when "001011111101110", -- t[6126] = 0
      "00000" when "001011111101111", -- t[6127] = 0
      "00000" when "001011111110000", -- t[6128] = 0
      "00000" when "001011111110001", -- t[6129] = 0
      "00000" when "001011111110010", -- t[6130] = 0
      "00000" when "001011111110011", -- t[6131] = 0
      "00000" when "001011111110100", -- t[6132] = 0
      "00000" when "001011111110101", -- t[6133] = 0
      "00000" when "001011111110110", -- t[6134] = 0
      "00000" when "001011111110111", -- t[6135] = 0
      "00000" when "001011111111000", -- t[6136] = 0
      "00000" when "001011111111001", -- t[6137] = 0
      "00000" when "001011111111010", -- t[6138] = 0
      "00000" when "001011111111011", -- t[6139] = 0
      "00000" when "001011111111100", -- t[6140] = 0
      "00000" when "001011111111101", -- t[6141] = 0
      "00000" when "001011111111110", -- t[6142] = 0
      "00000" when "001011111111111", -- t[6143] = 0
      "00000" when "001100000000000", -- t[6144] = 0
      "00000" when "001100000000001", -- t[6145] = 0
      "00000" when "001100000000010", -- t[6146] = 0
      "00000" when "001100000000011", -- t[6147] = 0
      "00000" when "001100000000100", -- t[6148] = 0
      "00000" when "001100000000101", -- t[6149] = 0
      "00000" when "001100000000110", -- t[6150] = 0
      "00000" when "001100000000111", -- t[6151] = 0
      "00000" when "001100000001000", -- t[6152] = 0
      "00000" when "001100000001001", -- t[6153] = 0
      "00000" when "001100000001010", -- t[6154] = 0
      "00000" when "001100000001011", -- t[6155] = 0
      "00000" when "001100000001100", -- t[6156] = 0
      "00000" when "001100000001101", -- t[6157] = 0
      "00000" when "001100000001110", -- t[6158] = 0
      "00000" when "001100000001111", -- t[6159] = 0
      "00000" when "001100000010000", -- t[6160] = 0
      "00000" when "001100000010001", -- t[6161] = 0
      "00000" when "001100000010010", -- t[6162] = 0
      "00000" when "001100000010011", -- t[6163] = 0
      "00000" when "001100000010100", -- t[6164] = 0
      "00000" when "001100000010101", -- t[6165] = 0
      "00000" when "001100000010110", -- t[6166] = 0
      "00000" when "001100000010111", -- t[6167] = 0
      "00000" when "001100000011000", -- t[6168] = 0
      "00000" when "001100000011001", -- t[6169] = 0
      "00000" when "001100000011010", -- t[6170] = 0
      "00000" when "001100000011011", -- t[6171] = 0
      "00000" when "001100000011100", -- t[6172] = 0
      "00000" when "001100000011101", -- t[6173] = 0
      "00000" when "001100000011110", -- t[6174] = 0
      "00000" when "001100000011111", -- t[6175] = 0
      "00000" when "001100000100000", -- t[6176] = 0
      "00000" when "001100000100001", -- t[6177] = 0
      "00000" when "001100000100010", -- t[6178] = 0
      "00000" when "001100000100011", -- t[6179] = 0
      "00000" when "001100000100100", -- t[6180] = 0
      "00000" when "001100000100101", -- t[6181] = 0
      "00000" when "001100000100110", -- t[6182] = 0
      "00000" when "001100000100111", -- t[6183] = 0
      "00000" when "001100000101000", -- t[6184] = 0
      "00000" when "001100000101001", -- t[6185] = 0
      "00000" when "001100000101010", -- t[6186] = 0
      "00000" when "001100000101011", -- t[6187] = 0
      "00000" when "001100000101100", -- t[6188] = 0
      "00000" when "001100000101101", -- t[6189] = 0
      "00000" when "001100000101110", -- t[6190] = 0
      "00000" when "001100000101111", -- t[6191] = 0
      "00000" when "001100000110000", -- t[6192] = 0
      "00000" when "001100000110001", -- t[6193] = 0
      "00000" when "001100000110010", -- t[6194] = 0
      "00000" when "001100000110011", -- t[6195] = 0
      "00000" when "001100000110100", -- t[6196] = 0
      "00000" when "001100000110101", -- t[6197] = 0
      "00000" when "001100000110110", -- t[6198] = 0
      "00000" when "001100000110111", -- t[6199] = 0
      "00000" when "001100000111000", -- t[6200] = 0
      "00000" when "001100000111001", -- t[6201] = 0
      "00000" when "001100000111010", -- t[6202] = 0
      "00000" when "001100000111011", -- t[6203] = 0
      "00000" when "001100000111100", -- t[6204] = 0
      "00000" when "001100000111101", -- t[6205] = 0
      "00000" when "001100000111110", -- t[6206] = 0
      "00000" when "001100000111111", -- t[6207] = 0
      "00000" when "001100001000000", -- t[6208] = 0
      "00000" when "001100001000001", -- t[6209] = 0
      "00000" when "001100001000010", -- t[6210] = 0
      "00000" when "001100001000011", -- t[6211] = 0
      "00000" when "001100001000100", -- t[6212] = 0
      "00000" when "001100001000101", -- t[6213] = 0
      "00000" when "001100001000110", -- t[6214] = 0
      "00000" when "001100001000111", -- t[6215] = 0
      "00000" when "001100001001000", -- t[6216] = 0
      "00000" when "001100001001001", -- t[6217] = 0
      "00000" when "001100001001010", -- t[6218] = 0
      "00000" when "001100001001011", -- t[6219] = 0
      "00000" when "001100001001100", -- t[6220] = 0
      "00000" when "001100001001101", -- t[6221] = 0
      "00000" when "001100001001110", -- t[6222] = 0
      "00000" when "001100001001111", -- t[6223] = 0
      "00000" when "001100001010000", -- t[6224] = 0
      "00000" when "001100001010001", -- t[6225] = 0
      "00000" when "001100001010010", -- t[6226] = 0
      "00000" when "001100001010011", -- t[6227] = 0
      "00000" when "001100001010100", -- t[6228] = 0
      "00000" when "001100001010101", -- t[6229] = 0
      "00000" when "001100001010110", -- t[6230] = 0
      "00000" when "001100001010111", -- t[6231] = 0
      "00000" when "001100001011000", -- t[6232] = 0
      "00000" when "001100001011001", -- t[6233] = 0
      "00000" when "001100001011010", -- t[6234] = 0
      "00000" when "001100001011011", -- t[6235] = 0
      "00000" when "001100001011100", -- t[6236] = 0
      "00000" when "001100001011101", -- t[6237] = 0
      "00000" when "001100001011110", -- t[6238] = 0
      "00000" when "001100001011111", -- t[6239] = 0
      "00000" when "001100001100000", -- t[6240] = 0
      "00000" when "001100001100001", -- t[6241] = 0
      "00000" when "001100001100010", -- t[6242] = 0
      "00000" when "001100001100011", -- t[6243] = 0
      "00000" when "001100001100100", -- t[6244] = 0
      "00000" when "001100001100101", -- t[6245] = 0
      "00000" when "001100001100110", -- t[6246] = 0
      "00000" when "001100001100111", -- t[6247] = 0
      "00000" when "001100001101000", -- t[6248] = 0
      "00000" when "001100001101001", -- t[6249] = 0
      "00000" when "001100001101010", -- t[6250] = 0
      "00000" when "001100001101011", -- t[6251] = 0
      "00000" when "001100001101100", -- t[6252] = 0
      "00000" when "001100001101101", -- t[6253] = 0
      "00000" when "001100001101110", -- t[6254] = 0
      "00000" when "001100001101111", -- t[6255] = 0
      "00000" when "001100001110000", -- t[6256] = 0
      "00000" when "001100001110001", -- t[6257] = 0
      "00000" when "001100001110010", -- t[6258] = 0
      "00000" when "001100001110011", -- t[6259] = 0
      "00000" when "001100001110100", -- t[6260] = 0
      "00000" when "001100001110101", -- t[6261] = 0
      "00000" when "001100001110110", -- t[6262] = 0
      "00000" when "001100001110111", -- t[6263] = 0
      "00000" when "001100001111000", -- t[6264] = 0
      "00000" when "001100001111001", -- t[6265] = 0
      "00000" when "001100001111010", -- t[6266] = 0
      "00000" when "001100001111011", -- t[6267] = 0
      "00000" when "001100001111100", -- t[6268] = 0
      "00000" when "001100001111101", -- t[6269] = 0
      "00000" when "001100001111110", -- t[6270] = 0
      "00000" when "001100001111111", -- t[6271] = 0
      "00000" when "001100010000000", -- t[6272] = 0
      "00000" when "001100010000001", -- t[6273] = 0
      "00000" when "001100010000010", -- t[6274] = 0
      "00000" when "001100010000011", -- t[6275] = 0
      "00000" when "001100010000100", -- t[6276] = 0
      "00000" when "001100010000101", -- t[6277] = 0
      "00000" when "001100010000110", -- t[6278] = 0
      "00000" when "001100010000111", -- t[6279] = 0
      "00000" when "001100010001000", -- t[6280] = 0
      "00000" when "001100010001001", -- t[6281] = 0
      "00000" when "001100010001010", -- t[6282] = 0
      "00000" when "001100010001011", -- t[6283] = 0
      "00000" when "001100010001100", -- t[6284] = 0
      "00000" when "001100010001101", -- t[6285] = 0
      "00000" when "001100010001110", -- t[6286] = 0
      "00000" when "001100010001111", -- t[6287] = 0
      "00000" when "001100010010000", -- t[6288] = 0
      "00000" when "001100010010001", -- t[6289] = 0
      "00000" when "001100010010010", -- t[6290] = 0
      "00000" when "001100010010011", -- t[6291] = 0
      "00000" when "001100010010100", -- t[6292] = 0
      "00000" when "001100010010101", -- t[6293] = 0
      "00000" when "001100010010110", -- t[6294] = 0
      "00000" when "001100010010111", -- t[6295] = 0
      "00000" when "001100010011000", -- t[6296] = 0
      "00000" when "001100010011001", -- t[6297] = 0
      "00000" when "001100010011010", -- t[6298] = 0
      "00000" when "001100010011011", -- t[6299] = 0
      "00000" when "001100010011100", -- t[6300] = 0
      "00000" when "001100010011101", -- t[6301] = 0
      "00000" when "001100010011110", -- t[6302] = 0
      "00000" when "001100010011111", -- t[6303] = 0
      "00000" when "001100010100000", -- t[6304] = 0
      "00000" when "001100010100001", -- t[6305] = 0
      "00000" when "001100010100010", -- t[6306] = 0
      "00000" when "001100010100011", -- t[6307] = 0
      "00000" when "001100010100100", -- t[6308] = 0
      "00000" when "001100010100101", -- t[6309] = 0
      "00000" when "001100010100110", -- t[6310] = 0
      "00000" when "001100010100111", -- t[6311] = 0
      "00000" when "001100010101000", -- t[6312] = 0
      "00000" when "001100010101001", -- t[6313] = 0
      "00000" when "001100010101010", -- t[6314] = 0
      "00000" when "001100010101011", -- t[6315] = 0
      "00000" when "001100010101100", -- t[6316] = 0
      "00000" when "001100010101101", -- t[6317] = 0
      "00000" when "001100010101110", -- t[6318] = 0
      "00000" when "001100010101111", -- t[6319] = 0
      "00000" when "001100010110000", -- t[6320] = 0
      "00000" when "001100010110001", -- t[6321] = 0
      "00000" when "001100010110010", -- t[6322] = 0
      "00000" when "001100010110011", -- t[6323] = 0
      "00000" when "001100010110100", -- t[6324] = 0
      "00000" when "001100010110101", -- t[6325] = 0
      "00000" when "001100010110110", -- t[6326] = 0
      "00000" when "001100010110111", -- t[6327] = 0
      "00000" when "001100010111000", -- t[6328] = 0
      "00000" when "001100010111001", -- t[6329] = 0
      "00000" when "001100010111010", -- t[6330] = 0
      "00000" when "001100010111011", -- t[6331] = 0
      "00000" when "001100010111100", -- t[6332] = 0
      "00000" when "001100010111101", -- t[6333] = 0
      "00000" when "001100010111110", -- t[6334] = 0
      "00000" when "001100010111111", -- t[6335] = 0
      "00000" when "001100011000000", -- t[6336] = 0
      "00000" when "001100011000001", -- t[6337] = 0
      "00000" when "001100011000010", -- t[6338] = 0
      "00000" when "001100011000011", -- t[6339] = 0
      "00000" when "001100011000100", -- t[6340] = 0
      "00000" when "001100011000101", -- t[6341] = 0
      "00000" when "001100011000110", -- t[6342] = 0
      "00000" when "001100011000111", -- t[6343] = 0
      "00000" when "001100011001000", -- t[6344] = 0
      "00000" when "001100011001001", -- t[6345] = 0
      "00000" when "001100011001010", -- t[6346] = 0
      "00000" when "001100011001011", -- t[6347] = 0
      "00000" when "001100011001100", -- t[6348] = 0
      "00000" when "001100011001101", -- t[6349] = 0
      "00000" when "001100011001110", -- t[6350] = 0
      "00000" when "001100011001111", -- t[6351] = 0
      "00000" when "001100011010000", -- t[6352] = 0
      "00000" when "001100011010001", -- t[6353] = 0
      "00000" when "001100011010010", -- t[6354] = 0
      "00000" when "001100011010011", -- t[6355] = 0
      "00000" when "001100011010100", -- t[6356] = 0
      "00000" when "001100011010101", -- t[6357] = 0
      "00000" when "001100011010110", -- t[6358] = 0
      "00000" when "001100011010111", -- t[6359] = 0
      "00000" when "001100011011000", -- t[6360] = 0
      "00000" when "001100011011001", -- t[6361] = 0
      "00000" when "001100011011010", -- t[6362] = 0
      "00000" when "001100011011011", -- t[6363] = 0
      "00000" when "001100011011100", -- t[6364] = 0
      "00000" when "001100011011101", -- t[6365] = 0
      "00000" when "001100011011110", -- t[6366] = 0
      "00000" when "001100011011111", -- t[6367] = 0
      "00000" when "001100011100000", -- t[6368] = 0
      "00000" when "001100011100001", -- t[6369] = 0
      "00000" when "001100011100010", -- t[6370] = 0
      "00000" when "001100011100011", -- t[6371] = 0
      "00000" when "001100011100100", -- t[6372] = 0
      "00000" when "001100011100101", -- t[6373] = 0
      "00000" when "001100011100110", -- t[6374] = 0
      "00000" when "001100011100111", -- t[6375] = 0
      "00000" when "001100011101000", -- t[6376] = 0
      "00000" when "001100011101001", -- t[6377] = 0
      "00000" when "001100011101010", -- t[6378] = 0
      "00000" when "001100011101011", -- t[6379] = 0
      "00000" when "001100011101100", -- t[6380] = 0
      "00000" when "001100011101101", -- t[6381] = 0
      "00000" when "001100011101110", -- t[6382] = 0
      "00000" when "001100011101111", -- t[6383] = 0
      "00000" when "001100011110000", -- t[6384] = 0
      "00000" when "001100011110001", -- t[6385] = 0
      "00000" when "001100011110010", -- t[6386] = 0
      "00000" when "001100011110011", -- t[6387] = 0
      "00000" when "001100011110100", -- t[6388] = 0
      "00000" when "001100011110101", -- t[6389] = 0
      "00000" when "001100011110110", -- t[6390] = 0
      "00000" when "001100011110111", -- t[6391] = 0
      "00000" when "001100011111000", -- t[6392] = 0
      "00000" when "001100011111001", -- t[6393] = 0
      "00000" when "001100011111010", -- t[6394] = 0
      "00000" when "001100011111011", -- t[6395] = 0
      "00000" when "001100011111100", -- t[6396] = 0
      "00000" when "001100011111101", -- t[6397] = 0
      "00000" when "001100011111110", -- t[6398] = 0
      "00000" when "001100011111111", -- t[6399] = 0
      "00000" when "001100100000000", -- t[6400] = 0
      "00000" when "001100100000001", -- t[6401] = 0
      "00000" when "001100100000010", -- t[6402] = 0
      "00000" when "001100100000011", -- t[6403] = 0
      "00000" when "001100100000100", -- t[6404] = 0
      "00000" when "001100100000101", -- t[6405] = 0
      "00000" when "001100100000110", -- t[6406] = 0
      "00000" when "001100100000111", -- t[6407] = 0
      "00000" when "001100100001000", -- t[6408] = 0
      "00000" when "001100100001001", -- t[6409] = 0
      "00000" when "001100100001010", -- t[6410] = 0
      "00000" when "001100100001011", -- t[6411] = 0
      "00000" when "001100100001100", -- t[6412] = 0
      "00000" when "001100100001101", -- t[6413] = 0
      "00000" when "001100100001110", -- t[6414] = 0
      "00000" when "001100100001111", -- t[6415] = 0
      "00000" when "001100100010000", -- t[6416] = 0
      "00000" when "001100100010001", -- t[6417] = 0
      "00000" when "001100100010010", -- t[6418] = 0
      "00000" when "001100100010011", -- t[6419] = 0
      "00000" when "001100100010100", -- t[6420] = 0
      "00000" when "001100100010101", -- t[6421] = 0
      "00000" when "001100100010110", -- t[6422] = 0
      "00000" when "001100100010111", -- t[6423] = 0
      "00000" when "001100100011000", -- t[6424] = 0
      "00000" when "001100100011001", -- t[6425] = 0
      "00000" when "001100100011010", -- t[6426] = 0
      "00000" when "001100100011011", -- t[6427] = 0
      "00000" when "001100100011100", -- t[6428] = 0
      "00000" when "001100100011101", -- t[6429] = 0
      "00000" when "001100100011110", -- t[6430] = 0
      "00000" when "001100100011111", -- t[6431] = 0
      "00000" when "001100100100000", -- t[6432] = 0
      "00000" when "001100100100001", -- t[6433] = 0
      "00000" when "001100100100010", -- t[6434] = 0
      "00000" when "001100100100011", -- t[6435] = 0
      "00000" when "001100100100100", -- t[6436] = 0
      "00000" when "001100100100101", -- t[6437] = 0
      "00000" when "001100100100110", -- t[6438] = 0
      "00000" when "001100100100111", -- t[6439] = 0
      "00000" when "001100100101000", -- t[6440] = 0
      "00000" when "001100100101001", -- t[6441] = 0
      "00000" when "001100100101010", -- t[6442] = 0
      "00000" when "001100100101011", -- t[6443] = 0
      "00000" when "001100100101100", -- t[6444] = 0
      "00000" when "001100100101101", -- t[6445] = 0
      "00000" when "001100100101110", -- t[6446] = 0
      "00000" when "001100100101111", -- t[6447] = 0
      "00000" when "001100100110000", -- t[6448] = 0
      "00000" when "001100100110001", -- t[6449] = 0
      "00000" when "001100100110010", -- t[6450] = 0
      "00000" when "001100100110011", -- t[6451] = 0
      "00000" when "001100100110100", -- t[6452] = 0
      "00000" when "001100100110101", -- t[6453] = 0
      "00000" when "001100100110110", -- t[6454] = 0
      "00000" when "001100100110111", -- t[6455] = 0
      "00000" when "001100100111000", -- t[6456] = 0
      "00000" when "001100100111001", -- t[6457] = 0
      "00000" when "001100100111010", -- t[6458] = 0
      "00000" when "001100100111011", -- t[6459] = 0
      "00000" when "001100100111100", -- t[6460] = 0
      "00000" when "001100100111101", -- t[6461] = 0
      "00000" when "001100100111110", -- t[6462] = 0
      "00000" when "001100100111111", -- t[6463] = 0
      "00000" when "001100101000000", -- t[6464] = 0
      "00000" when "001100101000001", -- t[6465] = 0
      "00000" when "001100101000010", -- t[6466] = 0
      "00000" when "001100101000011", -- t[6467] = 0
      "00000" when "001100101000100", -- t[6468] = 0
      "00000" when "001100101000101", -- t[6469] = 0
      "00000" when "001100101000110", -- t[6470] = 0
      "00000" when "001100101000111", -- t[6471] = 0
      "00000" when "001100101001000", -- t[6472] = 0
      "00000" when "001100101001001", -- t[6473] = 0
      "00000" when "001100101001010", -- t[6474] = 0
      "00000" when "001100101001011", -- t[6475] = 0
      "00000" when "001100101001100", -- t[6476] = 0
      "00000" when "001100101001101", -- t[6477] = 0
      "00000" when "001100101001110", -- t[6478] = 0
      "00000" when "001100101001111", -- t[6479] = 0
      "00000" when "001100101010000", -- t[6480] = 0
      "00000" when "001100101010001", -- t[6481] = 0
      "00000" when "001100101010010", -- t[6482] = 0
      "00000" when "001100101010011", -- t[6483] = 0
      "00000" when "001100101010100", -- t[6484] = 0
      "00000" when "001100101010101", -- t[6485] = 0
      "00000" when "001100101010110", -- t[6486] = 0
      "00000" when "001100101010111", -- t[6487] = 0
      "00000" when "001100101011000", -- t[6488] = 0
      "00000" when "001100101011001", -- t[6489] = 0
      "00000" when "001100101011010", -- t[6490] = 0
      "00000" when "001100101011011", -- t[6491] = 0
      "00000" when "001100101011100", -- t[6492] = 0
      "00000" when "001100101011101", -- t[6493] = 0
      "00000" when "001100101011110", -- t[6494] = 0
      "00000" when "001100101011111", -- t[6495] = 0
      "00000" when "001100101100000", -- t[6496] = 0
      "00000" when "001100101100001", -- t[6497] = 0
      "00000" when "001100101100010", -- t[6498] = 0
      "00000" when "001100101100011", -- t[6499] = 0
      "00000" when "001100101100100", -- t[6500] = 0
      "00000" when "001100101100101", -- t[6501] = 0
      "00000" when "001100101100110", -- t[6502] = 0
      "00000" when "001100101100111", -- t[6503] = 0
      "00000" when "001100101101000", -- t[6504] = 0
      "00000" when "001100101101001", -- t[6505] = 0
      "00000" when "001100101101010", -- t[6506] = 0
      "00000" when "001100101101011", -- t[6507] = 0
      "00000" when "001100101101100", -- t[6508] = 0
      "00000" when "001100101101101", -- t[6509] = 0
      "00000" when "001100101101110", -- t[6510] = 0
      "00000" when "001100101101111", -- t[6511] = 0
      "00000" when "001100101110000", -- t[6512] = 0
      "00000" when "001100101110001", -- t[6513] = 0
      "00000" when "001100101110010", -- t[6514] = 0
      "00000" when "001100101110011", -- t[6515] = 0
      "00000" when "001100101110100", -- t[6516] = 0
      "00000" when "001100101110101", -- t[6517] = 0
      "00000" when "001100101110110", -- t[6518] = 0
      "00000" when "001100101110111", -- t[6519] = 0
      "00000" when "001100101111000", -- t[6520] = 0
      "00000" when "001100101111001", -- t[6521] = 0
      "00000" when "001100101111010", -- t[6522] = 0
      "00000" when "001100101111011", -- t[6523] = 0
      "00000" when "001100101111100", -- t[6524] = 0
      "00000" when "001100101111101", -- t[6525] = 0
      "00000" when "001100101111110", -- t[6526] = 0
      "00000" when "001100101111111", -- t[6527] = 0
      "00000" when "001100110000000", -- t[6528] = 0
      "00000" when "001100110000001", -- t[6529] = 0
      "00000" when "001100110000010", -- t[6530] = 0
      "00000" when "001100110000011", -- t[6531] = 0
      "00000" when "001100110000100", -- t[6532] = 0
      "00000" when "001100110000101", -- t[6533] = 0
      "00000" when "001100110000110", -- t[6534] = 0
      "00000" when "001100110000111", -- t[6535] = 0
      "00000" when "001100110001000", -- t[6536] = 0
      "00000" when "001100110001001", -- t[6537] = 0
      "00000" when "001100110001010", -- t[6538] = 0
      "00000" when "001100110001011", -- t[6539] = 0
      "00000" when "001100110001100", -- t[6540] = 0
      "00000" when "001100110001101", -- t[6541] = 0
      "00000" when "001100110001110", -- t[6542] = 0
      "00000" when "001100110001111", -- t[6543] = 0
      "00000" when "001100110010000", -- t[6544] = 0
      "00000" when "001100110010001", -- t[6545] = 0
      "00000" when "001100110010010", -- t[6546] = 0
      "00000" when "001100110010011", -- t[6547] = 0
      "00000" when "001100110010100", -- t[6548] = 0
      "00000" when "001100110010101", -- t[6549] = 0
      "00000" when "001100110010110", -- t[6550] = 0
      "00000" when "001100110010111", -- t[6551] = 0
      "00000" when "001100110011000", -- t[6552] = 0
      "00000" when "001100110011001", -- t[6553] = 0
      "00000" when "001100110011010", -- t[6554] = 0
      "00000" when "001100110011011", -- t[6555] = 0
      "00000" when "001100110011100", -- t[6556] = 0
      "00000" when "001100110011101", -- t[6557] = 0
      "00000" when "001100110011110", -- t[6558] = 0
      "00000" when "001100110011111", -- t[6559] = 0
      "00000" when "001100110100000", -- t[6560] = 0
      "00000" when "001100110100001", -- t[6561] = 0
      "00000" when "001100110100010", -- t[6562] = 0
      "00000" when "001100110100011", -- t[6563] = 0
      "00000" when "001100110100100", -- t[6564] = 0
      "00000" when "001100110100101", -- t[6565] = 0
      "00000" when "001100110100110", -- t[6566] = 0
      "00000" when "001100110100111", -- t[6567] = 0
      "00000" when "001100110101000", -- t[6568] = 0
      "00000" when "001100110101001", -- t[6569] = 0
      "00000" when "001100110101010", -- t[6570] = 0
      "00000" when "001100110101011", -- t[6571] = 0
      "00000" when "001100110101100", -- t[6572] = 0
      "00000" when "001100110101101", -- t[6573] = 0
      "00000" when "001100110101110", -- t[6574] = 0
      "00000" when "001100110101111", -- t[6575] = 0
      "00000" when "001100110110000", -- t[6576] = 0
      "00000" when "001100110110001", -- t[6577] = 0
      "00000" when "001100110110010", -- t[6578] = 0
      "00000" when "001100110110011", -- t[6579] = 0
      "00000" when "001100110110100", -- t[6580] = 0
      "00000" when "001100110110101", -- t[6581] = 0
      "00000" when "001100110110110", -- t[6582] = 0
      "00000" when "001100110110111", -- t[6583] = 0
      "00000" when "001100110111000", -- t[6584] = 0
      "00000" when "001100110111001", -- t[6585] = 0
      "00000" when "001100110111010", -- t[6586] = 0
      "00000" when "001100110111011", -- t[6587] = 0
      "00000" when "001100110111100", -- t[6588] = 0
      "00000" when "001100110111101", -- t[6589] = 0
      "00000" when "001100110111110", -- t[6590] = 0
      "00000" when "001100110111111", -- t[6591] = 0
      "00000" when "001100111000000", -- t[6592] = 0
      "00000" when "001100111000001", -- t[6593] = 0
      "00000" when "001100111000010", -- t[6594] = 0
      "00000" when "001100111000011", -- t[6595] = 0
      "00000" when "001100111000100", -- t[6596] = 0
      "00000" when "001100111000101", -- t[6597] = 0
      "00000" when "001100111000110", -- t[6598] = 0
      "00000" when "001100111000111", -- t[6599] = 0
      "00000" when "001100111001000", -- t[6600] = 0
      "00000" when "001100111001001", -- t[6601] = 0
      "00000" when "001100111001010", -- t[6602] = 0
      "00000" when "001100111001011", -- t[6603] = 0
      "00000" when "001100111001100", -- t[6604] = 0
      "00000" when "001100111001101", -- t[6605] = 0
      "00000" when "001100111001110", -- t[6606] = 0
      "00000" when "001100111001111", -- t[6607] = 0
      "00000" when "001100111010000", -- t[6608] = 0
      "00000" when "001100111010001", -- t[6609] = 0
      "00000" when "001100111010010", -- t[6610] = 0
      "00000" when "001100111010011", -- t[6611] = 0
      "00000" when "001100111010100", -- t[6612] = 0
      "00000" when "001100111010101", -- t[6613] = 0
      "00000" when "001100111010110", -- t[6614] = 0
      "00000" when "001100111010111", -- t[6615] = 0
      "00000" when "001100111011000", -- t[6616] = 0
      "00000" when "001100111011001", -- t[6617] = 0
      "00000" when "001100111011010", -- t[6618] = 0
      "00000" when "001100111011011", -- t[6619] = 0
      "00000" when "001100111011100", -- t[6620] = 0
      "00000" when "001100111011101", -- t[6621] = 0
      "00000" when "001100111011110", -- t[6622] = 0
      "00000" when "001100111011111", -- t[6623] = 0
      "00000" when "001100111100000", -- t[6624] = 0
      "00000" when "001100111100001", -- t[6625] = 0
      "00000" when "001100111100010", -- t[6626] = 0
      "00000" when "001100111100011", -- t[6627] = 0
      "00000" when "001100111100100", -- t[6628] = 0
      "00000" when "001100111100101", -- t[6629] = 0
      "00000" when "001100111100110", -- t[6630] = 0
      "00000" when "001100111100111", -- t[6631] = 0
      "00000" when "001100111101000", -- t[6632] = 0
      "00000" when "001100111101001", -- t[6633] = 0
      "00000" when "001100111101010", -- t[6634] = 0
      "00000" when "001100111101011", -- t[6635] = 0
      "00000" when "001100111101100", -- t[6636] = 0
      "00000" when "001100111101101", -- t[6637] = 0
      "00000" when "001100111101110", -- t[6638] = 0
      "00000" when "001100111101111", -- t[6639] = 0
      "00000" when "001100111110000", -- t[6640] = 0
      "00000" when "001100111110001", -- t[6641] = 0
      "00000" when "001100111110010", -- t[6642] = 0
      "00000" when "001100111110011", -- t[6643] = 0
      "00000" when "001100111110100", -- t[6644] = 0
      "00000" when "001100111110101", -- t[6645] = 0
      "00000" when "001100111110110", -- t[6646] = 0
      "00000" when "001100111110111", -- t[6647] = 0
      "00000" when "001100111111000", -- t[6648] = 0
      "00000" when "001100111111001", -- t[6649] = 0
      "00000" when "001100111111010", -- t[6650] = 0
      "00000" when "001100111111011", -- t[6651] = 0
      "00000" when "001100111111100", -- t[6652] = 0
      "00000" when "001100111111101", -- t[6653] = 0
      "00000" when "001100111111110", -- t[6654] = 0
      "00000" when "001100111111111", -- t[6655] = 0
      "00000" when "001101000000000", -- t[6656] = 0
      "00000" when "001101000000001", -- t[6657] = 0
      "00000" when "001101000000010", -- t[6658] = 0
      "00000" when "001101000000011", -- t[6659] = 0
      "00000" when "001101000000100", -- t[6660] = 0
      "00000" when "001101000000101", -- t[6661] = 0
      "00000" when "001101000000110", -- t[6662] = 0
      "00000" when "001101000000111", -- t[6663] = 0
      "00000" when "001101000001000", -- t[6664] = 0
      "00000" when "001101000001001", -- t[6665] = 0
      "00000" when "001101000001010", -- t[6666] = 0
      "00000" when "001101000001011", -- t[6667] = 0
      "00000" when "001101000001100", -- t[6668] = 0
      "00000" when "001101000001101", -- t[6669] = 0
      "00000" when "001101000001110", -- t[6670] = 0
      "00000" when "001101000001111", -- t[6671] = 0
      "00000" when "001101000010000", -- t[6672] = 0
      "00000" when "001101000010001", -- t[6673] = 0
      "00000" when "001101000010010", -- t[6674] = 0
      "00000" when "001101000010011", -- t[6675] = 0
      "00000" when "001101000010100", -- t[6676] = 0
      "00000" when "001101000010101", -- t[6677] = 0
      "00000" when "001101000010110", -- t[6678] = 0
      "00000" when "001101000010111", -- t[6679] = 0
      "00000" when "001101000011000", -- t[6680] = 0
      "00000" when "001101000011001", -- t[6681] = 0
      "00000" when "001101000011010", -- t[6682] = 0
      "00000" when "001101000011011", -- t[6683] = 0
      "00000" when "001101000011100", -- t[6684] = 0
      "00000" when "001101000011101", -- t[6685] = 0
      "00000" when "001101000011110", -- t[6686] = 0
      "00000" when "001101000011111", -- t[6687] = 0
      "00000" when "001101000100000", -- t[6688] = 0
      "00000" when "001101000100001", -- t[6689] = 0
      "00000" when "001101000100010", -- t[6690] = 0
      "00000" when "001101000100011", -- t[6691] = 0
      "00000" when "001101000100100", -- t[6692] = 0
      "00000" when "001101000100101", -- t[6693] = 0
      "00000" when "001101000100110", -- t[6694] = 0
      "00000" when "001101000100111", -- t[6695] = 0
      "00000" when "001101000101000", -- t[6696] = 0
      "00000" when "001101000101001", -- t[6697] = 0
      "00000" when "001101000101010", -- t[6698] = 0
      "00000" when "001101000101011", -- t[6699] = 0
      "00000" when "001101000101100", -- t[6700] = 0
      "00000" when "001101000101101", -- t[6701] = 0
      "00000" when "001101000101110", -- t[6702] = 0
      "00000" when "001101000101111", -- t[6703] = 0
      "00000" when "001101000110000", -- t[6704] = 0
      "00000" when "001101000110001", -- t[6705] = 0
      "00000" when "001101000110010", -- t[6706] = 0
      "00000" when "001101000110011", -- t[6707] = 0
      "00000" when "001101000110100", -- t[6708] = 0
      "00000" when "001101000110101", -- t[6709] = 0
      "00000" when "001101000110110", -- t[6710] = 0
      "00000" when "001101000110111", -- t[6711] = 0
      "00000" when "001101000111000", -- t[6712] = 0
      "00000" when "001101000111001", -- t[6713] = 0
      "00000" when "001101000111010", -- t[6714] = 0
      "00000" when "001101000111011", -- t[6715] = 0
      "00000" when "001101000111100", -- t[6716] = 0
      "00000" when "001101000111101", -- t[6717] = 0
      "00000" when "001101000111110", -- t[6718] = 0
      "00000" when "001101000111111", -- t[6719] = 0
      "00000" when "001101001000000", -- t[6720] = 0
      "00000" when "001101001000001", -- t[6721] = 0
      "00000" when "001101001000010", -- t[6722] = 0
      "00000" when "001101001000011", -- t[6723] = 0
      "00000" when "001101001000100", -- t[6724] = 0
      "00000" when "001101001000101", -- t[6725] = 0
      "00000" when "001101001000110", -- t[6726] = 0
      "00000" when "001101001000111", -- t[6727] = 0
      "00000" when "001101001001000", -- t[6728] = 0
      "00000" when "001101001001001", -- t[6729] = 0
      "00000" when "001101001001010", -- t[6730] = 0
      "00000" when "001101001001011", -- t[6731] = 0
      "00000" when "001101001001100", -- t[6732] = 0
      "00000" when "001101001001101", -- t[6733] = 0
      "00000" when "001101001001110", -- t[6734] = 0
      "00000" when "001101001001111", -- t[6735] = 0
      "00000" when "001101001010000", -- t[6736] = 0
      "00000" when "001101001010001", -- t[6737] = 0
      "00000" when "001101001010010", -- t[6738] = 0
      "00000" when "001101001010011", -- t[6739] = 0
      "00000" when "001101001010100", -- t[6740] = 0
      "00000" when "001101001010101", -- t[6741] = 0
      "00000" when "001101001010110", -- t[6742] = 0
      "00000" when "001101001010111", -- t[6743] = 0
      "00000" when "001101001011000", -- t[6744] = 0
      "00000" when "001101001011001", -- t[6745] = 0
      "00000" when "001101001011010", -- t[6746] = 0
      "00000" when "001101001011011", -- t[6747] = 0
      "00000" when "001101001011100", -- t[6748] = 0
      "00000" when "001101001011101", -- t[6749] = 0
      "00000" when "001101001011110", -- t[6750] = 0
      "00000" when "001101001011111", -- t[6751] = 0
      "00000" when "001101001100000", -- t[6752] = 0
      "00000" when "001101001100001", -- t[6753] = 0
      "00000" when "001101001100010", -- t[6754] = 0
      "00000" when "001101001100011", -- t[6755] = 0
      "00000" when "001101001100100", -- t[6756] = 0
      "00000" when "001101001100101", -- t[6757] = 0
      "00000" when "001101001100110", -- t[6758] = 0
      "00000" when "001101001100111", -- t[6759] = 0
      "00000" when "001101001101000", -- t[6760] = 0
      "00000" when "001101001101001", -- t[6761] = 0
      "00000" when "001101001101010", -- t[6762] = 0
      "00000" when "001101001101011", -- t[6763] = 0
      "00000" when "001101001101100", -- t[6764] = 0
      "00000" when "001101001101101", -- t[6765] = 0
      "00000" when "001101001101110", -- t[6766] = 0
      "00000" when "001101001101111", -- t[6767] = 0
      "00000" when "001101001110000", -- t[6768] = 0
      "00000" when "001101001110001", -- t[6769] = 0
      "00000" when "001101001110010", -- t[6770] = 0
      "00000" when "001101001110011", -- t[6771] = 0
      "00000" when "001101001110100", -- t[6772] = 0
      "00000" when "001101001110101", -- t[6773] = 0
      "00000" when "001101001110110", -- t[6774] = 0
      "00000" when "001101001110111", -- t[6775] = 0
      "00000" when "001101001111000", -- t[6776] = 0
      "00000" when "001101001111001", -- t[6777] = 0
      "00000" when "001101001111010", -- t[6778] = 0
      "00000" when "001101001111011", -- t[6779] = 0
      "00000" when "001101001111100", -- t[6780] = 0
      "00000" when "001101001111101", -- t[6781] = 0
      "00000" when "001101001111110", -- t[6782] = 0
      "00000" when "001101001111111", -- t[6783] = 0
      "00000" when "001101010000000", -- t[6784] = 0
      "00000" when "001101010000001", -- t[6785] = 0
      "00000" when "001101010000010", -- t[6786] = 0
      "00000" when "001101010000011", -- t[6787] = 0
      "00000" when "001101010000100", -- t[6788] = 0
      "00000" when "001101010000101", -- t[6789] = 0
      "00000" when "001101010000110", -- t[6790] = 0
      "00000" when "001101010000111", -- t[6791] = 0
      "00000" when "001101010001000", -- t[6792] = 0
      "00000" when "001101010001001", -- t[6793] = 0
      "00000" when "001101010001010", -- t[6794] = 0
      "00000" when "001101010001011", -- t[6795] = 0
      "00000" when "001101010001100", -- t[6796] = 0
      "00000" when "001101010001101", -- t[6797] = 0
      "00000" when "001101010001110", -- t[6798] = 0
      "00000" when "001101010001111", -- t[6799] = 0
      "00000" when "001101010010000", -- t[6800] = 0
      "00000" when "001101010010001", -- t[6801] = 0
      "00000" when "001101010010010", -- t[6802] = 0
      "00000" when "001101010010011", -- t[6803] = 0
      "00000" when "001101010010100", -- t[6804] = 0
      "00000" when "001101010010101", -- t[6805] = 0
      "00000" when "001101010010110", -- t[6806] = 0
      "00000" when "001101010010111", -- t[6807] = 0
      "00000" when "001101010011000", -- t[6808] = 0
      "00000" when "001101010011001", -- t[6809] = 0
      "00000" when "001101010011010", -- t[6810] = 0
      "00000" when "001101010011011", -- t[6811] = 0
      "00000" when "001101010011100", -- t[6812] = 0
      "00000" when "001101010011101", -- t[6813] = 0
      "00000" when "001101010011110", -- t[6814] = 0
      "00000" when "001101010011111", -- t[6815] = 0
      "00000" when "001101010100000", -- t[6816] = 0
      "00000" when "001101010100001", -- t[6817] = 0
      "00000" when "001101010100010", -- t[6818] = 0
      "00000" when "001101010100011", -- t[6819] = 0
      "00000" when "001101010100100", -- t[6820] = 0
      "00000" when "001101010100101", -- t[6821] = 0
      "00000" when "001101010100110", -- t[6822] = 0
      "00000" when "001101010100111", -- t[6823] = 0
      "00000" when "001101010101000", -- t[6824] = 0
      "00000" when "001101010101001", -- t[6825] = 0
      "00000" when "001101010101010", -- t[6826] = 0
      "00000" when "001101010101011", -- t[6827] = 0
      "00000" when "001101010101100", -- t[6828] = 0
      "00000" when "001101010101101", -- t[6829] = 0
      "00000" when "001101010101110", -- t[6830] = 0
      "00000" when "001101010101111", -- t[6831] = 0
      "00000" when "001101010110000", -- t[6832] = 0
      "00000" when "001101010110001", -- t[6833] = 0
      "00000" when "001101010110010", -- t[6834] = 0
      "00000" when "001101010110011", -- t[6835] = 0
      "00000" when "001101010110100", -- t[6836] = 0
      "00000" when "001101010110101", -- t[6837] = 0
      "00000" when "001101010110110", -- t[6838] = 0
      "00000" when "001101010110111", -- t[6839] = 0
      "00000" when "001101010111000", -- t[6840] = 0
      "00000" when "001101010111001", -- t[6841] = 0
      "00000" when "001101010111010", -- t[6842] = 0
      "00000" when "001101010111011", -- t[6843] = 0
      "00000" when "001101010111100", -- t[6844] = 0
      "00000" when "001101010111101", -- t[6845] = 0
      "00000" when "001101010111110", -- t[6846] = 0
      "00000" when "001101010111111", -- t[6847] = 0
      "00000" when "001101011000000", -- t[6848] = 0
      "00000" when "001101011000001", -- t[6849] = 0
      "00000" when "001101011000010", -- t[6850] = 0
      "00000" when "001101011000011", -- t[6851] = 0
      "00000" when "001101011000100", -- t[6852] = 0
      "00000" when "001101011000101", -- t[6853] = 0
      "00000" when "001101011000110", -- t[6854] = 0
      "00000" when "001101011000111", -- t[6855] = 0
      "00000" when "001101011001000", -- t[6856] = 0
      "00000" when "001101011001001", -- t[6857] = 0
      "00000" when "001101011001010", -- t[6858] = 0
      "00000" when "001101011001011", -- t[6859] = 0
      "00000" when "001101011001100", -- t[6860] = 0
      "00000" when "001101011001101", -- t[6861] = 0
      "00000" when "001101011001110", -- t[6862] = 0
      "00000" when "001101011001111", -- t[6863] = 0
      "00000" when "001101011010000", -- t[6864] = 0
      "00000" when "001101011010001", -- t[6865] = 0
      "00000" when "001101011010010", -- t[6866] = 0
      "00000" when "001101011010011", -- t[6867] = 0
      "00000" when "001101011010100", -- t[6868] = 0
      "00000" when "001101011010101", -- t[6869] = 0
      "00000" when "001101011010110", -- t[6870] = 0
      "00000" when "001101011010111", -- t[6871] = 0
      "00000" when "001101011011000", -- t[6872] = 0
      "00000" when "001101011011001", -- t[6873] = 0
      "00000" when "001101011011010", -- t[6874] = 0
      "00000" when "001101011011011", -- t[6875] = 0
      "00000" when "001101011011100", -- t[6876] = 0
      "00000" when "001101011011101", -- t[6877] = 0
      "00000" when "001101011011110", -- t[6878] = 0
      "00000" when "001101011011111", -- t[6879] = 0
      "00000" when "001101011100000", -- t[6880] = 0
      "00000" when "001101011100001", -- t[6881] = 0
      "00000" when "001101011100010", -- t[6882] = 0
      "00000" when "001101011100011", -- t[6883] = 0
      "00000" when "001101011100100", -- t[6884] = 0
      "00000" when "001101011100101", -- t[6885] = 0
      "00000" when "001101011100110", -- t[6886] = 0
      "00000" when "001101011100111", -- t[6887] = 0
      "00000" when "001101011101000", -- t[6888] = 0
      "00000" when "001101011101001", -- t[6889] = 0
      "00000" when "001101011101010", -- t[6890] = 0
      "00000" when "001101011101011", -- t[6891] = 0
      "00000" when "001101011101100", -- t[6892] = 0
      "00000" when "001101011101101", -- t[6893] = 0
      "00000" when "001101011101110", -- t[6894] = 0
      "00000" when "001101011101111", -- t[6895] = 0
      "00000" when "001101011110000", -- t[6896] = 0
      "00000" when "001101011110001", -- t[6897] = 0
      "00000" when "001101011110010", -- t[6898] = 0
      "00000" when "001101011110011", -- t[6899] = 0
      "00000" when "001101011110100", -- t[6900] = 0
      "00000" when "001101011110101", -- t[6901] = 0
      "00000" when "001101011110110", -- t[6902] = 0
      "00000" when "001101011110111", -- t[6903] = 0
      "00000" when "001101011111000", -- t[6904] = 0
      "00000" when "001101011111001", -- t[6905] = 0
      "00000" when "001101011111010", -- t[6906] = 0
      "00000" when "001101011111011", -- t[6907] = 0
      "00000" when "001101011111100", -- t[6908] = 0
      "00000" when "001101011111101", -- t[6909] = 0
      "00000" when "001101011111110", -- t[6910] = 0
      "00000" when "001101011111111", -- t[6911] = 0
      "00000" when "001101100000000", -- t[6912] = 0
      "00000" when "001101100000001", -- t[6913] = 0
      "00000" when "001101100000010", -- t[6914] = 0
      "00000" when "001101100000011", -- t[6915] = 0
      "00000" when "001101100000100", -- t[6916] = 0
      "00000" when "001101100000101", -- t[6917] = 0
      "00000" when "001101100000110", -- t[6918] = 0
      "00000" when "001101100000111", -- t[6919] = 0
      "00000" when "001101100001000", -- t[6920] = 0
      "00000" when "001101100001001", -- t[6921] = 0
      "00000" when "001101100001010", -- t[6922] = 0
      "00000" when "001101100001011", -- t[6923] = 0
      "00000" when "001101100001100", -- t[6924] = 0
      "00000" when "001101100001101", -- t[6925] = 0
      "00000" when "001101100001110", -- t[6926] = 0
      "00000" when "001101100001111", -- t[6927] = 0
      "00000" when "001101100010000", -- t[6928] = 0
      "00000" when "001101100010001", -- t[6929] = 0
      "00000" when "001101100010010", -- t[6930] = 0
      "00000" when "001101100010011", -- t[6931] = 0
      "00000" when "001101100010100", -- t[6932] = 0
      "00000" when "001101100010101", -- t[6933] = 0
      "00000" when "001101100010110", -- t[6934] = 0
      "00000" when "001101100010111", -- t[6935] = 0
      "00000" when "001101100011000", -- t[6936] = 0
      "00000" when "001101100011001", -- t[6937] = 0
      "00000" when "001101100011010", -- t[6938] = 0
      "00000" when "001101100011011", -- t[6939] = 0
      "00000" when "001101100011100", -- t[6940] = 0
      "00000" when "001101100011101", -- t[6941] = 0
      "00000" when "001101100011110", -- t[6942] = 0
      "00000" when "001101100011111", -- t[6943] = 0
      "00000" when "001101100100000", -- t[6944] = 0
      "00000" when "001101100100001", -- t[6945] = 0
      "00000" when "001101100100010", -- t[6946] = 0
      "00000" when "001101100100011", -- t[6947] = 0
      "00000" when "001101100100100", -- t[6948] = 0
      "00000" when "001101100100101", -- t[6949] = 0
      "00000" when "001101100100110", -- t[6950] = 0
      "00000" when "001101100100111", -- t[6951] = 0
      "00000" when "001101100101000", -- t[6952] = 0
      "00000" when "001101100101001", -- t[6953] = 0
      "00000" when "001101100101010", -- t[6954] = 0
      "00000" when "001101100101011", -- t[6955] = 0
      "00000" when "001101100101100", -- t[6956] = 0
      "00000" when "001101100101101", -- t[6957] = 0
      "00000" when "001101100101110", -- t[6958] = 0
      "00000" when "001101100101111", -- t[6959] = 0
      "00000" when "001101100110000", -- t[6960] = 0
      "00000" when "001101100110001", -- t[6961] = 0
      "00000" when "001101100110010", -- t[6962] = 0
      "00000" when "001101100110011", -- t[6963] = 0
      "00000" when "001101100110100", -- t[6964] = 0
      "00000" when "001101100110101", -- t[6965] = 0
      "00000" when "001101100110110", -- t[6966] = 0
      "00000" when "001101100110111", -- t[6967] = 0
      "00000" when "001101100111000", -- t[6968] = 0
      "00000" when "001101100111001", -- t[6969] = 0
      "00000" when "001101100111010", -- t[6970] = 0
      "00000" when "001101100111011", -- t[6971] = 0
      "00000" when "001101100111100", -- t[6972] = 0
      "00000" when "001101100111101", -- t[6973] = 0
      "00000" when "001101100111110", -- t[6974] = 0
      "00000" when "001101100111111", -- t[6975] = 0
      "00000" when "001101101000000", -- t[6976] = 0
      "00000" when "001101101000001", -- t[6977] = 0
      "00000" when "001101101000010", -- t[6978] = 0
      "00000" when "001101101000011", -- t[6979] = 0
      "00000" when "001101101000100", -- t[6980] = 0
      "00000" when "001101101000101", -- t[6981] = 0
      "00000" when "001101101000110", -- t[6982] = 0
      "00000" when "001101101000111", -- t[6983] = 0
      "00000" when "001101101001000", -- t[6984] = 0
      "00000" when "001101101001001", -- t[6985] = 0
      "00000" when "001101101001010", -- t[6986] = 0
      "00000" when "001101101001011", -- t[6987] = 0
      "00000" when "001101101001100", -- t[6988] = 0
      "00000" when "001101101001101", -- t[6989] = 0
      "00000" when "001101101001110", -- t[6990] = 0
      "00000" when "001101101001111", -- t[6991] = 0
      "00000" when "001101101010000", -- t[6992] = 0
      "00000" when "001101101010001", -- t[6993] = 0
      "00000" when "001101101010010", -- t[6994] = 0
      "00000" when "001101101010011", -- t[6995] = 0
      "00000" when "001101101010100", -- t[6996] = 0
      "00000" when "001101101010101", -- t[6997] = 0
      "00000" when "001101101010110", -- t[6998] = 0
      "00000" when "001101101010111", -- t[6999] = 0
      "00000" when "001101101011000", -- t[7000] = 0
      "00000" when "001101101011001", -- t[7001] = 0
      "00000" when "001101101011010", -- t[7002] = 0
      "00000" when "001101101011011", -- t[7003] = 0
      "00000" when "001101101011100", -- t[7004] = 0
      "00000" when "001101101011101", -- t[7005] = 0
      "00000" when "001101101011110", -- t[7006] = 0
      "00000" when "001101101011111", -- t[7007] = 0
      "00000" when "001101101100000", -- t[7008] = 0
      "00000" when "001101101100001", -- t[7009] = 0
      "00000" when "001101101100010", -- t[7010] = 0
      "00000" when "001101101100011", -- t[7011] = 0
      "00000" when "001101101100100", -- t[7012] = 0
      "00000" when "001101101100101", -- t[7013] = 0
      "00000" when "001101101100110", -- t[7014] = 0
      "00000" when "001101101100111", -- t[7015] = 0
      "00000" when "001101101101000", -- t[7016] = 0
      "00000" when "001101101101001", -- t[7017] = 0
      "00000" when "001101101101010", -- t[7018] = 0
      "00000" when "001101101101011", -- t[7019] = 0
      "00000" when "001101101101100", -- t[7020] = 0
      "00000" when "001101101101101", -- t[7021] = 0
      "00000" when "001101101101110", -- t[7022] = 0
      "00000" when "001101101101111", -- t[7023] = 0
      "00000" when "001101101110000", -- t[7024] = 0
      "00000" when "001101101110001", -- t[7025] = 0
      "00000" when "001101101110010", -- t[7026] = 0
      "00000" when "001101101110011", -- t[7027] = 0
      "00000" when "001101101110100", -- t[7028] = 0
      "00000" when "001101101110101", -- t[7029] = 0
      "00000" when "001101101110110", -- t[7030] = 0
      "00000" when "001101101110111", -- t[7031] = 0
      "00000" when "001101101111000", -- t[7032] = 0
      "00000" when "001101101111001", -- t[7033] = 0
      "00000" when "001101101111010", -- t[7034] = 0
      "00000" when "001101101111011", -- t[7035] = 0
      "00000" when "001101101111100", -- t[7036] = 0
      "00000" when "001101101111101", -- t[7037] = 0
      "00000" when "001101101111110", -- t[7038] = 0
      "00000" when "001101101111111", -- t[7039] = 0
      "00000" when "001101110000000", -- t[7040] = 0
      "00000" when "001101110000001", -- t[7041] = 0
      "00000" when "001101110000010", -- t[7042] = 0
      "00000" when "001101110000011", -- t[7043] = 0
      "00000" when "001101110000100", -- t[7044] = 0
      "00000" when "001101110000101", -- t[7045] = 0
      "00000" when "001101110000110", -- t[7046] = 0
      "00000" when "001101110000111", -- t[7047] = 0
      "00000" when "001101110001000", -- t[7048] = 0
      "00000" when "001101110001001", -- t[7049] = 0
      "00000" when "001101110001010", -- t[7050] = 0
      "00000" when "001101110001011", -- t[7051] = 0
      "00000" when "001101110001100", -- t[7052] = 0
      "00000" when "001101110001101", -- t[7053] = 0
      "00000" when "001101110001110", -- t[7054] = 0
      "00000" when "001101110001111", -- t[7055] = 0
      "00000" when "001101110010000", -- t[7056] = 0
      "00000" when "001101110010001", -- t[7057] = 0
      "00000" when "001101110010010", -- t[7058] = 0
      "00000" when "001101110010011", -- t[7059] = 0
      "00000" when "001101110010100", -- t[7060] = 0
      "00000" when "001101110010101", -- t[7061] = 0
      "00000" when "001101110010110", -- t[7062] = 0
      "00000" when "001101110010111", -- t[7063] = 0
      "00000" when "001101110011000", -- t[7064] = 0
      "00000" when "001101110011001", -- t[7065] = 0
      "00000" when "001101110011010", -- t[7066] = 0
      "00000" when "001101110011011", -- t[7067] = 0
      "00000" when "001101110011100", -- t[7068] = 0
      "00000" when "001101110011101", -- t[7069] = 0
      "00000" when "001101110011110", -- t[7070] = 0
      "00000" when "001101110011111", -- t[7071] = 0
      "00000" when "001101110100000", -- t[7072] = 0
      "00000" when "001101110100001", -- t[7073] = 0
      "00000" when "001101110100010", -- t[7074] = 0
      "00000" when "001101110100011", -- t[7075] = 0
      "00000" when "001101110100100", -- t[7076] = 0
      "00000" when "001101110100101", -- t[7077] = 0
      "00000" when "001101110100110", -- t[7078] = 0
      "00000" when "001101110100111", -- t[7079] = 0
      "00000" when "001101110101000", -- t[7080] = 0
      "00000" when "001101110101001", -- t[7081] = 0
      "00000" when "001101110101010", -- t[7082] = 0
      "00000" when "001101110101011", -- t[7083] = 0
      "00000" when "001101110101100", -- t[7084] = 0
      "00000" when "001101110101101", -- t[7085] = 0
      "00000" when "001101110101110", -- t[7086] = 0
      "00000" when "001101110101111", -- t[7087] = 0
      "00000" when "001101110110000", -- t[7088] = 0
      "00000" when "001101110110001", -- t[7089] = 0
      "00000" when "001101110110010", -- t[7090] = 0
      "00000" when "001101110110011", -- t[7091] = 0
      "00000" when "001101110110100", -- t[7092] = 0
      "00000" when "001101110110101", -- t[7093] = 0
      "00000" when "001101110110110", -- t[7094] = 0
      "00000" when "001101110110111", -- t[7095] = 0
      "00000" when "001101110111000", -- t[7096] = 0
      "00000" when "001101110111001", -- t[7097] = 0
      "00000" when "001101110111010", -- t[7098] = 0
      "00000" when "001101110111011", -- t[7099] = 0
      "00000" when "001101110111100", -- t[7100] = 0
      "00000" when "001101110111101", -- t[7101] = 0
      "00000" when "001101110111110", -- t[7102] = 0
      "00000" when "001101110111111", -- t[7103] = 0
      "00000" when "001101111000000", -- t[7104] = 0
      "00000" when "001101111000001", -- t[7105] = 0
      "00000" when "001101111000010", -- t[7106] = 0
      "00000" when "001101111000011", -- t[7107] = 0
      "00000" when "001101111000100", -- t[7108] = 0
      "00001" when "001101111000101", -- t[7109] = 1
      "00001" when "001101111000110", -- t[7110] = 1
      "00001" when "001101111000111", -- t[7111] = 1
      "00001" when "001101111001000", -- t[7112] = 1
      "00001" when "001101111001001", -- t[7113] = 1
      "00001" when "001101111001010", -- t[7114] = 1
      "00001" when "001101111001011", -- t[7115] = 1
      "00001" when "001101111001100", -- t[7116] = 1
      "00001" when "001101111001101", -- t[7117] = 1
      "00001" when "001101111001110", -- t[7118] = 1
      "00001" when "001101111001111", -- t[7119] = 1
      "00001" when "001101111010000", -- t[7120] = 1
      "00001" when "001101111010001", -- t[7121] = 1
      "00001" when "001101111010010", -- t[7122] = 1
      "00001" when "001101111010011", -- t[7123] = 1
      "00001" when "001101111010100", -- t[7124] = 1
      "00001" when "001101111010101", -- t[7125] = 1
      "00001" when "001101111010110", -- t[7126] = 1
      "00001" when "001101111010111", -- t[7127] = 1
      "00001" when "001101111011000", -- t[7128] = 1
      "00001" when "001101111011001", -- t[7129] = 1
      "00001" when "001101111011010", -- t[7130] = 1
      "00001" when "001101111011011", -- t[7131] = 1
      "00001" when "001101111011100", -- t[7132] = 1
      "00001" when "001101111011101", -- t[7133] = 1
      "00001" when "001101111011110", -- t[7134] = 1
      "00001" when "001101111011111", -- t[7135] = 1
      "00001" when "001101111100000", -- t[7136] = 1
      "00001" when "001101111100001", -- t[7137] = 1
      "00001" when "001101111100010", -- t[7138] = 1
      "00001" when "001101111100011", -- t[7139] = 1
      "00001" when "001101111100100", -- t[7140] = 1
      "00001" when "001101111100101", -- t[7141] = 1
      "00001" when "001101111100110", -- t[7142] = 1
      "00001" when "001101111100111", -- t[7143] = 1
      "00001" when "001101111101000", -- t[7144] = 1
      "00001" when "001101111101001", -- t[7145] = 1
      "00001" when "001101111101010", -- t[7146] = 1
      "00001" when "001101111101011", -- t[7147] = 1
      "00001" when "001101111101100", -- t[7148] = 1
      "00001" when "001101111101101", -- t[7149] = 1
      "00001" when "001101111101110", -- t[7150] = 1
      "00001" when "001101111101111", -- t[7151] = 1
      "00001" when "001101111110000", -- t[7152] = 1
      "00001" when "001101111110001", -- t[7153] = 1
      "00001" when "001101111110010", -- t[7154] = 1
      "00001" when "001101111110011", -- t[7155] = 1
      "00001" when "001101111110100", -- t[7156] = 1
      "00001" when "001101111110101", -- t[7157] = 1
      "00001" when "001101111110110", -- t[7158] = 1
      "00001" when "001101111110111", -- t[7159] = 1
      "00001" when "001101111111000", -- t[7160] = 1
      "00001" when "001101111111001", -- t[7161] = 1
      "00001" when "001101111111010", -- t[7162] = 1
      "00001" when "001101111111011", -- t[7163] = 1
      "00001" when "001101111111100", -- t[7164] = 1
      "00001" when "001101111111101", -- t[7165] = 1
      "00001" when "001101111111110", -- t[7166] = 1
      "00001" when "001101111111111", -- t[7167] = 1
      "00001" when "001110000000000", -- t[7168] = 1
      "00001" when "001110000000001", -- t[7169] = 1
      "00001" when "001110000000010", -- t[7170] = 1
      "00001" when "001110000000011", -- t[7171] = 1
      "00001" when "001110000000100", -- t[7172] = 1
      "00001" when "001110000000101", -- t[7173] = 1
      "00001" when "001110000000110", -- t[7174] = 1
      "00001" when "001110000000111", -- t[7175] = 1
      "00001" when "001110000001000", -- t[7176] = 1
      "00001" when "001110000001001", -- t[7177] = 1
      "00001" when "001110000001010", -- t[7178] = 1
      "00001" when "001110000001011", -- t[7179] = 1
      "00001" when "001110000001100", -- t[7180] = 1
      "00001" when "001110000001101", -- t[7181] = 1
      "00001" when "001110000001110", -- t[7182] = 1
      "00001" when "001110000001111", -- t[7183] = 1
      "00001" when "001110000010000", -- t[7184] = 1
      "00001" when "001110000010001", -- t[7185] = 1
      "00001" when "001110000010010", -- t[7186] = 1
      "00001" when "001110000010011", -- t[7187] = 1
      "00001" when "001110000010100", -- t[7188] = 1
      "00001" when "001110000010101", -- t[7189] = 1
      "00001" when "001110000010110", -- t[7190] = 1
      "00001" when "001110000010111", -- t[7191] = 1
      "00001" when "001110000011000", -- t[7192] = 1
      "00001" when "001110000011001", -- t[7193] = 1
      "00001" when "001110000011010", -- t[7194] = 1
      "00001" when "001110000011011", -- t[7195] = 1
      "00001" when "001110000011100", -- t[7196] = 1
      "00001" when "001110000011101", -- t[7197] = 1
      "00001" when "001110000011110", -- t[7198] = 1
      "00001" when "001110000011111", -- t[7199] = 1
      "00001" when "001110000100000", -- t[7200] = 1
      "00001" when "001110000100001", -- t[7201] = 1
      "00001" when "001110000100010", -- t[7202] = 1
      "00001" when "001110000100011", -- t[7203] = 1
      "00001" when "001110000100100", -- t[7204] = 1
      "00001" when "001110000100101", -- t[7205] = 1
      "00001" when "001110000100110", -- t[7206] = 1
      "00001" when "001110000100111", -- t[7207] = 1
      "00001" when "001110000101000", -- t[7208] = 1
      "00001" when "001110000101001", -- t[7209] = 1
      "00001" when "001110000101010", -- t[7210] = 1
      "00001" when "001110000101011", -- t[7211] = 1
      "00001" when "001110000101100", -- t[7212] = 1
      "00001" when "001110000101101", -- t[7213] = 1
      "00001" when "001110000101110", -- t[7214] = 1
      "00001" when "001110000101111", -- t[7215] = 1
      "00001" when "001110000110000", -- t[7216] = 1
      "00001" when "001110000110001", -- t[7217] = 1
      "00001" when "001110000110010", -- t[7218] = 1
      "00001" when "001110000110011", -- t[7219] = 1
      "00001" when "001110000110100", -- t[7220] = 1
      "00001" when "001110000110101", -- t[7221] = 1
      "00001" when "001110000110110", -- t[7222] = 1
      "00001" when "001110000110111", -- t[7223] = 1
      "00001" when "001110000111000", -- t[7224] = 1
      "00001" when "001110000111001", -- t[7225] = 1
      "00001" when "001110000111010", -- t[7226] = 1
      "00001" when "001110000111011", -- t[7227] = 1
      "00001" when "001110000111100", -- t[7228] = 1
      "00001" when "001110000111101", -- t[7229] = 1
      "00001" when "001110000111110", -- t[7230] = 1
      "00001" when "001110000111111", -- t[7231] = 1
      "00001" when "001110001000000", -- t[7232] = 1
      "00001" when "001110001000001", -- t[7233] = 1
      "00001" when "001110001000010", -- t[7234] = 1
      "00001" when "001110001000011", -- t[7235] = 1
      "00001" when "001110001000100", -- t[7236] = 1
      "00001" when "001110001000101", -- t[7237] = 1
      "00001" when "001110001000110", -- t[7238] = 1
      "00001" when "001110001000111", -- t[7239] = 1
      "00001" when "001110001001000", -- t[7240] = 1
      "00001" when "001110001001001", -- t[7241] = 1
      "00001" when "001110001001010", -- t[7242] = 1
      "00001" when "001110001001011", -- t[7243] = 1
      "00001" when "001110001001100", -- t[7244] = 1
      "00001" when "001110001001101", -- t[7245] = 1
      "00001" when "001110001001110", -- t[7246] = 1
      "00001" when "001110001001111", -- t[7247] = 1
      "00001" when "001110001010000", -- t[7248] = 1
      "00001" when "001110001010001", -- t[7249] = 1
      "00001" when "001110001010010", -- t[7250] = 1
      "00001" when "001110001010011", -- t[7251] = 1
      "00001" when "001110001010100", -- t[7252] = 1
      "00001" when "001110001010101", -- t[7253] = 1
      "00001" when "001110001010110", -- t[7254] = 1
      "00001" when "001110001010111", -- t[7255] = 1
      "00001" when "001110001011000", -- t[7256] = 1
      "00001" when "001110001011001", -- t[7257] = 1
      "00001" when "001110001011010", -- t[7258] = 1
      "00001" when "001110001011011", -- t[7259] = 1
      "00001" when "001110001011100", -- t[7260] = 1
      "00001" when "001110001011101", -- t[7261] = 1
      "00001" when "001110001011110", -- t[7262] = 1
      "00001" when "001110001011111", -- t[7263] = 1
      "00001" when "001110001100000", -- t[7264] = 1
      "00001" when "001110001100001", -- t[7265] = 1
      "00001" when "001110001100010", -- t[7266] = 1
      "00001" when "001110001100011", -- t[7267] = 1
      "00001" when "001110001100100", -- t[7268] = 1
      "00001" when "001110001100101", -- t[7269] = 1
      "00001" when "001110001100110", -- t[7270] = 1
      "00001" when "001110001100111", -- t[7271] = 1
      "00001" when "001110001101000", -- t[7272] = 1
      "00001" when "001110001101001", -- t[7273] = 1
      "00001" when "001110001101010", -- t[7274] = 1
      "00001" when "001110001101011", -- t[7275] = 1
      "00001" when "001110001101100", -- t[7276] = 1
      "00001" when "001110001101101", -- t[7277] = 1
      "00001" when "001110001101110", -- t[7278] = 1
      "00001" when "001110001101111", -- t[7279] = 1
      "00001" when "001110001110000", -- t[7280] = 1
      "00001" when "001110001110001", -- t[7281] = 1
      "00001" when "001110001110010", -- t[7282] = 1
      "00001" when "001110001110011", -- t[7283] = 1
      "00001" when "001110001110100", -- t[7284] = 1
      "00001" when "001110001110101", -- t[7285] = 1
      "00001" when "001110001110110", -- t[7286] = 1
      "00001" when "001110001110111", -- t[7287] = 1
      "00001" when "001110001111000", -- t[7288] = 1
      "00001" when "001110001111001", -- t[7289] = 1
      "00001" when "001110001111010", -- t[7290] = 1
      "00001" when "001110001111011", -- t[7291] = 1
      "00001" when "001110001111100", -- t[7292] = 1
      "00001" when "001110001111101", -- t[7293] = 1
      "00001" when "001110001111110", -- t[7294] = 1
      "00001" when "001110001111111", -- t[7295] = 1
      "00001" when "001110010000000", -- t[7296] = 1
      "00001" when "001110010000001", -- t[7297] = 1
      "00001" when "001110010000010", -- t[7298] = 1
      "00001" when "001110010000011", -- t[7299] = 1
      "00001" when "001110010000100", -- t[7300] = 1
      "00001" when "001110010000101", -- t[7301] = 1
      "00001" when "001110010000110", -- t[7302] = 1
      "00001" when "001110010000111", -- t[7303] = 1
      "00001" when "001110010001000", -- t[7304] = 1
      "00001" when "001110010001001", -- t[7305] = 1
      "00001" when "001110010001010", -- t[7306] = 1
      "00001" when "001110010001011", -- t[7307] = 1
      "00001" when "001110010001100", -- t[7308] = 1
      "00001" when "001110010001101", -- t[7309] = 1
      "00001" when "001110010001110", -- t[7310] = 1
      "00001" when "001110010001111", -- t[7311] = 1
      "00001" when "001110010010000", -- t[7312] = 1
      "00001" when "001110010010001", -- t[7313] = 1
      "00001" when "001110010010010", -- t[7314] = 1
      "00001" when "001110010010011", -- t[7315] = 1
      "00001" when "001110010010100", -- t[7316] = 1
      "00001" when "001110010010101", -- t[7317] = 1
      "00001" when "001110010010110", -- t[7318] = 1
      "00001" when "001110010010111", -- t[7319] = 1
      "00001" when "001110010011000", -- t[7320] = 1
      "00001" when "001110010011001", -- t[7321] = 1
      "00001" when "001110010011010", -- t[7322] = 1
      "00001" when "001110010011011", -- t[7323] = 1
      "00001" when "001110010011100", -- t[7324] = 1
      "00001" when "001110010011101", -- t[7325] = 1
      "00001" when "001110010011110", -- t[7326] = 1
      "00001" when "001110010011111", -- t[7327] = 1
      "00001" when "001110010100000", -- t[7328] = 1
      "00001" when "001110010100001", -- t[7329] = 1
      "00001" when "001110010100010", -- t[7330] = 1
      "00001" when "001110010100011", -- t[7331] = 1
      "00001" when "001110010100100", -- t[7332] = 1
      "00001" when "001110010100101", -- t[7333] = 1
      "00001" when "001110010100110", -- t[7334] = 1
      "00001" when "001110010100111", -- t[7335] = 1
      "00001" when "001110010101000", -- t[7336] = 1
      "00001" when "001110010101001", -- t[7337] = 1
      "00001" when "001110010101010", -- t[7338] = 1
      "00001" when "001110010101011", -- t[7339] = 1
      "00001" when "001110010101100", -- t[7340] = 1
      "00001" when "001110010101101", -- t[7341] = 1
      "00001" when "001110010101110", -- t[7342] = 1
      "00001" when "001110010101111", -- t[7343] = 1
      "00001" when "001110010110000", -- t[7344] = 1
      "00001" when "001110010110001", -- t[7345] = 1
      "00001" when "001110010110010", -- t[7346] = 1
      "00001" when "001110010110011", -- t[7347] = 1
      "00001" when "001110010110100", -- t[7348] = 1
      "00001" when "001110010110101", -- t[7349] = 1
      "00001" when "001110010110110", -- t[7350] = 1
      "00001" when "001110010110111", -- t[7351] = 1
      "00001" when "001110010111000", -- t[7352] = 1
      "00001" when "001110010111001", -- t[7353] = 1
      "00001" when "001110010111010", -- t[7354] = 1
      "00001" when "001110010111011", -- t[7355] = 1
      "00001" when "001110010111100", -- t[7356] = 1
      "00001" when "001110010111101", -- t[7357] = 1
      "00001" when "001110010111110", -- t[7358] = 1
      "00001" when "001110010111111", -- t[7359] = 1
      "00001" when "001110011000000", -- t[7360] = 1
      "00001" when "001110011000001", -- t[7361] = 1
      "00001" when "001110011000010", -- t[7362] = 1
      "00001" when "001110011000011", -- t[7363] = 1
      "00001" when "001110011000100", -- t[7364] = 1
      "00001" when "001110011000101", -- t[7365] = 1
      "00001" when "001110011000110", -- t[7366] = 1
      "00001" when "001110011000111", -- t[7367] = 1
      "00001" when "001110011001000", -- t[7368] = 1
      "00001" when "001110011001001", -- t[7369] = 1
      "00001" when "001110011001010", -- t[7370] = 1
      "00001" when "001110011001011", -- t[7371] = 1
      "00001" when "001110011001100", -- t[7372] = 1
      "00001" when "001110011001101", -- t[7373] = 1
      "00001" when "001110011001110", -- t[7374] = 1
      "00001" when "001110011001111", -- t[7375] = 1
      "00001" when "001110011010000", -- t[7376] = 1
      "00001" when "001110011010001", -- t[7377] = 1
      "00001" when "001110011010010", -- t[7378] = 1
      "00001" when "001110011010011", -- t[7379] = 1
      "00001" when "001110011010100", -- t[7380] = 1
      "00001" when "001110011010101", -- t[7381] = 1
      "00001" when "001110011010110", -- t[7382] = 1
      "00001" when "001110011010111", -- t[7383] = 1
      "00001" when "001110011011000", -- t[7384] = 1
      "00001" when "001110011011001", -- t[7385] = 1
      "00001" when "001110011011010", -- t[7386] = 1
      "00001" when "001110011011011", -- t[7387] = 1
      "00001" when "001110011011100", -- t[7388] = 1
      "00001" when "001110011011101", -- t[7389] = 1
      "00001" when "001110011011110", -- t[7390] = 1
      "00001" when "001110011011111", -- t[7391] = 1
      "00001" when "001110011100000", -- t[7392] = 1
      "00001" when "001110011100001", -- t[7393] = 1
      "00001" when "001110011100010", -- t[7394] = 1
      "00001" when "001110011100011", -- t[7395] = 1
      "00001" when "001110011100100", -- t[7396] = 1
      "00001" when "001110011100101", -- t[7397] = 1
      "00001" when "001110011100110", -- t[7398] = 1
      "00001" when "001110011100111", -- t[7399] = 1
      "00001" when "001110011101000", -- t[7400] = 1
      "00001" when "001110011101001", -- t[7401] = 1
      "00001" when "001110011101010", -- t[7402] = 1
      "00001" when "001110011101011", -- t[7403] = 1
      "00001" when "001110011101100", -- t[7404] = 1
      "00001" when "001110011101101", -- t[7405] = 1
      "00001" when "001110011101110", -- t[7406] = 1
      "00001" when "001110011101111", -- t[7407] = 1
      "00001" when "001110011110000", -- t[7408] = 1
      "00001" when "001110011110001", -- t[7409] = 1
      "00001" when "001110011110010", -- t[7410] = 1
      "00001" when "001110011110011", -- t[7411] = 1
      "00001" when "001110011110100", -- t[7412] = 1
      "00001" when "001110011110101", -- t[7413] = 1
      "00001" when "001110011110110", -- t[7414] = 1
      "00001" when "001110011110111", -- t[7415] = 1
      "00001" when "001110011111000", -- t[7416] = 1
      "00001" when "001110011111001", -- t[7417] = 1
      "00001" when "001110011111010", -- t[7418] = 1
      "00001" when "001110011111011", -- t[7419] = 1
      "00001" when "001110011111100", -- t[7420] = 1
      "00001" when "001110011111101", -- t[7421] = 1
      "00001" when "001110011111110", -- t[7422] = 1
      "00001" when "001110011111111", -- t[7423] = 1
      "00001" when "001110100000000", -- t[7424] = 1
      "00001" when "001110100000001", -- t[7425] = 1
      "00001" when "001110100000010", -- t[7426] = 1
      "00001" when "001110100000011", -- t[7427] = 1
      "00001" when "001110100000100", -- t[7428] = 1
      "00001" when "001110100000101", -- t[7429] = 1
      "00001" when "001110100000110", -- t[7430] = 1
      "00001" when "001110100000111", -- t[7431] = 1
      "00001" when "001110100001000", -- t[7432] = 1
      "00001" when "001110100001001", -- t[7433] = 1
      "00001" when "001110100001010", -- t[7434] = 1
      "00001" when "001110100001011", -- t[7435] = 1
      "00001" when "001110100001100", -- t[7436] = 1
      "00001" when "001110100001101", -- t[7437] = 1
      "00001" when "001110100001110", -- t[7438] = 1
      "00001" when "001110100001111", -- t[7439] = 1
      "00001" when "001110100010000", -- t[7440] = 1
      "00001" when "001110100010001", -- t[7441] = 1
      "00001" when "001110100010010", -- t[7442] = 1
      "00001" when "001110100010011", -- t[7443] = 1
      "00001" when "001110100010100", -- t[7444] = 1
      "00001" when "001110100010101", -- t[7445] = 1
      "00001" when "001110100010110", -- t[7446] = 1
      "00001" when "001110100010111", -- t[7447] = 1
      "00001" when "001110100011000", -- t[7448] = 1
      "00001" when "001110100011001", -- t[7449] = 1
      "00001" when "001110100011010", -- t[7450] = 1
      "00001" when "001110100011011", -- t[7451] = 1
      "00001" when "001110100011100", -- t[7452] = 1
      "00001" when "001110100011101", -- t[7453] = 1
      "00001" when "001110100011110", -- t[7454] = 1
      "00001" when "001110100011111", -- t[7455] = 1
      "00001" when "001110100100000", -- t[7456] = 1
      "00001" when "001110100100001", -- t[7457] = 1
      "00001" when "001110100100010", -- t[7458] = 1
      "00001" when "001110100100011", -- t[7459] = 1
      "00001" when "001110100100100", -- t[7460] = 1
      "00001" when "001110100100101", -- t[7461] = 1
      "00001" when "001110100100110", -- t[7462] = 1
      "00001" when "001110100100111", -- t[7463] = 1
      "00001" when "001110100101000", -- t[7464] = 1
      "00001" when "001110100101001", -- t[7465] = 1
      "00001" when "001110100101010", -- t[7466] = 1
      "00001" when "001110100101011", -- t[7467] = 1
      "00001" when "001110100101100", -- t[7468] = 1
      "00001" when "001110100101101", -- t[7469] = 1
      "00001" when "001110100101110", -- t[7470] = 1
      "00001" when "001110100101111", -- t[7471] = 1
      "00001" when "001110100110000", -- t[7472] = 1
      "00001" when "001110100110001", -- t[7473] = 1
      "00001" when "001110100110010", -- t[7474] = 1
      "00001" when "001110100110011", -- t[7475] = 1
      "00001" when "001110100110100", -- t[7476] = 1
      "00001" when "001110100110101", -- t[7477] = 1
      "00001" when "001110100110110", -- t[7478] = 1
      "00001" when "001110100110111", -- t[7479] = 1
      "00001" when "001110100111000", -- t[7480] = 1
      "00001" when "001110100111001", -- t[7481] = 1
      "00001" when "001110100111010", -- t[7482] = 1
      "00001" when "001110100111011", -- t[7483] = 1
      "00001" when "001110100111100", -- t[7484] = 1
      "00001" when "001110100111101", -- t[7485] = 1
      "00001" when "001110100111110", -- t[7486] = 1
      "00001" when "001110100111111", -- t[7487] = 1
      "00001" when "001110101000000", -- t[7488] = 1
      "00001" when "001110101000001", -- t[7489] = 1
      "00001" when "001110101000010", -- t[7490] = 1
      "00001" when "001110101000011", -- t[7491] = 1
      "00001" when "001110101000100", -- t[7492] = 1
      "00001" when "001110101000101", -- t[7493] = 1
      "00001" when "001110101000110", -- t[7494] = 1
      "00001" when "001110101000111", -- t[7495] = 1
      "00001" when "001110101001000", -- t[7496] = 1
      "00001" when "001110101001001", -- t[7497] = 1
      "00001" when "001110101001010", -- t[7498] = 1
      "00001" when "001110101001011", -- t[7499] = 1
      "00001" when "001110101001100", -- t[7500] = 1
      "00001" when "001110101001101", -- t[7501] = 1
      "00001" when "001110101001110", -- t[7502] = 1
      "00001" when "001110101001111", -- t[7503] = 1
      "00001" when "001110101010000", -- t[7504] = 1
      "00001" when "001110101010001", -- t[7505] = 1
      "00001" when "001110101010010", -- t[7506] = 1
      "00001" when "001110101010011", -- t[7507] = 1
      "00001" when "001110101010100", -- t[7508] = 1
      "00001" when "001110101010101", -- t[7509] = 1
      "00001" when "001110101010110", -- t[7510] = 1
      "00001" when "001110101010111", -- t[7511] = 1
      "00001" when "001110101011000", -- t[7512] = 1
      "00001" when "001110101011001", -- t[7513] = 1
      "00001" when "001110101011010", -- t[7514] = 1
      "00001" when "001110101011011", -- t[7515] = 1
      "00001" when "001110101011100", -- t[7516] = 1
      "00001" when "001110101011101", -- t[7517] = 1
      "00001" when "001110101011110", -- t[7518] = 1
      "00001" when "001110101011111", -- t[7519] = 1
      "00001" when "001110101100000", -- t[7520] = 1
      "00001" when "001110101100001", -- t[7521] = 1
      "00001" when "001110101100010", -- t[7522] = 1
      "00001" when "001110101100011", -- t[7523] = 1
      "00001" when "001110101100100", -- t[7524] = 1
      "00001" when "001110101100101", -- t[7525] = 1
      "00001" when "001110101100110", -- t[7526] = 1
      "00001" when "001110101100111", -- t[7527] = 1
      "00001" when "001110101101000", -- t[7528] = 1
      "00001" when "001110101101001", -- t[7529] = 1
      "00001" when "001110101101010", -- t[7530] = 1
      "00001" when "001110101101011", -- t[7531] = 1
      "00001" when "001110101101100", -- t[7532] = 1
      "00001" when "001110101101101", -- t[7533] = 1
      "00001" when "001110101101110", -- t[7534] = 1
      "00001" when "001110101101111", -- t[7535] = 1
      "00001" when "001110101110000", -- t[7536] = 1
      "00001" when "001110101110001", -- t[7537] = 1
      "00001" when "001110101110010", -- t[7538] = 1
      "00001" when "001110101110011", -- t[7539] = 1
      "00001" when "001110101110100", -- t[7540] = 1
      "00001" when "001110101110101", -- t[7541] = 1
      "00001" when "001110101110110", -- t[7542] = 1
      "00001" when "001110101110111", -- t[7543] = 1
      "00001" when "001110101111000", -- t[7544] = 1
      "00001" when "001110101111001", -- t[7545] = 1
      "00001" when "001110101111010", -- t[7546] = 1
      "00001" when "001110101111011", -- t[7547] = 1
      "00001" when "001110101111100", -- t[7548] = 1
      "00001" when "001110101111101", -- t[7549] = 1
      "00001" when "001110101111110", -- t[7550] = 1
      "00001" when "001110101111111", -- t[7551] = 1
      "00001" when "001110110000000", -- t[7552] = 1
      "00001" when "001110110000001", -- t[7553] = 1
      "00001" when "001110110000010", -- t[7554] = 1
      "00001" when "001110110000011", -- t[7555] = 1
      "00001" when "001110110000100", -- t[7556] = 1
      "00001" when "001110110000101", -- t[7557] = 1
      "00001" when "001110110000110", -- t[7558] = 1
      "00001" when "001110110000111", -- t[7559] = 1
      "00001" when "001110110001000", -- t[7560] = 1
      "00001" when "001110110001001", -- t[7561] = 1
      "00001" when "001110110001010", -- t[7562] = 1
      "00001" when "001110110001011", -- t[7563] = 1
      "00001" when "001110110001100", -- t[7564] = 1
      "00001" when "001110110001101", -- t[7565] = 1
      "00001" when "001110110001110", -- t[7566] = 1
      "00001" when "001110110001111", -- t[7567] = 1
      "00001" when "001110110010000", -- t[7568] = 1
      "00001" when "001110110010001", -- t[7569] = 1
      "00001" when "001110110010010", -- t[7570] = 1
      "00001" when "001110110010011", -- t[7571] = 1
      "00001" when "001110110010100", -- t[7572] = 1
      "00001" when "001110110010101", -- t[7573] = 1
      "00001" when "001110110010110", -- t[7574] = 1
      "00001" when "001110110010111", -- t[7575] = 1
      "00001" when "001110110011000", -- t[7576] = 1
      "00001" when "001110110011001", -- t[7577] = 1
      "00001" when "001110110011010", -- t[7578] = 1
      "00001" when "001110110011011", -- t[7579] = 1
      "00001" when "001110110011100", -- t[7580] = 1
      "00001" when "001110110011101", -- t[7581] = 1
      "00001" when "001110110011110", -- t[7582] = 1
      "00001" when "001110110011111", -- t[7583] = 1
      "00001" when "001110110100000", -- t[7584] = 1
      "00001" when "001110110100001", -- t[7585] = 1
      "00001" when "001110110100010", -- t[7586] = 1
      "00001" when "001110110100011", -- t[7587] = 1
      "00001" when "001110110100100", -- t[7588] = 1
      "00001" when "001110110100101", -- t[7589] = 1
      "00001" when "001110110100110", -- t[7590] = 1
      "00001" when "001110110100111", -- t[7591] = 1
      "00001" when "001110110101000", -- t[7592] = 1
      "00001" when "001110110101001", -- t[7593] = 1
      "00001" when "001110110101010", -- t[7594] = 1
      "00001" when "001110110101011", -- t[7595] = 1
      "00001" when "001110110101100", -- t[7596] = 1
      "00001" when "001110110101101", -- t[7597] = 1
      "00001" when "001110110101110", -- t[7598] = 1
      "00001" when "001110110101111", -- t[7599] = 1
      "00001" when "001110110110000", -- t[7600] = 1
      "00001" when "001110110110001", -- t[7601] = 1
      "00001" when "001110110110010", -- t[7602] = 1
      "00001" when "001110110110011", -- t[7603] = 1
      "00001" when "001110110110100", -- t[7604] = 1
      "00001" when "001110110110101", -- t[7605] = 1
      "00001" when "001110110110110", -- t[7606] = 1
      "00001" when "001110110110111", -- t[7607] = 1
      "00001" when "001110110111000", -- t[7608] = 1
      "00001" when "001110110111001", -- t[7609] = 1
      "00001" when "001110110111010", -- t[7610] = 1
      "00001" when "001110110111011", -- t[7611] = 1
      "00001" when "001110110111100", -- t[7612] = 1
      "00001" when "001110110111101", -- t[7613] = 1
      "00001" when "001110110111110", -- t[7614] = 1
      "00001" when "001110110111111", -- t[7615] = 1
      "00001" when "001110111000000", -- t[7616] = 1
      "00001" when "001110111000001", -- t[7617] = 1
      "00001" when "001110111000010", -- t[7618] = 1
      "00001" when "001110111000011", -- t[7619] = 1
      "00001" when "001110111000100", -- t[7620] = 1
      "00001" when "001110111000101", -- t[7621] = 1
      "00001" when "001110111000110", -- t[7622] = 1
      "00001" when "001110111000111", -- t[7623] = 1
      "00001" when "001110111001000", -- t[7624] = 1
      "00001" when "001110111001001", -- t[7625] = 1
      "00001" when "001110111001010", -- t[7626] = 1
      "00001" when "001110111001011", -- t[7627] = 1
      "00001" when "001110111001100", -- t[7628] = 1
      "00001" when "001110111001101", -- t[7629] = 1
      "00001" when "001110111001110", -- t[7630] = 1
      "00001" when "001110111001111", -- t[7631] = 1
      "00001" when "001110111010000", -- t[7632] = 1
      "00001" when "001110111010001", -- t[7633] = 1
      "00001" when "001110111010010", -- t[7634] = 1
      "00001" when "001110111010011", -- t[7635] = 1
      "00001" when "001110111010100", -- t[7636] = 1
      "00001" when "001110111010101", -- t[7637] = 1
      "00001" when "001110111010110", -- t[7638] = 1
      "00001" when "001110111010111", -- t[7639] = 1
      "00001" when "001110111011000", -- t[7640] = 1
      "00001" when "001110111011001", -- t[7641] = 1
      "00001" when "001110111011010", -- t[7642] = 1
      "00001" when "001110111011011", -- t[7643] = 1
      "00001" when "001110111011100", -- t[7644] = 1
      "00001" when "001110111011101", -- t[7645] = 1
      "00001" when "001110111011110", -- t[7646] = 1
      "00001" when "001110111011111", -- t[7647] = 1
      "00001" when "001110111100000", -- t[7648] = 1
      "00001" when "001110111100001", -- t[7649] = 1
      "00001" when "001110111100010", -- t[7650] = 1
      "00001" when "001110111100011", -- t[7651] = 1
      "00001" when "001110111100100", -- t[7652] = 1
      "00001" when "001110111100101", -- t[7653] = 1
      "00001" when "001110111100110", -- t[7654] = 1
      "00001" when "001110111100111", -- t[7655] = 1
      "00001" when "001110111101000", -- t[7656] = 1
      "00001" when "001110111101001", -- t[7657] = 1
      "00001" when "001110111101010", -- t[7658] = 1
      "00001" when "001110111101011", -- t[7659] = 1
      "00001" when "001110111101100", -- t[7660] = 1
      "00001" when "001110111101101", -- t[7661] = 1
      "00001" when "001110111101110", -- t[7662] = 1
      "00001" when "001110111101111", -- t[7663] = 1
      "00001" when "001110111110000", -- t[7664] = 1
      "00001" when "001110111110001", -- t[7665] = 1
      "00001" when "001110111110010", -- t[7666] = 1
      "00001" when "001110111110011", -- t[7667] = 1
      "00001" when "001110111110100", -- t[7668] = 1
      "00001" when "001110111110101", -- t[7669] = 1
      "00001" when "001110111110110", -- t[7670] = 1
      "00001" when "001110111110111", -- t[7671] = 1
      "00001" when "001110111111000", -- t[7672] = 1
      "00001" when "001110111111001", -- t[7673] = 1
      "00001" when "001110111111010", -- t[7674] = 1
      "00001" when "001110111111011", -- t[7675] = 1
      "00001" when "001110111111100", -- t[7676] = 1
      "00001" when "001110111111101", -- t[7677] = 1
      "00001" when "001110111111110", -- t[7678] = 1
      "00001" when "001110111111111", -- t[7679] = 1
      "00001" when "001111000000000", -- t[7680] = 1
      "00001" when "001111000000001", -- t[7681] = 1
      "00001" when "001111000000010", -- t[7682] = 1
      "00001" when "001111000000011", -- t[7683] = 1
      "00001" when "001111000000100", -- t[7684] = 1
      "00001" when "001111000000101", -- t[7685] = 1
      "00001" when "001111000000110", -- t[7686] = 1
      "00001" when "001111000000111", -- t[7687] = 1
      "00001" when "001111000001000", -- t[7688] = 1
      "00001" when "001111000001001", -- t[7689] = 1
      "00001" when "001111000001010", -- t[7690] = 1
      "00001" when "001111000001011", -- t[7691] = 1
      "00001" when "001111000001100", -- t[7692] = 1
      "00001" when "001111000001101", -- t[7693] = 1
      "00001" when "001111000001110", -- t[7694] = 1
      "00001" when "001111000001111", -- t[7695] = 1
      "00001" when "001111000010000", -- t[7696] = 1
      "00001" when "001111000010001", -- t[7697] = 1
      "00001" when "001111000010010", -- t[7698] = 1
      "00001" when "001111000010011", -- t[7699] = 1
      "00001" when "001111000010100", -- t[7700] = 1
      "00001" when "001111000010101", -- t[7701] = 1
      "00001" when "001111000010110", -- t[7702] = 1
      "00001" when "001111000010111", -- t[7703] = 1
      "00001" when "001111000011000", -- t[7704] = 1
      "00001" when "001111000011001", -- t[7705] = 1
      "00001" when "001111000011010", -- t[7706] = 1
      "00001" when "001111000011011", -- t[7707] = 1
      "00001" when "001111000011100", -- t[7708] = 1
      "00001" when "001111000011101", -- t[7709] = 1
      "00001" when "001111000011110", -- t[7710] = 1
      "00001" when "001111000011111", -- t[7711] = 1
      "00001" when "001111000100000", -- t[7712] = 1
      "00001" when "001111000100001", -- t[7713] = 1
      "00001" when "001111000100010", -- t[7714] = 1
      "00001" when "001111000100011", -- t[7715] = 1
      "00001" when "001111000100100", -- t[7716] = 1
      "00001" when "001111000100101", -- t[7717] = 1
      "00001" when "001111000100110", -- t[7718] = 1
      "00001" when "001111000100111", -- t[7719] = 1
      "00001" when "001111000101000", -- t[7720] = 1
      "00001" when "001111000101001", -- t[7721] = 1
      "00001" when "001111000101010", -- t[7722] = 1
      "00001" when "001111000101011", -- t[7723] = 1
      "00001" when "001111000101100", -- t[7724] = 1
      "00001" when "001111000101101", -- t[7725] = 1
      "00001" when "001111000101110", -- t[7726] = 1
      "00001" when "001111000101111", -- t[7727] = 1
      "00001" when "001111000110000", -- t[7728] = 1
      "00001" when "001111000110001", -- t[7729] = 1
      "00001" when "001111000110010", -- t[7730] = 1
      "00001" when "001111000110011", -- t[7731] = 1
      "00001" when "001111000110100", -- t[7732] = 1
      "00001" when "001111000110101", -- t[7733] = 1
      "00001" when "001111000110110", -- t[7734] = 1
      "00001" when "001111000110111", -- t[7735] = 1
      "00001" when "001111000111000", -- t[7736] = 1
      "00001" when "001111000111001", -- t[7737] = 1
      "00001" when "001111000111010", -- t[7738] = 1
      "00001" when "001111000111011", -- t[7739] = 1
      "00001" when "001111000111100", -- t[7740] = 1
      "00001" when "001111000111101", -- t[7741] = 1
      "00001" when "001111000111110", -- t[7742] = 1
      "00001" when "001111000111111", -- t[7743] = 1
      "00001" when "001111001000000", -- t[7744] = 1
      "00001" when "001111001000001", -- t[7745] = 1
      "00001" when "001111001000010", -- t[7746] = 1
      "00001" when "001111001000011", -- t[7747] = 1
      "00001" when "001111001000100", -- t[7748] = 1
      "00001" when "001111001000101", -- t[7749] = 1
      "00001" when "001111001000110", -- t[7750] = 1
      "00001" when "001111001000111", -- t[7751] = 1
      "00001" when "001111001001000", -- t[7752] = 1
      "00001" when "001111001001001", -- t[7753] = 1
      "00001" when "001111001001010", -- t[7754] = 1
      "00001" when "001111001001011", -- t[7755] = 1
      "00001" when "001111001001100", -- t[7756] = 1
      "00001" when "001111001001101", -- t[7757] = 1
      "00001" when "001111001001110", -- t[7758] = 1
      "00001" when "001111001001111", -- t[7759] = 1
      "00001" when "001111001010000", -- t[7760] = 1
      "00001" when "001111001010001", -- t[7761] = 1
      "00001" when "001111001010010", -- t[7762] = 1
      "00001" when "001111001010011", -- t[7763] = 1
      "00001" when "001111001010100", -- t[7764] = 1
      "00001" when "001111001010101", -- t[7765] = 1
      "00001" when "001111001010110", -- t[7766] = 1
      "00001" when "001111001010111", -- t[7767] = 1
      "00001" when "001111001011000", -- t[7768] = 1
      "00001" when "001111001011001", -- t[7769] = 1
      "00001" when "001111001011010", -- t[7770] = 1
      "00001" when "001111001011011", -- t[7771] = 1
      "00001" when "001111001011100", -- t[7772] = 1
      "00001" when "001111001011101", -- t[7773] = 1
      "00001" when "001111001011110", -- t[7774] = 1
      "00001" when "001111001011111", -- t[7775] = 1
      "00001" when "001111001100000", -- t[7776] = 1
      "00001" when "001111001100001", -- t[7777] = 1
      "00001" when "001111001100010", -- t[7778] = 1
      "00001" when "001111001100011", -- t[7779] = 1
      "00001" when "001111001100100", -- t[7780] = 1
      "00001" when "001111001100101", -- t[7781] = 1
      "00001" when "001111001100110", -- t[7782] = 1
      "00001" when "001111001100111", -- t[7783] = 1
      "00001" when "001111001101000", -- t[7784] = 1
      "00001" when "001111001101001", -- t[7785] = 1
      "00001" when "001111001101010", -- t[7786] = 1
      "00001" when "001111001101011", -- t[7787] = 1
      "00001" when "001111001101100", -- t[7788] = 1
      "00001" when "001111001101101", -- t[7789] = 1
      "00001" when "001111001101110", -- t[7790] = 1
      "00001" when "001111001101111", -- t[7791] = 1
      "00001" when "001111001110000", -- t[7792] = 1
      "00001" when "001111001110001", -- t[7793] = 1
      "00001" when "001111001110010", -- t[7794] = 1
      "00001" when "001111001110011", -- t[7795] = 1
      "00001" when "001111001110100", -- t[7796] = 1
      "00001" when "001111001110101", -- t[7797] = 1
      "00001" when "001111001110110", -- t[7798] = 1
      "00001" when "001111001110111", -- t[7799] = 1
      "00001" when "001111001111000", -- t[7800] = 1
      "00001" when "001111001111001", -- t[7801] = 1
      "00001" when "001111001111010", -- t[7802] = 1
      "00001" when "001111001111011", -- t[7803] = 1
      "00001" when "001111001111100", -- t[7804] = 1
      "00001" when "001111001111101", -- t[7805] = 1
      "00001" when "001111001111110", -- t[7806] = 1
      "00001" when "001111001111111", -- t[7807] = 1
      "00001" when "001111010000000", -- t[7808] = 1
      "00001" when "001111010000001", -- t[7809] = 1
      "00001" when "001111010000010", -- t[7810] = 1
      "00001" when "001111010000011", -- t[7811] = 1
      "00001" when "001111010000100", -- t[7812] = 1
      "00001" when "001111010000101", -- t[7813] = 1
      "00001" when "001111010000110", -- t[7814] = 1
      "00001" when "001111010000111", -- t[7815] = 1
      "00001" when "001111010001000", -- t[7816] = 1
      "00001" when "001111010001001", -- t[7817] = 1
      "00001" when "001111010001010", -- t[7818] = 1
      "00001" when "001111010001011", -- t[7819] = 1
      "00001" when "001111010001100", -- t[7820] = 1
      "00001" when "001111010001101", -- t[7821] = 1
      "00001" when "001111010001110", -- t[7822] = 1
      "00001" when "001111010001111", -- t[7823] = 1
      "00001" when "001111010010000", -- t[7824] = 1
      "00001" when "001111010010001", -- t[7825] = 1
      "00001" when "001111010010010", -- t[7826] = 1
      "00001" when "001111010010011", -- t[7827] = 1
      "00001" when "001111010010100", -- t[7828] = 1
      "00001" when "001111010010101", -- t[7829] = 1
      "00001" when "001111010010110", -- t[7830] = 1
      "00001" when "001111010010111", -- t[7831] = 1
      "00001" when "001111010011000", -- t[7832] = 1
      "00001" when "001111010011001", -- t[7833] = 1
      "00001" when "001111010011010", -- t[7834] = 1
      "00001" when "001111010011011", -- t[7835] = 1
      "00001" when "001111010011100", -- t[7836] = 1
      "00001" when "001111010011101", -- t[7837] = 1
      "00001" when "001111010011110", -- t[7838] = 1
      "00001" when "001111010011111", -- t[7839] = 1
      "00001" when "001111010100000", -- t[7840] = 1
      "00001" when "001111010100001", -- t[7841] = 1
      "00001" when "001111010100010", -- t[7842] = 1
      "00001" when "001111010100011", -- t[7843] = 1
      "00001" when "001111010100100", -- t[7844] = 1
      "00001" when "001111010100101", -- t[7845] = 1
      "00001" when "001111010100110", -- t[7846] = 1
      "00001" when "001111010100111", -- t[7847] = 1
      "00001" when "001111010101000", -- t[7848] = 1
      "00001" when "001111010101001", -- t[7849] = 1
      "00001" when "001111010101010", -- t[7850] = 1
      "00001" when "001111010101011", -- t[7851] = 1
      "00001" when "001111010101100", -- t[7852] = 1
      "00001" when "001111010101101", -- t[7853] = 1
      "00001" when "001111010101110", -- t[7854] = 1
      "00001" when "001111010101111", -- t[7855] = 1
      "00001" when "001111010110000", -- t[7856] = 1
      "00001" when "001111010110001", -- t[7857] = 1
      "00001" when "001111010110010", -- t[7858] = 1
      "00001" when "001111010110011", -- t[7859] = 1
      "00001" when "001111010110100", -- t[7860] = 1
      "00001" when "001111010110101", -- t[7861] = 1
      "00001" when "001111010110110", -- t[7862] = 1
      "00001" when "001111010110111", -- t[7863] = 1
      "00001" when "001111010111000", -- t[7864] = 1
      "00001" when "001111010111001", -- t[7865] = 1
      "00001" when "001111010111010", -- t[7866] = 1
      "00001" when "001111010111011", -- t[7867] = 1
      "00001" when "001111010111100", -- t[7868] = 1
      "00001" when "001111010111101", -- t[7869] = 1
      "00001" when "001111010111110", -- t[7870] = 1
      "00001" when "001111010111111", -- t[7871] = 1
      "00001" when "001111011000000", -- t[7872] = 1
      "00001" when "001111011000001", -- t[7873] = 1
      "00001" when "001111011000010", -- t[7874] = 1
      "00001" when "001111011000011", -- t[7875] = 1
      "00001" when "001111011000100", -- t[7876] = 1
      "00001" when "001111011000101", -- t[7877] = 1
      "00001" when "001111011000110", -- t[7878] = 1
      "00001" when "001111011000111", -- t[7879] = 1
      "00001" when "001111011001000", -- t[7880] = 1
      "00001" when "001111011001001", -- t[7881] = 1
      "00001" when "001111011001010", -- t[7882] = 1
      "00001" when "001111011001011", -- t[7883] = 1
      "00001" when "001111011001100", -- t[7884] = 1
      "00001" when "001111011001101", -- t[7885] = 1
      "00001" when "001111011001110", -- t[7886] = 1
      "00001" when "001111011001111", -- t[7887] = 1
      "00001" when "001111011010000", -- t[7888] = 1
      "00001" when "001111011010001", -- t[7889] = 1
      "00001" when "001111011010010", -- t[7890] = 1
      "00001" when "001111011010011", -- t[7891] = 1
      "00001" when "001111011010100", -- t[7892] = 1
      "00001" when "001111011010101", -- t[7893] = 1
      "00001" when "001111011010110", -- t[7894] = 1
      "00001" when "001111011010111", -- t[7895] = 1
      "00001" when "001111011011000", -- t[7896] = 1
      "00001" when "001111011011001", -- t[7897] = 1
      "00001" when "001111011011010", -- t[7898] = 1
      "00001" when "001111011011011", -- t[7899] = 1
      "00001" when "001111011011100", -- t[7900] = 1
      "00001" when "001111011011101", -- t[7901] = 1
      "00001" when "001111011011110", -- t[7902] = 1
      "00001" when "001111011011111", -- t[7903] = 1
      "00001" when "001111011100000", -- t[7904] = 1
      "00001" when "001111011100001", -- t[7905] = 1
      "00001" when "001111011100010", -- t[7906] = 1
      "00001" when "001111011100011", -- t[7907] = 1
      "00001" when "001111011100100", -- t[7908] = 1
      "00001" when "001111011100101", -- t[7909] = 1
      "00001" when "001111011100110", -- t[7910] = 1
      "00001" when "001111011100111", -- t[7911] = 1
      "00001" when "001111011101000", -- t[7912] = 1
      "00001" when "001111011101001", -- t[7913] = 1
      "00001" when "001111011101010", -- t[7914] = 1
      "00001" when "001111011101011", -- t[7915] = 1
      "00001" when "001111011101100", -- t[7916] = 1
      "00001" when "001111011101101", -- t[7917] = 1
      "00001" when "001111011101110", -- t[7918] = 1
      "00001" when "001111011101111", -- t[7919] = 1
      "00001" when "001111011110000", -- t[7920] = 1
      "00001" when "001111011110001", -- t[7921] = 1
      "00001" when "001111011110010", -- t[7922] = 1
      "00001" when "001111011110011", -- t[7923] = 1
      "00001" when "001111011110100", -- t[7924] = 1
      "00001" when "001111011110101", -- t[7925] = 1
      "00001" when "001111011110110", -- t[7926] = 1
      "00001" when "001111011110111", -- t[7927] = 1
      "00001" when "001111011111000", -- t[7928] = 1
      "00001" when "001111011111001", -- t[7929] = 1
      "00001" when "001111011111010", -- t[7930] = 1
      "00001" when "001111011111011", -- t[7931] = 1
      "00001" when "001111011111100", -- t[7932] = 1
      "00001" when "001111011111101", -- t[7933] = 1
      "00001" when "001111011111110", -- t[7934] = 1
      "00001" when "001111011111111", -- t[7935] = 1
      "00001" when "001111100000000", -- t[7936] = 1
      "00001" when "001111100000001", -- t[7937] = 1
      "00001" when "001111100000010", -- t[7938] = 1
      "00001" when "001111100000011", -- t[7939] = 1
      "00001" when "001111100000100", -- t[7940] = 1
      "00001" when "001111100000101", -- t[7941] = 1
      "00001" when "001111100000110", -- t[7942] = 1
      "00001" when "001111100000111", -- t[7943] = 1
      "00001" when "001111100001000", -- t[7944] = 1
      "00001" when "001111100001001", -- t[7945] = 1
      "00001" when "001111100001010", -- t[7946] = 1
      "00001" when "001111100001011", -- t[7947] = 1
      "00001" when "001111100001100", -- t[7948] = 1
      "00001" when "001111100001101", -- t[7949] = 1
      "00001" when "001111100001110", -- t[7950] = 1
      "00001" when "001111100001111", -- t[7951] = 1
      "00001" when "001111100010000", -- t[7952] = 1
      "00001" when "001111100010001", -- t[7953] = 1
      "00001" when "001111100010010", -- t[7954] = 1
      "00001" when "001111100010011", -- t[7955] = 1
      "00001" when "001111100010100", -- t[7956] = 1
      "00001" when "001111100010101", -- t[7957] = 1
      "00001" when "001111100010110", -- t[7958] = 1
      "00001" when "001111100010111", -- t[7959] = 1
      "00001" when "001111100011000", -- t[7960] = 1
      "00001" when "001111100011001", -- t[7961] = 1
      "00001" when "001111100011010", -- t[7962] = 1
      "00001" when "001111100011011", -- t[7963] = 1
      "00001" when "001111100011100", -- t[7964] = 1
      "00001" when "001111100011101", -- t[7965] = 1
      "00001" when "001111100011110", -- t[7966] = 1
      "00001" when "001111100011111", -- t[7967] = 1
      "00001" when "001111100100000", -- t[7968] = 1
      "00001" when "001111100100001", -- t[7969] = 1
      "00001" when "001111100100010", -- t[7970] = 1
      "00001" when "001111100100011", -- t[7971] = 1
      "00001" when "001111100100100", -- t[7972] = 1
      "00001" when "001111100100101", -- t[7973] = 1
      "00001" when "001111100100110", -- t[7974] = 1
      "00001" when "001111100100111", -- t[7975] = 1
      "00001" when "001111100101000", -- t[7976] = 1
      "00001" when "001111100101001", -- t[7977] = 1
      "00001" when "001111100101010", -- t[7978] = 1
      "00001" when "001111100101011", -- t[7979] = 1
      "00001" when "001111100101100", -- t[7980] = 1
      "00001" when "001111100101101", -- t[7981] = 1
      "00001" when "001111100101110", -- t[7982] = 1
      "00001" when "001111100101111", -- t[7983] = 1
      "00001" when "001111100110000", -- t[7984] = 1
      "00001" when "001111100110001", -- t[7985] = 1
      "00001" when "001111100110010", -- t[7986] = 1
      "00001" when "001111100110011", -- t[7987] = 1
      "00001" when "001111100110100", -- t[7988] = 1
      "00001" when "001111100110101", -- t[7989] = 1
      "00001" when "001111100110110", -- t[7990] = 1
      "00001" when "001111100110111", -- t[7991] = 1
      "00001" when "001111100111000", -- t[7992] = 1
      "00001" when "001111100111001", -- t[7993] = 1
      "00001" when "001111100111010", -- t[7994] = 1
      "00001" when "001111100111011", -- t[7995] = 1
      "00001" when "001111100111100", -- t[7996] = 1
      "00001" when "001111100111101", -- t[7997] = 1
      "00001" when "001111100111110", -- t[7998] = 1
      "00001" when "001111100111111", -- t[7999] = 1
      "00001" when "001111101000000", -- t[8000] = 1
      "00001" when "001111101000001", -- t[8001] = 1
      "00001" when "001111101000010", -- t[8002] = 1
      "00001" when "001111101000011", -- t[8003] = 1
      "00001" when "001111101000100", -- t[8004] = 1
      "00001" when "001111101000101", -- t[8005] = 1
      "00001" when "001111101000110", -- t[8006] = 1
      "00001" when "001111101000111", -- t[8007] = 1
      "00001" when "001111101001000", -- t[8008] = 1
      "00001" when "001111101001001", -- t[8009] = 1
      "00001" when "001111101001010", -- t[8010] = 1
      "00001" when "001111101001011", -- t[8011] = 1
      "00001" when "001111101001100", -- t[8012] = 1
      "00001" when "001111101001101", -- t[8013] = 1
      "00001" when "001111101001110", -- t[8014] = 1
      "00001" when "001111101001111", -- t[8015] = 1
      "00001" when "001111101010000", -- t[8016] = 1
      "00001" when "001111101010001", -- t[8017] = 1
      "00001" when "001111101010010", -- t[8018] = 1
      "00001" when "001111101010011", -- t[8019] = 1
      "00001" when "001111101010100", -- t[8020] = 1
      "00001" when "001111101010101", -- t[8021] = 1
      "00001" when "001111101010110", -- t[8022] = 1
      "00001" when "001111101010111", -- t[8023] = 1
      "00001" when "001111101011000", -- t[8024] = 1
      "00001" when "001111101011001", -- t[8025] = 1
      "00001" when "001111101011010", -- t[8026] = 1
      "00001" when "001111101011011", -- t[8027] = 1
      "00001" when "001111101011100", -- t[8028] = 1
      "00001" when "001111101011101", -- t[8029] = 1
      "00001" when "001111101011110", -- t[8030] = 1
      "00001" when "001111101011111", -- t[8031] = 1
      "00001" when "001111101100000", -- t[8032] = 1
      "00001" when "001111101100001", -- t[8033] = 1
      "00001" when "001111101100010", -- t[8034] = 1
      "00001" when "001111101100011", -- t[8035] = 1
      "00001" when "001111101100100", -- t[8036] = 1
      "00001" when "001111101100101", -- t[8037] = 1
      "00001" when "001111101100110", -- t[8038] = 1
      "00001" when "001111101100111", -- t[8039] = 1
      "00001" when "001111101101000", -- t[8040] = 1
      "00001" when "001111101101001", -- t[8041] = 1
      "00001" when "001111101101010", -- t[8042] = 1
      "00001" when "001111101101011", -- t[8043] = 1
      "00001" when "001111101101100", -- t[8044] = 1
      "00001" when "001111101101101", -- t[8045] = 1
      "00001" when "001111101101110", -- t[8046] = 1
      "00001" when "001111101101111", -- t[8047] = 1
      "00001" when "001111101110000", -- t[8048] = 1
      "00001" when "001111101110001", -- t[8049] = 1
      "00001" when "001111101110010", -- t[8050] = 1
      "00001" when "001111101110011", -- t[8051] = 1
      "00001" when "001111101110100", -- t[8052] = 1
      "00001" when "001111101110101", -- t[8053] = 1
      "00001" when "001111101110110", -- t[8054] = 1
      "00001" when "001111101110111", -- t[8055] = 1
      "00001" when "001111101111000", -- t[8056] = 1
      "00001" when "001111101111001", -- t[8057] = 1
      "00001" when "001111101111010", -- t[8058] = 1
      "00001" when "001111101111011", -- t[8059] = 1
      "00001" when "001111101111100", -- t[8060] = 1
      "00001" when "001111101111101", -- t[8061] = 1
      "00001" when "001111101111110", -- t[8062] = 1
      "00001" when "001111101111111", -- t[8063] = 1
      "00001" when "001111110000000", -- t[8064] = 1
      "00001" when "001111110000001", -- t[8065] = 1
      "00001" when "001111110000010", -- t[8066] = 1
      "00001" when "001111110000011", -- t[8067] = 1
      "00001" when "001111110000100", -- t[8068] = 1
      "00001" when "001111110000101", -- t[8069] = 1
      "00001" when "001111110000110", -- t[8070] = 1
      "00001" when "001111110000111", -- t[8071] = 1
      "00001" when "001111110001000", -- t[8072] = 1
      "00001" when "001111110001001", -- t[8073] = 1
      "00001" when "001111110001010", -- t[8074] = 1
      "00001" when "001111110001011", -- t[8075] = 1
      "00001" when "001111110001100", -- t[8076] = 1
      "00001" when "001111110001101", -- t[8077] = 1
      "00001" when "001111110001110", -- t[8078] = 1
      "00001" when "001111110001111", -- t[8079] = 1
      "00001" when "001111110010000", -- t[8080] = 1
      "00001" when "001111110010001", -- t[8081] = 1
      "00001" when "001111110010010", -- t[8082] = 1
      "00001" when "001111110010011", -- t[8083] = 1
      "00001" when "001111110010100", -- t[8084] = 1
      "00001" when "001111110010101", -- t[8085] = 1
      "00001" when "001111110010110", -- t[8086] = 1
      "00001" when "001111110010111", -- t[8087] = 1
      "00001" when "001111110011000", -- t[8088] = 1
      "00001" when "001111110011001", -- t[8089] = 1
      "00001" when "001111110011010", -- t[8090] = 1
      "00001" when "001111110011011", -- t[8091] = 1
      "00001" when "001111110011100", -- t[8092] = 1
      "00001" when "001111110011101", -- t[8093] = 1
      "00001" when "001111110011110", -- t[8094] = 1
      "00001" when "001111110011111", -- t[8095] = 1
      "00001" when "001111110100000", -- t[8096] = 1
      "00001" when "001111110100001", -- t[8097] = 1
      "00001" when "001111110100010", -- t[8098] = 1
      "00001" when "001111110100011", -- t[8099] = 1
      "00001" when "001111110100100", -- t[8100] = 1
      "00001" when "001111110100101", -- t[8101] = 1
      "00001" when "001111110100110", -- t[8102] = 1
      "00001" when "001111110100111", -- t[8103] = 1
      "00001" when "001111110101000", -- t[8104] = 1
      "00001" when "001111110101001", -- t[8105] = 1
      "00001" when "001111110101010", -- t[8106] = 1
      "00001" when "001111110101011", -- t[8107] = 1
      "00001" when "001111110101100", -- t[8108] = 1
      "00001" when "001111110101101", -- t[8109] = 1
      "00001" when "001111110101110", -- t[8110] = 1
      "00001" when "001111110101111", -- t[8111] = 1
      "00001" when "001111110110000", -- t[8112] = 1
      "00001" when "001111110110001", -- t[8113] = 1
      "00001" when "001111110110010", -- t[8114] = 1
      "00001" when "001111110110011", -- t[8115] = 1
      "00001" when "001111110110100", -- t[8116] = 1
      "00001" when "001111110110101", -- t[8117] = 1
      "00001" when "001111110110110", -- t[8118] = 1
      "00001" when "001111110110111", -- t[8119] = 1
      "00001" when "001111110111000", -- t[8120] = 1
      "00001" when "001111110111001", -- t[8121] = 1
      "00001" when "001111110111010", -- t[8122] = 1
      "00001" when "001111110111011", -- t[8123] = 1
      "00001" when "001111110111100", -- t[8124] = 1
      "00001" when "001111110111101", -- t[8125] = 1
      "00001" when "001111110111110", -- t[8126] = 1
      "00001" when "001111110111111", -- t[8127] = 1
      "00001" when "001111111000000", -- t[8128] = 1
      "00001" when "001111111000001", -- t[8129] = 1
      "00001" when "001111111000010", -- t[8130] = 1
      "00001" when "001111111000011", -- t[8131] = 1
      "00001" when "001111111000100", -- t[8132] = 1
      "00001" when "001111111000101", -- t[8133] = 1
      "00001" when "001111111000110", -- t[8134] = 1
      "00001" when "001111111000111", -- t[8135] = 1
      "00001" when "001111111001000", -- t[8136] = 1
      "00001" when "001111111001001", -- t[8137] = 1
      "00001" when "001111111001010", -- t[8138] = 1
      "00001" when "001111111001011", -- t[8139] = 1
      "00001" when "001111111001100", -- t[8140] = 1
      "00001" when "001111111001101", -- t[8141] = 1
      "00001" when "001111111001110", -- t[8142] = 1
      "00001" when "001111111001111", -- t[8143] = 1
      "00001" when "001111111010000", -- t[8144] = 1
      "00001" when "001111111010001", -- t[8145] = 1
      "00001" when "001111111010010", -- t[8146] = 1
      "00001" when "001111111010011", -- t[8147] = 1
      "00001" when "001111111010100", -- t[8148] = 1
      "00001" when "001111111010101", -- t[8149] = 1
      "00001" when "001111111010110", -- t[8150] = 1
      "00001" when "001111111010111", -- t[8151] = 1
      "00001" when "001111111011000", -- t[8152] = 1
      "00001" when "001111111011001", -- t[8153] = 1
      "00001" when "001111111011010", -- t[8154] = 1
      "00001" when "001111111011011", -- t[8155] = 1
      "00001" when "001111111011100", -- t[8156] = 1
      "00001" when "001111111011101", -- t[8157] = 1
      "00001" when "001111111011110", -- t[8158] = 1
      "00001" when "001111111011111", -- t[8159] = 1
      "00001" when "001111111100000", -- t[8160] = 1
      "00001" when "001111111100001", -- t[8161] = 1
      "00001" when "001111111100010", -- t[8162] = 1
      "00001" when "001111111100011", -- t[8163] = 1
      "00001" when "001111111100100", -- t[8164] = 1
      "00001" when "001111111100101", -- t[8165] = 1
      "00001" when "001111111100110", -- t[8166] = 1
      "00001" when "001111111100111", -- t[8167] = 1
      "00001" when "001111111101000", -- t[8168] = 1
      "00001" when "001111111101001", -- t[8169] = 1
      "00001" when "001111111101010", -- t[8170] = 1
      "00001" when "001111111101011", -- t[8171] = 1
      "00001" when "001111111101100", -- t[8172] = 1
      "00001" when "001111111101101", -- t[8173] = 1
      "00001" when "001111111101110", -- t[8174] = 1
      "00001" when "001111111101111", -- t[8175] = 1
      "00001" when "001111111110000", -- t[8176] = 1
      "00001" when "001111111110001", -- t[8177] = 1
      "00001" when "001111111110010", -- t[8178] = 1
      "00001" when "001111111110011", -- t[8179] = 1
      "00001" when "001111111110100", -- t[8180] = 1
      "00001" when "001111111110101", -- t[8181] = 1
      "00001" when "001111111110110", -- t[8182] = 1
      "00001" when "001111111110111", -- t[8183] = 1
      "00001" when "001111111111000", -- t[8184] = 1
      "00001" when "001111111111001", -- t[8185] = 1
      "00001" when "001111111111010", -- t[8186] = 1
      "00001" when "001111111111011", -- t[8187] = 1
      "00001" when "001111111111100", -- t[8188] = 1
      "00001" when "001111111111101", -- t[8189] = 1
      "00001" when "001111111111110", -- t[8190] = 1
      "00001" when "001111111111111", -- t[8191] = 1
      "00001" when "010000000000000", -- t[8192] = 1
      "00001" when "010000000000001", -- t[8193] = 1
      "00001" when "010000000000010", -- t[8194] = 1
      "00001" when "010000000000011", -- t[8195] = 1
      "00001" when "010000000000100", -- t[8196] = 1
      "00001" when "010000000000101", -- t[8197] = 1
      "00001" when "010000000000110", -- t[8198] = 1
      "00001" when "010000000000111", -- t[8199] = 1
      "00001" when "010000000001000", -- t[8200] = 1
      "00001" when "010000000001001", -- t[8201] = 1
      "00001" when "010000000001010", -- t[8202] = 1
      "00001" when "010000000001011", -- t[8203] = 1
      "00001" when "010000000001100", -- t[8204] = 1
      "00001" when "010000000001101", -- t[8205] = 1
      "00001" when "010000000001110", -- t[8206] = 1
      "00001" when "010000000001111", -- t[8207] = 1
      "00001" when "010000000010000", -- t[8208] = 1
      "00001" when "010000000010001", -- t[8209] = 1
      "00001" when "010000000010010", -- t[8210] = 1
      "00001" when "010000000010011", -- t[8211] = 1
      "00001" when "010000000010100", -- t[8212] = 1
      "00001" when "010000000010101", -- t[8213] = 1
      "00001" when "010000000010110", -- t[8214] = 1
      "00001" when "010000000010111", -- t[8215] = 1
      "00001" when "010000000011000", -- t[8216] = 1
      "00001" when "010000000011001", -- t[8217] = 1
      "00001" when "010000000011010", -- t[8218] = 1
      "00001" when "010000000011011", -- t[8219] = 1
      "00001" when "010000000011100", -- t[8220] = 1
      "00001" when "010000000011101", -- t[8221] = 1
      "00001" when "010000000011110", -- t[8222] = 1
      "00001" when "010000000011111", -- t[8223] = 1
      "00001" when "010000000100000", -- t[8224] = 1
      "00001" when "010000000100001", -- t[8225] = 1
      "00001" when "010000000100010", -- t[8226] = 1
      "00001" when "010000000100011", -- t[8227] = 1
      "00001" when "010000000100100", -- t[8228] = 1
      "00001" when "010000000100101", -- t[8229] = 1
      "00001" when "010000000100110", -- t[8230] = 1
      "00001" when "010000000100111", -- t[8231] = 1
      "00001" when "010000000101000", -- t[8232] = 1
      "00001" when "010000000101001", -- t[8233] = 1
      "00001" when "010000000101010", -- t[8234] = 1
      "00001" when "010000000101011", -- t[8235] = 1
      "00001" when "010000000101100", -- t[8236] = 1
      "00001" when "010000000101101", -- t[8237] = 1
      "00001" when "010000000101110", -- t[8238] = 1
      "00001" when "010000000101111", -- t[8239] = 1
      "00001" when "010000000110000", -- t[8240] = 1
      "00001" when "010000000110001", -- t[8241] = 1
      "00001" when "010000000110010", -- t[8242] = 1
      "00001" when "010000000110011", -- t[8243] = 1
      "00001" when "010000000110100", -- t[8244] = 1
      "00001" when "010000000110101", -- t[8245] = 1
      "00001" when "010000000110110", -- t[8246] = 1
      "00001" when "010000000110111", -- t[8247] = 1
      "00001" when "010000000111000", -- t[8248] = 1
      "00001" when "010000000111001", -- t[8249] = 1
      "00001" when "010000000111010", -- t[8250] = 1
      "00001" when "010000000111011", -- t[8251] = 1
      "00001" when "010000000111100", -- t[8252] = 1
      "00001" when "010000000111101", -- t[8253] = 1
      "00001" when "010000000111110", -- t[8254] = 1
      "00001" when "010000000111111", -- t[8255] = 1
      "00001" when "010000001000000", -- t[8256] = 1
      "00001" when "010000001000001", -- t[8257] = 1
      "00001" when "010000001000010", -- t[8258] = 1
      "00001" when "010000001000011", -- t[8259] = 1
      "00001" when "010000001000100", -- t[8260] = 1
      "00001" when "010000001000101", -- t[8261] = 1
      "00001" when "010000001000110", -- t[8262] = 1
      "00001" when "010000001000111", -- t[8263] = 1
      "00001" when "010000001001000", -- t[8264] = 1
      "00001" when "010000001001001", -- t[8265] = 1
      "00001" when "010000001001010", -- t[8266] = 1
      "00001" when "010000001001011", -- t[8267] = 1
      "00001" when "010000001001100", -- t[8268] = 1
      "00001" when "010000001001101", -- t[8269] = 1
      "00001" when "010000001001110", -- t[8270] = 1
      "00001" when "010000001001111", -- t[8271] = 1
      "00001" when "010000001010000", -- t[8272] = 1
      "00001" when "010000001010001", -- t[8273] = 1
      "00001" when "010000001010010", -- t[8274] = 1
      "00001" when "010000001010011", -- t[8275] = 1
      "00001" when "010000001010100", -- t[8276] = 1
      "00001" when "010000001010101", -- t[8277] = 1
      "00001" when "010000001010110", -- t[8278] = 1
      "00001" when "010000001010111", -- t[8279] = 1
      "00001" when "010000001011000", -- t[8280] = 1
      "00001" when "010000001011001", -- t[8281] = 1
      "00001" when "010000001011010", -- t[8282] = 1
      "00001" when "010000001011011", -- t[8283] = 1
      "00001" when "010000001011100", -- t[8284] = 1
      "00001" when "010000001011101", -- t[8285] = 1
      "00001" when "010000001011110", -- t[8286] = 1
      "00001" when "010000001011111", -- t[8287] = 1
      "00001" when "010000001100000", -- t[8288] = 1
      "00001" when "010000001100001", -- t[8289] = 1
      "00001" when "010000001100010", -- t[8290] = 1
      "00001" when "010000001100011", -- t[8291] = 1
      "00001" when "010000001100100", -- t[8292] = 1
      "00001" when "010000001100101", -- t[8293] = 1
      "00001" when "010000001100110", -- t[8294] = 1
      "00001" when "010000001100111", -- t[8295] = 1
      "00001" when "010000001101000", -- t[8296] = 1
      "00001" when "010000001101001", -- t[8297] = 1
      "00001" when "010000001101010", -- t[8298] = 1
      "00001" when "010000001101011", -- t[8299] = 1
      "00001" when "010000001101100", -- t[8300] = 1
      "00001" when "010000001101101", -- t[8301] = 1
      "00001" when "010000001101110", -- t[8302] = 1
      "00001" when "010000001101111", -- t[8303] = 1
      "00001" when "010000001110000", -- t[8304] = 1
      "00001" when "010000001110001", -- t[8305] = 1
      "00001" when "010000001110010", -- t[8306] = 1
      "00001" when "010000001110011", -- t[8307] = 1
      "00001" when "010000001110100", -- t[8308] = 1
      "00001" when "010000001110101", -- t[8309] = 1
      "00001" when "010000001110110", -- t[8310] = 1
      "00001" when "010000001110111", -- t[8311] = 1
      "00001" when "010000001111000", -- t[8312] = 1
      "00001" when "010000001111001", -- t[8313] = 1
      "00001" when "010000001111010", -- t[8314] = 1
      "00001" when "010000001111011", -- t[8315] = 1
      "00001" when "010000001111100", -- t[8316] = 1
      "00001" when "010000001111101", -- t[8317] = 1
      "00001" when "010000001111110", -- t[8318] = 1
      "00001" when "010000001111111", -- t[8319] = 1
      "00001" when "010000010000000", -- t[8320] = 1
      "00001" when "010000010000001", -- t[8321] = 1
      "00001" when "010000010000010", -- t[8322] = 1
      "00001" when "010000010000011", -- t[8323] = 1
      "00001" when "010000010000100", -- t[8324] = 1
      "00001" when "010000010000101", -- t[8325] = 1
      "00001" when "010000010000110", -- t[8326] = 1
      "00001" when "010000010000111", -- t[8327] = 1
      "00001" when "010000010001000", -- t[8328] = 1
      "00001" when "010000010001001", -- t[8329] = 1
      "00001" when "010000010001010", -- t[8330] = 1
      "00001" when "010000010001011", -- t[8331] = 1
      "00001" when "010000010001100", -- t[8332] = 1
      "00001" when "010000010001101", -- t[8333] = 1
      "00001" when "010000010001110", -- t[8334] = 1
      "00001" when "010000010001111", -- t[8335] = 1
      "00001" when "010000010010000", -- t[8336] = 1
      "00001" when "010000010010001", -- t[8337] = 1
      "00001" when "010000010010010", -- t[8338] = 1
      "00001" when "010000010010011", -- t[8339] = 1
      "00001" when "010000010010100", -- t[8340] = 1
      "00001" when "010000010010101", -- t[8341] = 1
      "00001" when "010000010010110", -- t[8342] = 1
      "00001" when "010000010010111", -- t[8343] = 1
      "00001" when "010000010011000", -- t[8344] = 1
      "00001" when "010000010011001", -- t[8345] = 1
      "00001" when "010000010011010", -- t[8346] = 1
      "00001" when "010000010011011", -- t[8347] = 1
      "00001" when "010000010011100", -- t[8348] = 1
      "00001" when "010000010011101", -- t[8349] = 1
      "00001" when "010000010011110", -- t[8350] = 1
      "00001" when "010000010011111", -- t[8351] = 1
      "00001" when "010000010100000", -- t[8352] = 1
      "00001" when "010000010100001", -- t[8353] = 1
      "00001" when "010000010100010", -- t[8354] = 1
      "00001" when "010000010100011", -- t[8355] = 1
      "00001" when "010000010100100", -- t[8356] = 1
      "00001" when "010000010100101", -- t[8357] = 1
      "00001" when "010000010100110", -- t[8358] = 1
      "00001" when "010000010100111", -- t[8359] = 1
      "00001" when "010000010101000", -- t[8360] = 1
      "00001" when "010000010101001", -- t[8361] = 1
      "00001" when "010000010101010", -- t[8362] = 1
      "00001" when "010000010101011", -- t[8363] = 1
      "00001" when "010000010101100", -- t[8364] = 1
      "00001" when "010000010101101", -- t[8365] = 1
      "00001" when "010000010101110", -- t[8366] = 1
      "00001" when "010000010101111", -- t[8367] = 1
      "00001" when "010000010110000", -- t[8368] = 1
      "00001" when "010000010110001", -- t[8369] = 1
      "00001" when "010000010110010", -- t[8370] = 1
      "00001" when "010000010110011", -- t[8371] = 1
      "00001" when "010000010110100", -- t[8372] = 1
      "00001" when "010000010110101", -- t[8373] = 1
      "00001" when "010000010110110", -- t[8374] = 1
      "00001" when "010000010110111", -- t[8375] = 1
      "00001" when "010000010111000", -- t[8376] = 1
      "00001" when "010000010111001", -- t[8377] = 1
      "00001" when "010000010111010", -- t[8378] = 1
      "00001" when "010000010111011", -- t[8379] = 1
      "00001" when "010000010111100", -- t[8380] = 1
      "00001" when "010000010111101", -- t[8381] = 1
      "00001" when "010000010111110", -- t[8382] = 1
      "00001" when "010000010111111", -- t[8383] = 1
      "00001" when "010000011000000", -- t[8384] = 1
      "00001" when "010000011000001", -- t[8385] = 1
      "00001" when "010000011000010", -- t[8386] = 1
      "00001" when "010000011000011", -- t[8387] = 1
      "00001" when "010000011000100", -- t[8388] = 1
      "00001" when "010000011000101", -- t[8389] = 1
      "00001" when "010000011000110", -- t[8390] = 1
      "00001" when "010000011000111", -- t[8391] = 1
      "00001" when "010000011001000", -- t[8392] = 1
      "00001" when "010000011001001", -- t[8393] = 1
      "00001" when "010000011001010", -- t[8394] = 1
      "00001" when "010000011001011", -- t[8395] = 1
      "00001" when "010000011001100", -- t[8396] = 1
      "00001" when "010000011001101", -- t[8397] = 1
      "00001" when "010000011001110", -- t[8398] = 1
      "00001" when "010000011001111", -- t[8399] = 1
      "00001" when "010000011010000", -- t[8400] = 1
      "00001" when "010000011010001", -- t[8401] = 1
      "00001" when "010000011010010", -- t[8402] = 1
      "00001" when "010000011010011", -- t[8403] = 1
      "00001" when "010000011010100", -- t[8404] = 1
      "00001" when "010000011010101", -- t[8405] = 1
      "00001" when "010000011010110", -- t[8406] = 1
      "00001" when "010000011010111", -- t[8407] = 1
      "00001" when "010000011011000", -- t[8408] = 1
      "00001" when "010000011011001", -- t[8409] = 1
      "00001" when "010000011011010", -- t[8410] = 1
      "00001" when "010000011011011", -- t[8411] = 1
      "00001" when "010000011011100", -- t[8412] = 1
      "00001" when "010000011011101", -- t[8413] = 1
      "00001" when "010000011011110", -- t[8414] = 1
      "00001" when "010000011011111", -- t[8415] = 1
      "00001" when "010000011100000", -- t[8416] = 1
      "00001" when "010000011100001", -- t[8417] = 1
      "00001" when "010000011100010", -- t[8418] = 1
      "00001" when "010000011100011", -- t[8419] = 1
      "00001" when "010000011100100", -- t[8420] = 1
      "00001" when "010000011100101", -- t[8421] = 1
      "00001" when "010000011100110", -- t[8422] = 1
      "00001" when "010000011100111", -- t[8423] = 1
      "00001" when "010000011101000", -- t[8424] = 1
      "00001" when "010000011101001", -- t[8425] = 1
      "00001" when "010000011101010", -- t[8426] = 1
      "00001" when "010000011101011", -- t[8427] = 1
      "00001" when "010000011101100", -- t[8428] = 1
      "00001" when "010000011101101", -- t[8429] = 1
      "00001" when "010000011101110", -- t[8430] = 1
      "00001" when "010000011101111", -- t[8431] = 1
      "00001" when "010000011110000", -- t[8432] = 1
      "00001" when "010000011110001", -- t[8433] = 1
      "00001" when "010000011110010", -- t[8434] = 1
      "00001" when "010000011110011", -- t[8435] = 1
      "00001" when "010000011110100", -- t[8436] = 1
      "00001" when "010000011110101", -- t[8437] = 1
      "00001" when "010000011110110", -- t[8438] = 1
      "00001" when "010000011110111", -- t[8439] = 1
      "00001" when "010000011111000", -- t[8440] = 1
      "00001" when "010000011111001", -- t[8441] = 1
      "00001" when "010000011111010", -- t[8442] = 1
      "00001" when "010000011111011", -- t[8443] = 1
      "00001" when "010000011111100", -- t[8444] = 1
      "00001" when "010000011111101", -- t[8445] = 1
      "00001" when "010000011111110", -- t[8446] = 1
      "00001" when "010000011111111", -- t[8447] = 1
      "00001" when "010000100000000", -- t[8448] = 1
      "00001" when "010000100000001", -- t[8449] = 1
      "00001" when "010000100000010", -- t[8450] = 1
      "00001" when "010000100000011", -- t[8451] = 1
      "00001" when "010000100000100", -- t[8452] = 1
      "00001" when "010000100000101", -- t[8453] = 1
      "00001" when "010000100000110", -- t[8454] = 1
      "00001" when "010000100000111", -- t[8455] = 1
      "00001" when "010000100001000", -- t[8456] = 1
      "00001" when "010000100001001", -- t[8457] = 1
      "00001" when "010000100001010", -- t[8458] = 1
      "00001" when "010000100001011", -- t[8459] = 1
      "00001" when "010000100001100", -- t[8460] = 1
      "00001" when "010000100001101", -- t[8461] = 1
      "00001" when "010000100001110", -- t[8462] = 1
      "00001" when "010000100001111", -- t[8463] = 1
      "00001" when "010000100010000", -- t[8464] = 1
      "00001" when "010000100010001", -- t[8465] = 1
      "00001" when "010000100010010", -- t[8466] = 1
      "00001" when "010000100010011", -- t[8467] = 1
      "00001" when "010000100010100", -- t[8468] = 1
      "00001" when "010000100010101", -- t[8469] = 1
      "00001" when "010000100010110", -- t[8470] = 1
      "00001" when "010000100010111", -- t[8471] = 1
      "00001" when "010000100011000", -- t[8472] = 1
      "00001" when "010000100011001", -- t[8473] = 1
      "00001" when "010000100011010", -- t[8474] = 1
      "00001" when "010000100011011", -- t[8475] = 1
      "00001" when "010000100011100", -- t[8476] = 1
      "00001" when "010000100011101", -- t[8477] = 1
      "00001" when "010000100011110", -- t[8478] = 1
      "00001" when "010000100011111", -- t[8479] = 1
      "00001" when "010000100100000", -- t[8480] = 1
      "00001" when "010000100100001", -- t[8481] = 1
      "00001" when "010000100100010", -- t[8482] = 1
      "00001" when "010000100100011", -- t[8483] = 1
      "00001" when "010000100100100", -- t[8484] = 1
      "00001" when "010000100100101", -- t[8485] = 1
      "00001" when "010000100100110", -- t[8486] = 1
      "00001" when "010000100100111", -- t[8487] = 1
      "00001" when "010000100101000", -- t[8488] = 1
      "00001" when "010000100101001", -- t[8489] = 1
      "00001" when "010000100101010", -- t[8490] = 1
      "00001" when "010000100101011", -- t[8491] = 1
      "00001" when "010000100101100", -- t[8492] = 1
      "00001" when "010000100101101", -- t[8493] = 1
      "00001" when "010000100101110", -- t[8494] = 1
      "00001" when "010000100101111", -- t[8495] = 1
      "00001" when "010000100110000", -- t[8496] = 1
      "00001" when "010000100110001", -- t[8497] = 1
      "00001" when "010000100110010", -- t[8498] = 1
      "00001" when "010000100110011", -- t[8499] = 1
      "00001" when "010000100110100", -- t[8500] = 1
      "00001" when "010000100110101", -- t[8501] = 1
      "00001" when "010000100110110", -- t[8502] = 1
      "00001" when "010000100110111", -- t[8503] = 1
      "00001" when "010000100111000", -- t[8504] = 1
      "00001" when "010000100111001", -- t[8505] = 1
      "00001" when "010000100111010", -- t[8506] = 1
      "00001" when "010000100111011", -- t[8507] = 1
      "00001" when "010000100111100", -- t[8508] = 1
      "00001" when "010000100111101", -- t[8509] = 1
      "00001" when "010000100111110", -- t[8510] = 1
      "00001" when "010000100111111", -- t[8511] = 1
      "00001" when "010000101000000", -- t[8512] = 1
      "00001" when "010000101000001", -- t[8513] = 1
      "00001" when "010000101000010", -- t[8514] = 1
      "00001" when "010000101000011", -- t[8515] = 1
      "00001" when "010000101000100", -- t[8516] = 1
      "00001" when "010000101000101", -- t[8517] = 1
      "00001" when "010000101000110", -- t[8518] = 1
      "00001" when "010000101000111", -- t[8519] = 1
      "00001" when "010000101001000", -- t[8520] = 1
      "00001" when "010000101001001", -- t[8521] = 1
      "00001" when "010000101001010", -- t[8522] = 1
      "00001" when "010000101001011", -- t[8523] = 1
      "00001" when "010000101001100", -- t[8524] = 1
      "00001" when "010000101001101", -- t[8525] = 1
      "00001" when "010000101001110", -- t[8526] = 1
      "00001" when "010000101001111", -- t[8527] = 1
      "00001" when "010000101010000", -- t[8528] = 1
      "00001" when "010000101010001", -- t[8529] = 1
      "00001" when "010000101010010", -- t[8530] = 1
      "00001" when "010000101010011", -- t[8531] = 1
      "00001" when "010000101010100", -- t[8532] = 1
      "00001" when "010000101010101", -- t[8533] = 1
      "00001" when "010000101010110", -- t[8534] = 1
      "00001" when "010000101010111", -- t[8535] = 1
      "00001" when "010000101011000", -- t[8536] = 1
      "00001" when "010000101011001", -- t[8537] = 1
      "00001" when "010000101011010", -- t[8538] = 1
      "00001" when "010000101011011", -- t[8539] = 1
      "00001" when "010000101011100", -- t[8540] = 1
      "00001" when "010000101011101", -- t[8541] = 1
      "00001" when "010000101011110", -- t[8542] = 1
      "00001" when "010000101011111", -- t[8543] = 1
      "00001" when "010000101100000", -- t[8544] = 1
      "00001" when "010000101100001", -- t[8545] = 1
      "00001" when "010000101100010", -- t[8546] = 1
      "00001" when "010000101100011", -- t[8547] = 1
      "00001" when "010000101100100", -- t[8548] = 1
      "00001" when "010000101100101", -- t[8549] = 1
      "00001" when "010000101100110", -- t[8550] = 1
      "00001" when "010000101100111", -- t[8551] = 1
      "00001" when "010000101101000", -- t[8552] = 1
      "00001" when "010000101101001", -- t[8553] = 1
      "00001" when "010000101101010", -- t[8554] = 1
      "00001" when "010000101101011", -- t[8555] = 1
      "00001" when "010000101101100", -- t[8556] = 1
      "00001" when "010000101101101", -- t[8557] = 1
      "00001" when "010000101101110", -- t[8558] = 1
      "00001" when "010000101101111", -- t[8559] = 1
      "00001" when "010000101110000", -- t[8560] = 1
      "00001" when "010000101110001", -- t[8561] = 1
      "00001" when "010000101110010", -- t[8562] = 1
      "00001" when "010000101110011", -- t[8563] = 1
      "00001" when "010000101110100", -- t[8564] = 1
      "00001" when "010000101110101", -- t[8565] = 1
      "00001" when "010000101110110", -- t[8566] = 1
      "00001" when "010000101110111", -- t[8567] = 1
      "00001" when "010000101111000", -- t[8568] = 1
      "00001" when "010000101111001", -- t[8569] = 1
      "00001" when "010000101111010", -- t[8570] = 1
      "00001" when "010000101111011", -- t[8571] = 1
      "00001" when "010000101111100", -- t[8572] = 1
      "00001" when "010000101111101", -- t[8573] = 1
      "00001" when "010000101111110", -- t[8574] = 1
      "00001" when "010000101111111", -- t[8575] = 1
      "00001" when "010000110000000", -- t[8576] = 1
      "00001" when "010000110000001", -- t[8577] = 1
      "00001" when "010000110000010", -- t[8578] = 1
      "00001" when "010000110000011", -- t[8579] = 1
      "00001" when "010000110000100", -- t[8580] = 1
      "00001" when "010000110000101", -- t[8581] = 1
      "00001" when "010000110000110", -- t[8582] = 1
      "00001" when "010000110000111", -- t[8583] = 1
      "00001" when "010000110001000", -- t[8584] = 1
      "00001" when "010000110001001", -- t[8585] = 1
      "00001" when "010000110001010", -- t[8586] = 1
      "00001" when "010000110001011", -- t[8587] = 1
      "00001" when "010000110001100", -- t[8588] = 1
      "00001" when "010000110001101", -- t[8589] = 1
      "00001" when "010000110001110", -- t[8590] = 1
      "00001" when "010000110001111", -- t[8591] = 1
      "00001" when "010000110010000", -- t[8592] = 1
      "00001" when "010000110010001", -- t[8593] = 1
      "00001" when "010000110010010", -- t[8594] = 1
      "00001" when "010000110010011", -- t[8595] = 1
      "00001" when "010000110010100", -- t[8596] = 1
      "00001" when "010000110010101", -- t[8597] = 1
      "00001" when "010000110010110", -- t[8598] = 1
      "00001" when "010000110010111", -- t[8599] = 1
      "00001" when "010000110011000", -- t[8600] = 1
      "00001" when "010000110011001", -- t[8601] = 1
      "00001" when "010000110011010", -- t[8602] = 1
      "00001" when "010000110011011", -- t[8603] = 1
      "00001" when "010000110011100", -- t[8604] = 1
      "00001" when "010000110011101", -- t[8605] = 1
      "00001" when "010000110011110", -- t[8606] = 1
      "00001" when "010000110011111", -- t[8607] = 1
      "00001" when "010000110100000", -- t[8608] = 1
      "00001" when "010000110100001", -- t[8609] = 1
      "00001" when "010000110100010", -- t[8610] = 1
      "00001" when "010000110100011", -- t[8611] = 1
      "00001" when "010000110100100", -- t[8612] = 1
      "00001" when "010000110100101", -- t[8613] = 1
      "00001" when "010000110100110", -- t[8614] = 1
      "00001" when "010000110100111", -- t[8615] = 1
      "00001" when "010000110101000", -- t[8616] = 1
      "00001" when "010000110101001", -- t[8617] = 1
      "00001" when "010000110101010", -- t[8618] = 1
      "00001" when "010000110101011", -- t[8619] = 1
      "00001" when "010000110101100", -- t[8620] = 1
      "00001" when "010000110101101", -- t[8621] = 1
      "00001" when "010000110101110", -- t[8622] = 1
      "00001" when "010000110101111", -- t[8623] = 1
      "00001" when "010000110110000", -- t[8624] = 1
      "00001" when "010000110110001", -- t[8625] = 1
      "00001" when "010000110110010", -- t[8626] = 1
      "00001" when "010000110110011", -- t[8627] = 1
      "00001" when "010000110110100", -- t[8628] = 1
      "00001" when "010000110110101", -- t[8629] = 1
      "00001" when "010000110110110", -- t[8630] = 1
      "00001" when "010000110110111", -- t[8631] = 1
      "00001" when "010000110111000", -- t[8632] = 1
      "00001" when "010000110111001", -- t[8633] = 1
      "00001" when "010000110111010", -- t[8634] = 1
      "00001" when "010000110111011", -- t[8635] = 1
      "00001" when "010000110111100", -- t[8636] = 1
      "00001" when "010000110111101", -- t[8637] = 1
      "00001" when "010000110111110", -- t[8638] = 1
      "00001" when "010000110111111", -- t[8639] = 1
      "00001" when "010000111000000", -- t[8640] = 1
      "00001" when "010000111000001", -- t[8641] = 1
      "00001" when "010000111000010", -- t[8642] = 1
      "00001" when "010000111000011", -- t[8643] = 1
      "00001" when "010000111000100", -- t[8644] = 1
      "00001" when "010000111000101", -- t[8645] = 1
      "00001" when "010000111000110", -- t[8646] = 1
      "00001" when "010000111000111", -- t[8647] = 1
      "00001" when "010000111001000", -- t[8648] = 1
      "00001" when "010000111001001", -- t[8649] = 1
      "00001" when "010000111001010", -- t[8650] = 1
      "00001" when "010000111001011", -- t[8651] = 1
      "00001" when "010000111001100", -- t[8652] = 1
      "00001" when "010000111001101", -- t[8653] = 1
      "00001" when "010000111001110", -- t[8654] = 1
      "00001" when "010000111001111", -- t[8655] = 1
      "00001" when "010000111010000", -- t[8656] = 1
      "00001" when "010000111010001", -- t[8657] = 1
      "00001" when "010000111010010", -- t[8658] = 1
      "00001" when "010000111010011", -- t[8659] = 1
      "00001" when "010000111010100", -- t[8660] = 1
      "00001" when "010000111010101", -- t[8661] = 1
      "00001" when "010000111010110", -- t[8662] = 1
      "00001" when "010000111010111", -- t[8663] = 1
      "00001" when "010000111011000", -- t[8664] = 1
      "00001" when "010000111011001", -- t[8665] = 1
      "00001" when "010000111011010", -- t[8666] = 1
      "00001" when "010000111011011", -- t[8667] = 1
      "00001" when "010000111011100", -- t[8668] = 1
      "00001" when "010000111011101", -- t[8669] = 1
      "00001" when "010000111011110", -- t[8670] = 1
      "00001" when "010000111011111", -- t[8671] = 1
      "00001" when "010000111100000", -- t[8672] = 1
      "00001" when "010000111100001", -- t[8673] = 1
      "00001" when "010000111100010", -- t[8674] = 1
      "00001" when "010000111100011", -- t[8675] = 1
      "00001" when "010000111100100", -- t[8676] = 1
      "00001" when "010000111100101", -- t[8677] = 1
      "00001" when "010000111100110", -- t[8678] = 1
      "00001" when "010000111100111", -- t[8679] = 1
      "00001" when "010000111101000", -- t[8680] = 1
      "00001" when "010000111101001", -- t[8681] = 1
      "00001" when "010000111101010", -- t[8682] = 1
      "00001" when "010000111101011", -- t[8683] = 1
      "00001" when "010000111101100", -- t[8684] = 1
      "00001" when "010000111101101", -- t[8685] = 1
      "00001" when "010000111101110", -- t[8686] = 1
      "00001" when "010000111101111", -- t[8687] = 1
      "00001" when "010000111110000", -- t[8688] = 1
      "00001" when "010000111110001", -- t[8689] = 1
      "00001" when "010000111110010", -- t[8690] = 1
      "00001" when "010000111110011", -- t[8691] = 1
      "00001" when "010000111110100", -- t[8692] = 1
      "00001" when "010000111110101", -- t[8693] = 1
      "00001" when "010000111110110", -- t[8694] = 1
      "00001" when "010000111110111", -- t[8695] = 1
      "00001" when "010000111111000", -- t[8696] = 1
      "00001" when "010000111111001", -- t[8697] = 1
      "00001" when "010000111111010", -- t[8698] = 1
      "00001" when "010000111111011", -- t[8699] = 1
      "00001" when "010000111111100", -- t[8700] = 1
      "00001" when "010000111111101", -- t[8701] = 1
      "00001" when "010000111111110", -- t[8702] = 1
      "00001" when "010000111111111", -- t[8703] = 1
      "00001" when "010001000000000", -- t[8704] = 1
      "00001" when "010001000000001", -- t[8705] = 1
      "00001" when "010001000000010", -- t[8706] = 1
      "00001" when "010001000000011", -- t[8707] = 1
      "00001" when "010001000000100", -- t[8708] = 1
      "00001" when "010001000000101", -- t[8709] = 1
      "00001" when "010001000000110", -- t[8710] = 1
      "00001" when "010001000000111", -- t[8711] = 1
      "00001" when "010001000001000", -- t[8712] = 1
      "00001" when "010001000001001", -- t[8713] = 1
      "00001" when "010001000001010", -- t[8714] = 1
      "00001" when "010001000001011", -- t[8715] = 1
      "00001" when "010001000001100", -- t[8716] = 1
      "00001" when "010001000001101", -- t[8717] = 1
      "00001" when "010001000001110", -- t[8718] = 1
      "00001" when "010001000001111", -- t[8719] = 1
      "00001" when "010001000010000", -- t[8720] = 1
      "00001" when "010001000010001", -- t[8721] = 1
      "00001" when "010001000010010", -- t[8722] = 1
      "00001" when "010001000010011", -- t[8723] = 1
      "00001" when "010001000010100", -- t[8724] = 1
      "00001" when "010001000010101", -- t[8725] = 1
      "00001" when "010001000010110", -- t[8726] = 1
      "00001" when "010001000010111", -- t[8727] = 1
      "00001" when "010001000011000", -- t[8728] = 1
      "00001" when "010001000011001", -- t[8729] = 1
      "00001" when "010001000011010", -- t[8730] = 1
      "00001" when "010001000011011", -- t[8731] = 1
      "00001" when "010001000011100", -- t[8732] = 1
      "00001" when "010001000011101", -- t[8733] = 1
      "00001" when "010001000011110", -- t[8734] = 1
      "00001" when "010001000011111", -- t[8735] = 1
      "00001" when "010001000100000", -- t[8736] = 1
      "00001" when "010001000100001", -- t[8737] = 1
      "00001" when "010001000100010", -- t[8738] = 1
      "00001" when "010001000100011", -- t[8739] = 1
      "00001" when "010001000100100", -- t[8740] = 1
      "00001" when "010001000100101", -- t[8741] = 1
      "00001" when "010001000100110", -- t[8742] = 1
      "00001" when "010001000100111", -- t[8743] = 1
      "00001" when "010001000101000", -- t[8744] = 1
      "00001" when "010001000101001", -- t[8745] = 1
      "00001" when "010001000101010", -- t[8746] = 1
      "00001" when "010001000101011", -- t[8747] = 1
      "00001" when "010001000101100", -- t[8748] = 1
      "00001" when "010001000101101", -- t[8749] = 1
      "00001" when "010001000101110", -- t[8750] = 1
      "00001" when "010001000101111", -- t[8751] = 1
      "00001" when "010001000110000", -- t[8752] = 1
      "00001" when "010001000110001", -- t[8753] = 1
      "00001" when "010001000110010", -- t[8754] = 1
      "00001" when "010001000110011", -- t[8755] = 1
      "00001" when "010001000110100", -- t[8756] = 1
      "00001" when "010001000110101", -- t[8757] = 1
      "00001" when "010001000110110", -- t[8758] = 1
      "00001" when "010001000110111", -- t[8759] = 1
      "00001" when "010001000111000", -- t[8760] = 1
      "00001" when "010001000111001", -- t[8761] = 1
      "00001" when "010001000111010", -- t[8762] = 1
      "00001" when "010001000111011", -- t[8763] = 1
      "00001" when "010001000111100", -- t[8764] = 1
      "00001" when "010001000111101", -- t[8765] = 1
      "00001" when "010001000111110", -- t[8766] = 1
      "00001" when "010001000111111", -- t[8767] = 1
      "00001" when "010001001000000", -- t[8768] = 1
      "00001" when "010001001000001", -- t[8769] = 1
      "00001" when "010001001000010", -- t[8770] = 1
      "00001" when "010001001000011", -- t[8771] = 1
      "00001" when "010001001000100", -- t[8772] = 1
      "00001" when "010001001000101", -- t[8773] = 1
      "00001" when "010001001000110", -- t[8774] = 1
      "00001" when "010001001000111", -- t[8775] = 1
      "00001" when "010001001001000", -- t[8776] = 1
      "00001" when "010001001001001", -- t[8777] = 1
      "00001" when "010001001001010", -- t[8778] = 1
      "00001" when "010001001001011", -- t[8779] = 1
      "00001" when "010001001001100", -- t[8780] = 1
      "00001" when "010001001001101", -- t[8781] = 1
      "00001" when "010001001001110", -- t[8782] = 1
      "00001" when "010001001001111", -- t[8783] = 1
      "00001" when "010001001010000", -- t[8784] = 1
      "00001" when "010001001010001", -- t[8785] = 1
      "00001" when "010001001010010", -- t[8786] = 1
      "00001" when "010001001010011", -- t[8787] = 1
      "00001" when "010001001010100", -- t[8788] = 1
      "00001" when "010001001010101", -- t[8789] = 1
      "00001" when "010001001010110", -- t[8790] = 1
      "00001" when "010001001010111", -- t[8791] = 1
      "00001" when "010001001011000", -- t[8792] = 1
      "00001" when "010001001011001", -- t[8793] = 1
      "00001" when "010001001011010", -- t[8794] = 1
      "00001" when "010001001011011", -- t[8795] = 1
      "00001" when "010001001011100", -- t[8796] = 1
      "00001" when "010001001011101", -- t[8797] = 1
      "00001" when "010001001011110", -- t[8798] = 1
      "00001" when "010001001011111", -- t[8799] = 1
      "00001" when "010001001100000", -- t[8800] = 1
      "00001" when "010001001100001", -- t[8801] = 1
      "00001" when "010001001100010", -- t[8802] = 1
      "00001" when "010001001100011", -- t[8803] = 1
      "00001" when "010001001100100", -- t[8804] = 1
      "00001" when "010001001100101", -- t[8805] = 1
      "00001" when "010001001100110", -- t[8806] = 1
      "00001" when "010001001100111", -- t[8807] = 1
      "00001" when "010001001101000", -- t[8808] = 1
      "00001" when "010001001101001", -- t[8809] = 1
      "00001" when "010001001101010", -- t[8810] = 1
      "00001" when "010001001101011", -- t[8811] = 1
      "00001" when "010001001101100", -- t[8812] = 1
      "00001" when "010001001101101", -- t[8813] = 1
      "00001" when "010001001101110", -- t[8814] = 1
      "00001" when "010001001101111", -- t[8815] = 1
      "00001" when "010001001110000", -- t[8816] = 1
      "00001" when "010001001110001", -- t[8817] = 1
      "00001" when "010001001110010", -- t[8818] = 1
      "00001" when "010001001110011", -- t[8819] = 1
      "00001" when "010001001110100", -- t[8820] = 1
      "00001" when "010001001110101", -- t[8821] = 1
      "00001" when "010001001110110", -- t[8822] = 1
      "00001" when "010001001110111", -- t[8823] = 1
      "00001" when "010001001111000", -- t[8824] = 1
      "00001" when "010001001111001", -- t[8825] = 1
      "00001" when "010001001111010", -- t[8826] = 1
      "00001" when "010001001111011", -- t[8827] = 1
      "00001" when "010001001111100", -- t[8828] = 1
      "00001" when "010001001111101", -- t[8829] = 1
      "00001" when "010001001111110", -- t[8830] = 1
      "00001" when "010001001111111", -- t[8831] = 1
      "00001" when "010001010000000", -- t[8832] = 1
      "00001" when "010001010000001", -- t[8833] = 1
      "00001" when "010001010000010", -- t[8834] = 1
      "00001" when "010001010000011", -- t[8835] = 1
      "00001" when "010001010000100", -- t[8836] = 1
      "00001" when "010001010000101", -- t[8837] = 1
      "00001" when "010001010000110", -- t[8838] = 1
      "00001" when "010001010000111", -- t[8839] = 1
      "00001" when "010001010001000", -- t[8840] = 1
      "00001" when "010001010001001", -- t[8841] = 1
      "00001" when "010001010001010", -- t[8842] = 1
      "00001" when "010001010001011", -- t[8843] = 1
      "00001" when "010001010001100", -- t[8844] = 1
      "00001" when "010001010001101", -- t[8845] = 1
      "00001" when "010001010001110", -- t[8846] = 1
      "00001" when "010001010001111", -- t[8847] = 1
      "00001" when "010001010010000", -- t[8848] = 1
      "00001" when "010001010010001", -- t[8849] = 1
      "00001" when "010001010010010", -- t[8850] = 1
      "00001" when "010001010010011", -- t[8851] = 1
      "00001" when "010001010010100", -- t[8852] = 1
      "00001" when "010001010010101", -- t[8853] = 1
      "00001" when "010001010010110", -- t[8854] = 1
      "00001" when "010001010010111", -- t[8855] = 1
      "00001" when "010001010011000", -- t[8856] = 1
      "00001" when "010001010011001", -- t[8857] = 1
      "00001" when "010001010011010", -- t[8858] = 1
      "00001" when "010001010011011", -- t[8859] = 1
      "00001" when "010001010011100", -- t[8860] = 1
      "00001" when "010001010011101", -- t[8861] = 1
      "00001" when "010001010011110", -- t[8862] = 1
      "00001" when "010001010011111", -- t[8863] = 1
      "00001" when "010001010100000", -- t[8864] = 1
      "00001" when "010001010100001", -- t[8865] = 1
      "00001" when "010001010100010", -- t[8866] = 1
      "00001" when "010001010100011", -- t[8867] = 1
      "00001" when "010001010100100", -- t[8868] = 1
      "00001" when "010001010100101", -- t[8869] = 1
      "00001" when "010001010100110", -- t[8870] = 1
      "00001" when "010001010100111", -- t[8871] = 1
      "00001" when "010001010101000", -- t[8872] = 1
      "00001" when "010001010101001", -- t[8873] = 1
      "00001" when "010001010101010", -- t[8874] = 1
      "00001" when "010001010101011", -- t[8875] = 1
      "00001" when "010001010101100", -- t[8876] = 1
      "00001" when "010001010101101", -- t[8877] = 1
      "00001" when "010001010101110", -- t[8878] = 1
      "00001" when "010001010101111", -- t[8879] = 1
      "00001" when "010001010110000", -- t[8880] = 1
      "00001" when "010001010110001", -- t[8881] = 1
      "00001" when "010001010110010", -- t[8882] = 1
      "00001" when "010001010110011", -- t[8883] = 1
      "00001" when "010001010110100", -- t[8884] = 1
      "00001" when "010001010110101", -- t[8885] = 1
      "00001" when "010001010110110", -- t[8886] = 1
      "00001" when "010001010110111", -- t[8887] = 1
      "00001" when "010001010111000", -- t[8888] = 1
      "00001" when "010001010111001", -- t[8889] = 1
      "00001" when "010001010111010", -- t[8890] = 1
      "00001" when "010001010111011", -- t[8891] = 1
      "00001" when "010001010111100", -- t[8892] = 1
      "00001" when "010001010111101", -- t[8893] = 1
      "00001" when "010001010111110", -- t[8894] = 1
      "00001" when "010001010111111", -- t[8895] = 1
      "00001" when "010001011000000", -- t[8896] = 1
      "00001" when "010001011000001", -- t[8897] = 1
      "00001" when "010001011000010", -- t[8898] = 1
      "00001" when "010001011000011", -- t[8899] = 1
      "00001" when "010001011000100", -- t[8900] = 1
      "00001" when "010001011000101", -- t[8901] = 1
      "00001" when "010001011000110", -- t[8902] = 1
      "00001" when "010001011000111", -- t[8903] = 1
      "00001" when "010001011001000", -- t[8904] = 1
      "00001" when "010001011001001", -- t[8905] = 1
      "00001" when "010001011001010", -- t[8906] = 1
      "00001" when "010001011001011", -- t[8907] = 1
      "00001" when "010001011001100", -- t[8908] = 1
      "00001" when "010001011001101", -- t[8909] = 1
      "00001" when "010001011001110", -- t[8910] = 1
      "00001" when "010001011001111", -- t[8911] = 1
      "00001" when "010001011010000", -- t[8912] = 1
      "00001" when "010001011010001", -- t[8913] = 1
      "00001" when "010001011010010", -- t[8914] = 1
      "00001" when "010001011010011", -- t[8915] = 1
      "00001" when "010001011010100", -- t[8916] = 1
      "00001" when "010001011010101", -- t[8917] = 1
      "00001" when "010001011010110", -- t[8918] = 1
      "00001" when "010001011010111", -- t[8919] = 1
      "00001" when "010001011011000", -- t[8920] = 1
      "00001" when "010001011011001", -- t[8921] = 1
      "00001" when "010001011011010", -- t[8922] = 1
      "00001" when "010001011011011", -- t[8923] = 1
      "00001" when "010001011011100", -- t[8924] = 1
      "00001" when "010001011011101", -- t[8925] = 1
      "00001" when "010001011011110", -- t[8926] = 1
      "00001" when "010001011011111", -- t[8927] = 1
      "00001" when "010001011100000", -- t[8928] = 1
      "00001" when "010001011100001", -- t[8929] = 1
      "00001" when "010001011100010", -- t[8930] = 1
      "00001" when "010001011100011", -- t[8931] = 1
      "00001" when "010001011100100", -- t[8932] = 1
      "00001" when "010001011100101", -- t[8933] = 1
      "00001" when "010001011100110", -- t[8934] = 1
      "00001" when "010001011100111", -- t[8935] = 1
      "00001" when "010001011101000", -- t[8936] = 1
      "00001" when "010001011101001", -- t[8937] = 1
      "00001" when "010001011101010", -- t[8938] = 1
      "00001" when "010001011101011", -- t[8939] = 1
      "00001" when "010001011101100", -- t[8940] = 1
      "00001" when "010001011101101", -- t[8941] = 1
      "00001" when "010001011101110", -- t[8942] = 1
      "00001" when "010001011101111", -- t[8943] = 1
      "00001" when "010001011110000", -- t[8944] = 1
      "00001" when "010001011110001", -- t[8945] = 1
      "00001" when "010001011110010", -- t[8946] = 1
      "00001" when "010001011110011", -- t[8947] = 1
      "00001" when "010001011110100", -- t[8948] = 1
      "00001" when "010001011110101", -- t[8949] = 1
      "00001" when "010001011110110", -- t[8950] = 1
      "00001" when "010001011110111", -- t[8951] = 1
      "00001" when "010001011111000", -- t[8952] = 1
      "00001" when "010001011111001", -- t[8953] = 1
      "00001" when "010001011111010", -- t[8954] = 1
      "00001" when "010001011111011", -- t[8955] = 1
      "00001" when "010001011111100", -- t[8956] = 1
      "00001" when "010001011111101", -- t[8957] = 1
      "00001" when "010001011111110", -- t[8958] = 1
      "00001" when "010001011111111", -- t[8959] = 1
      "00001" when "010001100000000", -- t[8960] = 1
      "00001" when "010001100000001", -- t[8961] = 1
      "00001" when "010001100000010", -- t[8962] = 1
      "00001" when "010001100000011", -- t[8963] = 1
      "00001" when "010001100000100", -- t[8964] = 1
      "00001" when "010001100000101", -- t[8965] = 1
      "00001" when "010001100000110", -- t[8966] = 1
      "00001" when "010001100000111", -- t[8967] = 1
      "00001" when "010001100001000", -- t[8968] = 1
      "00001" when "010001100001001", -- t[8969] = 1
      "00001" when "010001100001010", -- t[8970] = 1
      "00001" when "010001100001011", -- t[8971] = 1
      "00001" when "010001100001100", -- t[8972] = 1
      "00001" when "010001100001101", -- t[8973] = 1
      "00001" when "010001100001110", -- t[8974] = 1
      "00001" when "010001100001111", -- t[8975] = 1
      "00001" when "010001100010000", -- t[8976] = 1
      "00001" when "010001100010001", -- t[8977] = 1
      "00001" when "010001100010010", -- t[8978] = 1
      "00001" when "010001100010011", -- t[8979] = 1
      "00001" when "010001100010100", -- t[8980] = 1
      "00001" when "010001100010101", -- t[8981] = 1
      "00001" when "010001100010110", -- t[8982] = 1
      "00001" when "010001100010111", -- t[8983] = 1
      "00001" when "010001100011000", -- t[8984] = 1
      "00001" when "010001100011001", -- t[8985] = 1
      "00001" when "010001100011010", -- t[8986] = 1
      "00001" when "010001100011011", -- t[8987] = 1
      "00001" when "010001100011100", -- t[8988] = 1
      "00001" when "010001100011101", -- t[8989] = 1
      "00001" when "010001100011110", -- t[8990] = 1
      "00001" when "010001100011111", -- t[8991] = 1
      "00001" when "010001100100000", -- t[8992] = 1
      "00001" when "010001100100001", -- t[8993] = 1
      "00001" when "010001100100010", -- t[8994] = 1
      "00001" when "010001100100011", -- t[8995] = 1
      "00001" when "010001100100100", -- t[8996] = 1
      "00001" when "010001100100101", -- t[8997] = 1
      "00001" when "010001100100110", -- t[8998] = 1
      "00001" when "010001100100111", -- t[8999] = 1
      "00001" when "010001100101000", -- t[9000] = 1
      "00001" when "010001100101001", -- t[9001] = 1
      "00001" when "010001100101010", -- t[9002] = 1
      "00001" when "010001100101011", -- t[9003] = 1
      "00001" when "010001100101100", -- t[9004] = 1
      "00001" when "010001100101101", -- t[9005] = 1
      "00001" when "010001100101110", -- t[9006] = 1
      "00001" when "010001100101111", -- t[9007] = 1
      "00001" when "010001100110000", -- t[9008] = 1
      "00001" when "010001100110001", -- t[9009] = 1
      "00001" when "010001100110010", -- t[9010] = 1
      "00001" when "010001100110011", -- t[9011] = 1
      "00001" when "010001100110100", -- t[9012] = 1
      "00001" when "010001100110101", -- t[9013] = 1
      "00001" when "010001100110110", -- t[9014] = 1
      "00001" when "010001100110111", -- t[9015] = 1
      "00001" when "010001100111000", -- t[9016] = 1
      "00001" when "010001100111001", -- t[9017] = 1
      "00001" when "010001100111010", -- t[9018] = 1
      "00001" when "010001100111011", -- t[9019] = 1
      "00001" when "010001100111100", -- t[9020] = 1
      "00001" when "010001100111101", -- t[9021] = 1
      "00001" when "010001100111110", -- t[9022] = 1
      "00001" when "010001100111111", -- t[9023] = 1
      "00001" when "010001101000000", -- t[9024] = 1
      "00001" when "010001101000001", -- t[9025] = 1
      "00001" when "010001101000010", -- t[9026] = 1
      "00001" when "010001101000011", -- t[9027] = 1
      "00001" when "010001101000100", -- t[9028] = 1
      "00001" when "010001101000101", -- t[9029] = 1
      "00001" when "010001101000110", -- t[9030] = 1
      "00001" when "010001101000111", -- t[9031] = 1
      "00001" when "010001101001000", -- t[9032] = 1
      "00001" when "010001101001001", -- t[9033] = 1
      "00001" when "010001101001010", -- t[9034] = 1
      "00001" when "010001101001011", -- t[9035] = 1
      "00001" when "010001101001100", -- t[9036] = 1
      "00001" when "010001101001101", -- t[9037] = 1
      "00001" when "010001101001110", -- t[9038] = 1
      "00001" when "010001101001111", -- t[9039] = 1
      "00001" when "010001101010000", -- t[9040] = 1
      "00001" when "010001101010001", -- t[9041] = 1
      "00001" when "010001101010010", -- t[9042] = 1
      "00001" when "010001101010011", -- t[9043] = 1
      "00001" when "010001101010100", -- t[9044] = 1
      "00001" when "010001101010101", -- t[9045] = 1
      "00001" when "010001101010110", -- t[9046] = 1
      "00001" when "010001101010111", -- t[9047] = 1
      "00001" when "010001101011000", -- t[9048] = 1
      "00001" when "010001101011001", -- t[9049] = 1
      "00001" when "010001101011010", -- t[9050] = 1
      "00001" when "010001101011011", -- t[9051] = 1
      "00001" when "010001101011100", -- t[9052] = 1
      "00001" when "010001101011101", -- t[9053] = 1
      "00001" when "010001101011110", -- t[9054] = 1
      "00001" when "010001101011111", -- t[9055] = 1
      "00001" when "010001101100000", -- t[9056] = 1
      "00001" when "010001101100001", -- t[9057] = 1
      "00001" when "010001101100010", -- t[9058] = 1
      "00001" when "010001101100011", -- t[9059] = 1
      "00001" when "010001101100100", -- t[9060] = 1
      "00001" when "010001101100101", -- t[9061] = 1
      "00001" when "010001101100110", -- t[9062] = 1
      "00001" when "010001101100111", -- t[9063] = 1
      "00001" when "010001101101000", -- t[9064] = 1
      "00001" when "010001101101001", -- t[9065] = 1
      "00001" when "010001101101010", -- t[9066] = 1
      "00001" when "010001101101011", -- t[9067] = 1
      "00001" when "010001101101100", -- t[9068] = 1
      "00001" when "010001101101101", -- t[9069] = 1
      "00001" when "010001101101110", -- t[9070] = 1
      "00001" when "010001101101111", -- t[9071] = 1
      "00001" when "010001101110000", -- t[9072] = 1
      "00001" when "010001101110001", -- t[9073] = 1
      "00001" when "010001101110010", -- t[9074] = 1
      "00001" when "010001101110011", -- t[9075] = 1
      "00001" when "010001101110100", -- t[9076] = 1
      "00001" when "010001101110101", -- t[9077] = 1
      "00001" when "010001101110110", -- t[9078] = 1
      "00001" when "010001101110111", -- t[9079] = 1
      "00001" when "010001101111000", -- t[9080] = 1
      "00001" when "010001101111001", -- t[9081] = 1
      "00001" when "010001101111010", -- t[9082] = 1
      "00001" when "010001101111011", -- t[9083] = 1
      "00001" when "010001101111100", -- t[9084] = 1
      "00001" when "010001101111101", -- t[9085] = 1
      "00001" when "010001101111110", -- t[9086] = 1
      "00001" when "010001101111111", -- t[9087] = 1
      "00001" when "010001110000000", -- t[9088] = 1
      "00001" when "010001110000001", -- t[9089] = 1
      "00001" when "010001110000010", -- t[9090] = 1
      "00001" when "010001110000011", -- t[9091] = 1
      "00001" when "010001110000100", -- t[9092] = 1
      "00001" when "010001110000101", -- t[9093] = 1
      "00001" when "010001110000110", -- t[9094] = 1
      "00001" when "010001110000111", -- t[9095] = 1
      "00001" when "010001110001000", -- t[9096] = 1
      "00001" when "010001110001001", -- t[9097] = 1
      "00001" when "010001110001010", -- t[9098] = 1
      "00001" when "010001110001011", -- t[9099] = 1
      "00001" when "010001110001100", -- t[9100] = 1
      "00001" when "010001110001101", -- t[9101] = 1
      "00001" when "010001110001110", -- t[9102] = 1
      "00001" when "010001110001111", -- t[9103] = 1
      "00001" when "010001110010000", -- t[9104] = 1
      "00001" when "010001110010001", -- t[9105] = 1
      "00001" when "010001110010010", -- t[9106] = 1
      "00001" when "010001110010011", -- t[9107] = 1
      "00001" when "010001110010100", -- t[9108] = 1
      "00001" when "010001110010101", -- t[9109] = 1
      "00001" when "010001110010110", -- t[9110] = 1
      "00001" when "010001110010111", -- t[9111] = 1
      "00001" when "010001110011000", -- t[9112] = 1
      "00001" when "010001110011001", -- t[9113] = 1
      "00001" when "010001110011010", -- t[9114] = 1
      "00001" when "010001110011011", -- t[9115] = 1
      "00001" when "010001110011100", -- t[9116] = 1
      "00001" when "010001110011101", -- t[9117] = 1
      "00001" when "010001110011110", -- t[9118] = 1
      "00001" when "010001110011111", -- t[9119] = 1
      "00001" when "010001110100000", -- t[9120] = 1
      "00001" when "010001110100001", -- t[9121] = 1
      "00001" when "010001110100010", -- t[9122] = 1
      "00001" when "010001110100011", -- t[9123] = 1
      "00001" when "010001110100100", -- t[9124] = 1
      "00001" when "010001110100101", -- t[9125] = 1
      "00001" when "010001110100110", -- t[9126] = 1
      "00001" when "010001110100111", -- t[9127] = 1
      "00001" when "010001110101000", -- t[9128] = 1
      "00001" when "010001110101001", -- t[9129] = 1
      "00001" when "010001110101010", -- t[9130] = 1
      "00001" when "010001110101011", -- t[9131] = 1
      "00001" when "010001110101100", -- t[9132] = 1
      "00001" when "010001110101101", -- t[9133] = 1
      "00001" when "010001110101110", -- t[9134] = 1
      "00001" when "010001110101111", -- t[9135] = 1
      "00001" when "010001110110000", -- t[9136] = 1
      "00001" when "010001110110001", -- t[9137] = 1
      "00001" when "010001110110010", -- t[9138] = 1
      "00001" when "010001110110011", -- t[9139] = 1
      "00001" when "010001110110100", -- t[9140] = 1
      "00001" when "010001110110101", -- t[9141] = 1
      "00001" when "010001110110110", -- t[9142] = 1
      "00001" when "010001110110111", -- t[9143] = 1
      "00001" when "010001110111000", -- t[9144] = 1
      "00001" when "010001110111001", -- t[9145] = 1
      "00001" when "010001110111010", -- t[9146] = 1
      "00001" when "010001110111011", -- t[9147] = 1
      "00001" when "010001110111100", -- t[9148] = 1
      "00001" when "010001110111101", -- t[9149] = 1
      "00001" when "010001110111110", -- t[9150] = 1
      "00001" when "010001110111111", -- t[9151] = 1
      "00001" when "010001111000000", -- t[9152] = 1
      "00001" when "010001111000001", -- t[9153] = 1
      "00001" when "010001111000010", -- t[9154] = 1
      "00001" when "010001111000011", -- t[9155] = 1
      "00001" when "010001111000100", -- t[9156] = 1
      "00001" when "010001111000101", -- t[9157] = 1
      "00001" when "010001111000110", -- t[9158] = 1
      "00001" when "010001111000111", -- t[9159] = 1
      "00001" when "010001111001000", -- t[9160] = 1
      "00001" when "010001111001001", -- t[9161] = 1
      "00001" when "010001111001010", -- t[9162] = 1
      "00001" when "010001111001011", -- t[9163] = 1
      "00001" when "010001111001100", -- t[9164] = 1
      "00001" when "010001111001101", -- t[9165] = 1
      "00001" when "010001111001110", -- t[9166] = 1
      "00001" when "010001111001111", -- t[9167] = 1
      "00001" when "010001111010000", -- t[9168] = 1
      "00001" when "010001111010001", -- t[9169] = 1
      "00001" when "010001111010010", -- t[9170] = 1
      "00001" when "010001111010011", -- t[9171] = 1
      "00001" when "010001111010100", -- t[9172] = 1
      "00001" when "010001111010101", -- t[9173] = 1
      "00001" when "010001111010110", -- t[9174] = 1
      "00001" when "010001111010111", -- t[9175] = 1
      "00001" when "010001111011000", -- t[9176] = 1
      "00001" when "010001111011001", -- t[9177] = 1
      "00001" when "010001111011010", -- t[9178] = 1
      "00001" when "010001111011011", -- t[9179] = 1
      "00001" when "010001111011100", -- t[9180] = 1
      "00001" when "010001111011101", -- t[9181] = 1
      "00001" when "010001111011110", -- t[9182] = 1
      "00001" when "010001111011111", -- t[9183] = 1
      "00001" when "010001111100000", -- t[9184] = 1
      "00001" when "010001111100001", -- t[9185] = 1
      "00001" when "010001111100010", -- t[9186] = 1
      "00001" when "010001111100011", -- t[9187] = 1
      "00001" when "010001111100100", -- t[9188] = 1
      "00001" when "010001111100101", -- t[9189] = 1
      "00001" when "010001111100110", -- t[9190] = 1
      "00001" when "010001111100111", -- t[9191] = 1
      "00001" when "010001111101000", -- t[9192] = 1
      "00001" when "010001111101001", -- t[9193] = 1
      "00001" when "010001111101010", -- t[9194] = 1
      "00001" when "010001111101011", -- t[9195] = 1
      "00001" when "010001111101100", -- t[9196] = 1
      "00001" when "010001111101101", -- t[9197] = 1
      "00001" when "010001111101110", -- t[9198] = 1
      "00001" when "010001111101111", -- t[9199] = 1
      "00001" when "010001111110000", -- t[9200] = 1
      "00001" when "010001111110001", -- t[9201] = 1
      "00001" when "010001111110010", -- t[9202] = 1
      "00001" when "010001111110011", -- t[9203] = 1
      "00001" when "010001111110100", -- t[9204] = 1
      "00001" when "010001111110101", -- t[9205] = 1
      "00001" when "010001111110110", -- t[9206] = 1
      "00001" when "010001111110111", -- t[9207] = 1
      "00001" when "010001111111000", -- t[9208] = 1
      "00001" when "010001111111001", -- t[9209] = 1
      "00001" when "010001111111010", -- t[9210] = 1
      "00001" when "010001111111011", -- t[9211] = 1
      "00001" when "010001111111100", -- t[9212] = 1
      "00001" when "010001111111101", -- t[9213] = 1
      "00001" when "010001111111110", -- t[9214] = 1
      "00001" when "010001111111111", -- t[9215] = 1
      "00001" when "010010000000000", -- t[9216] = 1
      "00001" when "010010000000001", -- t[9217] = 1
      "00001" when "010010000000010", -- t[9218] = 1
      "00001" when "010010000000011", -- t[9219] = 1
      "00001" when "010010000000100", -- t[9220] = 1
      "00001" when "010010000000101", -- t[9221] = 1
      "00001" when "010010000000110", -- t[9222] = 1
      "00001" when "010010000000111", -- t[9223] = 1
      "00001" when "010010000001000", -- t[9224] = 1
      "00001" when "010010000001001", -- t[9225] = 1
      "00001" when "010010000001010", -- t[9226] = 1
      "00001" when "010010000001011", -- t[9227] = 1
      "00001" when "010010000001100", -- t[9228] = 1
      "00001" when "010010000001101", -- t[9229] = 1
      "00001" when "010010000001110", -- t[9230] = 1
      "00001" when "010010000001111", -- t[9231] = 1
      "00001" when "010010000010000", -- t[9232] = 1
      "00001" when "010010000010001", -- t[9233] = 1
      "00001" when "010010000010010", -- t[9234] = 1
      "00001" when "010010000010011", -- t[9235] = 1
      "00001" when "010010000010100", -- t[9236] = 1
      "00001" when "010010000010101", -- t[9237] = 1
      "00001" when "010010000010110", -- t[9238] = 1
      "00001" when "010010000010111", -- t[9239] = 1
      "00001" when "010010000011000", -- t[9240] = 1
      "00001" when "010010000011001", -- t[9241] = 1
      "00001" when "010010000011010", -- t[9242] = 1
      "00001" when "010010000011011", -- t[9243] = 1
      "00001" when "010010000011100", -- t[9244] = 1
      "00001" when "010010000011101", -- t[9245] = 1
      "00001" when "010010000011110", -- t[9246] = 1
      "00001" when "010010000011111", -- t[9247] = 1
      "00001" when "010010000100000", -- t[9248] = 1
      "00001" when "010010000100001", -- t[9249] = 1
      "00001" when "010010000100010", -- t[9250] = 1
      "00001" when "010010000100011", -- t[9251] = 1
      "00001" when "010010000100100", -- t[9252] = 1
      "00001" when "010010000100101", -- t[9253] = 1
      "00001" when "010010000100110", -- t[9254] = 1
      "00001" when "010010000100111", -- t[9255] = 1
      "00001" when "010010000101000", -- t[9256] = 1
      "00001" when "010010000101001", -- t[9257] = 1
      "00001" when "010010000101010", -- t[9258] = 1
      "00001" when "010010000101011", -- t[9259] = 1
      "00001" when "010010000101100", -- t[9260] = 1
      "00001" when "010010000101101", -- t[9261] = 1
      "00001" when "010010000101110", -- t[9262] = 1
      "00001" when "010010000101111", -- t[9263] = 1
      "00001" when "010010000110000", -- t[9264] = 1
      "00001" when "010010000110001", -- t[9265] = 1
      "00001" when "010010000110010", -- t[9266] = 1
      "00001" when "010010000110011", -- t[9267] = 1
      "00001" when "010010000110100", -- t[9268] = 1
      "00001" when "010010000110101", -- t[9269] = 1
      "00001" when "010010000110110", -- t[9270] = 1
      "00001" when "010010000110111", -- t[9271] = 1
      "00001" when "010010000111000", -- t[9272] = 1
      "00001" when "010010000111001", -- t[9273] = 1
      "00001" when "010010000111010", -- t[9274] = 1
      "00001" when "010010000111011", -- t[9275] = 1
      "00001" when "010010000111100", -- t[9276] = 1
      "00001" when "010010000111101", -- t[9277] = 1
      "00001" when "010010000111110", -- t[9278] = 1
      "00001" when "010010000111111", -- t[9279] = 1
      "00001" when "010010001000000", -- t[9280] = 1
      "00001" when "010010001000001", -- t[9281] = 1
      "00001" when "010010001000010", -- t[9282] = 1
      "00001" when "010010001000011", -- t[9283] = 1
      "00001" when "010010001000100", -- t[9284] = 1
      "00001" when "010010001000101", -- t[9285] = 1
      "00001" when "010010001000110", -- t[9286] = 1
      "00001" when "010010001000111", -- t[9287] = 1
      "00001" when "010010001001000", -- t[9288] = 1
      "00001" when "010010001001001", -- t[9289] = 1
      "00001" when "010010001001010", -- t[9290] = 1
      "00001" when "010010001001011", -- t[9291] = 1
      "00001" when "010010001001100", -- t[9292] = 1
      "00001" when "010010001001101", -- t[9293] = 1
      "00001" when "010010001001110", -- t[9294] = 1
      "00001" when "010010001001111", -- t[9295] = 1
      "00001" when "010010001010000", -- t[9296] = 1
      "00001" when "010010001010001", -- t[9297] = 1
      "00001" when "010010001010010", -- t[9298] = 1
      "00001" when "010010001010011", -- t[9299] = 1
      "00001" when "010010001010100", -- t[9300] = 1
      "00001" when "010010001010101", -- t[9301] = 1
      "00001" when "010010001010110", -- t[9302] = 1
      "00001" when "010010001010111", -- t[9303] = 1
      "00001" when "010010001011000", -- t[9304] = 1
      "00001" when "010010001011001", -- t[9305] = 1
      "00001" when "010010001011010", -- t[9306] = 1
      "00001" when "010010001011011", -- t[9307] = 1
      "00001" when "010010001011100", -- t[9308] = 1
      "00001" when "010010001011101", -- t[9309] = 1
      "00001" when "010010001011110", -- t[9310] = 1
      "00001" when "010010001011111", -- t[9311] = 1
      "00001" when "010010001100000", -- t[9312] = 1
      "00001" when "010010001100001", -- t[9313] = 1
      "00001" when "010010001100010", -- t[9314] = 1
      "00001" when "010010001100011", -- t[9315] = 1
      "00001" when "010010001100100", -- t[9316] = 1
      "00001" when "010010001100101", -- t[9317] = 1
      "00001" when "010010001100110", -- t[9318] = 1
      "00001" when "010010001100111", -- t[9319] = 1
      "00001" when "010010001101000", -- t[9320] = 1
      "00001" when "010010001101001", -- t[9321] = 1
      "00001" when "010010001101010", -- t[9322] = 1
      "00001" when "010010001101011", -- t[9323] = 1
      "00001" when "010010001101100", -- t[9324] = 1
      "00001" when "010010001101101", -- t[9325] = 1
      "00001" when "010010001101110", -- t[9326] = 1
      "00001" when "010010001101111", -- t[9327] = 1
      "00001" when "010010001110000", -- t[9328] = 1
      "00001" when "010010001110001", -- t[9329] = 1
      "00001" when "010010001110010", -- t[9330] = 1
      "00001" when "010010001110011", -- t[9331] = 1
      "00001" when "010010001110100", -- t[9332] = 1
      "00001" when "010010001110101", -- t[9333] = 1
      "00001" when "010010001110110", -- t[9334] = 1
      "00001" when "010010001110111", -- t[9335] = 1
      "00001" when "010010001111000", -- t[9336] = 1
      "00001" when "010010001111001", -- t[9337] = 1
      "00001" when "010010001111010", -- t[9338] = 1
      "00001" when "010010001111011", -- t[9339] = 1
      "00001" when "010010001111100", -- t[9340] = 1
      "00001" when "010010001111101", -- t[9341] = 1
      "00001" when "010010001111110", -- t[9342] = 1
      "00001" when "010010001111111", -- t[9343] = 1
      "00001" when "010010010000000", -- t[9344] = 1
      "00001" when "010010010000001", -- t[9345] = 1
      "00001" when "010010010000010", -- t[9346] = 1
      "00001" when "010010010000011", -- t[9347] = 1
      "00001" when "010010010000100", -- t[9348] = 1
      "00001" when "010010010000101", -- t[9349] = 1
      "00001" when "010010010000110", -- t[9350] = 1
      "00001" when "010010010000111", -- t[9351] = 1
      "00001" when "010010010001000", -- t[9352] = 1
      "00001" when "010010010001001", -- t[9353] = 1
      "00001" when "010010010001010", -- t[9354] = 1
      "00001" when "010010010001011", -- t[9355] = 1
      "00001" when "010010010001100", -- t[9356] = 1
      "00001" when "010010010001101", -- t[9357] = 1
      "00001" when "010010010001110", -- t[9358] = 1
      "00001" when "010010010001111", -- t[9359] = 1
      "00001" when "010010010010000", -- t[9360] = 1
      "00001" when "010010010010001", -- t[9361] = 1
      "00001" when "010010010010010", -- t[9362] = 1
      "00001" when "010010010010011", -- t[9363] = 1
      "00001" when "010010010010100", -- t[9364] = 1
      "00001" when "010010010010101", -- t[9365] = 1
      "00001" when "010010010010110", -- t[9366] = 1
      "00001" when "010010010010111", -- t[9367] = 1
      "00001" when "010010010011000", -- t[9368] = 1
      "00001" when "010010010011001", -- t[9369] = 1
      "00001" when "010010010011010", -- t[9370] = 1
      "00001" when "010010010011011", -- t[9371] = 1
      "00001" when "010010010011100", -- t[9372] = 1
      "00001" when "010010010011101", -- t[9373] = 1
      "00001" when "010010010011110", -- t[9374] = 1
      "00001" when "010010010011111", -- t[9375] = 1
      "00001" when "010010010100000", -- t[9376] = 1
      "00001" when "010010010100001", -- t[9377] = 1
      "00001" when "010010010100010", -- t[9378] = 1
      "00001" when "010010010100011", -- t[9379] = 1
      "00001" when "010010010100100", -- t[9380] = 1
      "00001" when "010010010100101", -- t[9381] = 1
      "00001" when "010010010100110", -- t[9382] = 1
      "00001" when "010010010100111", -- t[9383] = 1
      "00001" when "010010010101000", -- t[9384] = 1
      "00001" when "010010010101001", -- t[9385] = 1
      "00001" when "010010010101010", -- t[9386] = 1
      "00001" when "010010010101011", -- t[9387] = 1
      "00001" when "010010010101100", -- t[9388] = 1
      "00001" when "010010010101101", -- t[9389] = 1
      "00001" when "010010010101110", -- t[9390] = 1
      "00001" when "010010010101111", -- t[9391] = 1
      "00001" when "010010010110000", -- t[9392] = 1
      "00001" when "010010010110001", -- t[9393] = 1
      "00001" when "010010010110010", -- t[9394] = 1
      "00001" when "010010010110011", -- t[9395] = 1
      "00001" when "010010010110100", -- t[9396] = 1
      "00001" when "010010010110101", -- t[9397] = 1
      "00001" when "010010010110110", -- t[9398] = 1
      "00001" when "010010010110111", -- t[9399] = 1
      "00001" when "010010010111000", -- t[9400] = 1
      "00001" when "010010010111001", -- t[9401] = 1
      "00001" when "010010010111010", -- t[9402] = 1
      "00001" when "010010010111011", -- t[9403] = 1
      "00001" when "010010010111100", -- t[9404] = 1
      "00001" when "010010010111101", -- t[9405] = 1
      "00001" when "010010010111110", -- t[9406] = 1
      "00001" when "010010010111111", -- t[9407] = 1
      "00001" when "010010011000000", -- t[9408] = 1
      "00001" when "010010011000001", -- t[9409] = 1
      "00001" when "010010011000010", -- t[9410] = 1
      "00001" when "010010011000011", -- t[9411] = 1
      "00001" when "010010011000100", -- t[9412] = 1
      "00001" when "010010011000101", -- t[9413] = 1
      "00001" when "010010011000110", -- t[9414] = 1
      "00001" when "010010011000111", -- t[9415] = 1
      "00001" when "010010011001000", -- t[9416] = 1
      "00001" when "010010011001001", -- t[9417] = 1
      "00001" when "010010011001010", -- t[9418] = 1
      "00001" when "010010011001011", -- t[9419] = 1
      "00001" when "010010011001100", -- t[9420] = 1
      "00001" when "010010011001101", -- t[9421] = 1
      "00001" when "010010011001110", -- t[9422] = 1
      "00001" when "010010011001111", -- t[9423] = 1
      "00001" when "010010011010000", -- t[9424] = 1
      "00001" when "010010011010001", -- t[9425] = 1
      "00001" when "010010011010010", -- t[9426] = 1
      "00001" when "010010011010011", -- t[9427] = 1
      "00001" when "010010011010100", -- t[9428] = 1
      "00001" when "010010011010101", -- t[9429] = 1
      "00001" when "010010011010110", -- t[9430] = 1
      "00001" when "010010011010111", -- t[9431] = 1
      "00001" when "010010011011000", -- t[9432] = 1
      "00001" when "010010011011001", -- t[9433] = 1
      "00001" when "010010011011010", -- t[9434] = 1
      "00001" when "010010011011011", -- t[9435] = 1
      "00001" when "010010011011100", -- t[9436] = 1
      "00001" when "010010011011101", -- t[9437] = 1
      "00001" when "010010011011110", -- t[9438] = 1
      "00001" when "010010011011111", -- t[9439] = 1
      "00001" when "010010011100000", -- t[9440] = 1
      "00001" when "010010011100001", -- t[9441] = 1
      "00001" when "010010011100010", -- t[9442] = 1
      "00001" when "010010011100011", -- t[9443] = 1
      "00001" when "010010011100100", -- t[9444] = 1
      "00001" when "010010011100101", -- t[9445] = 1
      "00001" when "010010011100110", -- t[9446] = 1
      "00001" when "010010011100111", -- t[9447] = 1
      "00001" when "010010011101000", -- t[9448] = 1
      "00001" when "010010011101001", -- t[9449] = 1
      "00001" when "010010011101010", -- t[9450] = 1
      "00001" when "010010011101011", -- t[9451] = 1
      "00001" when "010010011101100", -- t[9452] = 1
      "00001" when "010010011101101", -- t[9453] = 1
      "00001" when "010010011101110", -- t[9454] = 1
      "00001" when "010010011101111", -- t[9455] = 1
      "00001" when "010010011110000", -- t[9456] = 1
      "00001" when "010010011110001", -- t[9457] = 1
      "00001" when "010010011110010", -- t[9458] = 1
      "00001" when "010010011110011", -- t[9459] = 1
      "00001" when "010010011110100", -- t[9460] = 1
      "00001" when "010010011110101", -- t[9461] = 1
      "00001" when "010010011110110", -- t[9462] = 1
      "00001" when "010010011110111", -- t[9463] = 1
      "00001" when "010010011111000", -- t[9464] = 1
      "00001" when "010010011111001", -- t[9465] = 1
      "00001" when "010010011111010", -- t[9466] = 1
      "00001" when "010010011111011", -- t[9467] = 1
      "00001" when "010010011111100", -- t[9468] = 1
      "00001" when "010010011111101", -- t[9469] = 1
      "00001" when "010010011111110", -- t[9470] = 1
      "00001" when "010010011111111", -- t[9471] = 1
      "00001" when "010010100000000", -- t[9472] = 1
      "00001" when "010010100000001", -- t[9473] = 1
      "00001" when "010010100000010", -- t[9474] = 1
      "00001" when "010010100000011", -- t[9475] = 1
      "00001" when "010010100000100", -- t[9476] = 1
      "00001" when "010010100000101", -- t[9477] = 1
      "00001" when "010010100000110", -- t[9478] = 1
      "00001" when "010010100000111", -- t[9479] = 1
      "00001" when "010010100001000", -- t[9480] = 1
      "00001" when "010010100001001", -- t[9481] = 1
      "00001" when "010010100001010", -- t[9482] = 1
      "00001" when "010010100001011", -- t[9483] = 1
      "00001" when "010010100001100", -- t[9484] = 1
      "00001" when "010010100001101", -- t[9485] = 1
      "00001" when "010010100001110", -- t[9486] = 1
      "00001" when "010010100001111", -- t[9487] = 1
      "00001" when "010010100010000", -- t[9488] = 1
      "00001" when "010010100010001", -- t[9489] = 1
      "00001" when "010010100010010", -- t[9490] = 1
      "00001" when "010010100010011", -- t[9491] = 1
      "00001" when "010010100010100", -- t[9492] = 1
      "00001" when "010010100010101", -- t[9493] = 1
      "00001" when "010010100010110", -- t[9494] = 1
      "00001" when "010010100010111", -- t[9495] = 1
      "00001" when "010010100011000", -- t[9496] = 1
      "00001" when "010010100011001", -- t[9497] = 1
      "00001" when "010010100011010", -- t[9498] = 1
      "00001" when "010010100011011", -- t[9499] = 1
      "00001" when "010010100011100", -- t[9500] = 1
      "00001" when "010010100011101", -- t[9501] = 1
      "00001" when "010010100011110", -- t[9502] = 1
      "00001" when "010010100011111", -- t[9503] = 1
      "00001" when "010010100100000", -- t[9504] = 1
      "00001" when "010010100100001", -- t[9505] = 1
      "00001" when "010010100100010", -- t[9506] = 1
      "00001" when "010010100100011", -- t[9507] = 1
      "00001" when "010010100100100", -- t[9508] = 1
      "00001" when "010010100100101", -- t[9509] = 1
      "00001" when "010010100100110", -- t[9510] = 1
      "00001" when "010010100100111", -- t[9511] = 1
      "00001" when "010010100101000", -- t[9512] = 1
      "00001" when "010010100101001", -- t[9513] = 1
      "00001" when "010010100101010", -- t[9514] = 1
      "00001" when "010010100101011", -- t[9515] = 1
      "00001" when "010010100101100", -- t[9516] = 1
      "00001" when "010010100101101", -- t[9517] = 1
      "00001" when "010010100101110", -- t[9518] = 1
      "00001" when "010010100101111", -- t[9519] = 1
      "00001" when "010010100110000", -- t[9520] = 1
      "00001" when "010010100110001", -- t[9521] = 1
      "00001" when "010010100110010", -- t[9522] = 1
      "00001" when "010010100110011", -- t[9523] = 1
      "00001" when "010010100110100", -- t[9524] = 1
      "00001" when "010010100110101", -- t[9525] = 1
      "00001" when "010010100110110", -- t[9526] = 1
      "00001" when "010010100110111", -- t[9527] = 1
      "00001" when "010010100111000", -- t[9528] = 1
      "00001" when "010010100111001", -- t[9529] = 1
      "00001" when "010010100111010", -- t[9530] = 1
      "00001" when "010010100111011", -- t[9531] = 1
      "00001" when "010010100111100", -- t[9532] = 1
      "00001" when "010010100111101", -- t[9533] = 1
      "00001" when "010010100111110", -- t[9534] = 1
      "00001" when "010010100111111", -- t[9535] = 1
      "00001" when "010010101000000", -- t[9536] = 1
      "00001" when "010010101000001", -- t[9537] = 1
      "00001" when "010010101000010", -- t[9538] = 1
      "00001" when "010010101000011", -- t[9539] = 1
      "00001" when "010010101000100", -- t[9540] = 1
      "00001" when "010010101000101", -- t[9541] = 1
      "00001" when "010010101000110", -- t[9542] = 1
      "00001" when "010010101000111", -- t[9543] = 1
      "00001" when "010010101001000", -- t[9544] = 1
      "00001" when "010010101001001", -- t[9545] = 1
      "00001" when "010010101001010", -- t[9546] = 1
      "00001" when "010010101001011", -- t[9547] = 1
      "00001" when "010010101001100", -- t[9548] = 1
      "00001" when "010010101001101", -- t[9549] = 1
      "00001" when "010010101001110", -- t[9550] = 1
      "00001" when "010010101001111", -- t[9551] = 1
      "00001" when "010010101010000", -- t[9552] = 1
      "00001" when "010010101010001", -- t[9553] = 1
      "00001" when "010010101010010", -- t[9554] = 1
      "00001" when "010010101010011", -- t[9555] = 1
      "00001" when "010010101010100", -- t[9556] = 1
      "00001" when "010010101010101", -- t[9557] = 1
      "00001" when "010010101010110", -- t[9558] = 1
      "00001" when "010010101010111", -- t[9559] = 1
      "00001" when "010010101011000", -- t[9560] = 1
      "00001" when "010010101011001", -- t[9561] = 1
      "00001" when "010010101011010", -- t[9562] = 1
      "00001" when "010010101011011", -- t[9563] = 1
      "00001" when "010010101011100", -- t[9564] = 1
      "00001" when "010010101011101", -- t[9565] = 1
      "00001" when "010010101011110", -- t[9566] = 1
      "00001" when "010010101011111", -- t[9567] = 1
      "00001" when "010010101100000", -- t[9568] = 1
      "00001" when "010010101100001", -- t[9569] = 1
      "00001" when "010010101100010", -- t[9570] = 1
      "00001" when "010010101100011", -- t[9571] = 1
      "00001" when "010010101100100", -- t[9572] = 1
      "00001" when "010010101100101", -- t[9573] = 1
      "00001" when "010010101100110", -- t[9574] = 1
      "00001" when "010010101100111", -- t[9575] = 1
      "00001" when "010010101101000", -- t[9576] = 1
      "00001" when "010010101101001", -- t[9577] = 1
      "00001" when "010010101101010", -- t[9578] = 1
      "00001" when "010010101101011", -- t[9579] = 1
      "00001" when "010010101101100", -- t[9580] = 1
      "00001" when "010010101101101", -- t[9581] = 1
      "00001" when "010010101101110", -- t[9582] = 1
      "00001" when "010010101101111", -- t[9583] = 1
      "00001" when "010010101110000", -- t[9584] = 1
      "00001" when "010010101110001", -- t[9585] = 1
      "00001" when "010010101110010", -- t[9586] = 1
      "00001" when "010010101110011", -- t[9587] = 1
      "00001" when "010010101110100", -- t[9588] = 1
      "00001" when "010010101110101", -- t[9589] = 1
      "00001" when "010010101110110", -- t[9590] = 1
      "00001" when "010010101110111", -- t[9591] = 1
      "00001" when "010010101111000", -- t[9592] = 1
      "00001" when "010010101111001", -- t[9593] = 1
      "00001" when "010010101111010", -- t[9594] = 1
      "00001" when "010010101111011", -- t[9595] = 1
      "00001" when "010010101111100", -- t[9596] = 1
      "00001" when "010010101111101", -- t[9597] = 1
      "00001" when "010010101111110", -- t[9598] = 1
      "00001" when "010010101111111", -- t[9599] = 1
      "00001" when "010010110000000", -- t[9600] = 1
      "00001" when "010010110000001", -- t[9601] = 1
      "00001" when "010010110000010", -- t[9602] = 1
      "00001" when "010010110000011", -- t[9603] = 1
      "00001" when "010010110000100", -- t[9604] = 1
      "00001" when "010010110000101", -- t[9605] = 1
      "00001" when "010010110000110", -- t[9606] = 1
      "00001" when "010010110000111", -- t[9607] = 1
      "00001" when "010010110001000", -- t[9608] = 1
      "00001" when "010010110001001", -- t[9609] = 1
      "00001" when "010010110001010", -- t[9610] = 1
      "00001" when "010010110001011", -- t[9611] = 1
      "00001" when "010010110001100", -- t[9612] = 1
      "00001" when "010010110001101", -- t[9613] = 1
      "00001" when "010010110001110", -- t[9614] = 1
      "00001" when "010010110001111", -- t[9615] = 1
      "00001" when "010010110010000", -- t[9616] = 1
      "00001" when "010010110010001", -- t[9617] = 1
      "00001" when "010010110010010", -- t[9618] = 1
      "00001" when "010010110010011", -- t[9619] = 1
      "00001" when "010010110010100", -- t[9620] = 1
      "00001" when "010010110010101", -- t[9621] = 1
      "00001" when "010010110010110", -- t[9622] = 1
      "00001" when "010010110010111", -- t[9623] = 1
      "00001" when "010010110011000", -- t[9624] = 1
      "00001" when "010010110011001", -- t[9625] = 1
      "00001" when "010010110011010", -- t[9626] = 1
      "00001" when "010010110011011", -- t[9627] = 1
      "00001" when "010010110011100", -- t[9628] = 1
      "00001" when "010010110011101", -- t[9629] = 1
      "00001" when "010010110011110", -- t[9630] = 1
      "00001" when "010010110011111", -- t[9631] = 1
      "00001" when "010010110100000", -- t[9632] = 1
      "00001" when "010010110100001", -- t[9633] = 1
      "00001" when "010010110100010", -- t[9634] = 1
      "00001" when "010010110100011", -- t[9635] = 1
      "00001" when "010010110100100", -- t[9636] = 1
      "00001" when "010010110100101", -- t[9637] = 1
      "00001" when "010010110100110", -- t[9638] = 1
      "00001" when "010010110100111", -- t[9639] = 1
      "00001" when "010010110101000", -- t[9640] = 1
      "00001" when "010010110101001", -- t[9641] = 1
      "00001" when "010010110101010", -- t[9642] = 1
      "00001" when "010010110101011", -- t[9643] = 1
      "00001" when "010010110101100", -- t[9644] = 1
      "00001" when "010010110101101", -- t[9645] = 1
      "00001" when "010010110101110", -- t[9646] = 1
      "00001" when "010010110101111", -- t[9647] = 1
      "00001" when "010010110110000", -- t[9648] = 1
      "00001" when "010010110110001", -- t[9649] = 1
      "00001" when "010010110110010", -- t[9650] = 1
      "00001" when "010010110110011", -- t[9651] = 1
      "00001" when "010010110110100", -- t[9652] = 1
      "00001" when "010010110110101", -- t[9653] = 1
      "00001" when "010010110110110", -- t[9654] = 1
      "00001" when "010010110110111", -- t[9655] = 1
      "00001" when "010010110111000", -- t[9656] = 1
      "00001" when "010010110111001", -- t[9657] = 1
      "00001" when "010010110111010", -- t[9658] = 1
      "00001" when "010010110111011", -- t[9659] = 1
      "00001" when "010010110111100", -- t[9660] = 1
      "00001" when "010010110111101", -- t[9661] = 1
      "00001" when "010010110111110", -- t[9662] = 1
      "00001" when "010010110111111", -- t[9663] = 1
      "00001" when "010010111000000", -- t[9664] = 1
      "00001" when "010010111000001", -- t[9665] = 1
      "00001" when "010010111000010", -- t[9666] = 1
      "00001" when "010010111000011", -- t[9667] = 1
      "00001" when "010010111000100", -- t[9668] = 1
      "00001" when "010010111000101", -- t[9669] = 1
      "00001" when "010010111000110", -- t[9670] = 1
      "00001" when "010010111000111", -- t[9671] = 1
      "00001" when "010010111001000", -- t[9672] = 1
      "00001" when "010010111001001", -- t[9673] = 1
      "00001" when "010010111001010", -- t[9674] = 1
      "00001" when "010010111001011", -- t[9675] = 1
      "00001" when "010010111001100", -- t[9676] = 1
      "00001" when "010010111001101", -- t[9677] = 1
      "00001" when "010010111001110", -- t[9678] = 1
      "00001" when "010010111001111", -- t[9679] = 1
      "00001" when "010010111010000", -- t[9680] = 1
      "00001" when "010010111010001", -- t[9681] = 1
      "00001" when "010010111010010", -- t[9682] = 1
      "00001" when "010010111010011", -- t[9683] = 1
      "00001" when "010010111010100", -- t[9684] = 1
      "00001" when "010010111010101", -- t[9685] = 1
      "00001" when "010010111010110", -- t[9686] = 1
      "00001" when "010010111010111", -- t[9687] = 1
      "00001" when "010010111011000", -- t[9688] = 1
      "00001" when "010010111011001", -- t[9689] = 1
      "00001" when "010010111011010", -- t[9690] = 1
      "00001" when "010010111011011", -- t[9691] = 1
      "00001" when "010010111011100", -- t[9692] = 1
      "00001" when "010010111011101", -- t[9693] = 1
      "00001" when "010010111011110", -- t[9694] = 1
      "00001" when "010010111011111", -- t[9695] = 1
      "00001" when "010010111100000", -- t[9696] = 1
      "00001" when "010010111100001", -- t[9697] = 1
      "00001" when "010010111100010", -- t[9698] = 1
      "00001" when "010010111100011", -- t[9699] = 1
      "00001" when "010010111100100", -- t[9700] = 1
      "00001" when "010010111100101", -- t[9701] = 1
      "00001" when "010010111100110", -- t[9702] = 1
      "00001" when "010010111100111", -- t[9703] = 1
      "00001" when "010010111101000", -- t[9704] = 1
      "00001" when "010010111101001", -- t[9705] = 1
      "00001" when "010010111101010", -- t[9706] = 1
      "00001" when "010010111101011", -- t[9707] = 1
      "00001" when "010010111101100", -- t[9708] = 1
      "00001" when "010010111101101", -- t[9709] = 1
      "00001" when "010010111101110", -- t[9710] = 1
      "00001" when "010010111101111", -- t[9711] = 1
      "00001" when "010010111110000", -- t[9712] = 1
      "00001" when "010010111110001", -- t[9713] = 1
      "00001" when "010010111110010", -- t[9714] = 1
      "00001" when "010010111110011", -- t[9715] = 1
      "00001" when "010010111110100", -- t[9716] = 1
      "00001" when "010010111110101", -- t[9717] = 1
      "00001" when "010010111110110", -- t[9718] = 1
      "00001" when "010010111110111", -- t[9719] = 1
      "00001" when "010010111111000", -- t[9720] = 1
      "00001" when "010010111111001", -- t[9721] = 1
      "00001" when "010010111111010", -- t[9722] = 1
      "00001" when "010010111111011", -- t[9723] = 1
      "00001" when "010010111111100", -- t[9724] = 1
      "00001" when "010010111111101", -- t[9725] = 1
      "00001" when "010010111111110", -- t[9726] = 1
      "00001" when "010010111111111", -- t[9727] = 1
      "00001" when "010011000000000", -- t[9728] = 1
      "00001" when "010011000000001", -- t[9729] = 1
      "00001" when "010011000000010", -- t[9730] = 1
      "00001" when "010011000000011", -- t[9731] = 1
      "00001" when "010011000000100", -- t[9732] = 1
      "00001" when "010011000000101", -- t[9733] = 1
      "00001" when "010011000000110", -- t[9734] = 1
      "00001" when "010011000000111", -- t[9735] = 1
      "00001" when "010011000001000", -- t[9736] = 1
      "00001" when "010011000001001", -- t[9737] = 1
      "00001" when "010011000001010", -- t[9738] = 1
      "00001" when "010011000001011", -- t[9739] = 1
      "00001" when "010011000001100", -- t[9740] = 1
      "00001" when "010011000001101", -- t[9741] = 1
      "00001" when "010011000001110", -- t[9742] = 1
      "00001" when "010011000001111", -- t[9743] = 1
      "00001" when "010011000010000", -- t[9744] = 1
      "00001" when "010011000010001", -- t[9745] = 1
      "00001" when "010011000010010", -- t[9746] = 1
      "00001" when "010011000010011", -- t[9747] = 1
      "00001" when "010011000010100", -- t[9748] = 1
      "00001" when "010011000010101", -- t[9749] = 1
      "00001" when "010011000010110", -- t[9750] = 1
      "00001" when "010011000010111", -- t[9751] = 1
      "00001" when "010011000011000", -- t[9752] = 1
      "00001" when "010011000011001", -- t[9753] = 1
      "00001" when "010011000011010", -- t[9754] = 1
      "00001" when "010011000011011", -- t[9755] = 1
      "00001" when "010011000011100", -- t[9756] = 1
      "00001" when "010011000011101", -- t[9757] = 1
      "00001" when "010011000011110", -- t[9758] = 1
      "00001" when "010011000011111", -- t[9759] = 1
      "00001" when "010011000100000", -- t[9760] = 1
      "00001" when "010011000100001", -- t[9761] = 1
      "00001" when "010011000100010", -- t[9762] = 1
      "00001" when "010011000100011", -- t[9763] = 1
      "00001" when "010011000100100", -- t[9764] = 1
      "00001" when "010011000100101", -- t[9765] = 1
      "00001" when "010011000100110", -- t[9766] = 1
      "00001" when "010011000100111", -- t[9767] = 1
      "00001" when "010011000101000", -- t[9768] = 1
      "00001" when "010011000101001", -- t[9769] = 1
      "00001" when "010011000101010", -- t[9770] = 1
      "00001" when "010011000101011", -- t[9771] = 1
      "00001" when "010011000101100", -- t[9772] = 1
      "00001" when "010011000101101", -- t[9773] = 1
      "00001" when "010011000101110", -- t[9774] = 1
      "00001" when "010011000101111", -- t[9775] = 1
      "00001" when "010011000110000", -- t[9776] = 1
      "00001" when "010011000110001", -- t[9777] = 1
      "00001" when "010011000110010", -- t[9778] = 1
      "00001" when "010011000110011", -- t[9779] = 1
      "00001" when "010011000110100", -- t[9780] = 1
      "00001" when "010011000110101", -- t[9781] = 1
      "00001" when "010011000110110", -- t[9782] = 1
      "00001" when "010011000110111", -- t[9783] = 1
      "00001" when "010011000111000", -- t[9784] = 1
      "00001" when "010011000111001", -- t[9785] = 1
      "00001" when "010011000111010", -- t[9786] = 1
      "00001" when "010011000111011", -- t[9787] = 1
      "00001" when "010011000111100", -- t[9788] = 1
      "00001" when "010011000111101", -- t[9789] = 1
      "00001" when "010011000111110", -- t[9790] = 1
      "00001" when "010011000111111", -- t[9791] = 1
      "00001" when "010011001000000", -- t[9792] = 1
      "00001" when "010011001000001", -- t[9793] = 1
      "00001" when "010011001000010", -- t[9794] = 1
      "00001" when "010011001000011", -- t[9795] = 1
      "00001" when "010011001000100", -- t[9796] = 1
      "00001" when "010011001000101", -- t[9797] = 1
      "00001" when "010011001000110", -- t[9798] = 1
      "00001" when "010011001000111", -- t[9799] = 1
      "00001" when "010011001001000", -- t[9800] = 1
      "00001" when "010011001001001", -- t[9801] = 1
      "00001" when "010011001001010", -- t[9802] = 1
      "00001" when "010011001001011", -- t[9803] = 1
      "00001" when "010011001001100", -- t[9804] = 1
      "00001" when "010011001001101", -- t[9805] = 1
      "00001" when "010011001001110", -- t[9806] = 1
      "00001" when "010011001001111", -- t[9807] = 1
      "00001" when "010011001010000", -- t[9808] = 1
      "00001" when "010011001010001", -- t[9809] = 1
      "00001" when "010011001010010", -- t[9810] = 1
      "00001" when "010011001010011", -- t[9811] = 1
      "00001" when "010011001010100", -- t[9812] = 1
      "00001" when "010011001010101", -- t[9813] = 1
      "00001" when "010011001010110", -- t[9814] = 1
      "00001" when "010011001010111", -- t[9815] = 1
      "00001" when "010011001011000", -- t[9816] = 1
      "00001" when "010011001011001", -- t[9817] = 1
      "00001" when "010011001011010", -- t[9818] = 1
      "00001" when "010011001011011", -- t[9819] = 1
      "00001" when "010011001011100", -- t[9820] = 1
      "00001" when "010011001011101", -- t[9821] = 1
      "00001" when "010011001011110", -- t[9822] = 1
      "00001" when "010011001011111", -- t[9823] = 1
      "00001" when "010011001100000", -- t[9824] = 1
      "00001" when "010011001100001", -- t[9825] = 1
      "00001" when "010011001100010", -- t[9826] = 1
      "00001" when "010011001100011", -- t[9827] = 1
      "00001" when "010011001100100", -- t[9828] = 1
      "00001" when "010011001100101", -- t[9829] = 1
      "00001" when "010011001100110", -- t[9830] = 1
      "00001" when "010011001100111", -- t[9831] = 1
      "00001" when "010011001101000", -- t[9832] = 1
      "00001" when "010011001101001", -- t[9833] = 1
      "00001" when "010011001101010", -- t[9834] = 1
      "00001" when "010011001101011", -- t[9835] = 1
      "00001" when "010011001101100", -- t[9836] = 1
      "00001" when "010011001101101", -- t[9837] = 1
      "00001" when "010011001101110", -- t[9838] = 1
      "00001" when "010011001101111", -- t[9839] = 1
      "00001" when "010011001110000", -- t[9840] = 1
      "00001" when "010011001110001", -- t[9841] = 1
      "00001" when "010011001110010", -- t[9842] = 1
      "00001" when "010011001110011", -- t[9843] = 1
      "00001" when "010011001110100", -- t[9844] = 1
      "00001" when "010011001110101", -- t[9845] = 1
      "00001" when "010011001110110", -- t[9846] = 1
      "00001" when "010011001110111", -- t[9847] = 1
      "00001" when "010011001111000", -- t[9848] = 1
      "00001" when "010011001111001", -- t[9849] = 1
      "00001" when "010011001111010", -- t[9850] = 1
      "00001" when "010011001111011", -- t[9851] = 1
      "00001" when "010011001111100", -- t[9852] = 1
      "00001" when "010011001111101", -- t[9853] = 1
      "00001" when "010011001111110", -- t[9854] = 1
      "00001" when "010011001111111", -- t[9855] = 1
      "00001" when "010011010000000", -- t[9856] = 1
      "00001" when "010011010000001", -- t[9857] = 1
      "00001" when "010011010000010", -- t[9858] = 1
      "00001" when "010011010000011", -- t[9859] = 1
      "00001" when "010011010000100", -- t[9860] = 1
      "00001" when "010011010000101", -- t[9861] = 1
      "00001" when "010011010000110", -- t[9862] = 1
      "00001" when "010011010000111", -- t[9863] = 1
      "00001" when "010011010001000", -- t[9864] = 1
      "00001" when "010011010001001", -- t[9865] = 1
      "00001" when "010011010001010", -- t[9866] = 1
      "00001" when "010011010001011", -- t[9867] = 1
      "00001" when "010011010001100", -- t[9868] = 1
      "00001" when "010011010001101", -- t[9869] = 1
      "00001" when "010011010001110", -- t[9870] = 1
      "00001" when "010011010001111", -- t[9871] = 1
      "00001" when "010011010010000", -- t[9872] = 1
      "00001" when "010011010010001", -- t[9873] = 1
      "00001" when "010011010010010", -- t[9874] = 1
      "00001" when "010011010010011", -- t[9875] = 1
      "00001" when "010011010010100", -- t[9876] = 1
      "00001" when "010011010010101", -- t[9877] = 1
      "00001" when "010011010010110", -- t[9878] = 1
      "00001" when "010011010010111", -- t[9879] = 1
      "00001" when "010011010011000", -- t[9880] = 1
      "00001" when "010011010011001", -- t[9881] = 1
      "00001" when "010011010011010", -- t[9882] = 1
      "00001" when "010011010011011", -- t[9883] = 1
      "00001" when "010011010011100", -- t[9884] = 1
      "00001" when "010011010011101", -- t[9885] = 1
      "00001" when "010011010011110", -- t[9886] = 1
      "00001" when "010011010011111", -- t[9887] = 1
      "00001" when "010011010100000", -- t[9888] = 1
      "00001" when "010011010100001", -- t[9889] = 1
      "00001" when "010011010100010", -- t[9890] = 1
      "00001" when "010011010100011", -- t[9891] = 1
      "00001" when "010011010100100", -- t[9892] = 1
      "00001" when "010011010100101", -- t[9893] = 1
      "00001" when "010011010100110", -- t[9894] = 1
      "00001" when "010011010100111", -- t[9895] = 1
      "00001" when "010011010101000", -- t[9896] = 1
      "00001" when "010011010101001", -- t[9897] = 1
      "00001" when "010011010101010", -- t[9898] = 1
      "00001" when "010011010101011", -- t[9899] = 1
      "00001" when "010011010101100", -- t[9900] = 1
      "00001" when "010011010101101", -- t[9901] = 1
      "00001" when "010011010101110", -- t[9902] = 1
      "00001" when "010011010101111", -- t[9903] = 1
      "00001" when "010011010110000", -- t[9904] = 1
      "00001" when "010011010110001", -- t[9905] = 1
      "00001" when "010011010110010", -- t[9906] = 1
      "00001" when "010011010110011", -- t[9907] = 1
      "00001" when "010011010110100", -- t[9908] = 1
      "00001" when "010011010110101", -- t[9909] = 1
      "00001" when "010011010110110", -- t[9910] = 1
      "00001" when "010011010110111", -- t[9911] = 1
      "00001" when "010011010111000", -- t[9912] = 1
      "00001" when "010011010111001", -- t[9913] = 1
      "00001" when "010011010111010", -- t[9914] = 1
      "00001" when "010011010111011", -- t[9915] = 1
      "00001" when "010011010111100", -- t[9916] = 1
      "00001" when "010011010111101", -- t[9917] = 1
      "00001" when "010011010111110", -- t[9918] = 1
      "00001" when "010011010111111", -- t[9919] = 1
      "00001" when "010011011000000", -- t[9920] = 1
      "00001" when "010011011000001", -- t[9921] = 1
      "00001" when "010011011000010", -- t[9922] = 1
      "00001" when "010011011000011", -- t[9923] = 1
      "00001" when "010011011000100", -- t[9924] = 1
      "00001" when "010011011000101", -- t[9925] = 1
      "00001" when "010011011000110", -- t[9926] = 1
      "00001" when "010011011000111", -- t[9927] = 1
      "00001" when "010011011001000", -- t[9928] = 1
      "00001" when "010011011001001", -- t[9929] = 1
      "00001" when "010011011001010", -- t[9930] = 1
      "00001" when "010011011001011", -- t[9931] = 1
      "00001" when "010011011001100", -- t[9932] = 1
      "00001" when "010011011001101", -- t[9933] = 1
      "00001" when "010011011001110", -- t[9934] = 1
      "00001" when "010011011001111", -- t[9935] = 1
      "00001" when "010011011010000", -- t[9936] = 1
      "00001" when "010011011010001", -- t[9937] = 1
      "00001" when "010011011010010", -- t[9938] = 1
      "00001" when "010011011010011", -- t[9939] = 1
      "00001" when "010011011010100", -- t[9940] = 1
      "00001" when "010011011010101", -- t[9941] = 1
      "00001" when "010011011010110", -- t[9942] = 1
      "00001" when "010011011010111", -- t[9943] = 1
      "00001" when "010011011011000", -- t[9944] = 1
      "00001" when "010011011011001", -- t[9945] = 1
      "00001" when "010011011011010", -- t[9946] = 1
      "00001" when "010011011011011", -- t[9947] = 1
      "00001" when "010011011011100", -- t[9948] = 1
      "00001" when "010011011011101", -- t[9949] = 1
      "00001" when "010011011011110", -- t[9950] = 1
      "00001" when "010011011011111", -- t[9951] = 1
      "00001" when "010011011100000", -- t[9952] = 1
      "00001" when "010011011100001", -- t[9953] = 1
      "00001" when "010011011100010", -- t[9954] = 1
      "00001" when "010011011100011", -- t[9955] = 1
      "00001" when "010011011100100", -- t[9956] = 1
      "00001" when "010011011100101", -- t[9957] = 1
      "00001" when "010011011100110", -- t[9958] = 1
      "00001" when "010011011100111", -- t[9959] = 1
      "00001" when "010011011101000", -- t[9960] = 1
      "00001" when "010011011101001", -- t[9961] = 1
      "00001" when "010011011101010", -- t[9962] = 1
      "00001" when "010011011101011", -- t[9963] = 1
      "00001" when "010011011101100", -- t[9964] = 1
      "00001" when "010011011101101", -- t[9965] = 1
      "00001" when "010011011101110", -- t[9966] = 1
      "00001" when "010011011101111", -- t[9967] = 1
      "00001" when "010011011110000", -- t[9968] = 1
      "00001" when "010011011110001", -- t[9969] = 1
      "00001" when "010011011110010", -- t[9970] = 1
      "00001" when "010011011110011", -- t[9971] = 1
      "00001" when "010011011110100", -- t[9972] = 1
      "00001" when "010011011110101", -- t[9973] = 1
      "00001" when "010011011110110", -- t[9974] = 1
      "00001" when "010011011110111", -- t[9975] = 1
      "00001" when "010011011111000", -- t[9976] = 1
      "00001" when "010011011111001", -- t[9977] = 1
      "00001" when "010011011111010", -- t[9978] = 1
      "00001" when "010011011111011", -- t[9979] = 1
      "00001" when "010011011111100", -- t[9980] = 1
      "00001" when "010011011111101", -- t[9981] = 1
      "00001" when "010011011111110", -- t[9982] = 1
      "00001" when "010011011111111", -- t[9983] = 1
      "00001" when "010011100000000", -- t[9984] = 1
      "00001" when "010011100000001", -- t[9985] = 1
      "00001" when "010011100000010", -- t[9986] = 1
      "00001" when "010011100000011", -- t[9987] = 1
      "00001" when "010011100000100", -- t[9988] = 1
      "00001" when "010011100000101", -- t[9989] = 1
      "00001" when "010011100000110", -- t[9990] = 1
      "00001" when "010011100000111", -- t[9991] = 1
      "00001" when "010011100001000", -- t[9992] = 1
      "00001" when "010011100001001", -- t[9993] = 1
      "00001" when "010011100001010", -- t[9994] = 1
      "00001" when "010011100001011", -- t[9995] = 1
      "00001" when "010011100001100", -- t[9996] = 1
      "00001" when "010011100001101", -- t[9997] = 1
      "00001" when "010011100001110", -- t[9998] = 1
      "00001" when "010011100001111", -- t[9999] = 1
      "00001" when "010011100010000", -- t[10000] = 1
      "00001" when "010011100010001", -- t[10001] = 1
      "00001" when "010011100010010", -- t[10002] = 1
      "00001" when "010011100010011", -- t[10003] = 1
      "00001" when "010011100010100", -- t[10004] = 1
      "00001" when "010011100010101", -- t[10005] = 1
      "00001" when "010011100010110", -- t[10006] = 1
      "00001" when "010011100010111", -- t[10007] = 1
      "00001" when "010011100011000", -- t[10008] = 1
      "00001" when "010011100011001", -- t[10009] = 1
      "00001" when "010011100011010", -- t[10010] = 1
      "00001" when "010011100011011", -- t[10011] = 1
      "00001" when "010011100011100", -- t[10012] = 1
      "00001" when "010011100011101", -- t[10013] = 1
      "00001" when "010011100011110", -- t[10014] = 1
      "00001" when "010011100011111", -- t[10015] = 1
      "00001" when "010011100100000", -- t[10016] = 1
      "00001" when "010011100100001", -- t[10017] = 1
      "00001" when "010011100100010", -- t[10018] = 1
      "00001" when "010011100100011", -- t[10019] = 1
      "00001" when "010011100100100", -- t[10020] = 1
      "00001" when "010011100100101", -- t[10021] = 1
      "00001" when "010011100100110", -- t[10022] = 1
      "00001" when "010011100100111", -- t[10023] = 1
      "00001" when "010011100101000", -- t[10024] = 1
      "00001" when "010011100101001", -- t[10025] = 1
      "00001" when "010011100101010", -- t[10026] = 1
      "00001" when "010011100101011", -- t[10027] = 1
      "00001" when "010011100101100", -- t[10028] = 1
      "00001" when "010011100101101", -- t[10029] = 1
      "00001" when "010011100101110", -- t[10030] = 1
      "00001" when "010011100101111", -- t[10031] = 1
      "00001" when "010011100110000", -- t[10032] = 1
      "00001" when "010011100110001", -- t[10033] = 1
      "00001" when "010011100110010", -- t[10034] = 1
      "00001" when "010011100110011", -- t[10035] = 1
      "00001" when "010011100110100", -- t[10036] = 1
      "00001" when "010011100110101", -- t[10037] = 1
      "00001" when "010011100110110", -- t[10038] = 1
      "00001" when "010011100110111", -- t[10039] = 1
      "00001" when "010011100111000", -- t[10040] = 1
      "00001" when "010011100111001", -- t[10041] = 1
      "00001" when "010011100111010", -- t[10042] = 1
      "00001" when "010011100111011", -- t[10043] = 1
      "00001" when "010011100111100", -- t[10044] = 1
      "00001" when "010011100111101", -- t[10045] = 1
      "00001" when "010011100111110", -- t[10046] = 1
      "00001" when "010011100111111", -- t[10047] = 1
      "00001" when "010011101000000", -- t[10048] = 1
      "00001" when "010011101000001", -- t[10049] = 1
      "00001" when "010011101000010", -- t[10050] = 1
      "00001" when "010011101000011", -- t[10051] = 1
      "00001" when "010011101000100", -- t[10052] = 1
      "00001" when "010011101000101", -- t[10053] = 1
      "00001" when "010011101000110", -- t[10054] = 1
      "00001" when "010011101000111", -- t[10055] = 1
      "00001" when "010011101001000", -- t[10056] = 1
      "00001" when "010011101001001", -- t[10057] = 1
      "00001" when "010011101001010", -- t[10058] = 1
      "00001" when "010011101001011", -- t[10059] = 1
      "00001" when "010011101001100", -- t[10060] = 1
      "00001" when "010011101001101", -- t[10061] = 1
      "00001" when "010011101001110", -- t[10062] = 1
      "00001" when "010011101001111", -- t[10063] = 1
      "00001" when "010011101010000", -- t[10064] = 1
      "00001" when "010011101010001", -- t[10065] = 1
      "00001" when "010011101010010", -- t[10066] = 1
      "00001" when "010011101010011", -- t[10067] = 1
      "00001" when "010011101010100", -- t[10068] = 1
      "00001" when "010011101010101", -- t[10069] = 1
      "00001" when "010011101010110", -- t[10070] = 1
      "00001" when "010011101010111", -- t[10071] = 1
      "00001" when "010011101011000", -- t[10072] = 1
      "00001" when "010011101011001", -- t[10073] = 1
      "00001" when "010011101011010", -- t[10074] = 1
      "00001" when "010011101011011", -- t[10075] = 1
      "00001" when "010011101011100", -- t[10076] = 1
      "00001" when "010011101011101", -- t[10077] = 1
      "00001" when "010011101011110", -- t[10078] = 1
      "00001" when "010011101011111", -- t[10079] = 1
      "00001" when "010011101100000", -- t[10080] = 1
      "00001" when "010011101100001", -- t[10081] = 1
      "00001" when "010011101100010", -- t[10082] = 1
      "00001" when "010011101100011", -- t[10083] = 1
      "00001" when "010011101100100", -- t[10084] = 1
      "00001" when "010011101100101", -- t[10085] = 1
      "00001" when "010011101100110", -- t[10086] = 1
      "00001" when "010011101100111", -- t[10087] = 1
      "00001" when "010011101101000", -- t[10088] = 1
      "00001" when "010011101101001", -- t[10089] = 1
      "00001" when "010011101101010", -- t[10090] = 1
      "00001" when "010011101101011", -- t[10091] = 1
      "00001" when "010011101101100", -- t[10092] = 1
      "00001" when "010011101101101", -- t[10093] = 1
      "00001" when "010011101101110", -- t[10094] = 1
      "00001" when "010011101101111", -- t[10095] = 1
      "00001" when "010011101110000", -- t[10096] = 1
      "00001" when "010011101110001", -- t[10097] = 1
      "00001" when "010011101110010", -- t[10098] = 1
      "00001" when "010011101110011", -- t[10099] = 1
      "00001" when "010011101110100", -- t[10100] = 1
      "00001" when "010011101110101", -- t[10101] = 1
      "00001" when "010011101110110", -- t[10102] = 1
      "00001" when "010011101110111", -- t[10103] = 1
      "00001" when "010011101111000", -- t[10104] = 1
      "00001" when "010011101111001", -- t[10105] = 1
      "00001" when "010011101111010", -- t[10106] = 1
      "00001" when "010011101111011", -- t[10107] = 1
      "00001" when "010011101111100", -- t[10108] = 1
      "00001" when "010011101111101", -- t[10109] = 1
      "00001" when "010011101111110", -- t[10110] = 1
      "00001" when "010011101111111", -- t[10111] = 1
      "00001" when "010011110000000", -- t[10112] = 1
      "00001" when "010011110000001", -- t[10113] = 1
      "00001" when "010011110000010", -- t[10114] = 1
      "00001" when "010011110000011", -- t[10115] = 1
      "00001" when "010011110000100", -- t[10116] = 1
      "00001" when "010011110000101", -- t[10117] = 1
      "00001" when "010011110000110", -- t[10118] = 1
      "00001" when "010011110000111", -- t[10119] = 1
      "00001" when "010011110001000", -- t[10120] = 1
      "00001" when "010011110001001", -- t[10121] = 1
      "00001" when "010011110001010", -- t[10122] = 1
      "00001" when "010011110001011", -- t[10123] = 1
      "00001" when "010011110001100", -- t[10124] = 1
      "00001" when "010011110001101", -- t[10125] = 1
      "00001" when "010011110001110", -- t[10126] = 1
      "00001" when "010011110001111", -- t[10127] = 1
      "00001" when "010011110010000", -- t[10128] = 1
      "00001" when "010011110010001", -- t[10129] = 1
      "00001" when "010011110010010", -- t[10130] = 1
      "00001" when "010011110010011", -- t[10131] = 1
      "00001" when "010011110010100", -- t[10132] = 1
      "00001" when "010011110010101", -- t[10133] = 1
      "00001" when "010011110010110", -- t[10134] = 1
      "00001" when "010011110010111", -- t[10135] = 1
      "00001" when "010011110011000", -- t[10136] = 1
      "00001" when "010011110011001", -- t[10137] = 1
      "00001" when "010011110011010", -- t[10138] = 1
      "00001" when "010011110011011", -- t[10139] = 1
      "00001" when "010011110011100", -- t[10140] = 1
      "00001" when "010011110011101", -- t[10141] = 1
      "00001" when "010011110011110", -- t[10142] = 1
      "00001" when "010011110011111", -- t[10143] = 1
      "00001" when "010011110100000", -- t[10144] = 1
      "00001" when "010011110100001", -- t[10145] = 1
      "00001" when "010011110100010", -- t[10146] = 1
      "00001" when "010011110100011", -- t[10147] = 1
      "00001" when "010011110100100", -- t[10148] = 1
      "00001" when "010011110100101", -- t[10149] = 1
      "00001" when "010011110100110", -- t[10150] = 1
      "00001" when "010011110100111", -- t[10151] = 1
      "00001" when "010011110101000", -- t[10152] = 1
      "00001" when "010011110101001", -- t[10153] = 1
      "00001" when "010011110101010", -- t[10154] = 1
      "00001" when "010011110101011", -- t[10155] = 1
      "00001" when "010011110101100", -- t[10156] = 1
      "00001" when "010011110101101", -- t[10157] = 1
      "00001" when "010011110101110", -- t[10158] = 1
      "00001" when "010011110101111", -- t[10159] = 1
      "00001" when "010011110110000", -- t[10160] = 1
      "00001" when "010011110110001", -- t[10161] = 1
      "00001" when "010011110110010", -- t[10162] = 1
      "00001" when "010011110110011", -- t[10163] = 1
      "00001" when "010011110110100", -- t[10164] = 1
      "00001" when "010011110110101", -- t[10165] = 1
      "00001" when "010011110110110", -- t[10166] = 1
      "00001" when "010011110110111", -- t[10167] = 1
      "00001" when "010011110111000", -- t[10168] = 1
      "00001" when "010011110111001", -- t[10169] = 1
      "00001" when "010011110111010", -- t[10170] = 1
      "00001" when "010011110111011", -- t[10171] = 1
      "00001" when "010011110111100", -- t[10172] = 1
      "00001" when "010011110111101", -- t[10173] = 1
      "00001" when "010011110111110", -- t[10174] = 1
      "00001" when "010011110111111", -- t[10175] = 1
      "00001" when "010011111000000", -- t[10176] = 1
      "00001" when "010011111000001", -- t[10177] = 1
      "00001" when "010011111000010", -- t[10178] = 1
      "00001" when "010011111000011", -- t[10179] = 1
      "00001" when "010011111000100", -- t[10180] = 1
      "00001" when "010011111000101", -- t[10181] = 1
      "00001" when "010011111000110", -- t[10182] = 1
      "00001" when "010011111000111", -- t[10183] = 1
      "00001" when "010011111001000", -- t[10184] = 1
      "00001" when "010011111001001", -- t[10185] = 1
      "00001" when "010011111001010", -- t[10186] = 1
      "00001" when "010011111001011", -- t[10187] = 1
      "00001" when "010011111001100", -- t[10188] = 1
      "00001" when "010011111001101", -- t[10189] = 1
      "00001" when "010011111001110", -- t[10190] = 1
      "00001" when "010011111001111", -- t[10191] = 1
      "00001" when "010011111010000", -- t[10192] = 1
      "00001" when "010011111010001", -- t[10193] = 1
      "00001" when "010011111010010", -- t[10194] = 1
      "00001" when "010011111010011", -- t[10195] = 1
      "00001" when "010011111010100", -- t[10196] = 1
      "00001" when "010011111010101", -- t[10197] = 1
      "00001" when "010011111010110", -- t[10198] = 1
      "00001" when "010011111010111", -- t[10199] = 1
      "00001" when "010011111011000", -- t[10200] = 1
      "00001" when "010011111011001", -- t[10201] = 1
      "00001" when "010011111011010", -- t[10202] = 1
      "00001" when "010011111011011", -- t[10203] = 1
      "00001" when "010011111011100", -- t[10204] = 1
      "00001" when "010011111011101", -- t[10205] = 1
      "00001" when "010011111011110", -- t[10206] = 1
      "00001" when "010011111011111", -- t[10207] = 1
      "00001" when "010011111100000", -- t[10208] = 1
      "00001" when "010011111100001", -- t[10209] = 1
      "00001" when "010011111100010", -- t[10210] = 1
      "00001" when "010011111100011", -- t[10211] = 1
      "00001" when "010011111100100", -- t[10212] = 1
      "00001" when "010011111100101", -- t[10213] = 1
      "00001" when "010011111100110", -- t[10214] = 1
      "00001" when "010011111100111", -- t[10215] = 1
      "00001" when "010011111101000", -- t[10216] = 1
      "00001" when "010011111101001", -- t[10217] = 1
      "00001" when "010011111101010", -- t[10218] = 1
      "00001" when "010011111101011", -- t[10219] = 1
      "00001" when "010011111101100", -- t[10220] = 1
      "00001" when "010011111101101", -- t[10221] = 1
      "00001" when "010011111101110", -- t[10222] = 1
      "00001" when "010011111101111", -- t[10223] = 1
      "00001" when "010011111110000", -- t[10224] = 1
      "00001" when "010011111110001", -- t[10225] = 1
      "00001" when "010011111110010", -- t[10226] = 1
      "00001" when "010011111110011", -- t[10227] = 1
      "00001" when "010011111110100", -- t[10228] = 1
      "00001" when "010011111110101", -- t[10229] = 1
      "00001" when "010011111110110", -- t[10230] = 1
      "00001" when "010011111110111", -- t[10231] = 1
      "00001" when "010011111111000", -- t[10232] = 1
      "00001" when "010011111111001", -- t[10233] = 1
      "00001" when "010011111111010", -- t[10234] = 1
      "00001" when "010011111111011", -- t[10235] = 1
      "00001" when "010011111111100", -- t[10236] = 1
      "00001" when "010011111111101", -- t[10237] = 1
      "00001" when "010011111111110", -- t[10238] = 1
      "00001" when "010011111111111", -- t[10239] = 1
      "00001" when "010100000000000", -- t[10240] = 1
      "00001" when "010100000000001", -- t[10241] = 1
      "00001" when "010100000000010", -- t[10242] = 1
      "00001" when "010100000000011", -- t[10243] = 1
      "00001" when "010100000000100", -- t[10244] = 1
      "00001" when "010100000000101", -- t[10245] = 1
      "00001" when "010100000000110", -- t[10246] = 1
      "00001" when "010100000000111", -- t[10247] = 1
      "00001" when "010100000001000", -- t[10248] = 1
      "00001" when "010100000001001", -- t[10249] = 1
      "00001" when "010100000001010", -- t[10250] = 1
      "00001" when "010100000001011", -- t[10251] = 1
      "00001" when "010100000001100", -- t[10252] = 1
      "00001" when "010100000001101", -- t[10253] = 1
      "00001" when "010100000001110", -- t[10254] = 1
      "00001" when "010100000001111", -- t[10255] = 1
      "00001" when "010100000010000", -- t[10256] = 1
      "00001" when "010100000010001", -- t[10257] = 1
      "00001" when "010100000010010", -- t[10258] = 1
      "00001" when "010100000010011", -- t[10259] = 1
      "00001" when "010100000010100", -- t[10260] = 1
      "00001" when "010100000010101", -- t[10261] = 1
      "00001" when "010100000010110", -- t[10262] = 1
      "00001" when "010100000010111", -- t[10263] = 1
      "00001" when "010100000011000", -- t[10264] = 1
      "00001" when "010100000011001", -- t[10265] = 1
      "00001" when "010100000011010", -- t[10266] = 1
      "00001" when "010100000011011", -- t[10267] = 1
      "00001" when "010100000011100", -- t[10268] = 1
      "00001" when "010100000011101", -- t[10269] = 1
      "00001" when "010100000011110", -- t[10270] = 1
      "00001" when "010100000011111", -- t[10271] = 1
      "00001" when "010100000100000", -- t[10272] = 1
      "00001" when "010100000100001", -- t[10273] = 1
      "00001" when "010100000100010", -- t[10274] = 1
      "00001" when "010100000100011", -- t[10275] = 1
      "00001" when "010100000100100", -- t[10276] = 1
      "00001" when "010100000100101", -- t[10277] = 1
      "00001" when "010100000100110", -- t[10278] = 1
      "00001" when "010100000100111", -- t[10279] = 1
      "00001" when "010100000101000", -- t[10280] = 1
      "00001" when "010100000101001", -- t[10281] = 1
      "00001" when "010100000101010", -- t[10282] = 1
      "00001" when "010100000101011", -- t[10283] = 1
      "00001" when "010100000101100", -- t[10284] = 1
      "00001" when "010100000101101", -- t[10285] = 1
      "00001" when "010100000101110", -- t[10286] = 1
      "00001" when "010100000101111", -- t[10287] = 1
      "00001" when "010100000110000", -- t[10288] = 1
      "00001" when "010100000110001", -- t[10289] = 1
      "00001" when "010100000110010", -- t[10290] = 1
      "00001" when "010100000110011", -- t[10291] = 1
      "00001" when "010100000110100", -- t[10292] = 1
      "00001" when "010100000110101", -- t[10293] = 1
      "00001" when "010100000110110", -- t[10294] = 1
      "00001" when "010100000110111", -- t[10295] = 1
      "00001" when "010100000111000", -- t[10296] = 1
      "00001" when "010100000111001", -- t[10297] = 1
      "00001" when "010100000111010", -- t[10298] = 1
      "00001" when "010100000111011", -- t[10299] = 1
      "00001" when "010100000111100", -- t[10300] = 1
      "00001" when "010100000111101", -- t[10301] = 1
      "00001" when "010100000111110", -- t[10302] = 1
      "00001" when "010100000111111", -- t[10303] = 1
      "00001" when "010100001000000", -- t[10304] = 1
      "00001" when "010100001000001", -- t[10305] = 1
      "00001" when "010100001000010", -- t[10306] = 1
      "00001" when "010100001000011", -- t[10307] = 1
      "00001" when "010100001000100", -- t[10308] = 1
      "00001" when "010100001000101", -- t[10309] = 1
      "00001" when "010100001000110", -- t[10310] = 1
      "00001" when "010100001000111", -- t[10311] = 1
      "00001" when "010100001001000", -- t[10312] = 1
      "00001" when "010100001001001", -- t[10313] = 1
      "00001" when "010100001001010", -- t[10314] = 1
      "00001" when "010100001001011", -- t[10315] = 1
      "00001" when "010100001001100", -- t[10316] = 1
      "00001" when "010100001001101", -- t[10317] = 1
      "00001" when "010100001001110", -- t[10318] = 1
      "00001" when "010100001001111", -- t[10319] = 1
      "00001" when "010100001010000", -- t[10320] = 1
      "00001" when "010100001010001", -- t[10321] = 1
      "00001" when "010100001010010", -- t[10322] = 1
      "00001" when "010100001010011", -- t[10323] = 1
      "00001" when "010100001010100", -- t[10324] = 1
      "00001" when "010100001010101", -- t[10325] = 1
      "00001" when "010100001010110", -- t[10326] = 1
      "00001" when "010100001010111", -- t[10327] = 1
      "00001" when "010100001011000", -- t[10328] = 1
      "00001" when "010100001011001", -- t[10329] = 1
      "00001" when "010100001011010", -- t[10330] = 1
      "00001" when "010100001011011", -- t[10331] = 1
      "00001" when "010100001011100", -- t[10332] = 1
      "00001" when "010100001011101", -- t[10333] = 1
      "00001" when "010100001011110", -- t[10334] = 1
      "00001" when "010100001011111", -- t[10335] = 1
      "00001" when "010100001100000", -- t[10336] = 1
      "00001" when "010100001100001", -- t[10337] = 1
      "00001" when "010100001100010", -- t[10338] = 1
      "00001" when "010100001100011", -- t[10339] = 1
      "00001" when "010100001100100", -- t[10340] = 1
      "00001" when "010100001100101", -- t[10341] = 1
      "00001" when "010100001100110", -- t[10342] = 1
      "00001" when "010100001100111", -- t[10343] = 1
      "00001" when "010100001101000", -- t[10344] = 1
      "00001" when "010100001101001", -- t[10345] = 1
      "00001" when "010100001101010", -- t[10346] = 1
      "00001" when "010100001101011", -- t[10347] = 1
      "00001" when "010100001101100", -- t[10348] = 1
      "00001" when "010100001101101", -- t[10349] = 1
      "00001" when "010100001101110", -- t[10350] = 1
      "00001" when "010100001101111", -- t[10351] = 1
      "00001" when "010100001110000", -- t[10352] = 1
      "00001" when "010100001110001", -- t[10353] = 1
      "00001" when "010100001110010", -- t[10354] = 1
      "00010" when "010100001110011", -- t[10355] = 2
      "00010" when "010100001110100", -- t[10356] = 2
      "00010" when "010100001110101", -- t[10357] = 2
      "00010" when "010100001110110", -- t[10358] = 2
      "00010" when "010100001110111", -- t[10359] = 2
      "00010" when "010100001111000", -- t[10360] = 2
      "00010" when "010100001111001", -- t[10361] = 2
      "00010" when "010100001111010", -- t[10362] = 2
      "00010" when "010100001111011", -- t[10363] = 2
      "00010" when "010100001111100", -- t[10364] = 2
      "00010" when "010100001111101", -- t[10365] = 2
      "00010" when "010100001111110", -- t[10366] = 2
      "00010" when "010100001111111", -- t[10367] = 2
      "00010" when "010100010000000", -- t[10368] = 2
      "00010" when "010100010000001", -- t[10369] = 2
      "00010" when "010100010000010", -- t[10370] = 2
      "00010" when "010100010000011", -- t[10371] = 2
      "00010" when "010100010000100", -- t[10372] = 2
      "00010" when "010100010000101", -- t[10373] = 2
      "00010" when "010100010000110", -- t[10374] = 2
      "00010" when "010100010000111", -- t[10375] = 2
      "00010" when "010100010001000", -- t[10376] = 2
      "00010" when "010100010001001", -- t[10377] = 2
      "00010" when "010100010001010", -- t[10378] = 2
      "00010" when "010100010001011", -- t[10379] = 2
      "00010" when "010100010001100", -- t[10380] = 2
      "00010" when "010100010001101", -- t[10381] = 2
      "00010" when "010100010001110", -- t[10382] = 2
      "00010" when "010100010001111", -- t[10383] = 2
      "00010" when "010100010010000", -- t[10384] = 2
      "00010" when "010100010010001", -- t[10385] = 2
      "00010" when "010100010010010", -- t[10386] = 2
      "00010" when "010100010010011", -- t[10387] = 2
      "00010" when "010100010010100", -- t[10388] = 2
      "00010" when "010100010010101", -- t[10389] = 2
      "00010" when "010100010010110", -- t[10390] = 2
      "00010" when "010100010010111", -- t[10391] = 2
      "00010" when "010100010011000", -- t[10392] = 2
      "00010" when "010100010011001", -- t[10393] = 2
      "00010" when "010100010011010", -- t[10394] = 2
      "00010" when "010100010011011", -- t[10395] = 2
      "00010" when "010100010011100", -- t[10396] = 2
      "00010" when "010100010011101", -- t[10397] = 2
      "00010" when "010100010011110", -- t[10398] = 2
      "00010" when "010100010011111", -- t[10399] = 2
      "00010" when "010100010100000", -- t[10400] = 2
      "00010" when "010100010100001", -- t[10401] = 2
      "00010" when "010100010100010", -- t[10402] = 2
      "00010" when "010100010100011", -- t[10403] = 2
      "00010" when "010100010100100", -- t[10404] = 2
      "00010" when "010100010100101", -- t[10405] = 2
      "00010" when "010100010100110", -- t[10406] = 2
      "00010" when "010100010100111", -- t[10407] = 2
      "00010" when "010100010101000", -- t[10408] = 2
      "00010" when "010100010101001", -- t[10409] = 2
      "00010" when "010100010101010", -- t[10410] = 2
      "00010" when "010100010101011", -- t[10411] = 2
      "00010" when "010100010101100", -- t[10412] = 2
      "00010" when "010100010101101", -- t[10413] = 2
      "00010" when "010100010101110", -- t[10414] = 2
      "00010" when "010100010101111", -- t[10415] = 2
      "00010" when "010100010110000", -- t[10416] = 2
      "00010" when "010100010110001", -- t[10417] = 2
      "00010" when "010100010110010", -- t[10418] = 2
      "00010" when "010100010110011", -- t[10419] = 2
      "00010" when "010100010110100", -- t[10420] = 2
      "00010" when "010100010110101", -- t[10421] = 2
      "00010" when "010100010110110", -- t[10422] = 2
      "00010" when "010100010110111", -- t[10423] = 2
      "00010" when "010100010111000", -- t[10424] = 2
      "00010" when "010100010111001", -- t[10425] = 2
      "00010" when "010100010111010", -- t[10426] = 2
      "00010" when "010100010111011", -- t[10427] = 2
      "00010" when "010100010111100", -- t[10428] = 2
      "00010" when "010100010111101", -- t[10429] = 2
      "00010" when "010100010111110", -- t[10430] = 2
      "00010" when "010100010111111", -- t[10431] = 2
      "00010" when "010100011000000", -- t[10432] = 2
      "00010" when "010100011000001", -- t[10433] = 2
      "00010" when "010100011000010", -- t[10434] = 2
      "00010" when "010100011000011", -- t[10435] = 2
      "00010" when "010100011000100", -- t[10436] = 2
      "00010" when "010100011000101", -- t[10437] = 2
      "00010" when "010100011000110", -- t[10438] = 2
      "00010" when "010100011000111", -- t[10439] = 2
      "00010" when "010100011001000", -- t[10440] = 2
      "00010" when "010100011001001", -- t[10441] = 2
      "00010" when "010100011001010", -- t[10442] = 2
      "00010" when "010100011001011", -- t[10443] = 2
      "00010" when "010100011001100", -- t[10444] = 2
      "00010" when "010100011001101", -- t[10445] = 2
      "00010" when "010100011001110", -- t[10446] = 2
      "00010" when "010100011001111", -- t[10447] = 2
      "00010" when "010100011010000", -- t[10448] = 2
      "00010" when "010100011010001", -- t[10449] = 2
      "00010" when "010100011010010", -- t[10450] = 2
      "00010" when "010100011010011", -- t[10451] = 2
      "00010" when "010100011010100", -- t[10452] = 2
      "00010" when "010100011010101", -- t[10453] = 2
      "00010" when "010100011010110", -- t[10454] = 2
      "00010" when "010100011010111", -- t[10455] = 2
      "00010" when "010100011011000", -- t[10456] = 2
      "00010" when "010100011011001", -- t[10457] = 2
      "00010" when "010100011011010", -- t[10458] = 2
      "00010" when "010100011011011", -- t[10459] = 2
      "00010" when "010100011011100", -- t[10460] = 2
      "00010" when "010100011011101", -- t[10461] = 2
      "00010" when "010100011011110", -- t[10462] = 2
      "00010" when "010100011011111", -- t[10463] = 2
      "00010" when "010100011100000", -- t[10464] = 2
      "00010" when "010100011100001", -- t[10465] = 2
      "00010" when "010100011100010", -- t[10466] = 2
      "00010" when "010100011100011", -- t[10467] = 2
      "00010" when "010100011100100", -- t[10468] = 2
      "00010" when "010100011100101", -- t[10469] = 2
      "00010" when "010100011100110", -- t[10470] = 2
      "00010" when "010100011100111", -- t[10471] = 2
      "00010" when "010100011101000", -- t[10472] = 2
      "00010" when "010100011101001", -- t[10473] = 2
      "00010" when "010100011101010", -- t[10474] = 2
      "00010" when "010100011101011", -- t[10475] = 2
      "00010" when "010100011101100", -- t[10476] = 2
      "00010" when "010100011101101", -- t[10477] = 2
      "00010" when "010100011101110", -- t[10478] = 2
      "00010" when "010100011101111", -- t[10479] = 2
      "00010" when "010100011110000", -- t[10480] = 2
      "00010" when "010100011110001", -- t[10481] = 2
      "00010" when "010100011110010", -- t[10482] = 2
      "00010" when "010100011110011", -- t[10483] = 2
      "00010" when "010100011110100", -- t[10484] = 2
      "00010" when "010100011110101", -- t[10485] = 2
      "00010" when "010100011110110", -- t[10486] = 2
      "00010" when "010100011110111", -- t[10487] = 2
      "00010" when "010100011111000", -- t[10488] = 2
      "00010" when "010100011111001", -- t[10489] = 2
      "00010" when "010100011111010", -- t[10490] = 2
      "00010" when "010100011111011", -- t[10491] = 2
      "00010" when "010100011111100", -- t[10492] = 2
      "00010" when "010100011111101", -- t[10493] = 2
      "00010" when "010100011111110", -- t[10494] = 2
      "00010" when "010100011111111", -- t[10495] = 2
      "00010" when "010100100000000", -- t[10496] = 2
      "00010" when "010100100000001", -- t[10497] = 2
      "00010" when "010100100000010", -- t[10498] = 2
      "00010" when "010100100000011", -- t[10499] = 2
      "00010" when "010100100000100", -- t[10500] = 2
      "00010" when "010100100000101", -- t[10501] = 2
      "00010" when "010100100000110", -- t[10502] = 2
      "00010" when "010100100000111", -- t[10503] = 2
      "00010" when "010100100001000", -- t[10504] = 2
      "00010" when "010100100001001", -- t[10505] = 2
      "00010" when "010100100001010", -- t[10506] = 2
      "00010" when "010100100001011", -- t[10507] = 2
      "00010" when "010100100001100", -- t[10508] = 2
      "00010" when "010100100001101", -- t[10509] = 2
      "00010" when "010100100001110", -- t[10510] = 2
      "00010" when "010100100001111", -- t[10511] = 2
      "00010" when "010100100010000", -- t[10512] = 2
      "00010" when "010100100010001", -- t[10513] = 2
      "00010" when "010100100010010", -- t[10514] = 2
      "00010" when "010100100010011", -- t[10515] = 2
      "00010" when "010100100010100", -- t[10516] = 2
      "00010" when "010100100010101", -- t[10517] = 2
      "00010" when "010100100010110", -- t[10518] = 2
      "00010" when "010100100010111", -- t[10519] = 2
      "00010" when "010100100011000", -- t[10520] = 2
      "00010" when "010100100011001", -- t[10521] = 2
      "00010" when "010100100011010", -- t[10522] = 2
      "00010" when "010100100011011", -- t[10523] = 2
      "00010" when "010100100011100", -- t[10524] = 2
      "00010" when "010100100011101", -- t[10525] = 2
      "00010" when "010100100011110", -- t[10526] = 2
      "00010" when "010100100011111", -- t[10527] = 2
      "00010" when "010100100100000", -- t[10528] = 2
      "00010" when "010100100100001", -- t[10529] = 2
      "00010" when "010100100100010", -- t[10530] = 2
      "00010" when "010100100100011", -- t[10531] = 2
      "00010" when "010100100100100", -- t[10532] = 2
      "00010" when "010100100100101", -- t[10533] = 2
      "00010" when "010100100100110", -- t[10534] = 2
      "00010" when "010100100100111", -- t[10535] = 2
      "00010" when "010100100101000", -- t[10536] = 2
      "00010" when "010100100101001", -- t[10537] = 2
      "00010" when "010100100101010", -- t[10538] = 2
      "00010" when "010100100101011", -- t[10539] = 2
      "00010" when "010100100101100", -- t[10540] = 2
      "00010" when "010100100101101", -- t[10541] = 2
      "00010" when "010100100101110", -- t[10542] = 2
      "00010" when "010100100101111", -- t[10543] = 2
      "00010" when "010100100110000", -- t[10544] = 2
      "00010" when "010100100110001", -- t[10545] = 2
      "00010" when "010100100110010", -- t[10546] = 2
      "00010" when "010100100110011", -- t[10547] = 2
      "00010" when "010100100110100", -- t[10548] = 2
      "00010" when "010100100110101", -- t[10549] = 2
      "00010" when "010100100110110", -- t[10550] = 2
      "00010" when "010100100110111", -- t[10551] = 2
      "00010" when "010100100111000", -- t[10552] = 2
      "00010" when "010100100111001", -- t[10553] = 2
      "00010" when "010100100111010", -- t[10554] = 2
      "00010" when "010100100111011", -- t[10555] = 2
      "00010" when "010100100111100", -- t[10556] = 2
      "00010" when "010100100111101", -- t[10557] = 2
      "00010" when "010100100111110", -- t[10558] = 2
      "00010" when "010100100111111", -- t[10559] = 2
      "00010" when "010100101000000", -- t[10560] = 2
      "00010" when "010100101000001", -- t[10561] = 2
      "00010" when "010100101000010", -- t[10562] = 2
      "00010" when "010100101000011", -- t[10563] = 2
      "00010" when "010100101000100", -- t[10564] = 2
      "00010" when "010100101000101", -- t[10565] = 2
      "00010" when "010100101000110", -- t[10566] = 2
      "00010" when "010100101000111", -- t[10567] = 2
      "00010" when "010100101001000", -- t[10568] = 2
      "00010" when "010100101001001", -- t[10569] = 2
      "00010" when "010100101001010", -- t[10570] = 2
      "00010" when "010100101001011", -- t[10571] = 2
      "00010" when "010100101001100", -- t[10572] = 2
      "00010" when "010100101001101", -- t[10573] = 2
      "00010" when "010100101001110", -- t[10574] = 2
      "00010" when "010100101001111", -- t[10575] = 2
      "00010" when "010100101010000", -- t[10576] = 2
      "00010" when "010100101010001", -- t[10577] = 2
      "00010" when "010100101010010", -- t[10578] = 2
      "00010" when "010100101010011", -- t[10579] = 2
      "00010" when "010100101010100", -- t[10580] = 2
      "00010" when "010100101010101", -- t[10581] = 2
      "00010" when "010100101010110", -- t[10582] = 2
      "00010" when "010100101010111", -- t[10583] = 2
      "00010" when "010100101011000", -- t[10584] = 2
      "00010" when "010100101011001", -- t[10585] = 2
      "00010" when "010100101011010", -- t[10586] = 2
      "00010" when "010100101011011", -- t[10587] = 2
      "00010" when "010100101011100", -- t[10588] = 2
      "00010" when "010100101011101", -- t[10589] = 2
      "00010" when "010100101011110", -- t[10590] = 2
      "00010" when "010100101011111", -- t[10591] = 2
      "00010" when "010100101100000", -- t[10592] = 2
      "00010" when "010100101100001", -- t[10593] = 2
      "00010" when "010100101100010", -- t[10594] = 2
      "00010" when "010100101100011", -- t[10595] = 2
      "00010" when "010100101100100", -- t[10596] = 2
      "00010" when "010100101100101", -- t[10597] = 2
      "00010" when "010100101100110", -- t[10598] = 2
      "00010" when "010100101100111", -- t[10599] = 2
      "00010" when "010100101101000", -- t[10600] = 2
      "00010" when "010100101101001", -- t[10601] = 2
      "00010" when "010100101101010", -- t[10602] = 2
      "00010" when "010100101101011", -- t[10603] = 2
      "00010" when "010100101101100", -- t[10604] = 2
      "00010" when "010100101101101", -- t[10605] = 2
      "00010" when "010100101101110", -- t[10606] = 2
      "00010" when "010100101101111", -- t[10607] = 2
      "00010" when "010100101110000", -- t[10608] = 2
      "00010" when "010100101110001", -- t[10609] = 2
      "00010" when "010100101110010", -- t[10610] = 2
      "00010" when "010100101110011", -- t[10611] = 2
      "00010" when "010100101110100", -- t[10612] = 2
      "00010" when "010100101110101", -- t[10613] = 2
      "00010" when "010100101110110", -- t[10614] = 2
      "00010" when "010100101110111", -- t[10615] = 2
      "00010" when "010100101111000", -- t[10616] = 2
      "00010" when "010100101111001", -- t[10617] = 2
      "00010" when "010100101111010", -- t[10618] = 2
      "00010" when "010100101111011", -- t[10619] = 2
      "00010" when "010100101111100", -- t[10620] = 2
      "00010" when "010100101111101", -- t[10621] = 2
      "00010" when "010100101111110", -- t[10622] = 2
      "00010" when "010100101111111", -- t[10623] = 2
      "00010" when "010100110000000", -- t[10624] = 2
      "00010" when "010100110000001", -- t[10625] = 2
      "00010" when "010100110000010", -- t[10626] = 2
      "00010" when "010100110000011", -- t[10627] = 2
      "00010" when "010100110000100", -- t[10628] = 2
      "00010" when "010100110000101", -- t[10629] = 2
      "00010" when "010100110000110", -- t[10630] = 2
      "00010" when "010100110000111", -- t[10631] = 2
      "00010" when "010100110001000", -- t[10632] = 2
      "00010" when "010100110001001", -- t[10633] = 2
      "00010" when "010100110001010", -- t[10634] = 2
      "00010" when "010100110001011", -- t[10635] = 2
      "00010" when "010100110001100", -- t[10636] = 2
      "00010" when "010100110001101", -- t[10637] = 2
      "00010" when "010100110001110", -- t[10638] = 2
      "00010" when "010100110001111", -- t[10639] = 2
      "00010" when "010100110010000", -- t[10640] = 2
      "00010" when "010100110010001", -- t[10641] = 2
      "00010" when "010100110010010", -- t[10642] = 2
      "00010" when "010100110010011", -- t[10643] = 2
      "00010" when "010100110010100", -- t[10644] = 2
      "00010" when "010100110010101", -- t[10645] = 2
      "00010" when "010100110010110", -- t[10646] = 2
      "00010" when "010100110010111", -- t[10647] = 2
      "00010" when "010100110011000", -- t[10648] = 2
      "00010" when "010100110011001", -- t[10649] = 2
      "00010" when "010100110011010", -- t[10650] = 2
      "00010" when "010100110011011", -- t[10651] = 2
      "00010" when "010100110011100", -- t[10652] = 2
      "00010" when "010100110011101", -- t[10653] = 2
      "00010" when "010100110011110", -- t[10654] = 2
      "00010" when "010100110011111", -- t[10655] = 2
      "00010" when "010100110100000", -- t[10656] = 2
      "00010" when "010100110100001", -- t[10657] = 2
      "00010" when "010100110100010", -- t[10658] = 2
      "00010" when "010100110100011", -- t[10659] = 2
      "00010" when "010100110100100", -- t[10660] = 2
      "00010" when "010100110100101", -- t[10661] = 2
      "00010" when "010100110100110", -- t[10662] = 2
      "00010" when "010100110100111", -- t[10663] = 2
      "00010" when "010100110101000", -- t[10664] = 2
      "00010" when "010100110101001", -- t[10665] = 2
      "00010" when "010100110101010", -- t[10666] = 2
      "00010" when "010100110101011", -- t[10667] = 2
      "00010" when "010100110101100", -- t[10668] = 2
      "00010" when "010100110101101", -- t[10669] = 2
      "00010" when "010100110101110", -- t[10670] = 2
      "00010" when "010100110101111", -- t[10671] = 2
      "00010" when "010100110110000", -- t[10672] = 2
      "00010" when "010100110110001", -- t[10673] = 2
      "00010" when "010100110110010", -- t[10674] = 2
      "00010" when "010100110110011", -- t[10675] = 2
      "00010" when "010100110110100", -- t[10676] = 2
      "00010" when "010100110110101", -- t[10677] = 2
      "00010" when "010100110110110", -- t[10678] = 2
      "00010" when "010100110110111", -- t[10679] = 2
      "00010" when "010100110111000", -- t[10680] = 2
      "00010" when "010100110111001", -- t[10681] = 2
      "00010" when "010100110111010", -- t[10682] = 2
      "00010" when "010100110111011", -- t[10683] = 2
      "00010" when "010100110111100", -- t[10684] = 2
      "00010" when "010100110111101", -- t[10685] = 2
      "00010" when "010100110111110", -- t[10686] = 2
      "00010" when "010100110111111", -- t[10687] = 2
      "00010" when "010100111000000", -- t[10688] = 2
      "00010" when "010100111000001", -- t[10689] = 2
      "00010" when "010100111000010", -- t[10690] = 2
      "00010" when "010100111000011", -- t[10691] = 2
      "00010" when "010100111000100", -- t[10692] = 2
      "00010" when "010100111000101", -- t[10693] = 2
      "00010" when "010100111000110", -- t[10694] = 2
      "00010" when "010100111000111", -- t[10695] = 2
      "00010" when "010100111001000", -- t[10696] = 2
      "00010" when "010100111001001", -- t[10697] = 2
      "00010" when "010100111001010", -- t[10698] = 2
      "00010" when "010100111001011", -- t[10699] = 2
      "00010" when "010100111001100", -- t[10700] = 2
      "00010" when "010100111001101", -- t[10701] = 2
      "00010" when "010100111001110", -- t[10702] = 2
      "00010" when "010100111001111", -- t[10703] = 2
      "00010" when "010100111010000", -- t[10704] = 2
      "00010" when "010100111010001", -- t[10705] = 2
      "00010" when "010100111010010", -- t[10706] = 2
      "00010" when "010100111010011", -- t[10707] = 2
      "00010" when "010100111010100", -- t[10708] = 2
      "00010" when "010100111010101", -- t[10709] = 2
      "00010" when "010100111010110", -- t[10710] = 2
      "00010" when "010100111010111", -- t[10711] = 2
      "00010" when "010100111011000", -- t[10712] = 2
      "00010" when "010100111011001", -- t[10713] = 2
      "00010" when "010100111011010", -- t[10714] = 2
      "00010" when "010100111011011", -- t[10715] = 2
      "00010" when "010100111011100", -- t[10716] = 2
      "00010" when "010100111011101", -- t[10717] = 2
      "00010" when "010100111011110", -- t[10718] = 2
      "00010" when "010100111011111", -- t[10719] = 2
      "00010" when "010100111100000", -- t[10720] = 2
      "00010" when "010100111100001", -- t[10721] = 2
      "00010" when "010100111100010", -- t[10722] = 2
      "00010" when "010100111100011", -- t[10723] = 2
      "00010" when "010100111100100", -- t[10724] = 2
      "00010" when "010100111100101", -- t[10725] = 2
      "00010" when "010100111100110", -- t[10726] = 2
      "00010" when "010100111100111", -- t[10727] = 2
      "00010" when "010100111101000", -- t[10728] = 2
      "00010" when "010100111101001", -- t[10729] = 2
      "00010" when "010100111101010", -- t[10730] = 2
      "00010" when "010100111101011", -- t[10731] = 2
      "00010" when "010100111101100", -- t[10732] = 2
      "00010" when "010100111101101", -- t[10733] = 2
      "00010" when "010100111101110", -- t[10734] = 2
      "00010" when "010100111101111", -- t[10735] = 2
      "00010" when "010100111110000", -- t[10736] = 2
      "00010" when "010100111110001", -- t[10737] = 2
      "00010" when "010100111110010", -- t[10738] = 2
      "00010" when "010100111110011", -- t[10739] = 2
      "00010" when "010100111110100", -- t[10740] = 2
      "00010" when "010100111110101", -- t[10741] = 2
      "00010" when "010100111110110", -- t[10742] = 2
      "00010" when "010100111110111", -- t[10743] = 2
      "00010" when "010100111111000", -- t[10744] = 2
      "00010" when "010100111111001", -- t[10745] = 2
      "00010" when "010100111111010", -- t[10746] = 2
      "00010" when "010100111111011", -- t[10747] = 2
      "00010" when "010100111111100", -- t[10748] = 2
      "00010" when "010100111111101", -- t[10749] = 2
      "00010" when "010100111111110", -- t[10750] = 2
      "00010" when "010100111111111", -- t[10751] = 2
      "00010" when "010101000000000", -- t[10752] = 2
      "00010" when "010101000000001", -- t[10753] = 2
      "00010" when "010101000000010", -- t[10754] = 2
      "00010" when "010101000000011", -- t[10755] = 2
      "00010" when "010101000000100", -- t[10756] = 2
      "00010" when "010101000000101", -- t[10757] = 2
      "00010" when "010101000000110", -- t[10758] = 2
      "00010" when "010101000000111", -- t[10759] = 2
      "00010" when "010101000001000", -- t[10760] = 2
      "00010" when "010101000001001", -- t[10761] = 2
      "00010" when "010101000001010", -- t[10762] = 2
      "00010" when "010101000001011", -- t[10763] = 2
      "00010" when "010101000001100", -- t[10764] = 2
      "00010" when "010101000001101", -- t[10765] = 2
      "00010" when "010101000001110", -- t[10766] = 2
      "00010" when "010101000001111", -- t[10767] = 2
      "00010" when "010101000010000", -- t[10768] = 2
      "00010" when "010101000010001", -- t[10769] = 2
      "00010" when "010101000010010", -- t[10770] = 2
      "00010" when "010101000010011", -- t[10771] = 2
      "00010" when "010101000010100", -- t[10772] = 2
      "00010" when "010101000010101", -- t[10773] = 2
      "00010" when "010101000010110", -- t[10774] = 2
      "00010" when "010101000010111", -- t[10775] = 2
      "00010" when "010101000011000", -- t[10776] = 2
      "00010" when "010101000011001", -- t[10777] = 2
      "00010" when "010101000011010", -- t[10778] = 2
      "00010" when "010101000011011", -- t[10779] = 2
      "00010" when "010101000011100", -- t[10780] = 2
      "00010" when "010101000011101", -- t[10781] = 2
      "00010" when "010101000011110", -- t[10782] = 2
      "00010" when "010101000011111", -- t[10783] = 2
      "00010" when "010101000100000", -- t[10784] = 2
      "00010" when "010101000100001", -- t[10785] = 2
      "00010" when "010101000100010", -- t[10786] = 2
      "00010" when "010101000100011", -- t[10787] = 2
      "00010" when "010101000100100", -- t[10788] = 2
      "00010" when "010101000100101", -- t[10789] = 2
      "00010" when "010101000100110", -- t[10790] = 2
      "00010" when "010101000100111", -- t[10791] = 2
      "00010" when "010101000101000", -- t[10792] = 2
      "00010" when "010101000101001", -- t[10793] = 2
      "00010" when "010101000101010", -- t[10794] = 2
      "00010" when "010101000101011", -- t[10795] = 2
      "00010" when "010101000101100", -- t[10796] = 2
      "00010" when "010101000101101", -- t[10797] = 2
      "00010" when "010101000101110", -- t[10798] = 2
      "00010" when "010101000101111", -- t[10799] = 2
      "00010" when "010101000110000", -- t[10800] = 2
      "00010" when "010101000110001", -- t[10801] = 2
      "00010" when "010101000110010", -- t[10802] = 2
      "00010" when "010101000110011", -- t[10803] = 2
      "00010" when "010101000110100", -- t[10804] = 2
      "00010" when "010101000110101", -- t[10805] = 2
      "00010" when "010101000110110", -- t[10806] = 2
      "00010" when "010101000110111", -- t[10807] = 2
      "00010" when "010101000111000", -- t[10808] = 2
      "00010" when "010101000111001", -- t[10809] = 2
      "00010" when "010101000111010", -- t[10810] = 2
      "00010" when "010101000111011", -- t[10811] = 2
      "00010" when "010101000111100", -- t[10812] = 2
      "00010" when "010101000111101", -- t[10813] = 2
      "00010" when "010101000111110", -- t[10814] = 2
      "00010" when "010101000111111", -- t[10815] = 2
      "00010" when "010101001000000", -- t[10816] = 2
      "00010" when "010101001000001", -- t[10817] = 2
      "00010" when "010101001000010", -- t[10818] = 2
      "00010" when "010101001000011", -- t[10819] = 2
      "00010" when "010101001000100", -- t[10820] = 2
      "00010" when "010101001000101", -- t[10821] = 2
      "00010" when "010101001000110", -- t[10822] = 2
      "00010" when "010101001000111", -- t[10823] = 2
      "00010" when "010101001001000", -- t[10824] = 2
      "00010" when "010101001001001", -- t[10825] = 2
      "00010" when "010101001001010", -- t[10826] = 2
      "00010" when "010101001001011", -- t[10827] = 2
      "00010" when "010101001001100", -- t[10828] = 2
      "00010" when "010101001001101", -- t[10829] = 2
      "00010" when "010101001001110", -- t[10830] = 2
      "00010" when "010101001001111", -- t[10831] = 2
      "00010" when "010101001010000", -- t[10832] = 2
      "00010" when "010101001010001", -- t[10833] = 2
      "00010" when "010101001010010", -- t[10834] = 2
      "00010" when "010101001010011", -- t[10835] = 2
      "00010" when "010101001010100", -- t[10836] = 2
      "00010" when "010101001010101", -- t[10837] = 2
      "00010" when "010101001010110", -- t[10838] = 2
      "00010" when "010101001010111", -- t[10839] = 2
      "00010" when "010101001011000", -- t[10840] = 2
      "00010" when "010101001011001", -- t[10841] = 2
      "00010" when "010101001011010", -- t[10842] = 2
      "00010" when "010101001011011", -- t[10843] = 2
      "00010" when "010101001011100", -- t[10844] = 2
      "00010" when "010101001011101", -- t[10845] = 2
      "00010" when "010101001011110", -- t[10846] = 2
      "00010" when "010101001011111", -- t[10847] = 2
      "00010" when "010101001100000", -- t[10848] = 2
      "00010" when "010101001100001", -- t[10849] = 2
      "00010" when "010101001100010", -- t[10850] = 2
      "00010" when "010101001100011", -- t[10851] = 2
      "00010" when "010101001100100", -- t[10852] = 2
      "00010" when "010101001100101", -- t[10853] = 2
      "00010" when "010101001100110", -- t[10854] = 2
      "00010" when "010101001100111", -- t[10855] = 2
      "00010" when "010101001101000", -- t[10856] = 2
      "00010" when "010101001101001", -- t[10857] = 2
      "00010" when "010101001101010", -- t[10858] = 2
      "00010" when "010101001101011", -- t[10859] = 2
      "00010" when "010101001101100", -- t[10860] = 2
      "00010" when "010101001101101", -- t[10861] = 2
      "00010" when "010101001101110", -- t[10862] = 2
      "00010" when "010101001101111", -- t[10863] = 2
      "00010" when "010101001110000", -- t[10864] = 2
      "00010" when "010101001110001", -- t[10865] = 2
      "00010" when "010101001110010", -- t[10866] = 2
      "00010" when "010101001110011", -- t[10867] = 2
      "00010" when "010101001110100", -- t[10868] = 2
      "00010" when "010101001110101", -- t[10869] = 2
      "00010" when "010101001110110", -- t[10870] = 2
      "00010" when "010101001110111", -- t[10871] = 2
      "00010" when "010101001111000", -- t[10872] = 2
      "00010" when "010101001111001", -- t[10873] = 2
      "00010" when "010101001111010", -- t[10874] = 2
      "00010" when "010101001111011", -- t[10875] = 2
      "00010" when "010101001111100", -- t[10876] = 2
      "00010" when "010101001111101", -- t[10877] = 2
      "00010" when "010101001111110", -- t[10878] = 2
      "00010" when "010101001111111", -- t[10879] = 2
      "00010" when "010101010000000", -- t[10880] = 2
      "00010" when "010101010000001", -- t[10881] = 2
      "00010" when "010101010000010", -- t[10882] = 2
      "00010" when "010101010000011", -- t[10883] = 2
      "00010" when "010101010000100", -- t[10884] = 2
      "00010" when "010101010000101", -- t[10885] = 2
      "00010" when "010101010000110", -- t[10886] = 2
      "00010" when "010101010000111", -- t[10887] = 2
      "00010" when "010101010001000", -- t[10888] = 2
      "00010" when "010101010001001", -- t[10889] = 2
      "00010" when "010101010001010", -- t[10890] = 2
      "00010" when "010101010001011", -- t[10891] = 2
      "00010" when "010101010001100", -- t[10892] = 2
      "00010" when "010101010001101", -- t[10893] = 2
      "00010" when "010101010001110", -- t[10894] = 2
      "00010" when "010101010001111", -- t[10895] = 2
      "00010" when "010101010010000", -- t[10896] = 2
      "00010" when "010101010010001", -- t[10897] = 2
      "00010" when "010101010010010", -- t[10898] = 2
      "00010" when "010101010010011", -- t[10899] = 2
      "00010" when "010101010010100", -- t[10900] = 2
      "00010" when "010101010010101", -- t[10901] = 2
      "00010" when "010101010010110", -- t[10902] = 2
      "00010" when "010101010010111", -- t[10903] = 2
      "00010" when "010101010011000", -- t[10904] = 2
      "00010" when "010101010011001", -- t[10905] = 2
      "00010" when "010101010011010", -- t[10906] = 2
      "00010" when "010101010011011", -- t[10907] = 2
      "00010" when "010101010011100", -- t[10908] = 2
      "00010" when "010101010011101", -- t[10909] = 2
      "00010" when "010101010011110", -- t[10910] = 2
      "00010" when "010101010011111", -- t[10911] = 2
      "00010" when "010101010100000", -- t[10912] = 2
      "00010" when "010101010100001", -- t[10913] = 2
      "00010" when "010101010100010", -- t[10914] = 2
      "00010" when "010101010100011", -- t[10915] = 2
      "00010" when "010101010100100", -- t[10916] = 2
      "00010" when "010101010100101", -- t[10917] = 2
      "00010" when "010101010100110", -- t[10918] = 2
      "00010" when "010101010100111", -- t[10919] = 2
      "00010" when "010101010101000", -- t[10920] = 2
      "00010" when "010101010101001", -- t[10921] = 2
      "00010" when "010101010101010", -- t[10922] = 2
      "00010" when "010101010101011", -- t[10923] = 2
      "00010" when "010101010101100", -- t[10924] = 2
      "00010" when "010101010101101", -- t[10925] = 2
      "00010" when "010101010101110", -- t[10926] = 2
      "00010" when "010101010101111", -- t[10927] = 2
      "00010" when "010101010110000", -- t[10928] = 2
      "00010" when "010101010110001", -- t[10929] = 2
      "00010" when "010101010110010", -- t[10930] = 2
      "00010" when "010101010110011", -- t[10931] = 2
      "00010" when "010101010110100", -- t[10932] = 2
      "00010" when "010101010110101", -- t[10933] = 2
      "00010" when "010101010110110", -- t[10934] = 2
      "00010" when "010101010110111", -- t[10935] = 2
      "00010" when "010101010111000", -- t[10936] = 2
      "00010" when "010101010111001", -- t[10937] = 2
      "00010" when "010101010111010", -- t[10938] = 2
      "00010" when "010101010111011", -- t[10939] = 2
      "00010" when "010101010111100", -- t[10940] = 2
      "00010" when "010101010111101", -- t[10941] = 2
      "00010" when "010101010111110", -- t[10942] = 2
      "00010" when "010101010111111", -- t[10943] = 2
      "00010" when "010101011000000", -- t[10944] = 2
      "00010" when "010101011000001", -- t[10945] = 2
      "00010" when "010101011000010", -- t[10946] = 2
      "00010" when "010101011000011", -- t[10947] = 2
      "00010" when "010101011000100", -- t[10948] = 2
      "00010" when "010101011000101", -- t[10949] = 2
      "00010" when "010101011000110", -- t[10950] = 2
      "00010" when "010101011000111", -- t[10951] = 2
      "00010" when "010101011001000", -- t[10952] = 2
      "00010" when "010101011001001", -- t[10953] = 2
      "00010" when "010101011001010", -- t[10954] = 2
      "00010" when "010101011001011", -- t[10955] = 2
      "00010" when "010101011001100", -- t[10956] = 2
      "00010" when "010101011001101", -- t[10957] = 2
      "00010" when "010101011001110", -- t[10958] = 2
      "00010" when "010101011001111", -- t[10959] = 2
      "00010" when "010101011010000", -- t[10960] = 2
      "00010" when "010101011010001", -- t[10961] = 2
      "00010" when "010101011010010", -- t[10962] = 2
      "00010" when "010101011010011", -- t[10963] = 2
      "00010" when "010101011010100", -- t[10964] = 2
      "00010" when "010101011010101", -- t[10965] = 2
      "00010" when "010101011010110", -- t[10966] = 2
      "00010" when "010101011010111", -- t[10967] = 2
      "00010" when "010101011011000", -- t[10968] = 2
      "00010" when "010101011011001", -- t[10969] = 2
      "00010" when "010101011011010", -- t[10970] = 2
      "00010" when "010101011011011", -- t[10971] = 2
      "00010" when "010101011011100", -- t[10972] = 2
      "00010" when "010101011011101", -- t[10973] = 2
      "00010" when "010101011011110", -- t[10974] = 2
      "00010" when "010101011011111", -- t[10975] = 2
      "00010" when "010101011100000", -- t[10976] = 2
      "00010" when "010101011100001", -- t[10977] = 2
      "00010" when "010101011100010", -- t[10978] = 2
      "00010" when "010101011100011", -- t[10979] = 2
      "00010" when "010101011100100", -- t[10980] = 2
      "00010" when "010101011100101", -- t[10981] = 2
      "00010" when "010101011100110", -- t[10982] = 2
      "00010" when "010101011100111", -- t[10983] = 2
      "00010" when "010101011101000", -- t[10984] = 2
      "00010" when "010101011101001", -- t[10985] = 2
      "00010" when "010101011101010", -- t[10986] = 2
      "00010" when "010101011101011", -- t[10987] = 2
      "00010" when "010101011101100", -- t[10988] = 2
      "00010" when "010101011101101", -- t[10989] = 2
      "00010" when "010101011101110", -- t[10990] = 2
      "00010" when "010101011101111", -- t[10991] = 2
      "00010" when "010101011110000", -- t[10992] = 2
      "00010" when "010101011110001", -- t[10993] = 2
      "00010" when "010101011110010", -- t[10994] = 2
      "00010" when "010101011110011", -- t[10995] = 2
      "00010" when "010101011110100", -- t[10996] = 2
      "00010" when "010101011110101", -- t[10997] = 2
      "00010" when "010101011110110", -- t[10998] = 2
      "00010" when "010101011110111", -- t[10999] = 2
      "00010" when "010101011111000", -- t[11000] = 2
      "00010" when "010101011111001", -- t[11001] = 2
      "00010" when "010101011111010", -- t[11002] = 2
      "00010" when "010101011111011", -- t[11003] = 2
      "00010" when "010101011111100", -- t[11004] = 2
      "00010" when "010101011111101", -- t[11005] = 2
      "00010" when "010101011111110", -- t[11006] = 2
      "00010" when "010101011111111", -- t[11007] = 2
      "00010" when "010101100000000", -- t[11008] = 2
      "00010" when "010101100000001", -- t[11009] = 2
      "00010" when "010101100000010", -- t[11010] = 2
      "00010" when "010101100000011", -- t[11011] = 2
      "00010" when "010101100000100", -- t[11012] = 2
      "00010" when "010101100000101", -- t[11013] = 2
      "00010" when "010101100000110", -- t[11014] = 2
      "00010" when "010101100000111", -- t[11015] = 2
      "00010" when "010101100001000", -- t[11016] = 2
      "00010" when "010101100001001", -- t[11017] = 2
      "00010" when "010101100001010", -- t[11018] = 2
      "00010" when "010101100001011", -- t[11019] = 2
      "00010" when "010101100001100", -- t[11020] = 2
      "00010" when "010101100001101", -- t[11021] = 2
      "00010" when "010101100001110", -- t[11022] = 2
      "00010" when "010101100001111", -- t[11023] = 2
      "00010" when "010101100010000", -- t[11024] = 2
      "00010" when "010101100010001", -- t[11025] = 2
      "00010" when "010101100010010", -- t[11026] = 2
      "00010" when "010101100010011", -- t[11027] = 2
      "00010" when "010101100010100", -- t[11028] = 2
      "00010" when "010101100010101", -- t[11029] = 2
      "00010" when "010101100010110", -- t[11030] = 2
      "00010" when "010101100010111", -- t[11031] = 2
      "00010" when "010101100011000", -- t[11032] = 2
      "00010" when "010101100011001", -- t[11033] = 2
      "00010" when "010101100011010", -- t[11034] = 2
      "00010" when "010101100011011", -- t[11035] = 2
      "00010" when "010101100011100", -- t[11036] = 2
      "00010" when "010101100011101", -- t[11037] = 2
      "00010" when "010101100011110", -- t[11038] = 2
      "00010" when "010101100011111", -- t[11039] = 2
      "00010" when "010101100100000", -- t[11040] = 2
      "00010" when "010101100100001", -- t[11041] = 2
      "00010" when "010101100100010", -- t[11042] = 2
      "00010" when "010101100100011", -- t[11043] = 2
      "00010" when "010101100100100", -- t[11044] = 2
      "00010" when "010101100100101", -- t[11045] = 2
      "00010" when "010101100100110", -- t[11046] = 2
      "00010" when "010101100100111", -- t[11047] = 2
      "00010" when "010101100101000", -- t[11048] = 2
      "00010" when "010101100101001", -- t[11049] = 2
      "00010" when "010101100101010", -- t[11050] = 2
      "00010" when "010101100101011", -- t[11051] = 2
      "00010" when "010101100101100", -- t[11052] = 2
      "00010" when "010101100101101", -- t[11053] = 2
      "00010" when "010101100101110", -- t[11054] = 2
      "00010" when "010101100101111", -- t[11055] = 2
      "00010" when "010101100110000", -- t[11056] = 2
      "00010" when "010101100110001", -- t[11057] = 2
      "00010" when "010101100110010", -- t[11058] = 2
      "00010" when "010101100110011", -- t[11059] = 2
      "00010" when "010101100110100", -- t[11060] = 2
      "00010" when "010101100110101", -- t[11061] = 2
      "00010" when "010101100110110", -- t[11062] = 2
      "00010" when "010101100110111", -- t[11063] = 2
      "00010" when "010101100111000", -- t[11064] = 2
      "00010" when "010101100111001", -- t[11065] = 2
      "00010" when "010101100111010", -- t[11066] = 2
      "00010" when "010101100111011", -- t[11067] = 2
      "00010" when "010101100111100", -- t[11068] = 2
      "00010" when "010101100111101", -- t[11069] = 2
      "00010" when "010101100111110", -- t[11070] = 2
      "00010" when "010101100111111", -- t[11071] = 2
      "00010" when "010101101000000", -- t[11072] = 2
      "00010" when "010101101000001", -- t[11073] = 2
      "00010" when "010101101000010", -- t[11074] = 2
      "00010" when "010101101000011", -- t[11075] = 2
      "00010" when "010101101000100", -- t[11076] = 2
      "00010" when "010101101000101", -- t[11077] = 2
      "00010" when "010101101000110", -- t[11078] = 2
      "00010" when "010101101000111", -- t[11079] = 2
      "00010" when "010101101001000", -- t[11080] = 2
      "00010" when "010101101001001", -- t[11081] = 2
      "00010" when "010101101001010", -- t[11082] = 2
      "00010" when "010101101001011", -- t[11083] = 2
      "00010" when "010101101001100", -- t[11084] = 2
      "00010" when "010101101001101", -- t[11085] = 2
      "00010" when "010101101001110", -- t[11086] = 2
      "00010" when "010101101001111", -- t[11087] = 2
      "00010" when "010101101010000", -- t[11088] = 2
      "00010" when "010101101010001", -- t[11089] = 2
      "00010" when "010101101010010", -- t[11090] = 2
      "00010" when "010101101010011", -- t[11091] = 2
      "00010" when "010101101010100", -- t[11092] = 2
      "00010" when "010101101010101", -- t[11093] = 2
      "00010" when "010101101010110", -- t[11094] = 2
      "00010" when "010101101010111", -- t[11095] = 2
      "00010" when "010101101011000", -- t[11096] = 2
      "00010" when "010101101011001", -- t[11097] = 2
      "00010" when "010101101011010", -- t[11098] = 2
      "00010" when "010101101011011", -- t[11099] = 2
      "00010" when "010101101011100", -- t[11100] = 2
      "00010" when "010101101011101", -- t[11101] = 2
      "00010" when "010101101011110", -- t[11102] = 2
      "00010" when "010101101011111", -- t[11103] = 2
      "00010" when "010101101100000", -- t[11104] = 2
      "00010" when "010101101100001", -- t[11105] = 2
      "00010" when "010101101100010", -- t[11106] = 2
      "00010" when "010101101100011", -- t[11107] = 2
      "00010" when "010101101100100", -- t[11108] = 2
      "00010" when "010101101100101", -- t[11109] = 2
      "00010" when "010101101100110", -- t[11110] = 2
      "00010" when "010101101100111", -- t[11111] = 2
      "00010" when "010101101101000", -- t[11112] = 2
      "00010" when "010101101101001", -- t[11113] = 2
      "00010" when "010101101101010", -- t[11114] = 2
      "00010" when "010101101101011", -- t[11115] = 2
      "00010" when "010101101101100", -- t[11116] = 2
      "00010" when "010101101101101", -- t[11117] = 2
      "00010" when "010101101101110", -- t[11118] = 2
      "00010" when "010101101101111", -- t[11119] = 2
      "00010" when "010101101110000", -- t[11120] = 2
      "00010" when "010101101110001", -- t[11121] = 2
      "00010" when "010101101110010", -- t[11122] = 2
      "00010" when "010101101110011", -- t[11123] = 2
      "00010" when "010101101110100", -- t[11124] = 2
      "00010" when "010101101110101", -- t[11125] = 2
      "00010" when "010101101110110", -- t[11126] = 2
      "00010" when "010101101110111", -- t[11127] = 2
      "00010" when "010101101111000", -- t[11128] = 2
      "00010" when "010101101111001", -- t[11129] = 2
      "00010" when "010101101111010", -- t[11130] = 2
      "00010" when "010101101111011", -- t[11131] = 2
      "00010" when "010101101111100", -- t[11132] = 2
      "00010" when "010101101111101", -- t[11133] = 2
      "00010" when "010101101111110", -- t[11134] = 2
      "00010" when "010101101111111", -- t[11135] = 2
      "00010" when "010101110000000", -- t[11136] = 2
      "00010" when "010101110000001", -- t[11137] = 2
      "00010" when "010101110000010", -- t[11138] = 2
      "00010" when "010101110000011", -- t[11139] = 2
      "00010" when "010101110000100", -- t[11140] = 2
      "00010" when "010101110000101", -- t[11141] = 2
      "00010" when "010101110000110", -- t[11142] = 2
      "00010" when "010101110000111", -- t[11143] = 2
      "00010" when "010101110001000", -- t[11144] = 2
      "00010" when "010101110001001", -- t[11145] = 2
      "00010" when "010101110001010", -- t[11146] = 2
      "00010" when "010101110001011", -- t[11147] = 2
      "00010" when "010101110001100", -- t[11148] = 2
      "00010" when "010101110001101", -- t[11149] = 2
      "00010" when "010101110001110", -- t[11150] = 2
      "00010" when "010101110001111", -- t[11151] = 2
      "00010" when "010101110010000", -- t[11152] = 2
      "00010" when "010101110010001", -- t[11153] = 2
      "00010" when "010101110010010", -- t[11154] = 2
      "00010" when "010101110010011", -- t[11155] = 2
      "00010" when "010101110010100", -- t[11156] = 2
      "00010" when "010101110010101", -- t[11157] = 2
      "00010" when "010101110010110", -- t[11158] = 2
      "00010" when "010101110010111", -- t[11159] = 2
      "00010" when "010101110011000", -- t[11160] = 2
      "00010" when "010101110011001", -- t[11161] = 2
      "00010" when "010101110011010", -- t[11162] = 2
      "00010" when "010101110011011", -- t[11163] = 2
      "00010" when "010101110011100", -- t[11164] = 2
      "00010" when "010101110011101", -- t[11165] = 2
      "00010" when "010101110011110", -- t[11166] = 2
      "00010" when "010101110011111", -- t[11167] = 2
      "00010" when "010101110100000", -- t[11168] = 2
      "00010" when "010101110100001", -- t[11169] = 2
      "00010" when "010101110100010", -- t[11170] = 2
      "00010" when "010101110100011", -- t[11171] = 2
      "00010" when "010101110100100", -- t[11172] = 2
      "00010" when "010101110100101", -- t[11173] = 2
      "00010" when "010101110100110", -- t[11174] = 2
      "00010" when "010101110100111", -- t[11175] = 2
      "00010" when "010101110101000", -- t[11176] = 2
      "00010" when "010101110101001", -- t[11177] = 2
      "00010" when "010101110101010", -- t[11178] = 2
      "00010" when "010101110101011", -- t[11179] = 2
      "00010" when "010101110101100", -- t[11180] = 2
      "00010" when "010101110101101", -- t[11181] = 2
      "00010" when "010101110101110", -- t[11182] = 2
      "00010" when "010101110101111", -- t[11183] = 2
      "00010" when "010101110110000", -- t[11184] = 2
      "00010" when "010101110110001", -- t[11185] = 2
      "00010" when "010101110110010", -- t[11186] = 2
      "00010" when "010101110110011", -- t[11187] = 2
      "00010" when "010101110110100", -- t[11188] = 2
      "00010" when "010101110110101", -- t[11189] = 2
      "00010" when "010101110110110", -- t[11190] = 2
      "00010" when "010101110110111", -- t[11191] = 2
      "00010" when "010101110111000", -- t[11192] = 2
      "00010" when "010101110111001", -- t[11193] = 2
      "00010" when "010101110111010", -- t[11194] = 2
      "00010" when "010101110111011", -- t[11195] = 2
      "00010" when "010101110111100", -- t[11196] = 2
      "00010" when "010101110111101", -- t[11197] = 2
      "00010" when "010101110111110", -- t[11198] = 2
      "00010" when "010101110111111", -- t[11199] = 2
      "00010" when "010101111000000", -- t[11200] = 2
      "00010" when "010101111000001", -- t[11201] = 2
      "00010" when "010101111000010", -- t[11202] = 2
      "00010" when "010101111000011", -- t[11203] = 2
      "00010" when "010101111000100", -- t[11204] = 2
      "00010" when "010101111000101", -- t[11205] = 2
      "00010" when "010101111000110", -- t[11206] = 2
      "00010" when "010101111000111", -- t[11207] = 2
      "00010" when "010101111001000", -- t[11208] = 2
      "00010" when "010101111001001", -- t[11209] = 2
      "00010" when "010101111001010", -- t[11210] = 2
      "00010" when "010101111001011", -- t[11211] = 2
      "00010" when "010101111001100", -- t[11212] = 2
      "00010" when "010101111001101", -- t[11213] = 2
      "00010" when "010101111001110", -- t[11214] = 2
      "00010" when "010101111001111", -- t[11215] = 2
      "00010" when "010101111010000", -- t[11216] = 2
      "00010" when "010101111010001", -- t[11217] = 2
      "00010" when "010101111010010", -- t[11218] = 2
      "00010" when "010101111010011", -- t[11219] = 2
      "00010" when "010101111010100", -- t[11220] = 2
      "00010" when "010101111010101", -- t[11221] = 2
      "00010" when "010101111010110", -- t[11222] = 2
      "00010" when "010101111010111", -- t[11223] = 2
      "00010" when "010101111011000", -- t[11224] = 2
      "00010" when "010101111011001", -- t[11225] = 2
      "00010" when "010101111011010", -- t[11226] = 2
      "00010" when "010101111011011", -- t[11227] = 2
      "00010" when "010101111011100", -- t[11228] = 2
      "00010" when "010101111011101", -- t[11229] = 2
      "00010" when "010101111011110", -- t[11230] = 2
      "00010" when "010101111011111", -- t[11231] = 2
      "00010" when "010101111100000", -- t[11232] = 2
      "00010" when "010101111100001", -- t[11233] = 2
      "00010" when "010101111100010", -- t[11234] = 2
      "00010" when "010101111100011", -- t[11235] = 2
      "00010" when "010101111100100", -- t[11236] = 2
      "00010" when "010101111100101", -- t[11237] = 2
      "00010" when "010101111100110", -- t[11238] = 2
      "00010" when "010101111100111", -- t[11239] = 2
      "00010" when "010101111101000", -- t[11240] = 2
      "00010" when "010101111101001", -- t[11241] = 2
      "00010" when "010101111101010", -- t[11242] = 2
      "00010" when "010101111101011", -- t[11243] = 2
      "00010" when "010101111101100", -- t[11244] = 2
      "00010" when "010101111101101", -- t[11245] = 2
      "00010" when "010101111101110", -- t[11246] = 2
      "00010" when "010101111101111", -- t[11247] = 2
      "00010" when "010101111110000", -- t[11248] = 2
      "00010" when "010101111110001", -- t[11249] = 2
      "00010" when "010101111110010", -- t[11250] = 2
      "00010" when "010101111110011", -- t[11251] = 2
      "00010" when "010101111110100", -- t[11252] = 2
      "00010" when "010101111110101", -- t[11253] = 2
      "00010" when "010101111110110", -- t[11254] = 2
      "00010" when "010101111110111", -- t[11255] = 2
      "00010" when "010101111111000", -- t[11256] = 2
      "00010" when "010101111111001", -- t[11257] = 2
      "00010" when "010101111111010", -- t[11258] = 2
      "00010" when "010101111111011", -- t[11259] = 2
      "00010" when "010101111111100", -- t[11260] = 2
      "00010" when "010101111111101", -- t[11261] = 2
      "00010" when "010101111111110", -- t[11262] = 2
      "00010" when "010101111111111", -- t[11263] = 2
      "00010" when "010110000000000", -- t[11264] = 2
      "00010" when "010110000000001", -- t[11265] = 2
      "00010" when "010110000000010", -- t[11266] = 2
      "00010" when "010110000000011", -- t[11267] = 2
      "00010" when "010110000000100", -- t[11268] = 2
      "00010" when "010110000000101", -- t[11269] = 2
      "00010" when "010110000000110", -- t[11270] = 2
      "00010" when "010110000000111", -- t[11271] = 2
      "00010" when "010110000001000", -- t[11272] = 2
      "00010" when "010110000001001", -- t[11273] = 2
      "00010" when "010110000001010", -- t[11274] = 2
      "00010" when "010110000001011", -- t[11275] = 2
      "00010" when "010110000001100", -- t[11276] = 2
      "00010" when "010110000001101", -- t[11277] = 2
      "00010" when "010110000001110", -- t[11278] = 2
      "00010" when "010110000001111", -- t[11279] = 2
      "00010" when "010110000010000", -- t[11280] = 2
      "00010" when "010110000010001", -- t[11281] = 2
      "00010" when "010110000010010", -- t[11282] = 2
      "00010" when "010110000010011", -- t[11283] = 2
      "00010" when "010110000010100", -- t[11284] = 2
      "00010" when "010110000010101", -- t[11285] = 2
      "00010" when "010110000010110", -- t[11286] = 2
      "00010" when "010110000010111", -- t[11287] = 2
      "00010" when "010110000011000", -- t[11288] = 2
      "00010" when "010110000011001", -- t[11289] = 2
      "00010" when "010110000011010", -- t[11290] = 2
      "00010" when "010110000011011", -- t[11291] = 2
      "00010" when "010110000011100", -- t[11292] = 2
      "00010" when "010110000011101", -- t[11293] = 2
      "00010" when "010110000011110", -- t[11294] = 2
      "00010" when "010110000011111", -- t[11295] = 2
      "00010" when "010110000100000", -- t[11296] = 2
      "00010" when "010110000100001", -- t[11297] = 2
      "00010" when "010110000100010", -- t[11298] = 2
      "00010" when "010110000100011", -- t[11299] = 2
      "00010" when "010110000100100", -- t[11300] = 2
      "00010" when "010110000100101", -- t[11301] = 2
      "00010" when "010110000100110", -- t[11302] = 2
      "00010" when "010110000100111", -- t[11303] = 2
      "00010" when "010110000101000", -- t[11304] = 2
      "00010" when "010110000101001", -- t[11305] = 2
      "00010" when "010110000101010", -- t[11306] = 2
      "00010" when "010110000101011", -- t[11307] = 2
      "00010" when "010110000101100", -- t[11308] = 2
      "00010" when "010110000101101", -- t[11309] = 2
      "00010" when "010110000101110", -- t[11310] = 2
      "00010" when "010110000101111", -- t[11311] = 2
      "00010" when "010110000110000", -- t[11312] = 2
      "00010" when "010110000110001", -- t[11313] = 2
      "00010" when "010110000110010", -- t[11314] = 2
      "00010" when "010110000110011", -- t[11315] = 2
      "00010" when "010110000110100", -- t[11316] = 2
      "00010" when "010110000110101", -- t[11317] = 2
      "00010" when "010110000110110", -- t[11318] = 2
      "00010" when "010110000110111", -- t[11319] = 2
      "00010" when "010110000111000", -- t[11320] = 2
      "00010" when "010110000111001", -- t[11321] = 2
      "00010" when "010110000111010", -- t[11322] = 2
      "00010" when "010110000111011", -- t[11323] = 2
      "00010" when "010110000111100", -- t[11324] = 2
      "00010" when "010110000111101", -- t[11325] = 2
      "00010" when "010110000111110", -- t[11326] = 2
      "00010" when "010110000111111", -- t[11327] = 2
      "00010" when "010110001000000", -- t[11328] = 2
      "00010" when "010110001000001", -- t[11329] = 2
      "00010" when "010110001000010", -- t[11330] = 2
      "00010" when "010110001000011", -- t[11331] = 2
      "00010" when "010110001000100", -- t[11332] = 2
      "00010" when "010110001000101", -- t[11333] = 2
      "00010" when "010110001000110", -- t[11334] = 2
      "00010" when "010110001000111", -- t[11335] = 2
      "00010" when "010110001001000", -- t[11336] = 2
      "00010" when "010110001001001", -- t[11337] = 2
      "00010" when "010110001001010", -- t[11338] = 2
      "00010" when "010110001001011", -- t[11339] = 2
      "00010" when "010110001001100", -- t[11340] = 2
      "00010" when "010110001001101", -- t[11341] = 2
      "00010" when "010110001001110", -- t[11342] = 2
      "00010" when "010110001001111", -- t[11343] = 2
      "00010" when "010110001010000", -- t[11344] = 2
      "00010" when "010110001010001", -- t[11345] = 2
      "00010" when "010110001010010", -- t[11346] = 2
      "00010" when "010110001010011", -- t[11347] = 2
      "00010" when "010110001010100", -- t[11348] = 2
      "00010" when "010110001010101", -- t[11349] = 2
      "00010" when "010110001010110", -- t[11350] = 2
      "00010" when "010110001010111", -- t[11351] = 2
      "00010" when "010110001011000", -- t[11352] = 2
      "00010" when "010110001011001", -- t[11353] = 2
      "00010" when "010110001011010", -- t[11354] = 2
      "00010" when "010110001011011", -- t[11355] = 2
      "00010" when "010110001011100", -- t[11356] = 2
      "00010" when "010110001011101", -- t[11357] = 2
      "00010" when "010110001011110", -- t[11358] = 2
      "00010" when "010110001011111", -- t[11359] = 2
      "00010" when "010110001100000", -- t[11360] = 2
      "00010" when "010110001100001", -- t[11361] = 2
      "00010" when "010110001100010", -- t[11362] = 2
      "00010" when "010110001100011", -- t[11363] = 2
      "00010" when "010110001100100", -- t[11364] = 2
      "00010" when "010110001100101", -- t[11365] = 2
      "00010" when "010110001100110", -- t[11366] = 2
      "00010" when "010110001100111", -- t[11367] = 2
      "00010" when "010110001101000", -- t[11368] = 2
      "00010" when "010110001101001", -- t[11369] = 2
      "00010" when "010110001101010", -- t[11370] = 2
      "00010" when "010110001101011", -- t[11371] = 2
      "00010" when "010110001101100", -- t[11372] = 2
      "00010" when "010110001101101", -- t[11373] = 2
      "00010" when "010110001101110", -- t[11374] = 2
      "00010" when "010110001101111", -- t[11375] = 2
      "00010" when "010110001110000", -- t[11376] = 2
      "00010" when "010110001110001", -- t[11377] = 2
      "00010" when "010110001110010", -- t[11378] = 2
      "00010" when "010110001110011", -- t[11379] = 2
      "00010" when "010110001110100", -- t[11380] = 2
      "00010" when "010110001110101", -- t[11381] = 2
      "00010" when "010110001110110", -- t[11382] = 2
      "00010" when "010110001110111", -- t[11383] = 2
      "00010" when "010110001111000", -- t[11384] = 2
      "00010" when "010110001111001", -- t[11385] = 2
      "00010" when "010110001111010", -- t[11386] = 2
      "00010" when "010110001111011", -- t[11387] = 2
      "00010" when "010110001111100", -- t[11388] = 2
      "00010" when "010110001111101", -- t[11389] = 2
      "00010" when "010110001111110", -- t[11390] = 2
      "00010" when "010110001111111", -- t[11391] = 2
      "00010" when "010110010000000", -- t[11392] = 2
      "00010" when "010110010000001", -- t[11393] = 2
      "00010" when "010110010000010", -- t[11394] = 2
      "00010" when "010110010000011", -- t[11395] = 2
      "00010" when "010110010000100", -- t[11396] = 2
      "00010" when "010110010000101", -- t[11397] = 2
      "00010" when "010110010000110", -- t[11398] = 2
      "00010" when "010110010000111", -- t[11399] = 2
      "00010" when "010110010001000", -- t[11400] = 2
      "00010" when "010110010001001", -- t[11401] = 2
      "00010" when "010110010001010", -- t[11402] = 2
      "00010" when "010110010001011", -- t[11403] = 2
      "00010" when "010110010001100", -- t[11404] = 2
      "00010" when "010110010001101", -- t[11405] = 2
      "00010" when "010110010001110", -- t[11406] = 2
      "00010" when "010110010001111", -- t[11407] = 2
      "00010" when "010110010010000", -- t[11408] = 2
      "00010" when "010110010010001", -- t[11409] = 2
      "00010" when "010110010010010", -- t[11410] = 2
      "00010" when "010110010010011", -- t[11411] = 2
      "00010" when "010110010010100", -- t[11412] = 2
      "00010" when "010110010010101", -- t[11413] = 2
      "00010" when "010110010010110", -- t[11414] = 2
      "00010" when "010110010010111", -- t[11415] = 2
      "00010" when "010110010011000", -- t[11416] = 2
      "00010" when "010110010011001", -- t[11417] = 2
      "00010" when "010110010011010", -- t[11418] = 2
      "00010" when "010110010011011", -- t[11419] = 2
      "00010" when "010110010011100", -- t[11420] = 2
      "00010" when "010110010011101", -- t[11421] = 2
      "00010" when "010110010011110", -- t[11422] = 2
      "00010" when "010110010011111", -- t[11423] = 2
      "00010" when "010110010100000", -- t[11424] = 2
      "00010" when "010110010100001", -- t[11425] = 2
      "00010" when "010110010100010", -- t[11426] = 2
      "00010" when "010110010100011", -- t[11427] = 2
      "00010" when "010110010100100", -- t[11428] = 2
      "00010" when "010110010100101", -- t[11429] = 2
      "00010" when "010110010100110", -- t[11430] = 2
      "00010" when "010110010100111", -- t[11431] = 2
      "00010" when "010110010101000", -- t[11432] = 2
      "00010" when "010110010101001", -- t[11433] = 2
      "00010" when "010110010101010", -- t[11434] = 2
      "00010" when "010110010101011", -- t[11435] = 2
      "00010" when "010110010101100", -- t[11436] = 2
      "00010" when "010110010101101", -- t[11437] = 2
      "00010" when "010110010101110", -- t[11438] = 2
      "00010" when "010110010101111", -- t[11439] = 2
      "00010" when "010110010110000", -- t[11440] = 2
      "00010" when "010110010110001", -- t[11441] = 2
      "00010" when "010110010110010", -- t[11442] = 2
      "00010" when "010110010110011", -- t[11443] = 2
      "00010" when "010110010110100", -- t[11444] = 2
      "00010" when "010110010110101", -- t[11445] = 2
      "00010" when "010110010110110", -- t[11446] = 2
      "00010" when "010110010110111", -- t[11447] = 2
      "00010" when "010110010111000", -- t[11448] = 2
      "00010" when "010110010111001", -- t[11449] = 2
      "00010" when "010110010111010", -- t[11450] = 2
      "00010" when "010110010111011", -- t[11451] = 2
      "00010" when "010110010111100", -- t[11452] = 2
      "00010" when "010110010111101", -- t[11453] = 2
      "00010" when "010110010111110", -- t[11454] = 2
      "00010" when "010110010111111", -- t[11455] = 2
      "00010" when "010110011000000", -- t[11456] = 2
      "00010" when "010110011000001", -- t[11457] = 2
      "00010" when "010110011000010", -- t[11458] = 2
      "00010" when "010110011000011", -- t[11459] = 2
      "00010" when "010110011000100", -- t[11460] = 2
      "00010" when "010110011000101", -- t[11461] = 2
      "00010" when "010110011000110", -- t[11462] = 2
      "00010" when "010110011000111", -- t[11463] = 2
      "00010" when "010110011001000", -- t[11464] = 2
      "00010" when "010110011001001", -- t[11465] = 2
      "00010" when "010110011001010", -- t[11466] = 2
      "00010" when "010110011001011", -- t[11467] = 2
      "00010" when "010110011001100", -- t[11468] = 2
      "00010" when "010110011001101", -- t[11469] = 2
      "00010" when "010110011001110", -- t[11470] = 2
      "00010" when "010110011001111", -- t[11471] = 2
      "00010" when "010110011010000", -- t[11472] = 2
      "00010" when "010110011010001", -- t[11473] = 2
      "00010" when "010110011010010", -- t[11474] = 2
      "00010" when "010110011010011", -- t[11475] = 2
      "00010" when "010110011010100", -- t[11476] = 2
      "00010" when "010110011010101", -- t[11477] = 2
      "00010" when "010110011010110", -- t[11478] = 2
      "00010" when "010110011010111", -- t[11479] = 2
      "00010" when "010110011011000", -- t[11480] = 2
      "00010" when "010110011011001", -- t[11481] = 2
      "00010" when "010110011011010", -- t[11482] = 2
      "00010" when "010110011011011", -- t[11483] = 2
      "00010" when "010110011011100", -- t[11484] = 2
      "00010" when "010110011011101", -- t[11485] = 2
      "00010" when "010110011011110", -- t[11486] = 2
      "00010" when "010110011011111", -- t[11487] = 2
      "00010" when "010110011100000", -- t[11488] = 2
      "00010" when "010110011100001", -- t[11489] = 2
      "00010" when "010110011100010", -- t[11490] = 2
      "00010" when "010110011100011", -- t[11491] = 2
      "00010" when "010110011100100", -- t[11492] = 2
      "00010" when "010110011100101", -- t[11493] = 2
      "00010" when "010110011100110", -- t[11494] = 2
      "00010" when "010110011100111", -- t[11495] = 2
      "00010" when "010110011101000", -- t[11496] = 2
      "00010" when "010110011101001", -- t[11497] = 2
      "00010" when "010110011101010", -- t[11498] = 2
      "00010" when "010110011101011", -- t[11499] = 2
      "00010" when "010110011101100", -- t[11500] = 2
      "00010" when "010110011101101", -- t[11501] = 2
      "00010" when "010110011101110", -- t[11502] = 2
      "00010" when "010110011101111", -- t[11503] = 2
      "00010" when "010110011110000", -- t[11504] = 2
      "00010" when "010110011110001", -- t[11505] = 2
      "00010" when "010110011110010", -- t[11506] = 2
      "00010" when "010110011110011", -- t[11507] = 2
      "00010" when "010110011110100", -- t[11508] = 2
      "00010" when "010110011110101", -- t[11509] = 2
      "00010" when "010110011110110", -- t[11510] = 2
      "00010" when "010110011110111", -- t[11511] = 2
      "00010" when "010110011111000", -- t[11512] = 2
      "00010" when "010110011111001", -- t[11513] = 2
      "00010" when "010110011111010", -- t[11514] = 2
      "00010" when "010110011111011", -- t[11515] = 2
      "00010" when "010110011111100", -- t[11516] = 2
      "00010" when "010110011111101", -- t[11517] = 2
      "00010" when "010110011111110", -- t[11518] = 2
      "00010" when "010110011111111", -- t[11519] = 2
      "00010" when "010110100000000", -- t[11520] = 2
      "00010" when "010110100000001", -- t[11521] = 2
      "00010" when "010110100000010", -- t[11522] = 2
      "00010" when "010110100000011", -- t[11523] = 2
      "00010" when "010110100000100", -- t[11524] = 2
      "00010" when "010110100000101", -- t[11525] = 2
      "00010" when "010110100000110", -- t[11526] = 2
      "00010" when "010110100000111", -- t[11527] = 2
      "00010" when "010110100001000", -- t[11528] = 2
      "00010" when "010110100001001", -- t[11529] = 2
      "00010" when "010110100001010", -- t[11530] = 2
      "00010" when "010110100001011", -- t[11531] = 2
      "00010" when "010110100001100", -- t[11532] = 2
      "00010" when "010110100001101", -- t[11533] = 2
      "00010" when "010110100001110", -- t[11534] = 2
      "00010" when "010110100001111", -- t[11535] = 2
      "00010" when "010110100010000", -- t[11536] = 2
      "00010" when "010110100010001", -- t[11537] = 2
      "00010" when "010110100010010", -- t[11538] = 2
      "00010" when "010110100010011", -- t[11539] = 2
      "00010" when "010110100010100", -- t[11540] = 2
      "00010" when "010110100010101", -- t[11541] = 2
      "00010" when "010110100010110", -- t[11542] = 2
      "00010" when "010110100010111", -- t[11543] = 2
      "00010" when "010110100011000", -- t[11544] = 2
      "00010" when "010110100011001", -- t[11545] = 2
      "00010" when "010110100011010", -- t[11546] = 2
      "00010" when "010110100011011", -- t[11547] = 2
      "00010" when "010110100011100", -- t[11548] = 2
      "00010" when "010110100011101", -- t[11549] = 2
      "00010" when "010110100011110", -- t[11550] = 2
      "00010" when "010110100011111", -- t[11551] = 2
      "00010" when "010110100100000", -- t[11552] = 2
      "00010" when "010110100100001", -- t[11553] = 2
      "00010" when "010110100100010", -- t[11554] = 2
      "00010" when "010110100100011", -- t[11555] = 2
      "00010" when "010110100100100", -- t[11556] = 2
      "00010" when "010110100100101", -- t[11557] = 2
      "00010" when "010110100100110", -- t[11558] = 2
      "00010" when "010110100100111", -- t[11559] = 2
      "00010" when "010110100101000", -- t[11560] = 2
      "00010" when "010110100101001", -- t[11561] = 2
      "00010" when "010110100101010", -- t[11562] = 2
      "00010" when "010110100101011", -- t[11563] = 2
      "00010" when "010110100101100", -- t[11564] = 2
      "00010" when "010110100101101", -- t[11565] = 2
      "00010" when "010110100101110", -- t[11566] = 2
      "00010" when "010110100101111", -- t[11567] = 2
      "00010" when "010110100110000", -- t[11568] = 2
      "00010" when "010110100110001", -- t[11569] = 2
      "00010" when "010110100110010", -- t[11570] = 2
      "00010" when "010110100110011", -- t[11571] = 2
      "00010" when "010110100110100", -- t[11572] = 2
      "00010" when "010110100110101", -- t[11573] = 2
      "00010" when "010110100110110", -- t[11574] = 2
      "00010" when "010110100110111", -- t[11575] = 2
      "00010" when "010110100111000", -- t[11576] = 2
      "00010" when "010110100111001", -- t[11577] = 2
      "00010" when "010110100111010", -- t[11578] = 2
      "00010" when "010110100111011", -- t[11579] = 2
      "00010" when "010110100111100", -- t[11580] = 2
      "00010" when "010110100111101", -- t[11581] = 2
      "00010" when "010110100111110", -- t[11582] = 2
      "00010" when "010110100111111", -- t[11583] = 2
      "00010" when "010110101000000", -- t[11584] = 2
      "00010" when "010110101000001", -- t[11585] = 2
      "00010" when "010110101000010", -- t[11586] = 2
      "00010" when "010110101000011", -- t[11587] = 2
      "00010" when "010110101000100", -- t[11588] = 2
      "00010" when "010110101000101", -- t[11589] = 2
      "00010" when "010110101000110", -- t[11590] = 2
      "00010" when "010110101000111", -- t[11591] = 2
      "00010" when "010110101001000", -- t[11592] = 2
      "00010" when "010110101001001", -- t[11593] = 2
      "00010" when "010110101001010", -- t[11594] = 2
      "00010" when "010110101001011", -- t[11595] = 2
      "00010" when "010110101001100", -- t[11596] = 2
      "00010" when "010110101001101", -- t[11597] = 2
      "00010" when "010110101001110", -- t[11598] = 2
      "00010" when "010110101001111", -- t[11599] = 2
      "00010" when "010110101010000", -- t[11600] = 2
      "00010" when "010110101010001", -- t[11601] = 2
      "00010" when "010110101010010", -- t[11602] = 2
      "00010" when "010110101010011", -- t[11603] = 2
      "00010" when "010110101010100", -- t[11604] = 2
      "00010" when "010110101010101", -- t[11605] = 2
      "00010" when "010110101010110", -- t[11606] = 2
      "00010" when "010110101010111", -- t[11607] = 2
      "00010" when "010110101011000", -- t[11608] = 2
      "00010" when "010110101011001", -- t[11609] = 2
      "00010" when "010110101011010", -- t[11610] = 2
      "00010" when "010110101011011", -- t[11611] = 2
      "00010" when "010110101011100", -- t[11612] = 2
      "00010" when "010110101011101", -- t[11613] = 2
      "00010" when "010110101011110", -- t[11614] = 2
      "00010" when "010110101011111", -- t[11615] = 2
      "00010" when "010110101100000", -- t[11616] = 2
      "00010" when "010110101100001", -- t[11617] = 2
      "00010" when "010110101100010", -- t[11618] = 2
      "00010" when "010110101100011", -- t[11619] = 2
      "00010" when "010110101100100", -- t[11620] = 2
      "00010" when "010110101100101", -- t[11621] = 2
      "00010" when "010110101100110", -- t[11622] = 2
      "00010" when "010110101100111", -- t[11623] = 2
      "00010" when "010110101101000", -- t[11624] = 2
      "00010" when "010110101101001", -- t[11625] = 2
      "00010" when "010110101101010", -- t[11626] = 2
      "00010" when "010110101101011", -- t[11627] = 2
      "00010" when "010110101101100", -- t[11628] = 2
      "00010" when "010110101101101", -- t[11629] = 2
      "00010" when "010110101101110", -- t[11630] = 2
      "00010" when "010110101101111", -- t[11631] = 2
      "00010" when "010110101110000", -- t[11632] = 2
      "00010" when "010110101110001", -- t[11633] = 2
      "00010" when "010110101110010", -- t[11634] = 2
      "00010" when "010110101110011", -- t[11635] = 2
      "00010" when "010110101110100", -- t[11636] = 2
      "00010" when "010110101110101", -- t[11637] = 2
      "00010" when "010110101110110", -- t[11638] = 2
      "00010" when "010110101110111", -- t[11639] = 2
      "00010" when "010110101111000", -- t[11640] = 2
      "00010" when "010110101111001", -- t[11641] = 2
      "00010" when "010110101111010", -- t[11642] = 2
      "00010" when "010110101111011", -- t[11643] = 2
      "00010" when "010110101111100", -- t[11644] = 2
      "00010" when "010110101111101", -- t[11645] = 2
      "00010" when "010110101111110", -- t[11646] = 2
      "00010" when "010110101111111", -- t[11647] = 2
      "00010" when "010110110000000", -- t[11648] = 2
      "00010" when "010110110000001", -- t[11649] = 2
      "00010" when "010110110000010", -- t[11650] = 2
      "00010" when "010110110000011", -- t[11651] = 2
      "00010" when "010110110000100", -- t[11652] = 2
      "00010" when "010110110000101", -- t[11653] = 2
      "00010" when "010110110000110", -- t[11654] = 2
      "00010" when "010110110000111", -- t[11655] = 2
      "00010" when "010110110001000", -- t[11656] = 2
      "00010" when "010110110001001", -- t[11657] = 2
      "00010" when "010110110001010", -- t[11658] = 2
      "00010" when "010110110001011", -- t[11659] = 2
      "00010" when "010110110001100", -- t[11660] = 2
      "00010" when "010110110001101", -- t[11661] = 2
      "00010" when "010110110001110", -- t[11662] = 2
      "00010" when "010110110001111", -- t[11663] = 2
      "00010" when "010110110010000", -- t[11664] = 2
      "00010" when "010110110010001", -- t[11665] = 2
      "00010" when "010110110010010", -- t[11666] = 2
      "00010" when "010110110010011", -- t[11667] = 2
      "00010" when "010110110010100", -- t[11668] = 2
      "00010" when "010110110010101", -- t[11669] = 2
      "00010" when "010110110010110", -- t[11670] = 2
      "00010" when "010110110010111", -- t[11671] = 2
      "00010" when "010110110011000", -- t[11672] = 2
      "00010" when "010110110011001", -- t[11673] = 2
      "00010" when "010110110011010", -- t[11674] = 2
      "00010" when "010110110011011", -- t[11675] = 2
      "00010" when "010110110011100", -- t[11676] = 2
      "00010" when "010110110011101", -- t[11677] = 2
      "00010" when "010110110011110", -- t[11678] = 2
      "00010" when "010110110011111", -- t[11679] = 2
      "00010" when "010110110100000", -- t[11680] = 2
      "00010" when "010110110100001", -- t[11681] = 2
      "00010" when "010110110100010", -- t[11682] = 2
      "00010" when "010110110100011", -- t[11683] = 2
      "00010" when "010110110100100", -- t[11684] = 2
      "00010" when "010110110100101", -- t[11685] = 2
      "00010" when "010110110100110", -- t[11686] = 2
      "00010" when "010110110100111", -- t[11687] = 2
      "00010" when "010110110101000", -- t[11688] = 2
      "00010" when "010110110101001", -- t[11689] = 2
      "00010" when "010110110101010", -- t[11690] = 2
      "00010" when "010110110101011", -- t[11691] = 2
      "00010" when "010110110101100", -- t[11692] = 2
      "00010" when "010110110101101", -- t[11693] = 2
      "00010" when "010110110101110", -- t[11694] = 2
      "00010" when "010110110101111", -- t[11695] = 2
      "00010" when "010110110110000", -- t[11696] = 2
      "00010" when "010110110110001", -- t[11697] = 2
      "00010" when "010110110110010", -- t[11698] = 2
      "00010" when "010110110110011", -- t[11699] = 2
      "00010" when "010110110110100", -- t[11700] = 2
      "00010" when "010110110110101", -- t[11701] = 2
      "00010" when "010110110110110", -- t[11702] = 2
      "00010" when "010110110110111", -- t[11703] = 2
      "00010" when "010110110111000", -- t[11704] = 2
      "00010" when "010110110111001", -- t[11705] = 2
      "00010" when "010110110111010", -- t[11706] = 2
      "00010" when "010110110111011", -- t[11707] = 2
      "00010" when "010110110111100", -- t[11708] = 2
      "00010" when "010110110111101", -- t[11709] = 2
      "00010" when "010110110111110", -- t[11710] = 2
      "00010" when "010110110111111", -- t[11711] = 2
      "00010" when "010110111000000", -- t[11712] = 2
      "00010" when "010110111000001", -- t[11713] = 2
      "00010" when "010110111000010", -- t[11714] = 2
      "00010" when "010110111000011", -- t[11715] = 2
      "00010" when "010110111000100", -- t[11716] = 2
      "00010" when "010110111000101", -- t[11717] = 2
      "00010" when "010110111000110", -- t[11718] = 2
      "00010" when "010110111000111", -- t[11719] = 2
      "00010" when "010110111001000", -- t[11720] = 2
      "00010" when "010110111001001", -- t[11721] = 2
      "00010" when "010110111001010", -- t[11722] = 2
      "00010" when "010110111001011", -- t[11723] = 2
      "00010" when "010110111001100", -- t[11724] = 2
      "00010" when "010110111001101", -- t[11725] = 2
      "00010" when "010110111001110", -- t[11726] = 2
      "00010" when "010110111001111", -- t[11727] = 2
      "00010" when "010110111010000", -- t[11728] = 2
      "00010" when "010110111010001", -- t[11729] = 2
      "00010" when "010110111010010", -- t[11730] = 2
      "00010" when "010110111010011", -- t[11731] = 2
      "00010" when "010110111010100", -- t[11732] = 2
      "00010" when "010110111010101", -- t[11733] = 2
      "00010" when "010110111010110", -- t[11734] = 2
      "00010" when "010110111010111", -- t[11735] = 2
      "00010" when "010110111011000", -- t[11736] = 2
      "00010" when "010110111011001", -- t[11737] = 2
      "00010" when "010110111011010", -- t[11738] = 2
      "00010" when "010110111011011", -- t[11739] = 2
      "00010" when "010110111011100", -- t[11740] = 2
      "00010" when "010110111011101", -- t[11741] = 2
      "00010" when "010110111011110", -- t[11742] = 2
      "00010" when "010110111011111", -- t[11743] = 2
      "00010" when "010110111100000", -- t[11744] = 2
      "00010" when "010110111100001", -- t[11745] = 2
      "00010" when "010110111100010", -- t[11746] = 2
      "00010" when "010110111100011", -- t[11747] = 2
      "00010" when "010110111100100", -- t[11748] = 2
      "00010" when "010110111100101", -- t[11749] = 2
      "00010" when "010110111100110", -- t[11750] = 2
      "00010" when "010110111100111", -- t[11751] = 2
      "00010" when "010110111101000", -- t[11752] = 2
      "00010" when "010110111101001", -- t[11753] = 2
      "00010" when "010110111101010", -- t[11754] = 2
      "00010" when "010110111101011", -- t[11755] = 2
      "00010" when "010110111101100", -- t[11756] = 2
      "00010" when "010110111101101", -- t[11757] = 2
      "00010" when "010110111101110", -- t[11758] = 2
      "00010" when "010110111101111", -- t[11759] = 2
      "00010" when "010110111110000", -- t[11760] = 2
      "00010" when "010110111110001", -- t[11761] = 2
      "00010" when "010110111110010", -- t[11762] = 2
      "00010" when "010110111110011", -- t[11763] = 2
      "00010" when "010110111110100", -- t[11764] = 2
      "00010" when "010110111110101", -- t[11765] = 2
      "00010" when "010110111110110", -- t[11766] = 2
      "00010" when "010110111110111", -- t[11767] = 2
      "00010" when "010110111111000", -- t[11768] = 2
      "00010" when "010110111111001", -- t[11769] = 2
      "00010" when "010110111111010", -- t[11770] = 2
      "00010" when "010110111111011", -- t[11771] = 2
      "00010" when "010110111111100", -- t[11772] = 2
      "00010" when "010110111111101", -- t[11773] = 2
      "00010" when "010110111111110", -- t[11774] = 2
      "00010" when "010110111111111", -- t[11775] = 2
      "00010" when "010111000000000", -- t[11776] = 2
      "00010" when "010111000000001", -- t[11777] = 2
      "00010" when "010111000000010", -- t[11778] = 2
      "00010" when "010111000000011", -- t[11779] = 2
      "00010" when "010111000000100", -- t[11780] = 2
      "00010" when "010111000000101", -- t[11781] = 2
      "00010" when "010111000000110", -- t[11782] = 2
      "00010" when "010111000000111", -- t[11783] = 2
      "00010" when "010111000001000", -- t[11784] = 2
      "00010" when "010111000001001", -- t[11785] = 2
      "00010" when "010111000001010", -- t[11786] = 2
      "00010" when "010111000001011", -- t[11787] = 2
      "00010" when "010111000001100", -- t[11788] = 2
      "00010" when "010111000001101", -- t[11789] = 2
      "00010" when "010111000001110", -- t[11790] = 2
      "00010" when "010111000001111", -- t[11791] = 2
      "00010" when "010111000010000", -- t[11792] = 2
      "00010" when "010111000010001", -- t[11793] = 2
      "00010" when "010111000010010", -- t[11794] = 2
      "00010" when "010111000010011", -- t[11795] = 2
      "00010" when "010111000010100", -- t[11796] = 2
      "00010" when "010111000010101", -- t[11797] = 2
      "00010" when "010111000010110", -- t[11798] = 2
      "00010" when "010111000010111", -- t[11799] = 2
      "00010" when "010111000011000", -- t[11800] = 2
      "00010" when "010111000011001", -- t[11801] = 2
      "00010" when "010111000011010", -- t[11802] = 2
      "00010" when "010111000011011", -- t[11803] = 2
      "00010" when "010111000011100", -- t[11804] = 2
      "00010" when "010111000011101", -- t[11805] = 2
      "00010" when "010111000011110", -- t[11806] = 2
      "00010" when "010111000011111", -- t[11807] = 2
      "00010" when "010111000100000", -- t[11808] = 2
      "00010" when "010111000100001", -- t[11809] = 2
      "00010" when "010111000100010", -- t[11810] = 2
      "00010" when "010111000100011", -- t[11811] = 2
      "00010" when "010111000100100", -- t[11812] = 2
      "00010" when "010111000100101", -- t[11813] = 2
      "00010" when "010111000100110", -- t[11814] = 2
      "00010" when "010111000100111", -- t[11815] = 2
      "00010" when "010111000101000", -- t[11816] = 2
      "00010" when "010111000101001", -- t[11817] = 2
      "00010" when "010111000101010", -- t[11818] = 2
      "00010" when "010111000101011", -- t[11819] = 2
      "00010" when "010111000101100", -- t[11820] = 2
      "00010" when "010111000101101", -- t[11821] = 2
      "00010" when "010111000101110", -- t[11822] = 2
      "00010" when "010111000101111", -- t[11823] = 2
      "00010" when "010111000110000", -- t[11824] = 2
      "00010" when "010111000110001", -- t[11825] = 2
      "00010" when "010111000110010", -- t[11826] = 2
      "00010" when "010111000110011", -- t[11827] = 2
      "00010" when "010111000110100", -- t[11828] = 2
      "00010" when "010111000110101", -- t[11829] = 2
      "00010" when "010111000110110", -- t[11830] = 2
      "00010" when "010111000110111", -- t[11831] = 2
      "00010" when "010111000111000", -- t[11832] = 2
      "00010" when "010111000111001", -- t[11833] = 2
      "00010" when "010111000111010", -- t[11834] = 2
      "00010" when "010111000111011", -- t[11835] = 2
      "00010" when "010111000111100", -- t[11836] = 2
      "00010" when "010111000111101", -- t[11837] = 2
      "00010" when "010111000111110", -- t[11838] = 2
      "00010" when "010111000111111", -- t[11839] = 2
      "00010" when "010111001000000", -- t[11840] = 2
      "00010" when "010111001000001", -- t[11841] = 2
      "00010" when "010111001000010", -- t[11842] = 2
      "00010" when "010111001000011", -- t[11843] = 2
      "00010" when "010111001000100", -- t[11844] = 2
      "00010" when "010111001000101", -- t[11845] = 2
      "00010" when "010111001000110", -- t[11846] = 2
      "00010" when "010111001000111", -- t[11847] = 2
      "00010" when "010111001001000", -- t[11848] = 2
      "00010" when "010111001001001", -- t[11849] = 2
      "00010" when "010111001001010", -- t[11850] = 2
      "00010" when "010111001001011", -- t[11851] = 2
      "00010" when "010111001001100", -- t[11852] = 2
      "00010" when "010111001001101", -- t[11853] = 2
      "00010" when "010111001001110", -- t[11854] = 2
      "00010" when "010111001001111", -- t[11855] = 2
      "00010" when "010111001010000", -- t[11856] = 2
      "00010" when "010111001010001", -- t[11857] = 2
      "00010" when "010111001010010", -- t[11858] = 2
      "00010" when "010111001010011", -- t[11859] = 2
      "00010" when "010111001010100", -- t[11860] = 2
      "00010" when "010111001010101", -- t[11861] = 2
      "00010" when "010111001010110", -- t[11862] = 2
      "00010" when "010111001010111", -- t[11863] = 2
      "00011" when "010111001011000", -- t[11864] = 3
      "00011" when "010111001011001", -- t[11865] = 3
      "00011" when "010111001011010", -- t[11866] = 3
      "00011" when "010111001011011", -- t[11867] = 3
      "00011" when "010111001011100", -- t[11868] = 3
      "00011" when "010111001011101", -- t[11869] = 3
      "00011" when "010111001011110", -- t[11870] = 3
      "00011" when "010111001011111", -- t[11871] = 3
      "00011" when "010111001100000", -- t[11872] = 3
      "00011" when "010111001100001", -- t[11873] = 3
      "00011" when "010111001100010", -- t[11874] = 3
      "00011" when "010111001100011", -- t[11875] = 3
      "00011" when "010111001100100", -- t[11876] = 3
      "00011" when "010111001100101", -- t[11877] = 3
      "00011" when "010111001100110", -- t[11878] = 3
      "00011" when "010111001100111", -- t[11879] = 3
      "00011" when "010111001101000", -- t[11880] = 3
      "00011" when "010111001101001", -- t[11881] = 3
      "00011" when "010111001101010", -- t[11882] = 3
      "00011" when "010111001101011", -- t[11883] = 3
      "00011" when "010111001101100", -- t[11884] = 3
      "00011" when "010111001101101", -- t[11885] = 3
      "00011" when "010111001101110", -- t[11886] = 3
      "00011" when "010111001101111", -- t[11887] = 3
      "00011" when "010111001110000", -- t[11888] = 3
      "00011" when "010111001110001", -- t[11889] = 3
      "00011" when "010111001110010", -- t[11890] = 3
      "00011" when "010111001110011", -- t[11891] = 3
      "00011" when "010111001110100", -- t[11892] = 3
      "00011" when "010111001110101", -- t[11893] = 3
      "00011" when "010111001110110", -- t[11894] = 3
      "00011" when "010111001110111", -- t[11895] = 3
      "00011" when "010111001111000", -- t[11896] = 3
      "00011" when "010111001111001", -- t[11897] = 3
      "00011" when "010111001111010", -- t[11898] = 3
      "00011" when "010111001111011", -- t[11899] = 3
      "00011" when "010111001111100", -- t[11900] = 3
      "00011" when "010111001111101", -- t[11901] = 3
      "00011" when "010111001111110", -- t[11902] = 3
      "00011" when "010111001111111", -- t[11903] = 3
      "00011" when "010111010000000", -- t[11904] = 3
      "00011" when "010111010000001", -- t[11905] = 3
      "00011" when "010111010000010", -- t[11906] = 3
      "00011" when "010111010000011", -- t[11907] = 3
      "00011" when "010111010000100", -- t[11908] = 3
      "00011" when "010111010000101", -- t[11909] = 3
      "00011" when "010111010000110", -- t[11910] = 3
      "00011" when "010111010000111", -- t[11911] = 3
      "00011" when "010111010001000", -- t[11912] = 3
      "00011" when "010111010001001", -- t[11913] = 3
      "00011" when "010111010001010", -- t[11914] = 3
      "00011" when "010111010001011", -- t[11915] = 3
      "00011" when "010111010001100", -- t[11916] = 3
      "00011" when "010111010001101", -- t[11917] = 3
      "00011" when "010111010001110", -- t[11918] = 3
      "00011" when "010111010001111", -- t[11919] = 3
      "00011" when "010111010010000", -- t[11920] = 3
      "00011" when "010111010010001", -- t[11921] = 3
      "00011" when "010111010010010", -- t[11922] = 3
      "00011" when "010111010010011", -- t[11923] = 3
      "00011" when "010111010010100", -- t[11924] = 3
      "00011" when "010111010010101", -- t[11925] = 3
      "00011" when "010111010010110", -- t[11926] = 3
      "00011" when "010111010010111", -- t[11927] = 3
      "00011" when "010111010011000", -- t[11928] = 3
      "00011" when "010111010011001", -- t[11929] = 3
      "00011" when "010111010011010", -- t[11930] = 3
      "00011" when "010111010011011", -- t[11931] = 3
      "00011" when "010111010011100", -- t[11932] = 3
      "00011" when "010111010011101", -- t[11933] = 3
      "00011" when "010111010011110", -- t[11934] = 3
      "00011" when "010111010011111", -- t[11935] = 3
      "00011" when "010111010100000", -- t[11936] = 3
      "00011" when "010111010100001", -- t[11937] = 3
      "00011" when "010111010100010", -- t[11938] = 3
      "00011" when "010111010100011", -- t[11939] = 3
      "00011" when "010111010100100", -- t[11940] = 3
      "00011" when "010111010100101", -- t[11941] = 3
      "00011" when "010111010100110", -- t[11942] = 3
      "00011" when "010111010100111", -- t[11943] = 3
      "00011" when "010111010101000", -- t[11944] = 3
      "00011" when "010111010101001", -- t[11945] = 3
      "00011" when "010111010101010", -- t[11946] = 3
      "00011" when "010111010101011", -- t[11947] = 3
      "00011" when "010111010101100", -- t[11948] = 3
      "00011" when "010111010101101", -- t[11949] = 3
      "00011" when "010111010101110", -- t[11950] = 3
      "00011" when "010111010101111", -- t[11951] = 3
      "00011" when "010111010110000", -- t[11952] = 3
      "00011" when "010111010110001", -- t[11953] = 3
      "00011" when "010111010110010", -- t[11954] = 3
      "00011" when "010111010110011", -- t[11955] = 3
      "00011" when "010111010110100", -- t[11956] = 3
      "00011" when "010111010110101", -- t[11957] = 3
      "00011" when "010111010110110", -- t[11958] = 3
      "00011" when "010111010110111", -- t[11959] = 3
      "00011" when "010111010111000", -- t[11960] = 3
      "00011" when "010111010111001", -- t[11961] = 3
      "00011" when "010111010111010", -- t[11962] = 3
      "00011" when "010111010111011", -- t[11963] = 3
      "00011" when "010111010111100", -- t[11964] = 3
      "00011" when "010111010111101", -- t[11965] = 3
      "00011" when "010111010111110", -- t[11966] = 3
      "00011" when "010111010111111", -- t[11967] = 3
      "00011" when "010111011000000", -- t[11968] = 3
      "00011" when "010111011000001", -- t[11969] = 3
      "00011" when "010111011000010", -- t[11970] = 3
      "00011" when "010111011000011", -- t[11971] = 3
      "00011" when "010111011000100", -- t[11972] = 3
      "00011" when "010111011000101", -- t[11973] = 3
      "00011" when "010111011000110", -- t[11974] = 3
      "00011" when "010111011000111", -- t[11975] = 3
      "00011" when "010111011001000", -- t[11976] = 3
      "00011" when "010111011001001", -- t[11977] = 3
      "00011" when "010111011001010", -- t[11978] = 3
      "00011" when "010111011001011", -- t[11979] = 3
      "00011" when "010111011001100", -- t[11980] = 3
      "00011" when "010111011001101", -- t[11981] = 3
      "00011" when "010111011001110", -- t[11982] = 3
      "00011" when "010111011001111", -- t[11983] = 3
      "00011" when "010111011010000", -- t[11984] = 3
      "00011" when "010111011010001", -- t[11985] = 3
      "00011" when "010111011010010", -- t[11986] = 3
      "00011" when "010111011010011", -- t[11987] = 3
      "00011" when "010111011010100", -- t[11988] = 3
      "00011" when "010111011010101", -- t[11989] = 3
      "00011" when "010111011010110", -- t[11990] = 3
      "00011" when "010111011010111", -- t[11991] = 3
      "00011" when "010111011011000", -- t[11992] = 3
      "00011" when "010111011011001", -- t[11993] = 3
      "00011" when "010111011011010", -- t[11994] = 3
      "00011" when "010111011011011", -- t[11995] = 3
      "00011" when "010111011011100", -- t[11996] = 3
      "00011" when "010111011011101", -- t[11997] = 3
      "00011" when "010111011011110", -- t[11998] = 3
      "00011" when "010111011011111", -- t[11999] = 3
      "00011" when "010111011100000", -- t[12000] = 3
      "00011" when "010111011100001", -- t[12001] = 3
      "00011" when "010111011100010", -- t[12002] = 3
      "00011" when "010111011100011", -- t[12003] = 3
      "00011" when "010111011100100", -- t[12004] = 3
      "00011" when "010111011100101", -- t[12005] = 3
      "00011" when "010111011100110", -- t[12006] = 3
      "00011" when "010111011100111", -- t[12007] = 3
      "00011" when "010111011101000", -- t[12008] = 3
      "00011" when "010111011101001", -- t[12009] = 3
      "00011" when "010111011101010", -- t[12010] = 3
      "00011" when "010111011101011", -- t[12011] = 3
      "00011" when "010111011101100", -- t[12012] = 3
      "00011" when "010111011101101", -- t[12013] = 3
      "00011" when "010111011101110", -- t[12014] = 3
      "00011" when "010111011101111", -- t[12015] = 3
      "00011" when "010111011110000", -- t[12016] = 3
      "00011" when "010111011110001", -- t[12017] = 3
      "00011" when "010111011110010", -- t[12018] = 3
      "00011" when "010111011110011", -- t[12019] = 3
      "00011" when "010111011110100", -- t[12020] = 3
      "00011" when "010111011110101", -- t[12021] = 3
      "00011" when "010111011110110", -- t[12022] = 3
      "00011" when "010111011110111", -- t[12023] = 3
      "00011" when "010111011111000", -- t[12024] = 3
      "00011" when "010111011111001", -- t[12025] = 3
      "00011" when "010111011111010", -- t[12026] = 3
      "00011" when "010111011111011", -- t[12027] = 3
      "00011" when "010111011111100", -- t[12028] = 3
      "00011" when "010111011111101", -- t[12029] = 3
      "00011" when "010111011111110", -- t[12030] = 3
      "00011" when "010111011111111", -- t[12031] = 3
      "00011" when "010111100000000", -- t[12032] = 3
      "00011" when "010111100000001", -- t[12033] = 3
      "00011" when "010111100000010", -- t[12034] = 3
      "00011" when "010111100000011", -- t[12035] = 3
      "00011" when "010111100000100", -- t[12036] = 3
      "00011" when "010111100000101", -- t[12037] = 3
      "00011" when "010111100000110", -- t[12038] = 3
      "00011" when "010111100000111", -- t[12039] = 3
      "00011" when "010111100001000", -- t[12040] = 3
      "00011" when "010111100001001", -- t[12041] = 3
      "00011" when "010111100001010", -- t[12042] = 3
      "00011" when "010111100001011", -- t[12043] = 3
      "00011" when "010111100001100", -- t[12044] = 3
      "00011" when "010111100001101", -- t[12045] = 3
      "00011" when "010111100001110", -- t[12046] = 3
      "00011" when "010111100001111", -- t[12047] = 3
      "00011" when "010111100010000", -- t[12048] = 3
      "00011" when "010111100010001", -- t[12049] = 3
      "00011" when "010111100010010", -- t[12050] = 3
      "00011" when "010111100010011", -- t[12051] = 3
      "00011" when "010111100010100", -- t[12052] = 3
      "00011" when "010111100010101", -- t[12053] = 3
      "00011" when "010111100010110", -- t[12054] = 3
      "00011" when "010111100010111", -- t[12055] = 3
      "00011" when "010111100011000", -- t[12056] = 3
      "00011" when "010111100011001", -- t[12057] = 3
      "00011" when "010111100011010", -- t[12058] = 3
      "00011" when "010111100011011", -- t[12059] = 3
      "00011" when "010111100011100", -- t[12060] = 3
      "00011" when "010111100011101", -- t[12061] = 3
      "00011" when "010111100011110", -- t[12062] = 3
      "00011" when "010111100011111", -- t[12063] = 3
      "00011" when "010111100100000", -- t[12064] = 3
      "00011" when "010111100100001", -- t[12065] = 3
      "00011" when "010111100100010", -- t[12066] = 3
      "00011" when "010111100100011", -- t[12067] = 3
      "00011" when "010111100100100", -- t[12068] = 3
      "00011" when "010111100100101", -- t[12069] = 3
      "00011" when "010111100100110", -- t[12070] = 3
      "00011" when "010111100100111", -- t[12071] = 3
      "00011" when "010111100101000", -- t[12072] = 3
      "00011" when "010111100101001", -- t[12073] = 3
      "00011" when "010111100101010", -- t[12074] = 3
      "00011" when "010111100101011", -- t[12075] = 3
      "00011" when "010111100101100", -- t[12076] = 3
      "00011" when "010111100101101", -- t[12077] = 3
      "00011" when "010111100101110", -- t[12078] = 3
      "00011" when "010111100101111", -- t[12079] = 3
      "00011" when "010111100110000", -- t[12080] = 3
      "00011" when "010111100110001", -- t[12081] = 3
      "00011" when "010111100110010", -- t[12082] = 3
      "00011" when "010111100110011", -- t[12083] = 3
      "00011" when "010111100110100", -- t[12084] = 3
      "00011" when "010111100110101", -- t[12085] = 3
      "00011" when "010111100110110", -- t[12086] = 3
      "00011" when "010111100110111", -- t[12087] = 3
      "00011" when "010111100111000", -- t[12088] = 3
      "00011" when "010111100111001", -- t[12089] = 3
      "00011" when "010111100111010", -- t[12090] = 3
      "00011" when "010111100111011", -- t[12091] = 3
      "00011" when "010111100111100", -- t[12092] = 3
      "00011" when "010111100111101", -- t[12093] = 3
      "00011" when "010111100111110", -- t[12094] = 3
      "00011" when "010111100111111", -- t[12095] = 3
      "00011" when "010111101000000", -- t[12096] = 3
      "00011" when "010111101000001", -- t[12097] = 3
      "00011" when "010111101000010", -- t[12098] = 3
      "00011" when "010111101000011", -- t[12099] = 3
      "00011" when "010111101000100", -- t[12100] = 3
      "00011" when "010111101000101", -- t[12101] = 3
      "00011" when "010111101000110", -- t[12102] = 3
      "00011" when "010111101000111", -- t[12103] = 3
      "00011" when "010111101001000", -- t[12104] = 3
      "00011" when "010111101001001", -- t[12105] = 3
      "00011" when "010111101001010", -- t[12106] = 3
      "00011" when "010111101001011", -- t[12107] = 3
      "00011" when "010111101001100", -- t[12108] = 3
      "00011" when "010111101001101", -- t[12109] = 3
      "00011" when "010111101001110", -- t[12110] = 3
      "00011" when "010111101001111", -- t[12111] = 3
      "00011" when "010111101010000", -- t[12112] = 3
      "00011" when "010111101010001", -- t[12113] = 3
      "00011" when "010111101010010", -- t[12114] = 3
      "00011" when "010111101010011", -- t[12115] = 3
      "00011" when "010111101010100", -- t[12116] = 3
      "00011" when "010111101010101", -- t[12117] = 3
      "00011" when "010111101010110", -- t[12118] = 3
      "00011" when "010111101010111", -- t[12119] = 3
      "00011" when "010111101011000", -- t[12120] = 3
      "00011" when "010111101011001", -- t[12121] = 3
      "00011" when "010111101011010", -- t[12122] = 3
      "00011" when "010111101011011", -- t[12123] = 3
      "00011" when "010111101011100", -- t[12124] = 3
      "00011" when "010111101011101", -- t[12125] = 3
      "00011" when "010111101011110", -- t[12126] = 3
      "00011" when "010111101011111", -- t[12127] = 3
      "00011" when "010111101100000", -- t[12128] = 3
      "00011" when "010111101100001", -- t[12129] = 3
      "00011" when "010111101100010", -- t[12130] = 3
      "00011" when "010111101100011", -- t[12131] = 3
      "00011" when "010111101100100", -- t[12132] = 3
      "00011" when "010111101100101", -- t[12133] = 3
      "00011" when "010111101100110", -- t[12134] = 3
      "00011" when "010111101100111", -- t[12135] = 3
      "00011" when "010111101101000", -- t[12136] = 3
      "00011" when "010111101101001", -- t[12137] = 3
      "00011" when "010111101101010", -- t[12138] = 3
      "00011" when "010111101101011", -- t[12139] = 3
      "00011" when "010111101101100", -- t[12140] = 3
      "00011" when "010111101101101", -- t[12141] = 3
      "00011" when "010111101101110", -- t[12142] = 3
      "00011" when "010111101101111", -- t[12143] = 3
      "00011" when "010111101110000", -- t[12144] = 3
      "00011" when "010111101110001", -- t[12145] = 3
      "00011" when "010111101110010", -- t[12146] = 3
      "00011" when "010111101110011", -- t[12147] = 3
      "00011" when "010111101110100", -- t[12148] = 3
      "00011" when "010111101110101", -- t[12149] = 3
      "00011" when "010111101110110", -- t[12150] = 3
      "00011" when "010111101110111", -- t[12151] = 3
      "00011" when "010111101111000", -- t[12152] = 3
      "00011" when "010111101111001", -- t[12153] = 3
      "00011" when "010111101111010", -- t[12154] = 3
      "00011" when "010111101111011", -- t[12155] = 3
      "00011" when "010111101111100", -- t[12156] = 3
      "00011" when "010111101111101", -- t[12157] = 3
      "00011" when "010111101111110", -- t[12158] = 3
      "00011" when "010111101111111", -- t[12159] = 3
      "00011" when "010111110000000", -- t[12160] = 3
      "00011" when "010111110000001", -- t[12161] = 3
      "00011" when "010111110000010", -- t[12162] = 3
      "00011" when "010111110000011", -- t[12163] = 3
      "00011" when "010111110000100", -- t[12164] = 3
      "00011" when "010111110000101", -- t[12165] = 3
      "00011" when "010111110000110", -- t[12166] = 3
      "00011" when "010111110000111", -- t[12167] = 3
      "00011" when "010111110001000", -- t[12168] = 3
      "00011" when "010111110001001", -- t[12169] = 3
      "00011" when "010111110001010", -- t[12170] = 3
      "00011" when "010111110001011", -- t[12171] = 3
      "00011" when "010111110001100", -- t[12172] = 3
      "00011" when "010111110001101", -- t[12173] = 3
      "00011" when "010111110001110", -- t[12174] = 3
      "00011" when "010111110001111", -- t[12175] = 3
      "00011" when "010111110010000", -- t[12176] = 3
      "00011" when "010111110010001", -- t[12177] = 3
      "00011" when "010111110010010", -- t[12178] = 3
      "00011" when "010111110010011", -- t[12179] = 3
      "00011" when "010111110010100", -- t[12180] = 3
      "00011" when "010111110010101", -- t[12181] = 3
      "00011" when "010111110010110", -- t[12182] = 3
      "00011" when "010111110010111", -- t[12183] = 3
      "00011" when "010111110011000", -- t[12184] = 3
      "00011" when "010111110011001", -- t[12185] = 3
      "00011" when "010111110011010", -- t[12186] = 3
      "00011" when "010111110011011", -- t[12187] = 3
      "00011" when "010111110011100", -- t[12188] = 3
      "00011" when "010111110011101", -- t[12189] = 3
      "00011" when "010111110011110", -- t[12190] = 3
      "00011" when "010111110011111", -- t[12191] = 3
      "00011" when "010111110100000", -- t[12192] = 3
      "00011" when "010111110100001", -- t[12193] = 3
      "00011" when "010111110100010", -- t[12194] = 3
      "00011" when "010111110100011", -- t[12195] = 3
      "00011" when "010111110100100", -- t[12196] = 3
      "00011" when "010111110100101", -- t[12197] = 3
      "00011" when "010111110100110", -- t[12198] = 3
      "00011" when "010111110100111", -- t[12199] = 3
      "00011" when "010111110101000", -- t[12200] = 3
      "00011" when "010111110101001", -- t[12201] = 3
      "00011" when "010111110101010", -- t[12202] = 3
      "00011" when "010111110101011", -- t[12203] = 3
      "00011" when "010111110101100", -- t[12204] = 3
      "00011" when "010111110101101", -- t[12205] = 3
      "00011" when "010111110101110", -- t[12206] = 3
      "00011" when "010111110101111", -- t[12207] = 3
      "00011" when "010111110110000", -- t[12208] = 3
      "00011" when "010111110110001", -- t[12209] = 3
      "00011" when "010111110110010", -- t[12210] = 3
      "00011" when "010111110110011", -- t[12211] = 3
      "00011" when "010111110110100", -- t[12212] = 3
      "00011" when "010111110110101", -- t[12213] = 3
      "00011" when "010111110110110", -- t[12214] = 3
      "00011" when "010111110110111", -- t[12215] = 3
      "00011" when "010111110111000", -- t[12216] = 3
      "00011" when "010111110111001", -- t[12217] = 3
      "00011" when "010111110111010", -- t[12218] = 3
      "00011" when "010111110111011", -- t[12219] = 3
      "00011" when "010111110111100", -- t[12220] = 3
      "00011" when "010111110111101", -- t[12221] = 3
      "00011" when "010111110111110", -- t[12222] = 3
      "00011" when "010111110111111", -- t[12223] = 3
      "00011" when "010111111000000", -- t[12224] = 3
      "00011" when "010111111000001", -- t[12225] = 3
      "00011" when "010111111000010", -- t[12226] = 3
      "00011" when "010111111000011", -- t[12227] = 3
      "00011" when "010111111000100", -- t[12228] = 3
      "00011" when "010111111000101", -- t[12229] = 3
      "00011" when "010111111000110", -- t[12230] = 3
      "00011" when "010111111000111", -- t[12231] = 3
      "00011" when "010111111001000", -- t[12232] = 3
      "00011" when "010111111001001", -- t[12233] = 3
      "00011" when "010111111001010", -- t[12234] = 3
      "00011" when "010111111001011", -- t[12235] = 3
      "00011" when "010111111001100", -- t[12236] = 3
      "00011" when "010111111001101", -- t[12237] = 3
      "00011" when "010111111001110", -- t[12238] = 3
      "00011" when "010111111001111", -- t[12239] = 3
      "00011" when "010111111010000", -- t[12240] = 3
      "00011" when "010111111010001", -- t[12241] = 3
      "00011" when "010111111010010", -- t[12242] = 3
      "00011" when "010111111010011", -- t[12243] = 3
      "00011" when "010111111010100", -- t[12244] = 3
      "00011" when "010111111010101", -- t[12245] = 3
      "00011" when "010111111010110", -- t[12246] = 3
      "00011" when "010111111010111", -- t[12247] = 3
      "00011" when "010111111011000", -- t[12248] = 3
      "00011" when "010111111011001", -- t[12249] = 3
      "00011" when "010111111011010", -- t[12250] = 3
      "00011" when "010111111011011", -- t[12251] = 3
      "00011" when "010111111011100", -- t[12252] = 3
      "00011" when "010111111011101", -- t[12253] = 3
      "00011" when "010111111011110", -- t[12254] = 3
      "00011" when "010111111011111", -- t[12255] = 3
      "00011" when "010111111100000", -- t[12256] = 3
      "00011" when "010111111100001", -- t[12257] = 3
      "00011" when "010111111100010", -- t[12258] = 3
      "00011" when "010111111100011", -- t[12259] = 3
      "00011" when "010111111100100", -- t[12260] = 3
      "00011" when "010111111100101", -- t[12261] = 3
      "00011" when "010111111100110", -- t[12262] = 3
      "00011" when "010111111100111", -- t[12263] = 3
      "00011" when "010111111101000", -- t[12264] = 3
      "00011" when "010111111101001", -- t[12265] = 3
      "00011" when "010111111101010", -- t[12266] = 3
      "00011" when "010111111101011", -- t[12267] = 3
      "00011" when "010111111101100", -- t[12268] = 3
      "00011" when "010111111101101", -- t[12269] = 3
      "00011" when "010111111101110", -- t[12270] = 3
      "00011" when "010111111101111", -- t[12271] = 3
      "00011" when "010111111110000", -- t[12272] = 3
      "00011" when "010111111110001", -- t[12273] = 3
      "00011" when "010111111110010", -- t[12274] = 3
      "00011" when "010111111110011", -- t[12275] = 3
      "00011" when "010111111110100", -- t[12276] = 3
      "00011" when "010111111110101", -- t[12277] = 3
      "00011" when "010111111110110", -- t[12278] = 3
      "00011" when "010111111110111", -- t[12279] = 3
      "00011" when "010111111111000", -- t[12280] = 3
      "00011" when "010111111111001", -- t[12281] = 3
      "00011" when "010111111111010", -- t[12282] = 3
      "00011" when "010111111111011", -- t[12283] = 3
      "00011" when "010111111111100", -- t[12284] = 3
      "00011" when "010111111111101", -- t[12285] = 3
      "00011" when "010111111111110", -- t[12286] = 3
      "00011" when "010111111111111", -- t[12287] = 3
      "00011" when "011000000000000", -- t[12288] = 3
      "00011" when "011000000000001", -- t[12289] = 3
      "00011" when "011000000000010", -- t[12290] = 3
      "00011" when "011000000000011", -- t[12291] = 3
      "00011" when "011000000000100", -- t[12292] = 3
      "00011" when "011000000000101", -- t[12293] = 3
      "00011" when "011000000000110", -- t[12294] = 3
      "00011" when "011000000000111", -- t[12295] = 3
      "00011" when "011000000001000", -- t[12296] = 3
      "00011" when "011000000001001", -- t[12297] = 3
      "00011" when "011000000001010", -- t[12298] = 3
      "00011" when "011000000001011", -- t[12299] = 3
      "00011" when "011000000001100", -- t[12300] = 3
      "00011" when "011000000001101", -- t[12301] = 3
      "00011" when "011000000001110", -- t[12302] = 3
      "00011" when "011000000001111", -- t[12303] = 3
      "00011" when "011000000010000", -- t[12304] = 3
      "00011" when "011000000010001", -- t[12305] = 3
      "00011" when "011000000010010", -- t[12306] = 3
      "00011" when "011000000010011", -- t[12307] = 3
      "00011" when "011000000010100", -- t[12308] = 3
      "00011" when "011000000010101", -- t[12309] = 3
      "00011" when "011000000010110", -- t[12310] = 3
      "00011" when "011000000010111", -- t[12311] = 3
      "00011" when "011000000011000", -- t[12312] = 3
      "00011" when "011000000011001", -- t[12313] = 3
      "00011" when "011000000011010", -- t[12314] = 3
      "00011" when "011000000011011", -- t[12315] = 3
      "00011" when "011000000011100", -- t[12316] = 3
      "00011" when "011000000011101", -- t[12317] = 3
      "00011" when "011000000011110", -- t[12318] = 3
      "00011" when "011000000011111", -- t[12319] = 3
      "00011" when "011000000100000", -- t[12320] = 3
      "00011" when "011000000100001", -- t[12321] = 3
      "00011" when "011000000100010", -- t[12322] = 3
      "00011" when "011000000100011", -- t[12323] = 3
      "00011" when "011000000100100", -- t[12324] = 3
      "00011" when "011000000100101", -- t[12325] = 3
      "00011" when "011000000100110", -- t[12326] = 3
      "00011" when "011000000100111", -- t[12327] = 3
      "00011" when "011000000101000", -- t[12328] = 3
      "00011" when "011000000101001", -- t[12329] = 3
      "00011" when "011000000101010", -- t[12330] = 3
      "00011" when "011000000101011", -- t[12331] = 3
      "00011" when "011000000101100", -- t[12332] = 3
      "00011" when "011000000101101", -- t[12333] = 3
      "00011" when "011000000101110", -- t[12334] = 3
      "00011" when "011000000101111", -- t[12335] = 3
      "00011" when "011000000110000", -- t[12336] = 3
      "00011" when "011000000110001", -- t[12337] = 3
      "00011" when "011000000110010", -- t[12338] = 3
      "00011" when "011000000110011", -- t[12339] = 3
      "00011" when "011000000110100", -- t[12340] = 3
      "00011" when "011000000110101", -- t[12341] = 3
      "00011" when "011000000110110", -- t[12342] = 3
      "00011" when "011000000110111", -- t[12343] = 3
      "00011" when "011000000111000", -- t[12344] = 3
      "00011" when "011000000111001", -- t[12345] = 3
      "00011" when "011000000111010", -- t[12346] = 3
      "00011" when "011000000111011", -- t[12347] = 3
      "00011" when "011000000111100", -- t[12348] = 3
      "00011" when "011000000111101", -- t[12349] = 3
      "00011" when "011000000111110", -- t[12350] = 3
      "00011" when "011000000111111", -- t[12351] = 3
      "00011" when "011000001000000", -- t[12352] = 3
      "00011" when "011000001000001", -- t[12353] = 3
      "00011" when "011000001000010", -- t[12354] = 3
      "00011" when "011000001000011", -- t[12355] = 3
      "00011" when "011000001000100", -- t[12356] = 3
      "00011" when "011000001000101", -- t[12357] = 3
      "00011" when "011000001000110", -- t[12358] = 3
      "00011" when "011000001000111", -- t[12359] = 3
      "00011" when "011000001001000", -- t[12360] = 3
      "00011" when "011000001001001", -- t[12361] = 3
      "00011" when "011000001001010", -- t[12362] = 3
      "00011" when "011000001001011", -- t[12363] = 3
      "00011" when "011000001001100", -- t[12364] = 3
      "00011" when "011000001001101", -- t[12365] = 3
      "00011" when "011000001001110", -- t[12366] = 3
      "00011" when "011000001001111", -- t[12367] = 3
      "00011" when "011000001010000", -- t[12368] = 3
      "00011" when "011000001010001", -- t[12369] = 3
      "00011" when "011000001010010", -- t[12370] = 3
      "00011" when "011000001010011", -- t[12371] = 3
      "00011" when "011000001010100", -- t[12372] = 3
      "00011" when "011000001010101", -- t[12373] = 3
      "00011" when "011000001010110", -- t[12374] = 3
      "00011" when "011000001010111", -- t[12375] = 3
      "00011" when "011000001011000", -- t[12376] = 3
      "00011" when "011000001011001", -- t[12377] = 3
      "00011" when "011000001011010", -- t[12378] = 3
      "00011" when "011000001011011", -- t[12379] = 3
      "00011" when "011000001011100", -- t[12380] = 3
      "00011" when "011000001011101", -- t[12381] = 3
      "00011" when "011000001011110", -- t[12382] = 3
      "00011" when "011000001011111", -- t[12383] = 3
      "00011" when "011000001100000", -- t[12384] = 3
      "00011" when "011000001100001", -- t[12385] = 3
      "00011" when "011000001100010", -- t[12386] = 3
      "00011" when "011000001100011", -- t[12387] = 3
      "00011" when "011000001100100", -- t[12388] = 3
      "00011" when "011000001100101", -- t[12389] = 3
      "00011" when "011000001100110", -- t[12390] = 3
      "00011" when "011000001100111", -- t[12391] = 3
      "00011" when "011000001101000", -- t[12392] = 3
      "00011" when "011000001101001", -- t[12393] = 3
      "00011" when "011000001101010", -- t[12394] = 3
      "00011" when "011000001101011", -- t[12395] = 3
      "00011" when "011000001101100", -- t[12396] = 3
      "00011" when "011000001101101", -- t[12397] = 3
      "00011" when "011000001101110", -- t[12398] = 3
      "00011" when "011000001101111", -- t[12399] = 3
      "00011" when "011000001110000", -- t[12400] = 3
      "00011" when "011000001110001", -- t[12401] = 3
      "00011" when "011000001110010", -- t[12402] = 3
      "00011" when "011000001110011", -- t[12403] = 3
      "00011" when "011000001110100", -- t[12404] = 3
      "00011" when "011000001110101", -- t[12405] = 3
      "00011" when "011000001110110", -- t[12406] = 3
      "00011" when "011000001110111", -- t[12407] = 3
      "00011" when "011000001111000", -- t[12408] = 3
      "00011" when "011000001111001", -- t[12409] = 3
      "00011" when "011000001111010", -- t[12410] = 3
      "00011" when "011000001111011", -- t[12411] = 3
      "00011" when "011000001111100", -- t[12412] = 3
      "00011" when "011000001111101", -- t[12413] = 3
      "00011" when "011000001111110", -- t[12414] = 3
      "00011" when "011000001111111", -- t[12415] = 3
      "00011" when "011000010000000", -- t[12416] = 3
      "00011" when "011000010000001", -- t[12417] = 3
      "00011" when "011000010000010", -- t[12418] = 3
      "00011" when "011000010000011", -- t[12419] = 3
      "00011" when "011000010000100", -- t[12420] = 3
      "00011" when "011000010000101", -- t[12421] = 3
      "00011" when "011000010000110", -- t[12422] = 3
      "00011" when "011000010000111", -- t[12423] = 3
      "00011" when "011000010001000", -- t[12424] = 3
      "00011" when "011000010001001", -- t[12425] = 3
      "00011" when "011000010001010", -- t[12426] = 3
      "00011" when "011000010001011", -- t[12427] = 3
      "00011" when "011000010001100", -- t[12428] = 3
      "00011" when "011000010001101", -- t[12429] = 3
      "00011" when "011000010001110", -- t[12430] = 3
      "00011" when "011000010001111", -- t[12431] = 3
      "00011" when "011000010010000", -- t[12432] = 3
      "00011" when "011000010010001", -- t[12433] = 3
      "00011" when "011000010010010", -- t[12434] = 3
      "00011" when "011000010010011", -- t[12435] = 3
      "00011" when "011000010010100", -- t[12436] = 3
      "00011" when "011000010010101", -- t[12437] = 3
      "00011" when "011000010010110", -- t[12438] = 3
      "00011" when "011000010010111", -- t[12439] = 3
      "00011" when "011000010011000", -- t[12440] = 3
      "00011" when "011000010011001", -- t[12441] = 3
      "00011" when "011000010011010", -- t[12442] = 3
      "00011" when "011000010011011", -- t[12443] = 3
      "00011" when "011000010011100", -- t[12444] = 3
      "00011" when "011000010011101", -- t[12445] = 3
      "00011" when "011000010011110", -- t[12446] = 3
      "00011" when "011000010011111", -- t[12447] = 3
      "00011" when "011000010100000", -- t[12448] = 3
      "00011" when "011000010100001", -- t[12449] = 3
      "00011" when "011000010100010", -- t[12450] = 3
      "00011" when "011000010100011", -- t[12451] = 3
      "00011" when "011000010100100", -- t[12452] = 3
      "00011" when "011000010100101", -- t[12453] = 3
      "00011" when "011000010100110", -- t[12454] = 3
      "00011" when "011000010100111", -- t[12455] = 3
      "00011" when "011000010101000", -- t[12456] = 3
      "00011" when "011000010101001", -- t[12457] = 3
      "00011" when "011000010101010", -- t[12458] = 3
      "00011" when "011000010101011", -- t[12459] = 3
      "00011" when "011000010101100", -- t[12460] = 3
      "00011" when "011000010101101", -- t[12461] = 3
      "00011" when "011000010101110", -- t[12462] = 3
      "00011" when "011000010101111", -- t[12463] = 3
      "00011" when "011000010110000", -- t[12464] = 3
      "00011" when "011000010110001", -- t[12465] = 3
      "00011" when "011000010110010", -- t[12466] = 3
      "00011" when "011000010110011", -- t[12467] = 3
      "00011" when "011000010110100", -- t[12468] = 3
      "00011" when "011000010110101", -- t[12469] = 3
      "00011" when "011000010110110", -- t[12470] = 3
      "00011" when "011000010110111", -- t[12471] = 3
      "00011" when "011000010111000", -- t[12472] = 3
      "00011" when "011000010111001", -- t[12473] = 3
      "00011" when "011000010111010", -- t[12474] = 3
      "00011" when "011000010111011", -- t[12475] = 3
      "00011" when "011000010111100", -- t[12476] = 3
      "00011" when "011000010111101", -- t[12477] = 3
      "00011" when "011000010111110", -- t[12478] = 3
      "00011" when "011000010111111", -- t[12479] = 3
      "00011" when "011000011000000", -- t[12480] = 3
      "00011" when "011000011000001", -- t[12481] = 3
      "00011" when "011000011000010", -- t[12482] = 3
      "00011" when "011000011000011", -- t[12483] = 3
      "00011" when "011000011000100", -- t[12484] = 3
      "00011" when "011000011000101", -- t[12485] = 3
      "00011" when "011000011000110", -- t[12486] = 3
      "00011" when "011000011000111", -- t[12487] = 3
      "00011" when "011000011001000", -- t[12488] = 3
      "00011" when "011000011001001", -- t[12489] = 3
      "00011" when "011000011001010", -- t[12490] = 3
      "00011" when "011000011001011", -- t[12491] = 3
      "00011" when "011000011001100", -- t[12492] = 3
      "00011" when "011000011001101", -- t[12493] = 3
      "00011" when "011000011001110", -- t[12494] = 3
      "00011" when "011000011001111", -- t[12495] = 3
      "00011" when "011000011010000", -- t[12496] = 3
      "00011" when "011000011010001", -- t[12497] = 3
      "00011" when "011000011010010", -- t[12498] = 3
      "00011" when "011000011010011", -- t[12499] = 3
      "00011" when "011000011010100", -- t[12500] = 3
      "00011" when "011000011010101", -- t[12501] = 3
      "00011" when "011000011010110", -- t[12502] = 3
      "00011" when "011000011010111", -- t[12503] = 3
      "00011" when "011000011011000", -- t[12504] = 3
      "00011" when "011000011011001", -- t[12505] = 3
      "00011" when "011000011011010", -- t[12506] = 3
      "00011" when "011000011011011", -- t[12507] = 3
      "00011" when "011000011011100", -- t[12508] = 3
      "00011" when "011000011011101", -- t[12509] = 3
      "00011" when "011000011011110", -- t[12510] = 3
      "00011" when "011000011011111", -- t[12511] = 3
      "00011" when "011000011100000", -- t[12512] = 3
      "00011" when "011000011100001", -- t[12513] = 3
      "00011" when "011000011100010", -- t[12514] = 3
      "00011" when "011000011100011", -- t[12515] = 3
      "00011" when "011000011100100", -- t[12516] = 3
      "00011" when "011000011100101", -- t[12517] = 3
      "00011" when "011000011100110", -- t[12518] = 3
      "00011" when "011000011100111", -- t[12519] = 3
      "00011" when "011000011101000", -- t[12520] = 3
      "00011" when "011000011101001", -- t[12521] = 3
      "00011" when "011000011101010", -- t[12522] = 3
      "00011" when "011000011101011", -- t[12523] = 3
      "00011" when "011000011101100", -- t[12524] = 3
      "00011" when "011000011101101", -- t[12525] = 3
      "00011" when "011000011101110", -- t[12526] = 3
      "00011" when "011000011101111", -- t[12527] = 3
      "00011" when "011000011110000", -- t[12528] = 3
      "00011" when "011000011110001", -- t[12529] = 3
      "00011" when "011000011110010", -- t[12530] = 3
      "00011" when "011000011110011", -- t[12531] = 3
      "00011" when "011000011110100", -- t[12532] = 3
      "00011" when "011000011110101", -- t[12533] = 3
      "00011" when "011000011110110", -- t[12534] = 3
      "00011" when "011000011110111", -- t[12535] = 3
      "00011" when "011000011111000", -- t[12536] = 3
      "00011" when "011000011111001", -- t[12537] = 3
      "00011" when "011000011111010", -- t[12538] = 3
      "00011" when "011000011111011", -- t[12539] = 3
      "00011" when "011000011111100", -- t[12540] = 3
      "00011" when "011000011111101", -- t[12541] = 3
      "00011" when "011000011111110", -- t[12542] = 3
      "00011" when "011000011111111", -- t[12543] = 3
      "00011" when "011000100000000", -- t[12544] = 3
      "00011" when "011000100000001", -- t[12545] = 3
      "00011" when "011000100000010", -- t[12546] = 3
      "00011" when "011000100000011", -- t[12547] = 3
      "00011" when "011000100000100", -- t[12548] = 3
      "00011" when "011000100000101", -- t[12549] = 3
      "00011" when "011000100000110", -- t[12550] = 3
      "00011" when "011000100000111", -- t[12551] = 3
      "00011" when "011000100001000", -- t[12552] = 3
      "00011" when "011000100001001", -- t[12553] = 3
      "00011" when "011000100001010", -- t[12554] = 3
      "00011" when "011000100001011", -- t[12555] = 3
      "00011" when "011000100001100", -- t[12556] = 3
      "00011" when "011000100001101", -- t[12557] = 3
      "00011" when "011000100001110", -- t[12558] = 3
      "00011" when "011000100001111", -- t[12559] = 3
      "00011" when "011000100010000", -- t[12560] = 3
      "00011" when "011000100010001", -- t[12561] = 3
      "00011" when "011000100010010", -- t[12562] = 3
      "00011" when "011000100010011", -- t[12563] = 3
      "00011" when "011000100010100", -- t[12564] = 3
      "00011" when "011000100010101", -- t[12565] = 3
      "00011" when "011000100010110", -- t[12566] = 3
      "00011" when "011000100010111", -- t[12567] = 3
      "00011" when "011000100011000", -- t[12568] = 3
      "00011" when "011000100011001", -- t[12569] = 3
      "00011" when "011000100011010", -- t[12570] = 3
      "00011" when "011000100011011", -- t[12571] = 3
      "00011" when "011000100011100", -- t[12572] = 3
      "00011" when "011000100011101", -- t[12573] = 3
      "00011" when "011000100011110", -- t[12574] = 3
      "00011" when "011000100011111", -- t[12575] = 3
      "00011" when "011000100100000", -- t[12576] = 3
      "00011" when "011000100100001", -- t[12577] = 3
      "00011" when "011000100100010", -- t[12578] = 3
      "00011" when "011000100100011", -- t[12579] = 3
      "00011" when "011000100100100", -- t[12580] = 3
      "00011" when "011000100100101", -- t[12581] = 3
      "00011" when "011000100100110", -- t[12582] = 3
      "00011" when "011000100100111", -- t[12583] = 3
      "00011" when "011000100101000", -- t[12584] = 3
      "00011" when "011000100101001", -- t[12585] = 3
      "00011" when "011000100101010", -- t[12586] = 3
      "00011" when "011000100101011", -- t[12587] = 3
      "00011" when "011000100101100", -- t[12588] = 3
      "00011" when "011000100101101", -- t[12589] = 3
      "00011" when "011000100101110", -- t[12590] = 3
      "00011" when "011000100101111", -- t[12591] = 3
      "00011" when "011000100110000", -- t[12592] = 3
      "00011" when "011000100110001", -- t[12593] = 3
      "00011" when "011000100110010", -- t[12594] = 3
      "00011" when "011000100110011", -- t[12595] = 3
      "00011" when "011000100110100", -- t[12596] = 3
      "00011" when "011000100110101", -- t[12597] = 3
      "00011" when "011000100110110", -- t[12598] = 3
      "00011" when "011000100110111", -- t[12599] = 3
      "00011" when "011000100111000", -- t[12600] = 3
      "00011" when "011000100111001", -- t[12601] = 3
      "00011" when "011000100111010", -- t[12602] = 3
      "00011" when "011000100111011", -- t[12603] = 3
      "00011" when "011000100111100", -- t[12604] = 3
      "00011" when "011000100111101", -- t[12605] = 3
      "00011" when "011000100111110", -- t[12606] = 3
      "00011" when "011000100111111", -- t[12607] = 3
      "00011" when "011000101000000", -- t[12608] = 3
      "00011" when "011000101000001", -- t[12609] = 3
      "00011" when "011000101000010", -- t[12610] = 3
      "00011" when "011000101000011", -- t[12611] = 3
      "00011" when "011000101000100", -- t[12612] = 3
      "00011" when "011000101000101", -- t[12613] = 3
      "00011" when "011000101000110", -- t[12614] = 3
      "00011" when "011000101000111", -- t[12615] = 3
      "00011" when "011000101001000", -- t[12616] = 3
      "00011" when "011000101001001", -- t[12617] = 3
      "00011" when "011000101001010", -- t[12618] = 3
      "00011" when "011000101001011", -- t[12619] = 3
      "00011" when "011000101001100", -- t[12620] = 3
      "00011" when "011000101001101", -- t[12621] = 3
      "00011" when "011000101001110", -- t[12622] = 3
      "00011" when "011000101001111", -- t[12623] = 3
      "00011" when "011000101010000", -- t[12624] = 3
      "00011" when "011000101010001", -- t[12625] = 3
      "00011" when "011000101010010", -- t[12626] = 3
      "00011" when "011000101010011", -- t[12627] = 3
      "00011" when "011000101010100", -- t[12628] = 3
      "00011" when "011000101010101", -- t[12629] = 3
      "00011" when "011000101010110", -- t[12630] = 3
      "00011" when "011000101010111", -- t[12631] = 3
      "00011" when "011000101011000", -- t[12632] = 3
      "00011" when "011000101011001", -- t[12633] = 3
      "00011" when "011000101011010", -- t[12634] = 3
      "00011" when "011000101011011", -- t[12635] = 3
      "00011" when "011000101011100", -- t[12636] = 3
      "00011" when "011000101011101", -- t[12637] = 3
      "00011" when "011000101011110", -- t[12638] = 3
      "00011" when "011000101011111", -- t[12639] = 3
      "00011" when "011000101100000", -- t[12640] = 3
      "00011" when "011000101100001", -- t[12641] = 3
      "00011" when "011000101100010", -- t[12642] = 3
      "00011" when "011000101100011", -- t[12643] = 3
      "00011" when "011000101100100", -- t[12644] = 3
      "00011" when "011000101100101", -- t[12645] = 3
      "00011" when "011000101100110", -- t[12646] = 3
      "00011" when "011000101100111", -- t[12647] = 3
      "00011" when "011000101101000", -- t[12648] = 3
      "00011" when "011000101101001", -- t[12649] = 3
      "00011" when "011000101101010", -- t[12650] = 3
      "00011" when "011000101101011", -- t[12651] = 3
      "00011" when "011000101101100", -- t[12652] = 3
      "00011" when "011000101101101", -- t[12653] = 3
      "00011" when "011000101101110", -- t[12654] = 3
      "00011" when "011000101101111", -- t[12655] = 3
      "00011" when "011000101110000", -- t[12656] = 3
      "00011" when "011000101110001", -- t[12657] = 3
      "00011" when "011000101110010", -- t[12658] = 3
      "00011" when "011000101110011", -- t[12659] = 3
      "00011" when "011000101110100", -- t[12660] = 3
      "00011" when "011000101110101", -- t[12661] = 3
      "00011" when "011000101110110", -- t[12662] = 3
      "00011" when "011000101110111", -- t[12663] = 3
      "00011" when "011000101111000", -- t[12664] = 3
      "00011" when "011000101111001", -- t[12665] = 3
      "00011" when "011000101111010", -- t[12666] = 3
      "00011" when "011000101111011", -- t[12667] = 3
      "00011" when "011000101111100", -- t[12668] = 3
      "00011" when "011000101111101", -- t[12669] = 3
      "00011" when "011000101111110", -- t[12670] = 3
      "00011" when "011000101111111", -- t[12671] = 3
      "00011" when "011000110000000", -- t[12672] = 3
      "00011" when "011000110000001", -- t[12673] = 3
      "00011" when "011000110000010", -- t[12674] = 3
      "00011" when "011000110000011", -- t[12675] = 3
      "00011" when "011000110000100", -- t[12676] = 3
      "00011" when "011000110000101", -- t[12677] = 3
      "00011" when "011000110000110", -- t[12678] = 3
      "00011" when "011000110000111", -- t[12679] = 3
      "00011" when "011000110001000", -- t[12680] = 3
      "00011" when "011000110001001", -- t[12681] = 3
      "00011" when "011000110001010", -- t[12682] = 3
      "00011" when "011000110001011", -- t[12683] = 3
      "00011" when "011000110001100", -- t[12684] = 3
      "00011" when "011000110001101", -- t[12685] = 3
      "00011" when "011000110001110", -- t[12686] = 3
      "00011" when "011000110001111", -- t[12687] = 3
      "00011" when "011000110010000", -- t[12688] = 3
      "00011" when "011000110010001", -- t[12689] = 3
      "00011" when "011000110010010", -- t[12690] = 3
      "00011" when "011000110010011", -- t[12691] = 3
      "00011" when "011000110010100", -- t[12692] = 3
      "00011" when "011000110010101", -- t[12693] = 3
      "00011" when "011000110010110", -- t[12694] = 3
      "00011" when "011000110010111", -- t[12695] = 3
      "00011" when "011000110011000", -- t[12696] = 3
      "00011" when "011000110011001", -- t[12697] = 3
      "00011" when "011000110011010", -- t[12698] = 3
      "00011" when "011000110011011", -- t[12699] = 3
      "00011" when "011000110011100", -- t[12700] = 3
      "00011" when "011000110011101", -- t[12701] = 3
      "00011" when "011000110011110", -- t[12702] = 3
      "00011" when "011000110011111", -- t[12703] = 3
      "00011" when "011000110100000", -- t[12704] = 3
      "00011" when "011000110100001", -- t[12705] = 3
      "00011" when "011000110100010", -- t[12706] = 3
      "00011" when "011000110100011", -- t[12707] = 3
      "00011" when "011000110100100", -- t[12708] = 3
      "00011" when "011000110100101", -- t[12709] = 3
      "00011" when "011000110100110", -- t[12710] = 3
      "00011" when "011000110100111", -- t[12711] = 3
      "00011" when "011000110101000", -- t[12712] = 3
      "00011" when "011000110101001", -- t[12713] = 3
      "00011" when "011000110101010", -- t[12714] = 3
      "00011" when "011000110101011", -- t[12715] = 3
      "00011" when "011000110101100", -- t[12716] = 3
      "00011" when "011000110101101", -- t[12717] = 3
      "00011" when "011000110101110", -- t[12718] = 3
      "00011" when "011000110101111", -- t[12719] = 3
      "00011" when "011000110110000", -- t[12720] = 3
      "00011" when "011000110110001", -- t[12721] = 3
      "00011" when "011000110110010", -- t[12722] = 3
      "00011" when "011000110110011", -- t[12723] = 3
      "00011" when "011000110110100", -- t[12724] = 3
      "00011" when "011000110110101", -- t[12725] = 3
      "00011" when "011000110110110", -- t[12726] = 3
      "00011" when "011000110110111", -- t[12727] = 3
      "00011" when "011000110111000", -- t[12728] = 3
      "00011" when "011000110111001", -- t[12729] = 3
      "00011" when "011000110111010", -- t[12730] = 3
      "00011" when "011000110111011", -- t[12731] = 3
      "00011" when "011000110111100", -- t[12732] = 3
      "00011" when "011000110111101", -- t[12733] = 3
      "00011" when "011000110111110", -- t[12734] = 3
      "00011" when "011000110111111", -- t[12735] = 3
      "00011" when "011000111000000", -- t[12736] = 3
      "00011" when "011000111000001", -- t[12737] = 3
      "00011" when "011000111000010", -- t[12738] = 3
      "00011" when "011000111000011", -- t[12739] = 3
      "00011" when "011000111000100", -- t[12740] = 3
      "00011" when "011000111000101", -- t[12741] = 3
      "00011" when "011000111000110", -- t[12742] = 3
      "00011" when "011000111000111", -- t[12743] = 3
      "00011" when "011000111001000", -- t[12744] = 3
      "00011" when "011000111001001", -- t[12745] = 3
      "00011" when "011000111001010", -- t[12746] = 3
      "00011" when "011000111001011", -- t[12747] = 3
      "00011" when "011000111001100", -- t[12748] = 3
      "00011" when "011000111001101", -- t[12749] = 3
      "00011" when "011000111001110", -- t[12750] = 3
      "00011" when "011000111001111", -- t[12751] = 3
      "00011" when "011000111010000", -- t[12752] = 3
      "00011" when "011000111010001", -- t[12753] = 3
      "00011" when "011000111010010", -- t[12754] = 3
      "00011" when "011000111010011", -- t[12755] = 3
      "00011" when "011000111010100", -- t[12756] = 3
      "00011" when "011000111010101", -- t[12757] = 3
      "00011" when "011000111010110", -- t[12758] = 3
      "00011" when "011000111010111", -- t[12759] = 3
      "00011" when "011000111011000", -- t[12760] = 3
      "00011" when "011000111011001", -- t[12761] = 3
      "00011" when "011000111011010", -- t[12762] = 3
      "00011" when "011000111011011", -- t[12763] = 3
      "00011" when "011000111011100", -- t[12764] = 3
      "00011" when "011000111011101", -- t[12765] = 3
      "00011" when "011000111011110", -- t[12766] = 3
      "00011" when "011000111011111", -- t[12767] = 3
      "00011" when "011000111100000", -- t[12768] = 3
      "00011" when "011000111100001", -- t[12769] = 3
      "00011" when "011000111100010", -- t[12770] = 3
      "00011" when "011000111100011", -- t[12771] = 3
      "00011" when "011000111100100", -- t[12772] = 3
      "00011" when "011000111100101", -- t[12773] = 3
      "00011" when "011000111100110", -- t[12774] = 3
      "00011" when "011000111100111", -- t[12775] = 3
      "00011" when "011000111101000", -- t[12776] = 3
      "00011" when "011000111101001", -- t[12777] = 3
      "00011" when "011000111101010", -- t[12778] = 3
      "00011" when "011000111101011", -- t[12779] = 3
      "00011" when "011000111101100", -- t[12780] = 3
      "00011" when "011000111101101", -- t[12781] = 3
      "00011" when "011000111101110", -- t[12782] = 3
      "00011" when "011000111101111", -- t[12783] = 3
      "00011" when "011000111110000", -- t[12784] = 3
      "00011" when "011000111110001", -- t[12785] = 3
      "00011" when "011000111110010", -- t[12786] = 3
      "00011" when "011000111110011", -- t[12787] = 3
      "00011" when "011000111110100", -- t[12788] = 3
      "00011" when "011000111110101", -- t[12789] = 3
      "00011" when "011000111110110", -- t[12790] = 3
      "00011" when "011000111110111", -- t[12791] = 3
      "00011" when "011000111111000", -- t[12792] = 3
      "00011" when "011000111111001", -- t[12793] = 3
      "00011" when "011000111111010", -- t[12794] = 3
      "00011" when "011000111111011", -- t[12795] = 3
      "00011" when "011000111111100", -- t[12796] = 3
      "00011" when "011000111111101", -- t[12797] = 3
      "00011" when "011000111111110", -- t[12798] = 3
      "00011" when "011000111111111", -- t[12799] = 3
      "00011" when "011001000000000", -- t[12800] = 3
      "00011" when "011001000000001", -- t[12801] = 3
      "00011" when "011001000000010", -- t[12802] = 3
      "00011" when "011001000000011", -- t[12803] = 3
      "00011" when "011001000000100", -- t[12804] = 3
      "00011" when "011001000000101", -- t[12805] = 3
      "00011" when "011001000000110", -- t[12806] = 3
      "00011" when "011001000000111", -- t[12807] = 3
      "00011" when "011001000001000", -- t[12808] = 3
      "00011" when "011001000001001", -- t[12809] = 3
      "00011" when "011001000001010", -- t[12810] = 3
      "00011" when "011001000001011", -- t[12811] = 3
      "00011" when "011001000001100", -- t[12812] = 3
      "00011" when "011001000001101", -- t[12813] = 3
      "00011" when "011001000001110", -- t[12814] = 3
      "00011" when "011001000001111", -- t[12815] = 3
      "00011" when "011001000010000", -- t[12816] = 3
      "00011" when "011001000010001", -- t[12817] = 3
      "00011" when "011001000010010", -- t[12818] = 3
      "00011" when "011001000010011", -- t[12819] = 3
      "00011" when "011001000010100", -- t[12820] = 3
      "00011" when "011001000010101", -- t[12821] = 3
      "00011" when "011001000010110", -- t[12822] = 3
      "00011" when "011001000010111", -- t[12823] = 3
      "00011" when "011001000011000", -- t[12824] = 3
      "00011" when "011001000011001", -- t[12825] = 3
      "00011" when "011001000011010", -- t[12826] = 3
      "00011" when "011001000011011", -- t[12827] = 3
      "00011" when "011001000011100", -- t[12828] = 3
      "00011" when "011001000011101", -- t[12829] = 3
      "00011" when "011001000011110", -- t[12830] = 3
      "00011" when "011001000011111", -- t[12831] = 3
      "00011" when "011001000100000", -- t[12832] = 3
      "00011" when "011001000100001", -- t[12833] = 3
      "00011" when "011001000100010", -- t[12834] = 3
      "00011" when "011001000100011", -- t[12835] = 3
      "00011" when "011001000100100", -- t[12836] = 3
      "00011" when "011001000100101", -- t[12837] = 3
      "00011" when "011001000100110", -- t[12838] = 3
      "00011" when "011001000100111", -- t[12839] = 3
      "00011" when "011001000101000", -- t[12840] = 3
      "00011" when "011001000101001", -- t[12841] = 3
      "00011" when "011001000101010", -- t[12842] = 3
      "00011" when "011001000101011", -- t[12843] = 3
      "00011" when "011001000101100", -- t[12844] = 3
      "00011" when "011001000101101", -- t[12845] = 3
      "00011" when "011001000101110", -- t[12846] = 3
      "00011" when "011001000101111", -- t[12847] = 3
      "00011" when "011001000110000", -- t[12848] = 3
      "00011" when "011001000110001", -- t[12849] = 3
      "00011" when "011001000110010", -- t[12850] = 3
      "00011" when "011001000110011", -- t[12851] = 3
      "00011" when "011001000110100", -- t[12852] = 3
      "00011" when "011001000110101", -- t[12853] = 3
      "00011" when "011001000110110", -- t[12854] = 3
      "00011" when "011001000110111", -- t[12855] = 3
      "00011" when "011001000111000", -- t[12856] = 3
      "00100" when "011001000111001", -- t[12857] = 4
      "00100" when "011001000111010", -- t[12858] = 4
      "00100" when "011001000111011", -- t[12859] = 4
      "00100" when "011001000111100", -- t[12860] = 4
      "00100" when "011001000111101", -- t[12861] = 4
      "00100" when "011001000111110", -- t[12862] = 4
      "00100" when "011001000111111", -- t[12863] = 4
      "00100" when "011001001000000", -- t[12864] = 4
      "00100" when "011001001000001", -- t[12865] = 4
      "00100" when "011001001000010", -- t[12866] = 4
      "00100" when "011001001000011", -- t[12867] = 4
      "00100" when "011001001000100", -- t[12868] = 4
      "00100" when "011001001000101", -- t[12869] = 4
      "00100" when "011001001000110", -- t[12870] = 4
      "00100" when "011001001000111", -- t[12871] = 4
      "00100" when "011001001001000", -- t[12872] = 4
      "00100" when "011001001001001", -- t[12873] = 4
      "00100" when "011001001001010", -- t[12874] = 4
      "00100" when "011001001001011", -- t[12875] = 4
      "00100" when "011001001001100", -- t[12876] = 4
      "00100" when "011001001001101", -- t[12877] = 4
      "00100" when "011001001001110", -- t[12878] = 4
      "00100" when "011001001001111", -- t[12879] = 4
      "00100" when "011001001010000", -- t[12880] = 4
      "00100" when "011001001010001", -- t[12881] = 4
      "00100" when "011001001010010", -- t[12882] = 4
      "00100" when "011001001010011", -- t[12883] = 4
      "00100" when "011001001010100", -- t[12884] = 4
      "00100" when "011001001010101", -- t[12885] = 4
      "00100" when "011001001010110", -- t[12886] = 4
      "00100" when "011001001010111", -- t[12887] = 4
      "00100" when "011001001011000", -- t[12888] = 4
      "00100" when "011001001011001", -- t[12889] = 4
      "00100" when "011001001011010", -- t[12890] = 4
      "00100" when "011001001011011", -- t[12891] = 4
      "00100" when "011001001011100", -- t[12892] = 4
      "00100" when "011001001011101", -- t[12893] = 4
      "00100" when "011001001011110", -- t[12894] = 4
      "00100" when "011001001011111", -- t[12895] = 4
      "00100" when "011001001100000", -- t[12896] = 4
      "00100" when "011001001100001", -- t[12897] = 4
      "00100" when "011001001100010", -- t[12898] = 4
      "00100" when "011001001100011", -- t[12899] = 4
      "00100" when "011001001100100", -- t[12900] = 4
      "00100" when "011001001100101", -- t[12901] = 4
      "00100" when "011001001100110", -- t[12902] = 4
      "00100" when "011001001100111", -- t[12903] = 4
      "00100" when "011001001101000", -- t[12904] = 4
      "00100" when "011001001101001", -- t[12905] = 4
      "00100" when "011001001101010", -- t[12906] = 4
      "00100" when "011001001101011", -- t[12907] = 4
      "00100" when "011001001101100", -- t[12908] = 4
      "00100" when "011001001101101", -- t[12909] = 4
      "00100" when "011001001101110", -- t[12910] = 4
      "00100" when "011001001101111", -- t[12911] = 4
      "00100" when "011001001110000", -- t[12912] = 4
      "00100" when "011001001110001", -- t[12913] = 4
      "00100" when "011001001110010", -- t[12914] = 4
      "00100" when "011001001110011", -- t[12915] = 4
      "00100" when "011001001110100", -- t[12916] = 4
      "00100" when "011001001110101", -- t[12917] = 4
      "00100" when "011001001110110", -- t[12918] = 4
      "00100" when "011001001110111", -- t[12919] = 4
      "00100" when "011001001111000", -- t[12920] = 4
      "00100" when "011001001111001", -- t[12921] = 4
      "00100" when "011001001111010", -- t[12922] = 4
      "00100" when "011001001111011", -- t[12923] = 4
      "00100" when "011001001111100", -- t[12924] = 4
      "00100" when "011001001111101", -- t[12925] = 4
      "00100" when "011001001111110", -- t[12926] = 4
      "00100" when "011001001111111", -- t[12927] = 4
      "00100" when "011001010000000", -- t[12928] = 4
      "00100" when "011001010000001", -- t[12929] = 4
      "00100" when "011001010000010", -- t[12930] = 4
      "00100" when "011001010000011", -- t[12931] = 4
      "00100" when "011001010000100", -- t[12932] = 4
      "00100" when "011001010000101", -- t[12933] = 4
      "00100" when "011001010000110", -- t[12934] = 4
      "00100" when "011001010000111", -- t[12935] = 4
      "00100" when "011001010001000", -- t[12936] = 4
      "00100" when "011001010001001", -- t[12937] = 4
      "00100" when "011001010001010", -- t[12938] = 4
      "00100" when "011001010001011", -- t[12939] = 4
      "00100" when "011001010001100", -- t[12940] = 4
      "00100" when "011001010001101", -- t[12941] = 4
      "00100" when "011001010001110", -- t[12942] = 4
      "00100" when "011001010001111", -- t[12943] = 4
      "00100" when "011001010010000", -- t[12944] = 4
      "00100" when "011001010010001", -- t[12945] = 4
      "00100" when "011001010010010", -- t[12946] = 4
      "00100" when "011001010010011", -- t[12947] = 4
      "00100" when "011001010010100", -- t[12948] = 4
      "00100" when "011001010010101", -- t[12949] = 4
      "00100" when "011001010010110", -- t[12950] = 4
      "00100" when "011001010010111", -- t[12951] = 4
      "00100" when "011001010011000", -- t[12952] = 4
      "00100" when "011001010011001", -- t[12953] = 4
      "00100" when "011001010011010", -- t[12954] = 4
      "00100" when "011001010011011", -- t[12955] = 4
      "00100" when "011001010011100", -- t[12956] = 4
      "00100" when "011001010011101", -- t[12957] = 4
      "00100" when "011001010011110", -- t[12958] = 4
      "00100" when "011001010011111", -- t[12959] = 4
      "00100" when "011001010100000", -- t[12960] = 4
      "00100" when "011001010100001", -- t[12961] = 4
      "00100" when "011001010100010", -- t[12962] = 4
      "00100" when "011001010100011", -- t[12963] = 4
      "00100" when "011001010100100", -- t[12964] = 4
      "00100" when "011001010100101", -- t[12965] = 4
      "00100" when "011001010100110", -- t[12966] = 4
      "00100" when "011001010100111", -- t[12967] = 4
      "00100" when "011001010101000", -- t[12968] = 4
      "00100" when "011001010101001", -- t[12969] = 4
      "00100" when "011001010101010", -- t[12970] = 4
      "00100" when "011001010101011", -- t[12971] = 4
      "00100" when "011001010101100", -- t[12972] = 4
      "00100" when "011001010101101", -- t[12973] = 4
      "00100" when "011001010101110", -- t[12974] = 4
      "00100" when "011001010101111", -- t[12975] = 4
      "00100" when "011001010110000", -- t[12976] = 4
      "00100" when "011001010110001", -- t[12977] = 4
      "00100" when "011001010110010", -- t[12978] = 4
      "00100" when "011001010110011", -- t[12979] = 4
      "00100" when "011001010110100", -- t[12980] = 4
      "00100" when "011001010110101", -- t[12981] = 4
      "00100" when "011001010110110", -- t[12982] = 4
      "00100" when "011001010110111", -- t[12983] = 4
      "00100" when "011001010111000", -- t[12984] = 4
      "00100" when "011001010111001", -- t[12985] = 4
      "00100" when "011001010111010", -- t[12986] = 4
      "00100" when "011001010111011", -- t[12987] = 4
      "00100" when "011001010111100", -- t[12988] = 4
      "00100" when "011001010111101", -- t[12989] = 4
      "00100" when "011001010111110", -- t[12990] = 4
      "00100" when "011001010111111", -- t[12991] = 4
      "00100" when "011001011000000", -- t[12992] = 4
      "00100" when "011001011000001", -- t[12993] = 4
      "00100" when "011001011000010", -- t[12994] = 4
      "00100" when "011001011000011", -- t[12995] = 4
      "00100" when "011001011000100", -- t[12996] = 4
      "00100" when "011001011000101", -- t[12997] = 4
      "00100" when "011001011000110", -- t[12998] = 4
      "00100" when "011001011000111", -- t[12999] = 4
      "00100" when "011001011001000", -- t[13000] = 4
      "00100" when "011001011001001", -- t[13001] = 4
      "00100" when "011001011001010", -- t[13002] = 4
      "00100" when "011001011001011", -- t[13003] = 4
      "00100" when "011001011001100", -- t[13004] = 4
      "00100" when "011001011001101", -- t[13005] = 4
      "00100" when "011001011001110", -- t[13006] = 4
      "00100" when "011001011001111", -- t[13007] = 4
      "00100" when "011001011010000", -- t[13008] = 4
      "00100" when "011001011010001", -- t[13009] = 4
      "00100" when "011001011010010", -- t[13010] = 4
      "00100" when "011001011010011", -- t[13011] = 4
      "00100" when "011001011010100", -- t[13012] = 4
      "00100" when "011001011010101", -- t[13013] = 4
      "00100" when "011001011010110", -- t[13014] = 4
      "00100" when "011001011010111", -- t[13015] = 4
      "00100" when "011001011011000", -- t[13016] = 4
      "00100" when "011001011011001", -- t[13017] = 4
      "00100" when "011001011011010", -- t[13018] = 4
      "00100" when "011001011011011", -- t[13019] = 4
      "00100" when "011001011011100", -- t[13020] = 4
      "00100" when "011001011011101", -- t[13021] = 4
      "00100" when "011001011011110", -- t[13022] = 4
      "00100" when "011001011011111", -- t[13023] = 4
      "00100" when "011001011100000", -- t[13024] = 4
      "00100" when "011001011100001", -- t[13025] = 4
      "00100" when "011001011100010", -- t[13026] = 4
      "00100" when "011001011100011", -- t[13027] = 4
      "00100" when "011001011100100", -- t[13028] = 4
      "00100" when "011001011100101", -- t[13029] = 4
      "00100" when "011001011100110", -- t[13030] = 4
      "00100" when "011001011100111", -- t[13031] = 4
      "00100" when "011001011101000", -- t[13032] = 4
      "00100" when "011001011101001", -- t[13033] = 4
      "00100" when "011001011101010", -- t[13034] = 4
      "00100" when "011001011101011", -- t[13035] = 4
      "00100" when "011001011101100", -- t[13036] = 4
      "00100" when "011001011101101", -- t[13037] = 4
      "00100" when "011001011101110", -- t[13038] = 4
      "00100" when "011001011101111", -- t[13039] = 4
      "00100" when "011001011110000", -- t[13040] = 4
      "00100" when "011001011110001", -- t[13041] = 4
      "00100" when "011001011110010", -- t[13042] = 4
      "00100" when "011001011110011", -- t[13043] = 4
      "00100" when "011001011110100", -- t[13044] = 4
      "00100" when "011001011110101", -- t[13045] = 4
      "00100" when "011001011110110", -- t[13046] = 4
      "00100" when "011001011110111", -- t[13047] = 4
      "00100" when "011001011111000", -- t[13048] = 4
      "00100" when "011001011111001", -- t[13049] = 4
      "00100" when "011001011111010", -- t[13050] = 4
      "00100" when "011001011111011", -- t[13051] = 4
      "00100" when "011001011111100", -- t[13052] = 4
      "00100" when "011001011111101", -- t[13053] = 4
      "00100" when "011001011111110", -- t[13054] = 4
      "00100" when "011001011111111", -- t[13055] = 4
      "00100" when "011001100000000", -- t[13056] = 4
      "00100" when "011001100000001", -- t[13057] = 4
      "00100" when "011001100000010", -- t[13058] = 4
      "00100" when "011001100000011", -- t[13059] = 4
      "00100" when "011001100000100", -- t[13060] = 4
      "00100" when "011001100000101", -- t[13061] = 4
      "00100" when "011001100000110", -- t[13062] = 4
      "00100" when "011001100000111", -- t[13063] = 4
      "00100" when "011001100001000", -- t[13064] = 4
      "00100" when "011001100001001", -- t[13065] = 4
      "00100" when "011001100001010", -- t[13066] = 4
      "00100" when "011001100001011", -- t[13067] = 4
      "00100" when "011001100001100", -- t[13068] = 4
      "00100" when "011001100001101", -- t[13069] = 4
      "00100" when "011001100001110", -- t[13070] = 4
      "00100" when "011001100001111", -- t[13071] = 4
      "00100" when "011001100010000", -- t[13072] = 4
      "00100" when "011001100010001", -- t[13073] = 4
      "00100" when "011001100010010", -- t[13074] = 4
      "00100" when "011001100010011", -- t[13075] = 4
      "00100" when "011001100010100", -- t[13076] = 4
      "00100" when "011001100010101", -- t[13077] = 4
      "00100" when "011001100010110", -- t[13078] = 4
      "00100" when "011001100010111", -- t[13079] = 4
      "00100" when "011001100011000", -- t[13080] = 4
      "00100" when "011001100011001", -- t[13081] = 4
      "00100" when "011001100011010", -- t[13082] = 4
      "00100" when "011001100011011", -- t[13083] = 4
      "00100" when "011001100011100", -- t[13084] = 4
      "00100" when "011001100011101", -- t[13085] = 4
      "00100" when "011001100011110", -- t[13086] = 4
      "00100" when "011001100011111", -- t[13087] = 4
      "00100" when "011001100100000", -- t[13088] = 4
      "00100" when "011001100100001", -- t[13089] = 4
      "00100" when "011001100100010", -- t[13090] = 4
      "00100" when "011001100100011", -- t[13091] = 4
      "00100" when "011001100100100", -- t[13092] = 4
      "00100" when "011001100100101", -- t[13093] = 4
      "00100" when "011001100100110", -- t[13094] = 4
      "00100" when "011001100100111", -- t[13095] = 4
      "00100" when "011001100101000", -- t[13096] = 4
      "00100" when "011001100101001", -- t[13097] = 4
      "00100" when "011001100101010", -- t[13098] = 4
      "00100" when "011001100101011", -- t[13099] = 4
      "00100" when "011001100101100", -- t[13100] = 4
      "00100" when "011001100101101", -- t[13101] = 4
      "00100" when "011001100101110", -- t[13102] = 4
      "00100" when "011001100101111", -- t[13103] = 4
      "00100" when "011001100110000", -- t[13104] = 4
      "00100" when "011001100110001", -- t[13105] = 4
      "00100" when "011001100110010", -- t[13106] = 4
      "00100" when "011001100110011", -- t[13107] = 4
      "00100" when "011001100110100", -- t[13108] = 4
      "00100" when "011001100110101", -- t[13109] = 4
      "00100" when "011001100110110", -- t[13110] = 4
      "00100" when "011001100110111", -- t[13111] = 4
      "00100" when "011001100111000", -- t[13112] = 4
      "00100" when "011001100111001", -- t[13113] = 4
      "00100" when "011001100111010", -- t[13114] = 4
      "00100" when "011001100111011", -- t[13115] = 4
      "00100" when "011001100111100", -- t[13116] = 4
      "00100" when "011001100111101", -- t[13117] = 4
      "00100" when "011001100111110", -- t[13118] = 4
      "00100" when "011001100111111", -- t[13119] = 4
      "00100" when "011001101000000", -- t[13120] = 4
      "00100" when "011001101000001", -- t[13121] = 4
      "00100" when "011001101000010", -- t[13122] = 4
      "00100" when "011001101000011", -- t[13123] = 4
      "00100" when "011001101000100", -- t[13124] = 4
      "00100" when "011001101000101", -- t[13125] = 4
      "00100" when "011001101000110", -- t[13126] = 4
      "00100" when "011001101000111", -- t[13127] = 4
      "00100" when "011001101001000", -- t[13128] = 4
      "00100" when "011001101001001", -- t[13129] = 4
      "00100" when "011001101001010", -- t[13130] = 4
      "00100" when "011001101001011", -- t[13131] = 4
      "00100" when "011001101001100", -- t[13132] = 4
      "00100" when "011001101001101", -- t[13133] = 4
      "00100" when "011001101001110", -- t[13134] = 4
      "00100" when "011001101001111", -- t[13135] = 4
      "00100" when "011001101010000", -- t[13136] = 4
      "00100" when "011001101010001", -- t[13137] = 4
      "00100" when "011001101010010", -- t[13138] = 4
      "00100" when "011001101010011", -- t[13139] = 4
      "00100" when "011001101010100", -- t[13140] = 4
      "00100" when "011001101010101", -- t[13141] = 4
      "00100" when "011001101010110", -- t[13142] = 4
      "00100" when "011001101010111", -- t[13143] = 4
      "00100" when "011001101011000", -- t[13144] = 4
      "00100" when "011001101011001", -- t[13145] = 4
      "00100" when "011001101011010", -- t[13146] = 4
      "00100" when "011001101011011", -- t[13147] = 4
      "00100" when "011001101011100", -- t[13148] = 4
      "00100" when "011001101011101", -- t[13149] = 4
      "00100" when "011001101011110", -- t[13150] = 4
      "00100" when "011001101011111", -- t[13151] = 4
      "00100" when "011001101100000", -- t[13152] = 4
      "00100" when "011001101100001", -- t[13153] = 4
      "00100" when "011001101100010", -- t[13154] = 4
      "00100" when "011001101100011", -- t[13155] = 4
      "00100" when "011001101100100", -- t[13156] = 4
      "00100" when "011001101100101", -- t[13157] = 4
      "00100" when "011001101100110", -- t[13158] = 4
      "00100" when "011001101100111", -- t[13159] = 4
      "00100" when "011001101101000", -- t[13160] = 4
      "00100" when "011001101101001", -- t[13161] = 4
      "00100" when "011001101101010", -- t[13162] = 4
      "00100" when "011001101101011", -- t[13163] = 4
      "00100" when "011001101101100", -- t[13164] = 4
      "00100" when "011001101101101", -- t[13165] = 4
      "00100" when "011001101101110", -- t[13166] = 4
      "00100" when "011001101101111", -- t[13167] = 4
      "00100" when "011001101110000", -- t[13168] = 4
      "00100" when "011001101110001", -- t[13169] = 4
      "00100" when "011001101110010", -- t[13170] = 4
      "00100" when "011001101110011", -- t[13171] = 4
      "00100" when "011001101110100", -- t[13172] = 4
      "00100" when "011001101110101", -- t[13173] = 4
      "00100" when "011001101110110", -- t[13174] = 4
      "00100" when "011001101110111", -- t[13175] = 4
      "00100" when "011001101111000", -- t[13176] = 4
      "00100" when "011001101111001", -- t[13177] = 4
      "00100" when "011001101111010", -- t[13178] = 4
      "00100" when "011001101111011", -- t[13179] = 4
      "00100" when "011001101111100", -- t[13180] = 4
      "00100" when "011001101111101", -- t[13181] = 4
      "00100" when "011001101111110", -- t[13182] = 4
      "00100" when "011001101111111", -- t[13183] = 4
      "00100" when "011001110000000", -- t[13184] = 4
      "00100" when "011001110000001", -- t[13185] = 4
      "00100" when "011001110000010", -- t[13186] = 4
      "00100" when "011001110000011", -- t[13187] = 4
      "00100" when "011001110000100", -- t[13188] = 4
      "00100" when "011001110000101", -- t[13189] = 4
      "00100" when "011001110000110", -- t[13190] = 4
      "00100" when "011001110000111", -- t[13191] = 4
      "00100" when "011001110001000", -- t[13192] = 4
      "00100" when "011001110001001", -- t[13193] = 4
      "00100" when "011001110001010", -- t[13194] = 4
      "00100" when "011001110001011", -- t[13195] = 4
      "00100" when "011001110001100", -- t[13196] = 4
      "00100" when "011001110001101", -- t[13197] = 4
      "00100" when "011001110001110", -- t[13198] = 4
      "00100" when "011001110001111", -- t[13199] = 4
      "00100" when "011001110010000", -- t[13200] = 4
      "00100" when "011001110010001", -- t[13201] = 4
      "00100" when "011001110010010", -- t[13202] = 4
      "00100" when "011001110010011", -- t[13203] = 4
      "00100" when "011001110010100", -- t[13204] = 4
      "00100" when "011001110010101", -- t[13205] = 4
      "00100" when "011001110010110", -- t[13206] = 4
      "00100" when "011001110010111", -- t[13207] = 4
      "00100" when "011001110011000", -- t[13208] = 4
      "00100" when "011001110011001", -- t[13209] = 4
      "00100" when "011001110011010", -- t[13210] = 4
      "00100" when "011001110011011", -- t[13211] = 4
      "00100" when "011001110011100", -- t[13212] = 4
      "00100" when "011001110011101", -- t[13213] = 4
      "00100" when "011001110011110", -- t[13214] = 4
      "00100" when "011001110011111", -- t[13215] = 4
      "00100" when "011001110100000", -- t[13216] = 4
      "00100" when "011001110100001", -- t[13217] = 4
      "00100" when "011001110100010", -- t[13218] = 4
      "00100" when "011001110100011", -- t[13219] = 4
      "00100" when "011001110100100", -- t[13220] = 4
      "00100" when "011001110100101", -- t[13221] = 4
      "00100" when "011001110100110", -- t[13222] = 4
      "00100" when "011001110100111", -- t[13223] = 4
      "00100" when "011001110101000", -- t[13224] = 4
      "00100" when "011001110101001", -- t[13225] = 4
      "00100" when "011001110101010", -- t[13226] = 4
      "00100" when "011001110101011", -- t[13227] = 4
      "00100" when "011001110101100", -- t[13228] = 4
      "00100" when "011001110101101", -- t[13229] = 4
      "00100" when "011001110101110", -- t[13230] = 4
      "00100" when "011001110101111", -- t[13231] = 4
      "00100" when "011001110110000", -- t[13232] = 4
      "00100" when "011001110110001", -- t[13233] = 4
      "00100" when "011001110110010", -- t[13234] = 4
      "00100" when "011001110110011", -- t[13235] = 4
      "00100" when "011001110110100", -- t[13236] = 4
      "00100" when "011001110110101", -- t[13237] = 4
      "00100" when "011001110110110", -- t[13238] = 4
      "00100" when "011001110110111", -- t[13239] = 4
      "00100" when "011001110111000", -- t[13240] = 4
      "00100" when "011001110111001", -- t[13241] = 4
      "00100" when "011001110111010", -- t[13242] = 4
      "00100" when "011001110111011", -- t[13243] = 4
      "00100" when "011001110111100", -- t[13244] = 4
      "00100" when "011001110111101", -- t[13245] = 4
      "00100" when "011001110111110", -- t[13246] = 4
      "00100" when "011001110111111", -- t[13247] = 4
      "00100" when "011001111000000", -- t[13248] = 4
      "00100" when "011001111000001", -- t[13249] = 4
      "00100" when "011001111000010", -- t[13250] = 4
      "00100" when "011001111000011", -- t[13251] = 4
      "00100" when "011001111000100", -- t[13252] = 4
      "00100" when "011001111000101", -- t[13253] = 4
      "00100" when "011001111000110", -- t[13254] = 4
      "00100" when "011001111000111", -- t[13255] = 4
      "00100" when "011001111001000", -- t[13256] = 4
      "00100" when "011001111001001", -- t[13257] = 4
      "00100" when "011001111001010", -- t[13258] = 4
      "00100" when "011001111001011", -- t[13259] = 4
      "00100" when "011001111001100", -- t[13260] = 4
      "00100" when "011001111001101", -- t[13261] = 4
      "00100" when "011001111001110", -- t[13262] = 4
      "00100" when "011001111001111", -- t[13263] = 4
      "00100" when "011001111010000", -- t[13264] = 4
      "00100" when "011001111010001", -- t[13265] = 4
      "00100" when "011001111010010", -- t[13266] = 4
      "00100" when "011001111010011", -- t[13267] = 4
      "00100" when "011001111010100", -- t[13268] = 4
      "00100" when "011001111010101", -- t[13269] = 4
      "00100" when "011001111010110", -- t[13270] = 4
      "00100" when "011001111010111", -- t[13271] = 4
      "00100" when "011001111011000", -- t[13272] = 4
      "00100" when "011001111011001", -- t[13273] = 4
      "00100" when "011001111011010", -- t[13274] = 4
      "00100" when "011001111011011", -- t[13275] = 4
      "00100" when "011001111011100", -- t[13276] = 4
      "00100" when "011001111011101", -- t[13277] = 4
      "00100" when "011001111011110", -- t[13278] = 4
      "00100" when "011001111011111", -- t[13279] = 4
      "00100" when "011001111100000", -- t[13280] = 4
      "00100" when "011001111100001", -- t[13281] = 4
      "00100" when "011001111100010", -- t[13282] = 4
      "00100" when "011001111100011", -- t[13283] = 4
      "00100" when "011001111100100", -- t[13284] = 4
      "00100" when "011001111100101", -- t[13285] = 4
      "00100" when "011001111100110", -- t[13286] = 4
      "00100" when "011001111100111", -- t[13287] = 4
      "00100" when "011001111101000", -- t[13288] = 4
      "00100" when "011001111101001", -- t[13289] = 4
      "00100" when "011001111101010", -- t[13290] = 4
      "00100" when "011001111101011", -- t[13291] = 4
      "00100" when "011001111101100", -- t[13292] = 4
      "00100" when "011001111101101", -- t[13293] = 4
      "00100" when "011001111101110", -- t[13294] = 4
      "00100" when "011001111101111", -- t[13295] = 4
      "00100" when "011001111110000", -- t[13296] = 4
      "00100" when "011001111110001", -- t[13297] = 4
      "00100" when "011001111110010", -- t[13298] = 4
      "00100" when "011001111110011", -- t[13299] = 4
      "00100" when "011001111110100", -- t[13300] = 4
      "00100" when "011001111110101", -- t[13301] = 4
      "00100" when "011001111110110", -- t[13302] = 4
      "00100" when "011001111110111", -- t[13303] = 4
      "00100" when "011001111111000", -- t[13304] = 4
      "00100" when "011001111111001", -- t[13305] = 4
      "00100" when "011001111111010", -- t[13306] = 4
      "00100" when "011001111111011", -- t[13307] = 4
      "00100" when "011001111111100", -- t[13308] = 4
      "00100" when "011001111111101", -- t[13309] = 4
      "00100" when "011001111111110", -- t[13310] = 4
      "00100" when "011001111111111", -- t[13311] = 4
      "00100" when "011010000000000", -- t[13312] = 4
      "00100" when "011010000000001", -- t[13313] = 4
      "00100" when "011010000000010", -- t[13314] = 4
      "00100" when "011010000000011", -- t[13315] = 4
      "00100" when "011010000000100", -- t[13316] = 4
      "00100" when "011010000000101", -- t[13317] = 4
      "00100" when "011010000000110", -- t[13318] = 4
      "00100" when "011010000000111", -- t[13319] = 4
      "00100" when "011010000001000", -- t[13320] = 4
      "00100" when "011010000001001", -- t[13321] = 4
      "00100" when "011010000001010", -- t[13322] = 4
      "00100" when "011010000001011", -- t[13323] = 4
      "00100" when "011010000001100", -- t[13324] = 4
      "00100" when "011010000001101", -- t[13325] = 4
      "00100" when "011010000001110", -- t[13326] = 4
      "00100" when "011010000001111", -- t[13327] = 4
      "00100" when "011010000010000", -- t[13328] = 4
      "00100" when "011010000010001", -- t[13329] = 4
      "00100" when "011010000010010", -- t[13330] = 4
      "00100" when "011010000010011", -- t[13331] = 4
      "00100" when "011010000010100", -- t[13332] = 4
      "00100" when "011010000010101", -- t[13333] = 4
      "00100" when "011010000010110", -- t[13334] = 4
      "00100" when "011010000010111", -- t[13335] = 4
      "00100" when "011010000011000", -- t[13336] = 4
      "00100" when "011010000011001", -- t[13337] = 4
      "00100" when "011010000011010", -- t[13338] = 4
      "00100" when "011010000011011", -- t[13339] = 4
      "00100" when "011010000011100", -- t[13340] = 4
      "00100" when "011010000011101", -- t[13341] = 4
      "00100" when "011010000011110", -- t[13342] = 4
      "00100" when "011010000011111", -- t[13343] = 4
      "00100" when "011010000100000", -- t[13344] = 4
      "00100" when "011010000100001", -- t[13345] = 4
      "00100" when "011010000100010", -- t[13346] = 4
      "00100" when "011010000100011", -- t[13347] = 4
      "00100" when "011010000100100", -- t[13348] = 4
      "00100" when "011010000100101", -- t[13349] = 4
      "00100" when "011010000100110", -- t[13350] = 4
      "00100" when "011010000100111", -- t[13351] = 4
      "00100" when "011010000101000", -- t[13352] = 4
      "00100" when "011010000101001", -- t[13353] = 4
      "00100" when "011010000101010", -- t[13354] = 4
      "00100" when "011010000101011", -- t[13355] = 4
      "00100" when "011010000101100", -- t[13356] = 4
      "00100" when "011010000101101", -- t[13357] = 4
      "00100" when "011010000101110", -- t[13358] = 4
      "00100" when "011010000101111", -- t[13359] = 4
      "00100" when "011010000110000", -- t[13360] = 4
      "00100" when "011010000110001", -- t[13361] = 4
      "00100" when "011010000110010", -- t[13362] = 4
      "00100" when "011010000110011", -- t[13363] = 4
      "00100" when "011010000110100", -- t[13364] = 4
      "00100" when "011010000110101", -- t[13365] = 4
      "00100" when "011010000110110", -- t[13366] = 4
      "00100" when "011010000110111", -- t[13367] = 4
      "00100" when "011010000111000", -- t[13368] = 4
      "00100" when "011010000111001", -- t[13369] = 4
      "00100" when "011010000111010", -- t[13370] = 4
      "00100" when "011010000111011", -- t[13371] = 4
      "00100" when "011010000111100", -- t[13372] = 4
      "00100" when "011010000111101", -- t[13373] = 4
      "00100" when "011010000111110", -- t[13374] = 4
      "00100" when "011010000111111", -- t[13375] = 4
      "00100" when "011010001000000", -- t[13376] = 4
      "00100" when "011010001000001", -- t[13377] = 4
      "00100" when "011010001000010", -- t[13378] = 4
      "00100" when "011010001000011", -- t[13379] = 4
      "00100" when "011010001000100", -- t[13380] = 4
      "00100" when "011010001000101", -- t[13381] = 4
      "00100" when "011010001000110", -- t[13382] = 4
      "00100" when "011010001000111", -- t[13383] = 4
      "00100" when "011010001001000", -- t[13384] = 4
      "00100" when "011010001001001", -- t[13385] = 4
      "00100" when "011010001001010", -- t[13386] = 4
      "00100" when "011010001001011", -- t[13387] = 4
      "00100" when "011010001001100", -- t[13388] = 4
      "00100" when "011010001001101", -- t[13389] = 4
      "00100" when "011010001001110", -- t[13390] = 4
      "00100" when "011010001001111", -- t[13391] = 4
      "00100" when "011010001010000", -- t[13392] = 4
      "00100" when "011010001010001", -- t[13393] = 4
      "00100" when "011010001010010", -- t[13394] = 4
      "00100" when "011010001010011", -- t[13395] = 4
      "00100" when "011010001010100", -- t[13396] = 4
      "00100" when "011010001010101", -- t[13397] = 4
      "00100" when "011010001010110", -- t[13398] = 4
      "00100" when "011010001010111", -- t[13399] = 4
      "00100" when "011010001011000", -- t[13400] = 4
      "00100" when "011010001011001", -- t[13401] = 4
      "00100" when "011010001011010", -- t[13402] = 4
      "00100" when "011010001011011", -- t[13403] = 4
      "00100" when "011010001011100", -- t[13404] = 4
      "00100" when "011010001011101", -- t[13405] = 4
      "00100" when "011010001011110", -- t[13406] = 4
      "00100" when "011010001011111", -- t[13407] = 4
      "00100" when "011010001100000", -- t[13408] = 4
      "00100" when "011010001100001", -- t[13409] = 4
      "00100" when "011010001100010", -- t[13410] = 4
      "00100" when "011010001100011", -- t[13411] = 4
      "00100" when "011010001100100", -- t[13412] = 4
      "00100" when "011010001100101", -- t[13413] = 4
      "00100" when "011010001100110", -- t[13414] = 4
      "00100" when "011010001100111", -- t[13415] = 4
      "00100" when "011010001101000", -- t[13416] = 4
      "00100" when "011010001101001", -- t[13417] = 4
      "00100" when "011010001101010", -- t[13418] = 4
      "00100" when "011010001101011", -- t[13419] = 4
      "00100" when "011010001101100", -- t[13420] = 4
      "00100" when "011010001101101", -- t[13421] = 4
      "00100" when "011010001101110", -- t[13422] = 4
      "00100" when "011010001101111", -- t[13423] = 4
      "00100" when "011010001110000", -- t[13424] = 4
      "00100" when "011010001110001", -- t[13425] = 4
      "00100" when "011010001110010", -- t[13426] = 4
      "00100" when "011010001110011", -- t[13427] = 4
      "00100" when "011010001110100", -- t[13428] = 4
      "00100" when "011010001110101", -- t[13429] = 4
      "00100" when "011010001110110", -- t[13430] = 4
      "00100" when "011010001110111", -- t[13431] = 4
      "00100" when "011010001111000", -- t[13432] = 4
      "00100" when "011010001111001", -- t[13433] = 4
      "00100" when "011010001111010", -- t[13434] = 4
      "00100" when "011010001111011", -- t[13435] = 4
      "00100" when "011010001111100", -- t[13436] = 4
      "00100" when "011010001111101", -- t[13437] = 4
      "00100" when "011010001111110", -- t[13438] = 4
      "00100" when "011010001111111", -- t[13439] = 4
      "00100" when "011010010000000", -- t[13440] = 4
      "00100" when "011010010000001", -- t[13441] = 4
      "00100" when "011010010000010", -- t[13442] = 4
      "00100" when "011010010000011", -- t[13443] = 4
      "00100" when "011010010000100", -- t[13444] = 4
      "00100" when "011010010000101", -- t[13445] = 4
      "00100" when "011010010000110", -- t[13446] = 4
      "00100" when "011010010000111", -- t[13447] = 4
      "00100" when "011010010001000", -- t[13448] = 4
      "00100" when "011010010001001", -- t[13449] = 4
      "00100" when "011010010001010", -- t[13450] = 4
      "00100" when "011010010001011", -- t[13451] = 4
      "00100" when "011010010001100", -- t[13452] = 4
      "00100" when "011010010001101", -- t[13453] = 4
      "00100" when "011010010001110", -- t[13454] = 4
      "00100" when "011010010001111", -- t[13455] = 4
      "00100" when "011010010010000", -- t[13456] = 4
      "00100" when "011010010010001", -- t[13457] = 4
      "00100" when "011010010010010", -- t[13458] = 4
      "00100" when "011010010010011", -- t[13459] = 4
      "00100" when "011010010010100", -- t[13460] = 4
      "00100" when "011010010010101", -- t[13461] = 4
      "00100" when "011010010010110", -- t[13462] = 4
      "00100" when "011010010010111", -- t[13463] = 4
      "00100" when "011010010011000", -- t[13464] = 4
      "00100" when "011010010011001", -- t[13465] = 4
      "00100" when "011010010011010", -- t[13466] = 4
      "00100" when "011010010011011", -- t[13467] = 4
      "00100" when "011010010011100", -- t[13468] = 4
      "00100" when "011010010011101", -- t[13469] = 4
      "00100" when "011010010011110", -- t[13470] = 4
      "00100" when "011010010011111", -- t[13471] = 4
      "00100" when "011010010100000", -- t[13472] = 4
      "00100" when "011010010100001", -- t[13473] = 4
      "00100" when "011010010100010", -- t[13474] = 4
      "00100" when "011010010100011", -- t[13475] = 4
      "00100" when "011010010100100", -- t[13476] = 4
      "00100" when "011010010100101", -- t[13477] = 4
      "00100" when "011010010100110", -- t[13478] = 4
      "00100" when "011010010100111", -- t[13479] = 4
      "00100" when "011010010101000", -- t[13480] = 4
      "00100" when "011010010101001", -- t[13481] = 4
      "00100" when "011010010101010", -- t[13482] = 4
      "00100" when "011010010101011", -- t[13483] = 4
      "00100" when "011010010101100", -- t[13484] = 4
      "00100" when "011010010101101", -- t[13485] = 4
      "00100" when "011010010101110", -- t[13486] = 4
      "00100" when "011010010101111", -- t[13487] = 4
      "00100" when "011010010110000", -- t[13488] = 4
      "00100" when "011010010110001", -- t[13489] = 4
      "00100" when "011010010110010", -- t[13490] = 4
      "00100" when "011010010110011", -- t[13491] = 4
      "00100" when "011010010110100", -- t[13492] = 4
      "00100" when "011010010110101", -- t[13493] = 4
      "00100" when "011010010110110", -- t[13494] = 4
      "00100" when "011010010110111", -- t[13495] = 4
      "00100" when "011010010111000", -- t[13496] = 4
      "00100" when "011010010111001", -- t[13497] = 4
      "00100" when "011010010111010", -- t[13498] = 4
      "00100" when "011010010111011", -- t[13499] = 4
      "00100" when "011010010111100", -- t[13500] = 4
      "00100" when "011010010111101", -- t[13501] = 4
      "00100" when "011010010111110", -- t[13502] = 4
      "00100" when "011010010111111", -- t[13503] = 4
      "00100" when "011010011000000", -- t[13504] = 4
      "00100" when "011010011000001", -- t[13505] = 4
      "00100" when "011010011000010", -- t[13506] = 4
      "00100" when "011010011000011", -- t[13507] = 4
      "00100" when "011010011000100", -- t[13508] = 4
      "00100" when "011010011000101", -- t[13509] = 4
      "00100" when "011010011000110", -- t[13510] = 4
      "00100" when "011010011000111", -- t[13511] = 4
      "00100" when "011010011001000", -- t[13512] = 4
      "00100" when "011010011001001", -- t[13513] = 4
      "00100" when "011010011001010", -- t[13514] = 4
      "00100" when "011010011001011", -- t[13515] = 4
      "00100" when "011010011001100", -- t[13516] = 4
      "00100" when "011010011001101", -- t[13517] = 4
      "00100" when "011010011001110", -- t[13518] = 4
      "00100" when "011010011001111", -- t[13519] = 4
      "00100" when "011010011010000", -- t[13520] = 4
      "00100" when "011010011010001", -- t[13521] = 4
      "00100" when "011010011010010", -- t[13522] = 4
      "00100" when "011010011010011", -- t[13523] = 4
      "00100" when "011010011010100", -- t[13524] = 4
      "00100" when "011010011010101", -- t[13525] = 4
      "00100" when "011010011010110", -- t[13526] = 4
      "00100" when "011010011010111", -- t[13527] = 4
      "00100" when "011010011011000", -- t[13528] = 4
      "00100" when "011010011011001", -- t[13529] = 4
      "00100" when "011010011011010", -- t[13530] = 4
      "00100" when "011010011011011", -- t[13531] = 4
      "00100" when "011010011011100", -- t[13532] = 4
      "00100" when "011010011011101", -- t[13533] = 4
      "00100" when "011010011011110", -- t[13534] = 4
      "00100" when "011010011011111", -- t[13535] = 4
      "00100" when "011010011100000", -- t[13536] = 4
      "00100" when "011010011100001", -- t[13537] = 4
      "00100" when "011010011100010", -- t[13538] = 4
      "00100" when "011010011100011", -- t[13539] = 4
      "00100" when "011010011100100", -- t[13540] = 4
      "00100" when "011010011100101", -- t[13541] = 4
      "00100" when "011010011100110", -- t[13542] = 4
      "00100" when "011010011100111", -- t[13543] = 4
      "00100" when "011010011101000", -- t[13544] = 4
      "00100" when "011010011101001", -- t[13545] = 4
      "00100" when "011010011101010", -- t[13546] = 4
      "00100" when "011010011101011", -- t[13547] = 4
      "00100" when "011010011101100", -- t[13548] = 4
      "00100" when "011010011101101", -- t[13549] = 4
      "00100" when "011010011101110", -- t[13550] = 4
      "00100" when "011010011101111", -- t[13551] = 4
      "00100" when "011010011110000", -- t[13552] = 4
      "00100" when "011010011110001", -- t[13553] = 4
      "00100" when "011010011110010", -- t[13554] = 4
      "00100" when "011010011110011", -- t[13555] = 4
      "00100" when "011010011110100", -- t[13556] = 4
      "00100" when "011010011110101", -- t[13557] = 4
      "00100" when "011010011110110", -- t[13558] = 4
      "00100" when "011010011110111", -- t[13559] = 4
      "00100" when "011010011111000", -- t[13560] = 4
      "00100" when "011010011111001", -- t[13561] = 4
      "00100" when "011010011111010", -- t[13562] = 4
      "00100" when "011010011111011", -- t[13563] = 4
      "00100" when "011010011111100", -- t[13564] = 4
      "00100" when "011010011111101", -- t[13565] = 4
      "00100" when "011010011111110", -- t[13566] = 4
      "00100" when "011010011111111", -- t[13567] = 4
      "00100" when "011010100000000", -- t[13568] = 4
      "00100" when "011010100000001", -- t[13569] = 4
      "00100" when "011010100000010", -- t[13570] = 4
      "00100" when "011010100000011", -- t[13571] = 4
      "00100" when "011010100000100", -- t[13572] = 4
      "00100" when "011010100000101", -- t[13573] = 4
      "00100" when "011010100000110", -- t[13574] = 4
      "00100" when "011010100000111", -- t[13575] = 4
      "00100" when "011010100001000", -- t[13576] = 4
      "00100" when "011010100001001", -- t[13577] = 4
      "00100" when "011010100001010", -- t[13578] = 4
      "00100" when "011010100001011", -- t[13579] = 4
      "00100" when "011010100001100", -- t[13580] = 4
      "00100" when "011010100001101", -- t[13581] = 4
      "00100" when "011010100001110", -- t[13582] = 4
      "00100" when "011010100001111", -- t[13583] = 4
      "00100" when "011010100010000", -- t[13584] = 4
      "00100" when "011010100010001", -- t[13585] = 4
      "00100" when "011010100010010", -- t[13586] = 4
      "00100" when "011010100010011", -- t[13587] = 4
      "00100" when "011010100010100", -- t[13588] = 4
      "00100" when "011010100010101", -- t[13589] = 4
      "00100" when "011010100010110", -- t[13590] = 4
      "00100" when "011010100010111", -- t[13591] = 4
      "00100" when "011010100011000", -- t[13592] = 4
      "00100" when "011010100011001", -- t[13593] = 4
      "00100" when "011010100011010", -- t[13594] = 4
      "00100" when "011010100011011", -- t[13595] = 4
      "00100" when "011010100011100", -- t[13596] = 4
      "00100" when "011010100011101", -- t[13597] = 4
      "00100" when "011010100011110", -- t[13598] = 4
      "00101" when "011010100011111", -- t[13599] = 5
      "00101" when "011010100100000", -- t[13600] = 5
      "00101" when "011010100100001", -- t[13601] = 5
      "00101" when "011010100100010", -- t[13602] = 5
      "00101" when "011010100100011", -- t[13603] = 5
      "00101" when "011010100100100", -- t[13604] = 5
      "00101" when "011010100100101", -- t[13605] = 5
      "00101" when "011010100100110", -- t[13606] = 5
      "00101" when "011010100100111", -- t[13607] = 5
      "00101" when "011010100101000", -- t[13608] = 5
      "00101" when "011010100101001", -- t[13609] = 5
      "00101" when "011010100101010", -- t[13610] = 5
      "00101" when "011010100101011", -- t[13611] = 5
      "00101" when "011010100101100", -- t[13612] = 5
      "00101" when "011010100101101", -- t[13613] = 5
      "00101" when "011010100101110", -- t[13614] = 5
      "00101" when "011010100101111", -- t[13615] = 5
      "00101" when "011010100110000", -- t[13616] = 5
      "00101" when "011010100110001", -- t[13617] = 5
      "00101" when "011010100110010", -- t[13618] = 5
      "00101" when "011010100110011", -- t[13619] = 5
      "00101" when "011010100110100", -- t[13620] = 5
      "00101" when "011010100110101", -- t[13621] = 5
      "00101" when "011010100110110", -- t[13622] = 5
      "00101" when "011010100110111", -- t[13623] = 5
      "00101" when "011010100111000", -- t[13624] = 5
      "00101" when "011010100111001", -- t[13625] = 5
      "00101" when "011010100111010", -- t[13626] = 5
      "00101" when "011010100111011", -- t[13627] = 5
      "00101" when "011010100111100", -- t[13628] = 5
      "00101" when "011010100111101", -- t[13629] = 5
      "00101" when "011010100111110", -- t[13630] = 5
      "00101" when "011010100111111", -- t[13631] = 5
      "00101" when "011010101000000", -- t[13632] = 5
      "00101" when "011010101000001", -- t[13633] = 5
      "00101" when "011010101000010", -- t[13634] = 5
      "00101" when "011010101000011", -- t[13635] = 5
      "00101" when "011010101000100", -- t[13636] = 5
      "00101" when "011010101000101", -- t[13637] = 5
      "00101" when "011010101000110", -- t[13638] = 5
      "00101" when "011010101000111", -- t[13639] = 5
      "00101" when "011010101001000", -- t[13640] = 5
      "00101" when "011010101001001", -- t[13641] = 5
      "00101" when "011010101001010", -- t[13642] = 5
      "00101" when "011010101001011", -- t[13643] = 5
      "00101" when "011010101001100", -- t[13644] = 5
      "00101" when "011010101001101", -- t[13645] = 5
      "00101" when "011010101001110", -- t[13646] = 5
      "00101" when "011010101001111", -- t[13647] = 5
      "00101" when "011010101010000", -- t[13648] = 5
      "00101" when "011010101010001", -- t[13649] = 5
      "00101" when "011010101010010", -- t[13650] = 5
      "00101" when "011010101010011", -- t[13651] = 5
      "00101" when "011010101010100", -- t[13652] = 5
      "00101" when "011010101010101", -- t[13653] = 5
      "00101" when "011010101010110", -- t[13654] = 5
      "00101" when "011010101010111", -- t[13655] = 5
      "00101" when "011010101011000", -- t[13656] = 5
      "00101" when "011010101011001", -- t[13657] = 5
      "00101" when "011010101011010", -- t[13658] = 5
      "00101" when "011010101011011", -- t[13659] = 5
      "00101" when "011010101011100", -- t[13660] = 5
      "00101" when "011010101011101", -- t[13661] = 5
      "00101" when "011010101011110", -- t[13662] = 5
      "00101" when "011010101011111", -- t[13663] = 5
      "00101" when "011010101100000", -- t[13664] = 5
      "00101" when "011010101100001", -- t[13665] = 5
      "00101" when "011010101100010", -- t[13666] = 5
      "00101" when "011010101100011", -- t[13667] = 5
      "00101" when "011010101100100", -- t[13668] = 5
      "00101" when "011010101100101", -- t[13669] = 5
      "00101" when "011010101100110", -- t[13670] = 5
      "00101" when "011010101100111", -- t[13671] = 5
      "00101" when "011010101101000", -- t[13672] = 5
      "00101" when "011010101101001", -- t[13673] = 5
      "00101" when "011010101101010", -- t[13674] = 5
      "00101" when "011010101101011", -- t[13675] = 5
      "00101" when "011010101101100", -- t[13676] = 5
      "00101" when "011010101101101", -- t[13677] = 5
      "00101" when "011010101101110", -- t[13678] = 5
      "00101" when "011010101101111", -- t[13679] = 5
      "00101" when "011010101110000", -- t[13680] = 5
      "00101" when "011010101110001", -- t[13681] = 5
      "00101" when "011010101110010", -- t[13682] = 5
      "00101" when "011010101110011", -- t[13683] = 5
      "00101" when "011010101110100", -- t[13684] = 5
      "00101" when "011010101110101", -- t[13685] = 5
      "00101" when "011010101110110", -- t[13686] = 5
      "00101" when "011010101110111", -- t[13687] = 5
      "00101" when "011010101111000", -- t[13688] = 5
      "00101" when "011010101111001", -- t[13689] = 5
      "00101" when "011010101111010", -- t[13690] = 5
      "00101" when "011010101111011", -- t[13691] = 5
      "00101" when "011010101111100", -- t[13692] = 5
      "00101" when "011010101111101", -- t[13693] = 5
      "00101" when "011010101111110", -- t[13694] = 5
      "00101" when "011010101111111", -- t[13695] = 5
      "00101" when "011010110000000", -- t[13696] = 5
      "00101" when "011010110000001", -- t[13697] = 5
      "00101" when "011010110000010", -- t[13698] = 5
      "00101" when "011010110000011", -- t[13699] = 5
      "00101" when "011010110000100", -- t[13700] = 5
      "00101" when "011010110000101", -- t[13701] = 5
      "00101" when "011010110000110", -- t[13702] = 5
      "00101" when "011010110000111", -- t[13703] = 5
      "00101" when "011010110001000", -- t[13704] = 5
      "00101" when "011010110001001", -- t[13705] = 5
      "00101" when "011010110001010", -- t[13706] = 5
      "00101" when "011010110001011", -- t[13707] = 5
      "00101" when "011010110001100", -- t[13708] = 5
      "00101" when "011010110001101", -- t[13709] = 5
      "00101" when "011010110001110", -- t[13710] = 5
      "00101" when "011010110001111", -- t[13711] = 5
      "00101" when "011010110010000", -- t[13712] = 5
      "00101" when "011010110010001", -- t[13713] = 5
      "00101" when "011010110010010", -- t[13714] = 5
      "00101" when "011010110010011", -- t[13715] = 5
      "00101" when "011010110010100", -- t[13716] = 5
      "00101" when "011010110010101", -- t[13717] = 5
      "00101" when "011010110010110", -- t[13718] = 5
      "00101" when "011010110010111", -- t[13719] = 5
      "00101" when "011010110011000", -- t[13720] = 5
      "00101" when "011010110011001", -- t[13721] = 5
      "00101" when "011010110011010", -- t[13722] = 5
      "00101" when "011010110011011", -- t[13723] = 5
      "00101" when "011010110011100", -- t[13724] = 5
      "00101" when "011010110011101", -- t[13725] = 5
      "00101" when "011010110011110", -- t[13726] = 5
      "00101" when "011010110011111", -- t[13727] = 5
      "00101" when "011010110100000", -- t[13728] = 5
      "00101" when "011010110100001", -- t[13729] = 5
      "00101" when "011010110100010", -- t[13730] = 5
      "00101" when "011010110100011", -- t[13731] = 5
      "00101" when "011010110100100", -- t[13732] = 5
      "00101" when "011010110100101", -- t[13733] = 5
      "00101" when "011010110100110", -- t[13734] = 5
      "00101" when "011010110100111", -- t[13735] = 5
      "00101" when "011010110101000", -- t[13736] = 5
      "00101" when "011010110101001", -- t[13737] = 5
      "00101" when "011010110101010", -- t[13738] = 5
      "00101" when "011010110101011", -- t[13739] = 5
      "00101" when "011010110101100", -- t[13740] = 5
      "00101" when "011010110101101", -- t[13741] = 5
      "00101" when "011010110101110", -- t[13742] = 5
      "00101" when "011010110101111", -- t[13743] = 5
      "00101" when "011010110110000", -- t[13744] = 5
      "00101" when "011010110110001", -- t[13745] = 5
      "00101" when "011010110110010", -- t[13746] = 5
      "00101" when "011010110110011", -- t[13747] = 5
      "00101" when "011010110110100", -- t[13748] = 5
      "00101" when "011010110110101", -- t[13749] = 5
      "00101" when "011010110110110", -- t[13750] = 5
      "00101" when "011010110110111", -- t[13751] = 5
      "00101" when "011010110111000", -- t[13752] = 5
      "00101" when "011010110111001", -- t[13753] = 5
      "00101" when "011010110111010", -- t[13754] = 5
      "00101" when "011010110111011", -- t[13755] = 5
      "00101" when "011010110111100", -- t[13756] = 5
      "00101" when "011010110111101", -- t[13757] = 5
      "00101" when "011010110111110", -- t[13758] = 5
      "00101" when "011010110111111", -- t[13759] = 5
      "00101" when "011010111000000", -- t[13760] = 5
      "00101" when "011010111000001", -- t[13761] = 5
      "00101" when "011010111000010", -- t[13762] = 5
      "00101" when "011010111000011", -- t[13763] = 5
      "00101" when "011010111000100", -- t[13764] = 5
      "00101" when "011010111000101", -- t[13765] = 5
      "00101" when "011010111000110", -- t[13766] = 5
      "00101" when "011010111000111", -- t[13767] = 5
      "00101" when "011010111001000", -- t[13768] = 5
      "00101" when "011010111001001", -- t[13769] = 5
      "00101" when "011010111001010", -- t[13770] = 5
      "00101" when "011010111001011", -- t[13771] = 5
      "00101" when "011010111001100", -- t[13772] = 5
      "00101" when "011010111001101", -- t[13773] = 5
      "00101" when "011010111001110", -- t[13774] = 5
      "00101" when "011010111001111", -- t[13775] = 5
      "00101" when "011010111010000", -- t[13776] = 5
      "00101" when "011010111010001", -- t[13777] = 5
      "00101" when "011010111010010", -- t[13778] = 5
      "00101" when "011010111010011", -- t[13779] = 5
      "00101" when "011010111010100", -- t[13780] = 5
      "00101" when "011010111010101", -- t[13781] = 5
      "00101" when "011010111010110", -- t[13782] = 5
      "00101" when "011010111010111", -- t[13783] = 5
      "00101" when "011010111011000", -- t[13784] = 5
      "00101" when "011010111011001", -- t[13785] = 5
      "00101" when "011010111011010", -- t[13786] = 5
      "00101" when "011010111011011", -- t[13787] = 5
      "00101" when "011010111011100", -- t[13788] = 5
      "00101" when "011010111011101", -- t[13789] = 5
      "00101" when "011010111011110", -- t[13790] = 5
      "00101" when "011010111011111", -- t[13791] = 5
      "00101" when "011010111100000", -- t[13792] = 5
      "00101" when "011010111100001", -- t[13793] = 5
      "00101" when "011010111100010", -- t[13794] = 5
      "00101" when "011010111100011", -- t[13795] = 5
      "00101" when "011010111100100", -- t[13796] = 5
      "00101" when "011010111100101", -- t[13797] = 5
      "00101" when "011010111100110", -- t[13798] = 5
      "00101" when "011010111100111", -- t[13799] = 5
      "00101" when "011010111101000", -- t[13800] = 5
      "00101" when "011010111101001", -- t[13801] = 5
      "00101" when "011010111101010", -- t[13802] = 5
      "00101" when "011010111101011", -- t[13803] = 5
      "00101" when "011010111101100", -- t[13804] = 5
      "00101" when "011010111101101", -- t[13805] = 5
      "00101" when "011010111101110", -- t[13806] = 5
      "00101" when "011010111101111", -- t[13807] = 5
      "00101" when "011010111110000", -- t[13808] = 5
      "00101" when "011010111110001", -- t[13809] = 5
      "00101" when "011010111110010", -- t[13810] = 5
      "00101" when "011010111110011", -- t[13811] = 5
      "00101" when "011010111110100", -- t[13812] = 5
      "00101" when "011010111110101", -- t[13813] = 5
      "00101" when "011010111110110", -- t[13814] = 5
      "00101" when "011010111110111", -- t[13815] = 5
      "00101" when "011010111111000", -- t[13816] = 5
      "00101" when "011010111111001", -- t[13817] = 5
      "00101" when "011010111111010", -- t[13818] = 5
      "00101" when "011010111111011", -- t[13819] = 5
      "00101" when "011010111111100", -- t[13820] = 5
      "00101" when "011010111111101", -- t[13821] = 5
      "00101" when "011010111111110", -- t[13822] = 5
      "00101" when "011010111111111", -- t[13823] = 5
      "00101" when "011011000000000", -- t[13824] = 5
      "00101" when "011011000000001", -- t[13825] = 5
      "00101" when "011011000000010", -- t[13826] = 5
      "00101" when "011011000000011", -- t[13827] = 5
      "00101" when "011011000000100", -- t[13828] = 5
      "00101" when "011011000000101", -- t[13829] = 5
      "00101" when "011011000000110", -- t[13830] = 5
      "00101" when "011011000000111", -- t[13831] = 5
      "00101" when "011011000001000", -- t[13832] = 5
      "00101" when "011011000001001", -- t[13833] = 5
      "00101" when "011011000001010", -- t[13834] = 5
      "00101" when "011011000001011", -- t[13835] = 5
      "00101" when "011011000001100", -- t[13836] = 5
      "00101" when "011011000001101", -- t[13837] = 5
      "00101" when "011011000001110", -- t[13838] = 5
      "00101" when "011011000001111", -- t[13839] = 5
      "00101" when "011011000010000", -- t[13840] = 5
      "00101" when "011011000010001", -- t[13841] = 5
      "00101" when "011011000010010", -- t[13842] = 5
      "00101" when "011011000010011", -- t[13843] = 5
      "00101" when "011011000010100", -- t[13844] = 5
      "00101" when "011011000010101", -- t[13845] = 5
      "00101" when "011011000010110", -- t[13846] = 5
      "00101" when "011011000010111", -- t[13847] = 5
      "00101" when "011011000011000", -- t[13848] = 5
      "00101" when "011011000011001", -- t[13849] = 5
      "00101" when "011011000011010", -- t[13850] = 5
      "00101" when "011011000011011", -- t[13851] = 5
      "00101" when "011011000011100", -- t[13852] = 5
      "00101" when "011011000011101", -- t[13853] = 5
      "00101" when "011011000011110", -- t[13854] = 5
      "00101" when "011011000011111", -- t[13855] = 5
      "00101" when "011011000100000", -- t[13856] = 5
      "00101" when "011011000100001", -- t[13857] = 5
      "00101" when "011011000100010", -- t[13858] = 5
      "00101" when "011011000100011", -- t[13859] = 5
      "00101" when "011011000100100", -- t[13860] = 5
      "00101" when "011011000100101", -- t[13861] = 5
      "00101" when "011011000100110", -- t[13862] = 5
      "00101" when "011011000100111", -- t[13863] = 5
      "00101" when "011011000101000", -- t[13864] = 5
      "00101" when "011011000101001", -- t[13865] = 5
      "00101" when "011011000101010", -- t[13866] = 5
      "00101" when "011011000101011", -- t[13867] = 5
      "00101" when "011011000101100", -- t[13868] = 5
      "00101" when "011011000101101", -- t[13869] = 5
      "00101" when "011011000101110", -- t[13870] = 5
      "00101" when "011011000101111", -- t[13871] = 5
      "00101" when "011011000110000", -- t[13872] = 5
      "00101" when "011011000110001", -- t[13873] = 5
      "00101" when "011011000110010", -- t[13874] = 5
      "00101" when "011011000110011", -- t[13875] = 5
      "00101" when "011011000110100", -- t[13876] = 5
      "00101" when "011011000110101", -- t[13877] = 5
      "00101" when "011011000110110", -- t[13878] = 5
      "00101" when "011011000110111", -- t[13879] = 5
      "00101" when "011011000111000", -- t[13880] = 5
      "00101" when "011011000111001", -- t[13881] = 5
      "00101" when "011011000111010", -- t[13882] = 5
      "00101" when "011011000111011", -- t[13883] = 5
      "00101" when "011011000111100", -- t[13884] = 5
      "00101" when "011011000111101", -- t[13885] = 5
      "00101" when "011011000111110", -- t[13886] = 5
      "00101" when "011011000111111", -- t[13887] = 5
      "00101" when "011011001000000", -- t[13888] = 5
      "00101" when "011011001000001", -- t[13889] = 5
      "00101" when "011011001000010", -- t[13890] = 5
      "00101" when "011011001000011", -- t[13891] = 5
      "00101" when "011011001000100", -- t[13892] = 5
      "00101" when "011011001000101", -- t[13893] = 5
      "00101" when "011011001000110", -- t[13894] = 5
      "00101" when "011011001000111", -- t[13895] = 5
      "00101" when "011011001001000", -- t[13896] = 5
      "00101" when "011011001001001", -- t[13897] = 5
      "00101" when "011011001001010", -- t[13898] = 5
      "00101" when "011011001001011", -- t[13899] = 5
      "00101" when "011011001001100", -- t[13900] = 5
      "00101" when "011011001001101", -- t[13901] = 5
      "00101" when "011011001001110", -- t[13902] = 5
      "00101" when "011011001001111", -- t[13903] = 5
      "00101" when "011011001010000", -- t[13904] = 5
      "00101" when "011011001010001", -- t[13905] = 5
      "00101" when "011011001010010", -- t[13906] = 5
      "00101" when "011011001010011", -- t[13907] = 5
      "00101" when "011011001010100", -- t[13908] = 5
      "00101" when "011011001010101", -- t[13909] = 5
      "00101" when "011011001010110", -- t[13910] = 5
      "00101" when "011011001010111", -- t[13911] = 5
      "00101" when "011011001011000", -- t[13912] = 5
      "00101" when "011011001011001", -- t[13913] = 5
      "00101" when "011011001011010", -- t[13914] = 5
      "00101" when "011011001011011", -- t[13915] = 5
      "00101" when "011011001011100", -- t[13916] = 5
      "00101" when "011011001011101", -- t[13917] = 5
      "00101" when "011011001011110", -- t[13918] = 5
      "00101" when "011011001011111", -- t[13919] = 5
      "00101" when "011011001100000", -- t[13920] = 5
      "00101" when "011011001100001", -- t[13921] = 5
      "00101" when "011011001100010", -- t[13922] = 5
      "00101" when "011011001100011", -- t[13923] = 5
      "00101" when "011011001100100", -- t[13924] = 5
      "00101" when "011011001100101", -- t[13925] = 5
      "00101" when "011011001100110", -- t[13926] = 5
      "00101" when "011011001100111", -- t[13927] = 5
      "00101" when "011011001101000", -- t[13928] = 5
      "00101" when "011011001101001", -- t[13929] = 5
      "00101" when "011011001101010", -- t[13930] = 5
      "00101" when "011011001101011", -- t[13931] = 5
      "00101" when "011011001101100", -- t[13932] = 5
      "00101" when "011011001101101", -- t[13933] = 5
      "00101" when "011011001101110", -- t[13934] = 5
      "00101" when "011011001101111", -- t[13935] = 5
      "00101" when "011011001110000", -- t[13936] = 5
      "00101" when "011011001110001", -- t[13937] = 5
      "00101" when "011011001110010", -- t[13938] = 5
      "00101" when "011011001110011", -- t[13939] = 5
      "00101" when "011011001110100", -- t[13940] = 5
      "00101" when "011011001110101", -- t[13941] = 5
      "00101" when "011011001110110", -- t[13942] = 5
      "00101" when "011011001110111", -- t[13943] = 5
      "00101" when "011011001111000", -- t[13944] = 5
      "00101" when "011011001111001", -- t[13945] = 5
      "00101" when "011011001111010", -- t[13946] = 5
      "00101" when "011011001111011", -- t[13947] = 5
      "00101" when "011011001111100", -- t[13948] = 5
      "00101" when "011011001111101", -- t[13949] = 5
      "00101" when "011011001111110", -- t[13950] = 5
      "00101" when "011011001111111", -- t[13951] = 5
      "00101" when "011011010000000", -- t[13952] = 5
      "00101" when "011011010000001", -- t[13953] = 5
      "00101" when "011011010000010", -- t[13954] = 5
      "00101" when "011011010000011", -- t[13955] = 5
      "00101" when "011011010000100", -- t[13956] = 5
      "00101" when "011011010000101", -- t[13957] = 5
      "00101" when "011011010000110", -- t[13958] = 5
      "00101" when "011011010000111", -- t[13959] = 5
      "00101" when "011011010001000", -- t[13960] = 5
      "00101" when "011011010001001", -- t[13961] = 5
      "00101" when "011011010001010", -- t[13962] = 5
      "00101" when "011011010001011", -- t[13963] = 5
      "00101" when "011011010001100", -- t[13964] = 5
      "00101" when "011011010001101", -- t[13965] = 5
      "00101" when "011011010001110", -- t[13966] = 5
      "00101" when "011011010001111", -- t[13967] = 5
      "00101" when "011011010010000", -- t[13968] = 5
      "00101" when "011011010010001", -- t[13969] = 5
      "00101" when "011011010010010", -- t[13970] = 5
      "00101" when "011011010010011", -- t[13971] = 5
      "00101" when "011011010010100", -- t[13972] = 5
      "00101" when "011011010010101", -- t[13973] = 5
      "00101" when "011011010010110", -- t[13974] = 5
      "00101" when "011011010010111", -- t[13975] = 5
      "00101" when "011011010011000", -- t[13976] = 5
      "00101" when "011011010011001", -- t[13977] = 5
      "00101" when "011011010011010", -- t[13978] = 5
      "00101" when "011011010011011", -- t[13979] = 5
      "00101" when "011011010011100", -- t[13980] = 5
      "00101" when "011011010011101", -- t[13981] = 5
      "00101" when "011011010011110", -- t[13982] = 5
      "00101" when "011011010011111", -- t[13983] = 5
      "00101" when "011011010100000", -- t[13984] = 5
      "00101" when "011011010100001", -- t[13985] = 5
      "00101" when "011011010100010", -- t[13986] = 5
      "00101" when "011011010100011", -- t[13987] = 5
      "00101" when "011011010100100", -- t[13988] = 5
      "00101" when "011011010100101", -- t[13989] = 5
      "00101" when "011011010100110", -- t[13990] = 5
      "00101" when "011011010100111", -- t[13991] = 5
      "00101" when "011011010101000", -- t[13992] = 5
      "00101" when "011011010101001", -- t[13993] = 5
      "00101" when "011011010101010", -- t[13994] = 5
      "00101" when "011011010101011", -- t[13995] = 5
      "00101" when "011011010101100", -- t[13996] = 5
      "00101" when "011011010101101", -- t[13997] = 5
      "00101" when "011011010101110", -- t[13998] = 5
      "00101" when "011011010101111", -- t[13999] = 5
      "00101" when "011011010110000", -- t[14000] = 5
      "00101" when "011011010110001", -- t[14001] = 5
      "00101" when "011011010110010", -- t[14002] = 5
      "00101" when "011011010110011", -- t[14003] = 5
      "00101" when "011011010110100", -- t[14004] = 5
      "00101" when "011011010110101", -- t[14005] = 5
      "00101" when "011011010110110", -- t[14006] = 5
      "00101" when "011011010110111", -- t[14007] = 5
      "00101" when "011011010111000", -- t[14008] = 5
      "00101" when "011011010111001", -- t[14009] = 5
      "00101" when "011011010111010", -- t[14010] = 5
      "00101" when "011011010111011", -- t[14011] = 5
      "00101" when "011011010111100", -- t[14012] = 5
      "00101" when "011011010111101", -- t[14013] = 5
      "00101" when "011011010111110", -- t[14014] = 5
      "00101" when "011011010111111", -- t[14015] = 5
      "00101" when "011011011000000", -- t[14016] = 5
      "00101" when "011011011000001", -- t[14017] = 5
      "00101" when "011011011000010", -- t[14018] = 5
      "00101" when "011011011000011", -- t[14019] = 5
      "00101" when "011011011000100", -- t[14020] = 5
      "00101" when "011011011000101", -- t[14021] = 5
      "00101" when "011011011000110", -- t[14022] = 5
      "00101" when "011011011000111", -- t[14023] = 5
      "00101" when "011011011001000", -- t[14024] = 5
      "00101" when "011011011001001", -- t[14025] = 5
      "00101" when "011011011001010", -- t[14026] = 5
      "00101" when "011011011001011", -- t[14027] = 5
      "00101" when "011011011001100", -- t[14028] = 5
      "00101" when "011011011001101", -- t[14029] = 5
      "00101" when "011011011001110", -- t[14030] = 5
      "00101" when "011011011001111", -- t[14031] = 5
      "00101" when "011011011010000", -- t[14032] = 5
      "00101" when "011011011010001", -- t[14033] = 5
      "00101" when "011011011010010", -- t[14034] = 5
      "00101" when "011011011010011", -- t[14035] = 5
      "00101" when "011011011010100", -- t[14036] = 5
      "00101" when "011011011010101", -- t[14037] = 5
      "00101" when "011011011010110", -- t[14038] = 5
      "00101" when "011011011010111", -- t[14039] = 5
      "00101" when "011011011011000", -- t[14040] = 5
      "00101" when "011011011011001", -- t[14041] = 5
      "00101" when "011011011011010", -- t[14042] = 5
      "00101" when "011011011011011", -- t[14043] = 5
      "00101" when "011011011011100", -- t[14044] = 5
      "00101" when "011011011011101", -- t[14045] = 5
      "00101" when "011011011011110", -- t[14046] = 5
      "00101" when "011011011011111", -- t[14047] = 5
      "00101" when "011011011100000", -- t[14048] = 5
      "00101" when "011011011100001", -- t[14049] = 5
      "00101" when "011011011100010", -- t[14050] = 5
      "00101" when "011011011100011", -- t[14051] = 5
      "00101" when "011011011100100", -- t[14052] = 5
      "00101" when "011011011100101", -- t[14053] = 5
      "00101" when "011011011100110", -- t[14054] = 5
      "00101" when "011011011100111", -- t[14055] = 5
      "00101" when "011011011101000", -- t[14056] = 5
      "00101" when "011011011101001", -- t[14057] = 5
      "00101" when "011011011101010", -- t[14058] = 5
      "00101" when "011011011101011", -- t[14059] = 5
      "00101" when "011011011101100", -- t[14060] = 5
      "00101" when "011011011101101", -- t[14061] = 5
      "00101" when "011011011101110", -- t[14062] = 5
      "00101" when "011011011101111", -- t[14063] = 5
      "00101" when "011011011110000", -- t[14064] = 5
      "00101" when "011011011110001", -- t[14065] = 5
      "00101" when "011011011110010", -- t[14066] = 5
      "00101" when "011011011110011", -- t[14067] = 5
      "00101" when "011011011110100", -- t[14068] = 5
      "00101" when "011011011110101", -- t[14069] = 5
      "00101" when "011011011110110", -- t[14070] = 5
      "00101" when "011011011110111", -- t[14071] = 5
      "00101" when "011011011111000", -- t[14072] = 5
      "00101" when "011011011111001", -- t[14073] = 5
      "00101" when "011011011111010", -- t[14074] = 5
      "00101" when "011011011111011", -- t[14075] = 5
      "00101" when "011011011111100", -- t[14076] = 5
      "00101" when "011011011111101", -- t[14077] = 5
      "00101" when "011011011111110", -- t[14078] = 5
      "00101" when "011011011111111", -- t[14079] = 5
      "00101" when "011011100000000", -- t[14080] = 5
      "00101" when "011011100000001", -- t[14081] = 5
      "00101" when "011011100000010", -- t[14082] = 5
      "00101" when "011011100000011", -- t[14083] = 5
      "00101" when "011011100000100", -- t[14084] = 5
      "00101" when "011011100000101", -- t[14085] = 5
      "00101" when "011011100000110", -- t[14086] = 5
      "00101" when "011011100000111", -- t[14087] = 5
      "00101" when "011011100001000", -- t[14088] = 5
      "00101" when "011011100001001", -- t[14089] = 5
      "00101" when "011011100001010", -- t[14090] = 5
      "00101" when "011011100001011", -- t[14091] = 5
      "00101" when "011011100001100", -- t[14092] = 5
      "00101" when "011011100001101", -- t[14093] = 5
      "00101" when "011011100001110", -- t[14094] = 5
      "00101" when "011011100001111", -- t[14095] = 5
      "00101" when "011011100010000", -- t[14096] = 5
      "00101" when "011011100010001", -- t[14097] = 5
      "00101" when "011011100010010", -- t[14098] = 5
      "00101" when "011011100010011", -- t[14099] = 5
      "00101" when "011011100010100", -- t[14100] = 5
      "00101" when "011011100010101", -- t[14101] = 5
      "00101" when "011011100010110", -- t[14102] = 5
      "00101" when "011011100010111", -- t[14103] = 5
      "00101" when "011011100011000", -- t[14104] = 5
      "00101" when "011011100011001", -- t[14105] = 5
      "00101" when "011011100011010", -- t[14106] = 5
      "00101" when "011011100011011", -- t[14107] = 5
      "00101" when "011011100011100", -- t[14108] = 5
      "00101" when "011011100011101", -- t[14109] = 5
      "00101" when "011011100011110", -- t[14110] = 5
      "00101" when "011011100011111", -- t[14111] = 5
      "00101" when "011011100100000", -- t[14112] = 5
      "00101" when "011011100100001", -- t[14113] = 5
      "00101" when "011011100100010", -- t[14114] = 5
      "00101" when "011011100100011", -- t[14115] = 5
      "00101" when "011011100100100", -- t[14116] = 5
      "00101" when "011011100100101", -- t[14117] = 5
      "00101" when "011011100100110", -- t[14118] = 5
      "00101" when "011011100100111", -- t[14119] = 5
      "00101" when "011011100101000", -- t[14120] = 5
      "00101" when "011011100101001", -- t[14121] = 5
      "00101" when "011011100101010", -- t[14122] = 5
      "00101" when "011011100101011", -- t[14123] = 5
      "00101" when "011011100101100", -- t[14124] = 5
      "00101" when "011011100101101", -- t[14125] = 5
      "00101" when "011011100101110", -- t[14126] = 5
      "00101" when "011011100101111", -- t[14127] = 5
      "00101" when "011011100110000", -- t[14128] = 5
      "00101" when "011011100110001", -- t[14129] = 5
      "00101" when "011011100110010", -- t[14130] = 5
      "00101" when "011011100110011", -- t[14131] = 5
      "00101" when "011011100110100", -- t[14132] = 5
      "00101" when "011011100110101", -- t[14133] = 5
      "00101" when "011011100110110", -- t[14134] = 5
      "00101" when "011011100110111", -- t[14135] = 5
      "00101" when "011011100111000", -- t[14136] = 5
      "00101" when "011011100111001", -- t[14137] = 5
      "00101" when "011011100111010", -- t[14138] = 5
      "00101" when "011011100111011", -- t[14139] = 5
      "00101" when "011011100111100", -- t[14140] = 5
      "00101" when "011011100111101", -- t[14141] = 5
      "00101" when "011011100111110", -- t[14142] = 5
      "00101" when "011011100111111", -- t[14143] = 5
      "00101" when "011011101000000", -- t[14144] = 5
      "00101" when "011011101000001", -- t[14145] = 5
      "00101" when "011011101000010", -- t[14146] = 5
      "00101" when "011011101000011", -- t[14147] = 5
      "00101" when "011011101000100", -- t[14148] = 5
      "00101" when "011011101000101", -- t[14149] = 5
      "00101" when "011011101000110", -- t[14150] = 5
      "00101" when "011011101000111", -- t[14151] = 5
      "00101" when "011011101001000", -- t[14152] = 5
      "00101" when "011011101001001", -- t[14153] = 5
      "00101" when "011011101001010", -- t[14154] = 5
      "00101" when "011011101001011", -- t[14155] = 5
      "00101" when "011011101001100", -- t[14156] = 5
      "00101" when "011011101001101", -- t[14157] = 5
      "00101" when "011011101001110", -- t[14158] = 5
      "00101" when "011011101001111", -- t[14159] = 5
      "00101" when "011011101010000", -- t[14160] = 5
      "00101" when "011011101010001", -- t[14161] = 5
      "00101" when "011011101010010", -- t[14162] = 5
      "00101" when "011011101010011", -- t[14163] = 5
      "00101" when "011011101010100", -- t[14164] = 5
      "00101" when "011011101010101", -- t[14165] = 5
      "00101" when "011011101010110", -- t[14166] = 5
      "00101" when "011011101010111", -- t[14167] = 5
      "00101" when "011011101011000", -- t[14168] = 5
      "00101" when "011011101011001", -- t[14169] = 5
      "00101" when "011011101011010", -- t[14170] = 5
      "00101" when "011011101011011", -- t[14171] = 5
      "00101" when "011011101011100", -- t[14172] = 5
      "00101" when "011011101011101", -- t[14173] = 5
      "00101" when "011011101011110", -- t[14174] = 5
      "00101" when "011011101011111", -- t[14175] = 5
      "00101" when "011011101100000", -- t[14176] = 5
      "00101" when "011011101100001", -- t[14177] = 5
      "00101" when "011011101100010", -- t[14178] = 5
      "00101" when "011011101100011", -- t[14179] = 5
      "00101" when "011011101100100", -- t[14180] = 5
      "00101" when "011011101100101", -- t[14181] = 5
      "00101" when "011011101100110", -- t[14182] = 5
      "00101" when "011011101100111", -- t[14183] = 5
      "00101" when "011011101101000", -- t[14184] = 5
      "00101" when "011011101101001", -- t[14185] = 5
      "00101" when "011011101101010", -- t[14186] = 5
      "00101" when "011011101101011", -- t[14187] = 5
      "00101" when "011011101101100", -- t[14188] = 5
      "00101" when "011011101101101", -- t[14189] = 5
      "00101" when "011011101101110", -- t[14190] = 5
      "00101" when "011011101101111", -- t[14191] = 5
      "00110" when "011011101110000", -- t[14192] = 6
      "00110" when "011011101110001", -- t[14193] = 6
      "00110" when "011011101110010", -- t[14194] = 6
      "00110" when "011011101110011", -- t[14195] = 6
      "00110" when "011011101110100", -- t[14196] = 6
      "00110" when "011011101110101", -- t[14197] = 6
      "00110" when "011011101110110", -- t[14198] = 6
      "00110" when "011011101110111", -- t[14199] = 6
      "00110" when "011011101111000", -- t[14200] = 6
      "00110" when "011011101111001", -- t[14201] = 6
      "00110" when "011011101111010", -- t[14202] = 6
      "00110" when "011011101111011", -- t[14203] = 6
      "00110" when "011011101111100", -- t[14204] = 6
      "00110" when "011011101111101", -- t[14205] = 6
      "00110" when "011011101111110", -- t[14206] = 6
      "00110" when "011011101111111", -- t[14207] = 6
      "00110" when "011011110000000", -- t[14208] = 6
      "00110" when "011011110000001", -- t[14209] = 6
      "00110" when "011011110000010", -- t[14210] = 6
      "00110" when "011011110000011", -- t[14211] = 6
      "00110" when "011011110000100", -- t[14212] = 6
      "00110" when "011011110000101", -- t[14213] = 6
      "00110" when "011011110000110", -- t[14214] = 6
      "00110" when "011011110000111", -- t[14215] = 6
      "00110" when "011011110001000", -- t[14216] = 6
      "00110" when "011011110001001", -- t[14217] = 6
      "00110" when "011011110001010", -- t[14218] = 6
      "00110" when "011011110001011", -- t[14219] = 6
      "00110" when "011011110001100", -- t[14220] = 6
      "00110" when "011011110001101", -- t[14221] = 6
      "00110" when "011011110001110", -- t[14222] = 6
      "00110" when "011011110001111", -- t[14223] = 6
      "00110" when "011011110010000", -- t[14224] = 6
      "00110" when "011011110010001", -- t[14225] = 6
      "00110" when "011011110010010", -- t[14226] = 6
      "00110" when "011011110010011", -- t[14227] = 6
      "00110" when "011011110010100", -- t[14228] = 6
      "00110" when "011011110010101", -- t[14229] = 6
      "00110" when "011011110010110", -- t[14230] = 6
      "00110" when "011011110010111", -- t[14231] = 6
      "00110" when "011011110011000", -- t[14232] = 6
      "00110" when "011011110011001", -- t[14233] = 6
      "00110" when "011011110011010", -- t[14234] = 6
      "00110" when "011011110011011", -- t[14235] = 6
      "00110" when "011011110011100", -- t[14236] = 6
      "00110" when "011011110011101", -- t[14237] = 6
      "00110" when "011011110011110", -- t[14238] = 6
      "00110" when "011011110011111", -- t[14239] = 6
      "00110" when "011011110100000", -- t[14240] = 6
      "00110" when "011011110100001", -- t[14241] = 6
      "00110" when "011011110100010", -- t[14242] = 6
      "00110" when "011011110100011", -- t[14243] = 6
      "00110" when "011011110100100", -- t[14244] = 6
      "00110" when "011011110100101", -- t[14245] = 6
      "00110" when "011011110100110", -- t[14246] = 6
      "00110" when "011011110100111", -- t[14247] = 6
      "00110" when "011011110101000", -- t[14248] = 6
      "00110" when "011011110101001", -- t[14249] = 6
      "00110" when "011011110101010", -- t[14250] = 6
      "00110" when "011011110101011", -- t[14251] = 6
      "00110" when "011011110101100", -- t[14252] = 6
      "00110" when "011011110101101", -- t[14253] = 6
      "00110" when "011011110101110", -- t[14254] = 6
      "00110" when "011011110101111", -- t[14255] = 6
      "00110" when "011011110110000", -- t[14256] = 6
      "00110" when "011011110110001", -- t[14257] = 6
      "00110" when "011011110110010", -- t[14258] = 6
      "00110" when "011011110110011", -- t[14259] = 6
      "00110" when "011011110110100", -- t[14260] = 6
      "00110" when "011011110110101", -- t[14261] = 6
      "00110" when "011011110110110", -- t[14262] = 6
      "00110" when "011011110110111", -- t[14263] = 6
      "00110" when "011011110111000", -- t[14264] = 6
      "00110" when "011011110111001", -- t[14265] = 6
      "00110" when "011011110111010", -- t[14266] = 6
      "00110" when "011011110111011", -- t[14267] = 6
      "00110" when "011011110111100", -- t[14268] = 6
      "00110" when "011011110111101", -- t[14269] = 6
      "00110" when "011011110111110", -- t[14270] = 6
      "00110" when "011011110111111", -- t[14271] = 6
      "00110" when "011011111000000", -- t[14272] = 6
      "00110" when "011011111000001", -- t[14273] = 6
      "00110" when "011011111000010", -- t[14274] = 6
      "00110" when "011011111000011", -- t[14275] = 6
      "00110" when "011011111000100", -- t[14276] = 6
      "00110" when "011011111000101", -- t[14277] = 6
      "00110" when "011011111000110", -- t[14278] = 6
      "00110" when "011011111000111", -- t[14279] = 6
      "00110" when "011011111001000", -- t[14280] = 6
      "00110" when "011011111001001", -- t[14281] = 6
      "00110" when "011011111001010", -- t[14282] = 6
      "00110" when "011011111001011", -- t[14283] = 6
      "00110" when "011011111001100", -- t[14284] = 6
      "00110" when "011011111001101", -- t[14285] = 6
      "00110" when "011011111001110", -- t[14286] = 6
      "00110" when "011011111001111", -- t[14287] = 6
      "00110" when "011011111010000", -- t[14288] = 6
      "00110" when "011011111010001", -- t[14289] = 6
      "00110" when "011011111010010", -- t[14290] = 6
      "00110" when "011011111010011", -- t[14291] = 6
      "00110" when "011011111010100", -- t[14292] = 6
      "00110" when "011011111010101", -- t[14293] = 6
      "00110" when "011011111010110", -- t[14294] = 6
      "00110" when "011011111010111", -- t[14295] = 6
      "00110" when "011011111011000", -- t[14296] = 6
      "00110" when "011011111011001", -- t[14297] = 6
      "00110" when "011011111011010", -- t[14298] = 6
      "00110" when "011011111011011", -- t[14299] = 6
      "00110" when "011011111011100", -- t[14300] = 6
      "00110" when "011011111011101", -- t[14301] = 6
      "00110" when "011011111011110", -- t[14302] = 6
      "00110" when "011011111011111", -- t[14303] = 6
      "00110" when "011011111100000", -- t[14304] = 6
      "00110" when "011011111100001", -- t[14305] = 6
      "00110" when "011011111100010", -- t[14306] = 6
      "00110" when "011011111100011", -- t[14307] = 6
      "00110" when "011011111100100", -- t[14308] = 6
      "00110" when "011011111100101", -- t[14309] = 6
      "00110" when "011011111100110", -- t[14310] = 6
      "00110" when "011011111100111", -- t[14311] = 6
      "00110" when "011011111101000", -- t[14312] = 6
      "00110" when "011011111101001", -- t[14313] = 6
      "00110" when "011011111101010", -- t[14314] = 6
      "00110" when "011011111101011", -- t[14315] = 6
      "00110" when "011011111101100", -- t[14316] = 6
      "00110" when "011011111101101", -- t[14317] = 6
      "00110" when "011011111101110", -- t[14318] = 6
      "00110" when "011011111101111", -- t[14319] = 6
      "00110" when "011011111110000", -- t[14320] = 6
      "00110" when "011011111110001", -- t[14321] = 6
      "00110" when "011011111110010", -- t[14322] = 6
      "00110" when "011011111110011", -- t[14323] = 6
      "00110" when "011011111110100", -- t[14324] = 6
      "00110" when "011011111110101", -- t[14325] = 6
      "00110" when "011011111110110", -- t[14326] = 6
      "00110" when "011011111110111", -- t[14327] = 6
      "00110" when "011011111111000", -- t[14328] = 6
      "00110" when "011011111111001", -- t[14329] = 6
      "00110" when "011011111111010", -- t[14330] = 6
      "00110" when "011011111111011", -- t[14331] = 6
      "00110" when "011011111111100", -- t[14332] = 6
      "00110" when "011011111111101", -- t[14333] = 6
      "00110" when "011011111111110", -- t[14334] = 6
      "00110" when "011011111111111", -- t[14335] = 6
      "00110" when "011100000000000", -- t[14336] = 6
      "00110" when "011100000000001", -- t[14337] = 6
      "00110" when "011100000000010", -- t[14338] = 6
      "00110" when "011100000000011", -- t[14339] = 6
      "00110" when "011100000000100", -- t[14340] = 6
      "00110" when "011100000000101", -- t[14341] = 6
      "00110" when "011100000000110", -- t[14342] = 6
      "00110" when "011100000000111", -- t[14343] = 6
      "00110" when "011100000001000", -- t[14344] = 6
      "00110" when "011100000001001", -- t[14345] = 6
      "00110" when "011100000001010", -- t[14346] = 6
      "00110" when "011100000001011", -- t[14347] = 6
      "00110" when "011100000001100", -- t[14348] = 6
      "00110" when "011100000001101", -- t[14349] = 6
      "00110" when "011100000001110", -- t[14350] = 6
      "00110" when "011100000001111", -- t[14351] = 6
      "00110" when "011100000010000", -- t[14352] = 6
      "00110" when "011100000010001", -- t[14353] = 6
      "00110" when "011100000010010", -- t[14354] = 6
      "00110" when "011100000010011", -- t[14355] = 6
      "00110" when "011100000010100", -- t[14356] = 6
      "00110" when "011100000010101", -- t[14357] = 6
      "00110" when "011100000010110", -- t[14358] = 6
      "00110" when "011100000010111", -- t[14359] = 6
      "00110" when "011100000011000", -- t[14360] = 6
      "00110" when "011100000011001", -- t[14361] = 6
      "00110" when "011100000011010", -- t[14362] = 6
      "00110" when "011100000011011", -- t[14363] = 6
      "00110" when "011100000011100", -- t[14364] = 6
      "00110" when "011100000011101", -- t[14365] = 6
      "00110" when "011100000011110", -- t[14366] = 6
      "00110" when "011100000011111", -- t[14367] = 6
      "00110" when "011100000100000", -- t[14368] = 6
      "00110" when "011100000100001", -- t[14369] = 6
      "00110" when "011100000100010", -- t[14370] = 6
      "00110" when "011100000100011", -- t[14371] = 6
      "00110" when "011100000100100", -- t[14372] = 6
      "00110" when "011100000100101", -- t[14373] = 6
      "00110" when "011100000100110", -- t[14374] = 6
      "00110" when "011100000100111", -- t[14375] = 6
      "00110" when "011100000101000", -- t[14376] = 6
      "00110" when "011100000101001", -- t[14377] = 6
      "00110" when "011100000101010", -- t[14378] = 6
      "00110" when "011100000101011", -- t[14379] = 6
      "00110" when "011100000101100", -- t[14380] = 6
      "00110" when "011100000101101", -- t[14381] = 6
      "00110" when "011100000101110", -- t[14382] = 6
      "00110" when "011100000101111", -- t[14383] = 6
      "00110" when "011100000110000", -- t[14384] = 6
      "00110" when "011100000110001", -- t[14385] = 6
      "00110" when "011100000110010", -- t[14386] = 6
      "00110" when "011100000110011", -- t[14387] = 6
      "00110" when "011100000110100", -- t[14388] = 6
      "00110" when "011100000110101", -- t[14389] = 6
      "00110" when "011100000110110", -- t[14390] = 6
      "00110" when "011100000110111", -- t[14391] = 6
      "00110" when "011100000111000", -- t[14392] = 6
      "00110" when "011100000111001", -- t[14393] = 6
      "00110" when "011100000111010", -- t[14394] = 6
      "00110" when "011100000111011", -- t[14395] = 6
      "00110" when "011100000111100", -- t[14396] = 6
      "00110" when "011100000111101", -- t[14397] = 6
      "00110" when "011100000111110", -- t[14398] = 6
      "00110" when "011100000111111", -- t[14399] = 6
      "00110" when "011100001000000", -- t[14400] = 6
      "00110" when "011100001000001", -- t[14401] = 6
      "00110" when "011100001000010", -- t[14402] = 6
      "00110" when "011100001000011", -- t[14403] = 6
      "00110" when "011100001000100", -- t[14404] = 6
      "00110" when "011100001000101", -- t[14405] = 6
      "00110" when "011100001000110", -- t[14406] = 6
      "00110" when "011100001000111", -- t[14407] = 6
      "00110" when "011100001001000", -- t[14408] = 6
      "00110" when "011100001001001", -- t[14409] = 6
      "00110" when "011100001001010", -- t[14410] = 6
      "00110" when "011100001001011", -- t[14411] = 6
      "00110" when "011100001001100", -- t[14412] = 6
      "00110" when "011100001001101", -- t[14413] = 6
      "00110" when "011100001001110", -- t[14414] = 6
      "00110" when "011100001001111", -- t[14415] = 6
      "00110" when "011100001010000", -- t[14416] = 6
      "00110" when "011100001010001", -- t[14417] = 6
      "00110" when "011100001010010", -- t[14418] = 6
      "00110" when "011100001010011", -- t[14419] = 6
      "00110" when "011100001010100", -- t[14420] = 6
      "00110" when "011100001010101", -- t[14421] = 6
      "00110" when "011100001010110", -- t[14422] = 6
      "00110" when "011100001010111", -- t[14423] = 6
      "00110" when "011100001011000", -- t[14424] = 6
      "00110" when "011100001011001", -- t[14425] = 6
      "00110" when "011100001011010", -- t[14426] = 6
      "00110" when "011100001011011", -- t[14427] = 6
      "00110" when "011100001011100", -- t[14428] = 6
      "00110" when "011100001011101", -- t[14429] = 6
      "00110" when "011100001011110", -- t[14430] = 6
      "00110" when "011100001011111", -- t[14431] = 6
      "00110" when "011100001100000", -- t[14432] = 6
      "00110" when "011100001100001", -- t[14433] = 6
      "00110" when "011100001100010", -- t[14434] = 6
      "00110" when "011100001100011", -- t[14435] = 6
      "00110" when "011100001100100", -- t[14436] = 6
      "00110" when "011100001100101", -- t[14437] = 6
      "00110" when "011100001100110", -- t[14438] = 6
      "00110" when "011100001100111", -- t[14439] = 6
      "00110" when "011100001101000", -- t[14440] = 6
      "00110" when "011100001101001", -- t[14441] = 6
      "00110" when "011100001101010", -- t[14442] = 6
      "00110" when "011100001101011", -- t[14443] = 6
      "00110" when "011100001101100", -- t[14444] = 6
      "00110" when "011100001101101", -- t[14445] = 6
      "00110" when "011100001101110", -- t[14446] = 6
      "00110" when "011100001101111", -- t[14447] = 6
      "00110" when "011100001110000", -- t[14448] = 6
      "00110" when "011100001110001", -- t[14449] = 6
      "00110" when "011100001110010", -- t[14450] = 6
      "00110" when "011100001110011", -- t[14451] = 6
      "00110" when "011100001110100", -- t[14452] = 6
      "00110" when "011100001110101", -- t[14453] = 6
      "00110" when "011100001110110", -- t[14454] = 6
      "00110" when "011100001110111", -- t[14455] = 6
      "00110" when "011100001111000", -- t[14456] = 6
      "00110" when "011100001111001", -- t[14457] = 6
      "00110" when "011100001111010", -- t[14458] = 6
      "00110" when "011100001111011", -- t[14459] = 6
      "00110" when "011100001111100", -- t[14460] = 6
      "00110" when "011100001111101", -- t[14461] = 6
      "00110" when "011100001111110", -- t[14462] = 6
      "00110" when "011100001111111", -- t[14463] = 6
      "00110" when "011100010000000", -- t[14464] = 6
      "00110" when "011100010000001", -- t[14465] = 6
      "00110" when "011100010000010", -- t[14466] = 6
      "00110" when "011100010000011", -- t[14467] = 6
      "00110" when "011100010000100", -- t[14468] = 6
      "00110" when "011100010000101", -- t[14469] = 6
      "00110" when "011100010000110", -- t[14470] = 6
      "00110" when "011100010000111", -- t[14471] = 6
      "00110" when "011100010001000", -- t[14472] = 6
      "00110" when "011100010001001", -- t[14473] = 6
      "00110" when "011100010001010", -- t[14474] = 6
      "00110" when "011100010001011", -- t[14475] = 6
      "00110" when "011100010001100", -- t[14476] = 6
      "00110" when "011100010001101", -- t[14477] = 6
      "00110" when "011100010001110", -- t[14478] = 6
      "00110" when "011100010001111", -- t[14479] = 6
      "00110" when "011100010010000", -- t[14480] = 6
      "00110" when "011100010010001", -- t[14481] = 6
      "00110" when "011100010010010", -- t[14482] = 6
      "00110" when "011100010010011", -- t[14483] = 6
      "00110" when "011100010010100", -- t[14484] = 6
      "00110" when "011100010010101", -- t[14485] = 6
      "00110" when "011100010010110", -- t[14486] = 6
      "00110" when "011100010010111", -- t[14487] = 6
      "00110" when "011100010011000", -- t[14488] = 6
      "00110" when "011100010011001", -- t[14489] = 6
      "00110" when "011100010011010", -- t[14490] = 6
      "00110" when "011100010011011", -- t[14491] = 6
      "00110" when "011100010011100", -- t[14492] = 6
      "00110" when "011100010011101", -- t[14493] = 6
      "00110" when "011100010011110", -- t[14494] = 6
      "00110" when "011100010011111", -- t[14495] = 6
      "00110" when "011100010100000", -- t[14496] = 6
      "00110" when "011100010100001", -- t[14497] = 6
      "00110" when "011100010100010", -- t[14498] = 6
      "00110" when "011100010100011", -- t[14499] = 6
      "00110" when "011100010100100", -- t[14500] = 6
      "00110" when "011100010100101", -- t[14501] = 6
      "00110" when "011100010100110", -- t[14502] = 6
      "00110" when "011100010100111", -- t[14503] = 6
      "00110" when "011100010101000", -- t[14504] = 6
      "00110" when "011100010101001", -- t[14505] = 6
      "00110" when "011100010101010", -- t[14506] = 6
      "00110" when "011100010101011", -- t[14507] = 6
      "00110" when "011100010101100", -- t[14508] = 6
      "00110" when "011100010101101", -- t[14509] = 6
      "00110" when "011100010101110", -- t[14510] = 6
      "00110" when "011100010101111", -- t[14511] = 6
      "00110" when "011100010110000", -- t[14512] = 6
      "00110" when "011100010110001", -- t[14513] = 6
      "00110" when "011100010110010", -- t[14514] = 6
      "00110" when "011100010110011", -- t[14515] = 6
      "00110" when "011100010110100", -- t[14516] = 6
      "00110" when "011100010110101", -- t[14517] = 6
      "00110" when "011100010110110", -- t[14518] = 6
      "00110" when "011100010110111", -- t[14519] = 6
      "00110" when "011100010111000", -- t[14520] = 6
      "00110" when "011100010111001", -- t[14521] = 6
      "00110" when "011100010111010", -- t[14522] = 6
      "00110" when "011100010111011", -- t[14523] = 6
      "00110" when "011100010111100", -- t[14524] = 6
      "00110" when "011100010111101", -- t[14525] = 6
      "00110" when "011100010111110", -- t[14526] = 6
      "00110" when "011100010111111", -- t[14527] = 6
      "00110" when "011100011000000", -- t[14528] = 6
      "00110" when "011100011000001", -- t[14529] = 6
      "00110" when "011100011000010", -- t[14530] = 6
      "00110" when "011100011000011", -- t[14531] = 6
      "00110" when "011100011000100", -- t[14532] = 6
      "00110" when "011100011000101", -- t[14533] = 6
      "00110" when "011100011000110", -- t[14534] = 6
      "00110" when "011100011000111", -- t[14535] = 6
      "00110" when "011100011001000", -- t[14536] = 6
      "00110" when "011100011001001", -- t[14537] = 6
      "00110" when "011100011001010", -- t[14538] = 6
      "00110" when "011100011001011", -- t[14539] = 6
      "00110" when "011100011001100", -- t[14540] = 6
      "00110" when "011100011001101", -- t[14541] = 6
      "00110" when "011100011001110", -- t[14542] = 6
      "00110" when "011100011001111", -- t[14543] = 6
      "00110" when "011100011010000", -- t[14544] = 6
      "00110" when "011100011010001", -- t[14545] = 6
      "00110" when "011100011010010", -- t[14546] = 6
      "00110" when "011100011010011", -- t[14547] = 6
      "00110" when "011100011010100", -- t[14548] = 6
      "00110" when "011100011010101", -- t[14549] = 6
      "00110" when "011100011010110", -- t[14550] = 6
      "00110" when "011100011010111", -- t[14551] = 6
      "00110" when "011100011011000", -- t[14552] = 6
      "00110" when "011100011011001", -- t[14553] = 6
      "00110" when "011100011011010", -- t[14554] = 6
      "00110" when "011100011011011", -- t[14555] = 6
      "00110" when "011100011011100", -- t[14556] = 6
      "00110" when "011100011011101", -- t[14557] = 6
      "00110" when "011100011011110", -- t[14558] = 6
      "00110" when "011100011011111", -- t[14559] = 6
      "00110" when "011100011100000", -- t[14560] = 6
      "00110" when "011100011100001", -- t[14561] = 6
      "00110" when "011100011100010", -- t[14562] = 6
      "00110" when "011100011100011", -- t[14563] = 6
      "00110" when "011100011100100", -- t[14564] = 6
      "00110" when "011100011100101", -- t[14565] = 6
      "00110" when "011100011100110", -- t[14566] = 6
      "00110" when "011100011100111", -- t[14567] = 6
      "00110" when "011100011101000", -- t[14568] = 6
      "00110" when "011100011101001", -- t[14569] = 6
      "00110" when "011100011101010", -- t[14570] = 6
      "00110" when "011100011101011", -- t[14571] = 6
      "00110" when "011100011101100", -- t[14572] = 6
      "00110" when "011100011101101", -- t[14573] = 6
      "00110" when "011100011101110", -- t[14574] = 6
      "00110" when "011100011101111", -- t[14575] = 6
      "00110" when "011100011110000", -- t[14576] = 6
      "00110" when "011100011110001", -- t[14577] = 6
      "00110" when "011100011110010", -- t[14578] = 6
      "00110" when "011100011110011", -- t[14579] = 6
      "00110" when "011100011110100", -- t[14580] = 6
      "00110" when "011100011110101", -- t[14581] = 6
      "00110" when "011100011110110", -- t[14582] = 6
      "00110" when "011100011110111", -- t[14583] = 6
      "00110" when "011100011111000", -- t[14584] = 6
      "00110" when "011100011111001", -- t[14585] = 6
      "00110" when "011100011111010", -- t[14586] = 6
      "00110" when "011100011111011", -- t[14587] = 6
      "00110" when "011100011111100", -- t[14588] = 6
      "00110" when "011100011111101", -- t[14589] = 6
      "00110" when "011100011111110", -- t[14590] = 6
      "00110" when "011100011111111", -- t[14591] = 6
      "00110" when "011100100000000", -- t[14592] = 6
      "00110" when "011100100000001", -- t[14593] = 6
      "00110" when "011100100000010", -- t[14594] = 6
      "00110" when "011100100000011", -- t[14595] = 6
      "00110" when "011100100000100", -- t[14596] = 6
      "00110" when "011100100000101", -- t[14597] = 6
      "00110" when "011100100000110", -- t[14598] = 6
      "00110" when "011100100000111", -- t[14599] = 6
      "00110" when "011100100001000", -- t[14600] = 6
      "00110" when "011100100001001", -- t[14601] = 6
      "00110" when "011100100001010", -- t[14602] = 6
      "00110" when "011100100001011", -- t[14603] = 6
      "00110" when "011100100001100", -- t[14604] = 6
      "00110" when "011100100001101", -- t[14605] = 6
      "00110" when "011100100001110", -- t[14606] = 6
      "00110" when "011100100001111", -- t[14607] = 6
      "00110" when "011100100010000", -- t[14608] = 6
      "00110" when "011100100010001", -- t[14609] = 6
      "00110" when "011100100010010", -- t[14610] = 6
      "00110" when "011100100010011", -- t[14611] = 6
      "00110" when "011100100010100", -- t[14612] = 6
      "00110" when "011100100010101", -- t[14613] = 6
      "00110" when "011100100010110", -- t[14614] = 6
      "00110" when "011100100010111", -- t[14615] = 6
      "00110" when "011100100011000", -- t[14616] = 6
      "00110" when "011100100011001", -- t[14617] = 6
      "00110" when "011100100011010", -- t[14618] = 6
      "00110" when "011100100011011", -- t[14619] = 6
      "00110" when "011100100011100", -- t[14620] = 6
      "00110" when "011100100011101", -- t[14621] = 6
      "00110" when "011100100011110", -- t[14622] = 6
      "00110" when "011100100011111", -- t[14623] = 6
      "00110" when "011100100100000", -- t[14624] = 6
      "00110" when "011100100100001", -- t[14625] = 6
      "00110" when "011100100100010", -- t[14626] = 6
      "00110" when "011100100100011", -- t[14627] = 6
      "00110" when "011100100100100", -- t[14628] = 6
      "00110" when "011100100100101", -- t[14629] = 6
      "00110" when "011100100100110", -- t[14630] = 6
      "00110" when "011100100100111", -- t[14631] = 6
      "00110" when "011100100101000", -- t[14632] = 6
      "00110" when "011100100101001", -- t[14633] = 6
      "00110" when "011100100101010", -- t[14634] = 6
      "00110" when "011100100101011", -- t[14635] = 6
      "00110" when "011100100101100", -- t[14636] = 6
      "00110" when "011100100101101", -- t[14637] = 6
      "00110" when "011100100101110", -- t[14638] = 6
      "00110" when "011100100101111", -- t[14639] = 6
      "00110" when "011100100110000", -- t[14640] = 6
      "00110" when "011100100110001", -- t[14641] = 6
      "00110" when "011100100110010", -- t[14642] = 6
      "00110" when "011100100110011", -- t[14643] = 6
      "00110" when "011100100110100", -- t[14644] = 6
      "00110" when "011100100110101", -- t[14645] = 6
      "00110" when "011100100110110", -- t[14646] = 6
      "00110" when "011100100110111", -- t[14647] = 6
      "00110" when "011100100111000", -- t[14648] = 6
      "00110" when "011100100111001", -- t[14649] = 6
      "00110" when "011100100111010", -- t[14650] = 6
      "00110" when "011100100111011", -- t[14651] = 6
      "00110" when "011100100111100", -- t[14652] = 6
      "00110" when "011100100111101", -- t[14653] = 6
      "00110" when "011100100111110", -- t[14654] = 6
      "00110" when "011100100111111", -- t[14655] = 6
      "00110" when "011100101000000", -- t[14656] = 6
      "00110" when "011100101000001", -- t[14657] = 6
      "00110" when "011100101000010", -- t[14658] = 6
      "00110" when "011100101000011", -- t[14659] = 6
      "00110" when "011100101000100", -- t[14660] = 6
      "00110" when "011100101000101", -- t[14661] = 6
      "00110" when "011100101000110", -- t[14662] = 6
      "00110" when "011100101000111", -- t[14663] = 6
      "00110" when "011100101001000", -- t[14664] = 6
      "00110" when "011100101001001", -- t[14665] = 6
      "00110" when "011100101001010", -- t[14666] = 6
      "00110" when "011100101001011", -- t[14667] = 6
      "00110" when "011100101001100", -- t[14668] = 6
      "00110" when "011100101001101", -- t[14669] = 6
      "00110" when "011100101001110", -- t[14670] = 6
      "00110" when "011100101001111", -- t[14671] = 6
      "00110" when "011100101010000", -- t[14672] = 6
      "00110" when "011100101010001", -- t[14673] = 6
      "00110" when "011100101010010", -- t[14674] = 6
      "00110" when "011100101010011", -- t[14675] = 6
      "00110" when "011100101010100", -- t[14676] = 6
      "00110" when "011100101010101", -- t[14677] = 6
      "00110" when "011100101010110", -- t[14678] = 6
      "00110" when "011100101010111", -- t[14679] = 6
      "00110" when "011100101011000", -- t[14680] = 6
      "00110" when "011100101011001", -- t[14681] = 6
      "00110" when "011100101011010", -- t[14682] = 6
      "00110" when "011100101011011", -- t[14683] = 6
      "00110" when "011100101011100", -- t[14684] = 6
      "00111" when "011100101011101", -- t[14685] = 7
      "00111" when "011100101011110", -- t[14686] = 7
      "00111" when "011100101011111", -- t[14687] = 7
      "00111" when "011100101100000", -- t[14688] = 7
      "00111" when "011100101100001", -- t[14689] = 7
      "00111" when "011100101100010", -- t[14690] = 7
      "00111" when "011100101100011", -- t[14691] = 7
      "00111" when "011100101100100", -- t[14692] = 7
      "00111" when "011100101100101", -- t[14693] = 7
      "00111" when "011100101100110", -- t[14694] = 7
      "00111" when "011100101100111", -- t[14695] = 7
      "00111" when "011100101101000", -- t[14696] = 7
      "00111" when "011100101101001", -- t[14697] = 7
      "00111" when "011100101101010", -- t[14698] = 7
      "00111" when "011100101101011", -- t[14699] = 7
      "00111" when "011100101101100", -- t[14700] = 7
      "00111" when "011100101101101", -- t[14701] = 7
      "00111" when "011100101101110", -- t[14702] = 7
      "00111" when "011100101101111", -- t[14703] = 7
      "00111" when "011100101110000", -- t[14704] = 7
      "00111" when "011100101110001", -- t[14705] = 7
      "00111" when "011100101110010", -- t[14706] = 7
      "00111" when "011100101110011", -- t[14707] = 7
      "00111" when "011100101110100", -- t[14708] = 7
      "00111" when "011100101110101", -- t[14709] = 7
      "00111" when "011100101110110", -- t[14710] = 7
      "00111" when "011100101110111", -- t[14711] = 7
      "00111" when "011100101111000", -- t[14712] = 7
      "00111" when "011100101111001", -- t[14713] = 7
      "00111" when "011100101111010", -- t[14714] = 7
      "00111" when "011100101111011", -- t[14715] = 7
      "00111" when "011100101111100", -- t[14716] = 7
      "00111" when "011100101111101", -- t[14717] = 7
      "00111" when "011100101111110", -- t[14718] = 7
      "00111" when "011100101111111", -- t[14719] = 7
      "00111" when "011100110000000", -- t[14720] = 7
      "00111" when "011100110000001", -- t[14721] = 7
      "00111" when "011100110000010", -- t[14722] = 7
      "00111" when "011100110000011", -- t[14723] = 7
      "00111" when "011100110000100", -- t[14724] = 7
      "00111" when "011100110000101", -- t[14725] = 7
      "00111" when "011100110000110", -- t[14726] = 7
      "00111" when "011100110000111", -- t[14727] = 7
      "00111" when "011100110001000", -- t[14728] = 7
      "00111" when "011100110001001", -- t[14729] = 7
      "00111" when "011100110001010", -- t[14730] = 7
      "00111" when "011100110001011", -- t[14731] = 7
      "00111" when "011100110001100", -- t[14732] = 7
      "00111" when "011100110001101", -- t[14733] = 7
      "00111" when "011100110001110", -- t[14734] = 7
      "00111" when "011100110001111", -- t[14735] = 7
      "00111" when "011100110010000", -- t[14736] = 7
      "00111" when "011100110010001", -- t[14737] = 7
      "00111" when "011100110010010", -- t[14738] = 7
      "00111" when "011100110010011", -- t[14739] = 7
      "00111" when "011100110010100", -- t[14740] = 7
      "00111" when "011100110010101", -- t[14741] = 7
      "00111" when "011100110010110", -- t[14742] = 7
      "00111" when "011100110010111", -- t[14743] = 7
      "00111" when "011100110011000", -- t[14744] = 7
      "00111" when "011100110011001", -- t[14745] = 7
      "00111" when "011100110011010", -- t[14746] = 7
      "00111" when "011100110011011", -- t[14747] = 7
      "00111" when "011100110011100", -- t[14748] = 7
      "00111" when "011100110011101", -- t[14749] = 7
      "00111" when "011100110011110", -- t[14750] = 7
      "00111" when "011100110011111", -- t[14751] = 7
      "00111" when "011100110100000", -- t[14752] = 7
      "00111" when "011100110100001", -- t[14753] = 7
      "00111" when "011100110100010", -- t[14754] = 7
      "00111" when "011100110100011", -- t[14755] = 7
      "00111" when "011100110100100", -- t[14756] = 7
      "00111" when "011100110100101", -- t[14757] = 7
      "00111" when "011100110100110", -- t[14758] = 7
      "00111" when "011100110100111", -- t[14759] = 7
      "00111" when "011100110101000", -- t[14760] = 7
      "00111" when "011100110101001", -- t[14761] = 7
      "00111" when "011100110101010", -- t[14762] = 7
      "00111" when "011100110101011", -- t[14763] = 7
      "00111" when "011100110101100", -- t[14764] = 7
      "00111" when "011100110101101", -- t[14765] = 7
      "00111" when "011100110101110", -- t[14766] = 7
      "00111" when "011100110101111", -- t[14767] = 7
      "00111" when "011100110110000", -- t[14768] = 7
      "00111" when "011100110110001", -- t[14769] = 7
      "00111" when "011100110110010", -- t[14770] = 7
      "00111" when "011100110110011", -- t[14771] = 7
      "00111" when "011100110110100", -- t[14772] = 7
      "00111" when "011100110110101", -- t[14773] = 7
      "00111" when "011100110110110", -- t[14774] = 7
      "00111" when "011100110110111", -- t[14775] = 7
      "00111" when "011100110111000", -- t[14776] = 7
      "00111" when "011100110111001", -- t[14777] = 7
      "00111" when "011100110111010", -- t[14778] = 7
      "00111" when "011100110111011", -- t[14779] = 7
      "00111" when "011100110111100", -- t[14780] = 7
      "00111" when "011100110111101", -- t[14781] = 7
      "00111" when "011100110111110", -- t[14782] = 7
      "00111" when "011100110111111", -- t[14783] = 7
      "00111" when "011100111000000", -- t[14784] = 7
      "00111" when "011100111000001", -- t[14785] = 7
      "00111" when "011100111000010", -- t[14786] = 7
      "00111" when "011100111000011", -- t[14787] = 7
      "00111" when "011100111000100", -- t[14788] = 7
      "00111" when "011100111000101", -- t[14789] = 7
      "00111" when "011100111000110", -- t[14790] = 7
      "00111" when "011100111000111", -- t[14791] = 7
      "00111" when "011100111001000", -- t[14792] = 7
      "00111" when "011100111001001", -- t[14793] = 7
      "00111" when "011100111001010", -- t[14794] = 7
      "00111" when "011100111001011", -- t[14795] = 7
      "00111" when "011100111001100", -- t[14796] = 7
      "00111" when "011100111001101", -- t[14797] = 7
      "00111" when "011100111001110", -- t[14798] = 7
      "00111" when "011100111001111", -- t[14799] = 7
      "00111" when "011100111010000", -- t[14800] = 7
      "00111" when "011100111010001", -- t[14801] = 7
      "00111" when "011100111010010", -- t[14802] = 7
      "00111" when "011100111010011", -- t[14803] = 7
      "00111" when "011100111010100", -- t[14804] = 7
      "00111" when "011100111010101", -- t[14805] = 7
      "00111" when "011100111010110", -- t[14806] = 7
      "00111" when "011100111010111", -- t[14807] = 7
      "00111" when "011100111011000", -- t[14808] = 7
      "00111" when "011100111011001", -- t[14809] = 7
      "00111" when "011100111011010", -- t[14810] = 7
      "00111" when "011100111011011", -- t[14811] = 7
      "00111" when "011100111011100", -- t[14812] = 7
      "00111" when "011100111011101", -- t[14813] = 7
      "00111" when "011100111011110", -- t[14814] = 7
      "00111" when "011100111011111", -- t[14815] = 7
      "00111" when "011100111100000", -- t[14816] = 7
      "00111" when "011100111100001", -- t[14817] = 7
      "00111" when "011100111100010", -- t[14818] = 7
      "00111" when "011100111100011", -- t[14819] = 7
      "00111" when "011100111100100", -- t[14820] = 7
      "00111" when "011100111100101", -- t[14821] = 7
      "00111" when "011100111100110", -- t[14822] = 7
      "00111" when "011100111100111", -- t[14823] = 7
      "00111" when "011100111101000", -- t[14824] = 7
      "00111" when "011100111101001", -- t[14825] = 7
      "00111" when "011100111101010", -- t[14826] = 7
      "00111" when "011100111101011", -- t[14827] = 7
      "00111" when "011100111101100", -- t[14828] = 7
      "00111" when "011100111101101", -- t[14829] = 7
      "00111" when "011100111101110", -- t[14830] = 7
      "00111" when "011100111101111", -- t[14831] = 7
      "00111" when "011100111110000", -- t[14832] = 7
      "00111" when "011100111110001", -- t[14833] = 7
      "00111" when "011100111110010", -- t[14834] = 7
      "00111" when "011100111110011", -- t[14835] = 7
      "00111" when "011100111110100", -- t[14836] = 7
      "00111" when "011100111110101", -- t[14837] = 7
      "00111" when "011100111110110", -- t[14838] = 7
      "00111" when "011100111110111", -- t[14839] = 7
      "00111" when "011100111111000", -- t[14840] = 7
      "00111" when "011100111111001", -- t[14841] = 7
      "00111" when "011100111111010", -- t[14842] = 7
      "00111" when "011100111111011", -- t[14843] = 7
      "00111" when "011100111111100", -- t[14844] = 7
      "00111" when "011100111111101", -- t[14845] = 7
      "00111" when "011100111111110", -- t[14846] = 7
      "00111" when "011100111111111", -- t[14847] = 7
      "00111" when "011101000000000", -- t[14848] = 7
      "00111" when "011101000000001", -- t[14849] = 7
      "00111" when "011101000000010", -- t[14850] = 7
      "00111" when "011101000000011", -- t[14851] = 7
      "00111" when "011101000000100", -- t[14852] = 7
      "00111" when "011101000000101", -- t[14853] = 7
      "00111" when "011101000000110", -- t[14854] = 7
      "00111" when "011101000000111", -- t[14855] = 7
      "00111" when "011101000001000", -- t[14856] = 7
      "00111" when "011101000001001", -- t[14857] = 7
      "00111" when "011101000001010", -- t[14858] = 7
      "00111" when "011101000001011", -- t[14859] = 7
      "00111" when "011101000001100", -- t[14860] = 7
      "00111" when "011101000001101", -- t[14861] = 7
      "00111" when "011101000001110", -- t[14862] = 7
      "00111" when "011101000001111", -- t[14863] = 7
      "00111" when "011101000010000", -- t[14864] = 7
      "00111" when "011101000010001", -- t[14865] = 7
      "00111" when "011101000010010", -- t[14866] = 7
      "00111" when "011101000010011", -- t[14867] = 7
      "00111" when "011101000010100", -- t[14868] = 7
      "00111" when "011101000010101", -- t[14869] = 7
      "00111" when "011101000010110", -- t[14870] = 7
      "00111" when "011101000010111", -- t[14871] = 7
      "00111" when "011101000011000", -- t[14872] = 7
      "00111" when "011101000011001", -- t[14873] = 7
      "00111" when "011101000011010", -- t[14874] = 7
      "00111" when "011101000011011", -- t[14875] = 7
      "00111" when "011101000011100", -- t[14876] = 7
      "00111" when "011101000011101", -- t[14877] = 7
      "00111" when "011101000011110", -- t[14878] = 7
      "00111" when "011101000011111", -- t[14879] = 7
      "00111" when "011101000100000", -- t[14880] = 7
      "00111" when "011101000100001", -- t[14881] = 7
      "00111" when "011101000100010", -- t[14882] = 7
      "00111" when "011101000100011", -- t[14883] = 7
      "00111" when "011101000100100", -- t[14884] = 7
      "00111" when "011101000100101", -- t[14885] = 7
      "00111" when "011101000100110", -- t[14886] = 7
      "00111" when "011101000100111", -- t[14887] = 7
      "00111" when "011101000101000", -- t[14888] = 7
      "00111" when "011101000101001", -- t[14889] = 7
      "00111" when "011101000101010", -- t[14890] = 7
      "00111" when "011101000101011", -- t[14891] = 7
      "00111" when "011101000101100", -- t[14892] = 7
      "00111" when "011101000101101", -- t[14893] = 7
      "00111" when "011101000101110", -- t[14894] = 7
      "00111" when "011101000101111", -- t[14895] = 7
      "00111" when "011101000110000", -- t[14896] = 7
      "00111" when "011101000110001", -- t[14897] = 7
      "00111" when "011101000110010", -- t[14898] = 7
      "00111" when "011101000110011", -- t[14899] = 7
      "00111" when "011101000110100", -- t[14900] = 7
      "00111" when "011101000110101", -- t[14901] = 7
      "00111" when "011101000110110", -- t[14902] = 7
      "00111" when "011101000110111", -- t[14903] = 7
      "00111" when "011101000111000", -- t[14904] = 7
      "00111" when "011101000111001", -- t[14905] = 7
      "00111" when "011101000111010", -- t[14906] = 7
      "00111" when "011101000111011", -- t[14907] = 7
      "00111" when "011101000111100", -- t[14908] = 7
      "00111" when "011101000111101", -- t[14909] = 7
      "00111" when "011101000111110", -- t[14910] = 7
      "00111" when "011101000111111", -- t[14911] = 7
      "00111" when "011101001000000", -- t[14912] = 7
      "00111" when "011101001000001", -- t[14913] = 7
      "00111" when "011101001000010", -- t[14914] = 7
      "00111" when "011101001000011", -- t[14915] = 7
      "00111" when "011101001000100", -- t[14916] = 7
      "00111" when "011101001000101", -- t[14917] = 7
      "00111" when "011101001000110", -- t[14918] = 7
      "00111" when "011101001000111", -- t[14919] = 7
      "00111" when "011101001001000", -- t[14920] = 7
      "00111" when "011101001001001", -- t[14921] = 7
      "00111" when "011101001001010", -- t[14922] = 7
      "00111" when "011101001001011", -- t[14923] = 7
      "00111" when "011101001001100", -- t[14924] = 7
      "00111" when "011101001001101", -- t[14925] = 7
      "00111" when "011101001001110", -- t[14926] = 7
      "00111" when "011101001001111", -- t[14927] = 7
      "00111" when "011101001010000", -- t[14928] = 7
      "00111" when "011101001010001", -- t[14929] = 7
      "00111" when "011101001010010", -- t[14930] = 7
      "00111" when "011101001010011", -- t[14931] = 7
      "00111" when "011101001010100", -- t[14932] = 7
      "00111" when "011101001010101", -- t[14933] = 7
      "00111" when "011101001010110", -- t[14934] = 7
      "00111" when "011101001010111", -- t[14935] = 7
      "00111" when "011101001011000", -- t[14936] = 7
      "00111" when "011101001011001", -- t[14937] = 7
      "00111" when "011101001011010", -- t[14938] = 7
      "00111" when "011101001011011", -- t[14939] = 7
      "00111" when "011101001011100", -- t[14940] = 7
      "00111" when "011101001011101", -- t[14941] = 7
      "00111" when "011101001011110", -- t[14942] = 7
      "00111" when "011101001011111", -- t[14943] = 7
      "00111" when "011101001100000", -- t[14944] = 7
      "00111" when "011101001100001", -- t[14945] = 7
      "00111" when "011101001100010", -- t[14946] = 7
      "00111" when "011101001100011", -- t[14947] = 7
      "00111" when "011101001100100", -- t[14948] = 7
      "00111" when "011101001100101", -- t[14949] = 7
      "00111" when "011101001100110", -- t[14950] = 7
      "00111" when "011101001100111", -- t[14951] = 7
      "00111" when "011101001101000", -- t[14952] = 7
      "00111" when "011101001101001", -- t[14953] = 7
      "00111" when "011101001101010", -- t[14954] = 7
      "00111" when "011101001101011", -- t[14955] = 7
      "00111" when "011101001101100", -- t[14956] = 7
      "00111" when "011101001101101", -- t[14957] = 7
      "00111" when "011101001101110", -- t[14958] = 7
      "00111" when "011101001101111", -- t[14959] = 7
      "00111" when "011101001110000", -- t[14960] = 7
      "00111" when "011101001110001", -- t[14961] = 7
      "00111" when "011101001110010", -- t[14962] = 7
      "00111" when "011101001110011", -- t[14963] = 7
      "00111" when "011101001110100", -- t[14964] = 7
      "00111" when "011101001110101", -- t[14965] = 7
      "00111" when "011101001110110", -- t[14966] = 7
      "00111" when "011101001110111", -- t[14967] = 7
      "00111" when "011101001111000", -- t[14968] = 7
      "00111" when "011101001111001", -- t[14969] = 7
      "00111" when "011101001111010", -- t[14970] = 7
      "00111" when "011101001111011", -- t[14971] = 7
      "00111" when "011101001111100", -- t[14972] = 7
      "00111" when "011101001111101", -- t[14973] = 7
      "00111" when "011101001111110", -- t[14974] = 7
      "00111" when "011101001111111", -- t[14975] = 7
      "00111" when "011101010000000", -- t[14976] = 7
      "00111" when "011101010000001", -- t[14977] = 7
      "00111" when "011101010000010", -- t[14978] = 7
      "00111" when "011101010000011", -- t[14979] = 7
      "00111" when "011101010000100", -- t[14980] = 7
      "00111" when "011101010000101", -- t[14981] = 7
      "00111" when "011101010000110", -- t[14982] = 7
      "00111" when "011101010000111", -- t[14983] = 7
      "00111" when "011101010001000", -- t[14984] = 7
      "00111" when "011101010001001", -- t[14985] = 7
      "00111" when "011101010001010", -- t[14986] = 7
      "00111" when "011101010001011", -- t[14987] = 7
      "00111" when "011101010001100", -- t[14988] = 7
      "00111" when "011101010001101", -- t[14989] = 7
      "00111" when "011101010001110", -- t[14990] = 7
      "00111" when "011101010001111", -- t[14991] = 7
      "00111" when "011101010010000", -- t[14992] = 7
      "00111" when "011101010010001", -- t[14993] = 7
      "00111" when "011101010010010", -- t[14994] = 7
      "00111" when "011101010010011", -- t[14995] = 7
      "00111" when "011101010010100", -- t[14996] = 7
      "00111" when "011101010010101", -- t[14997] = 7
      "00111" when "011101010010110", -- t[14998] = 7
      "00111" when "011101010010111", -- t[14999] = 7
      "00111" when "011101010011000", -- t[15000] = 7
      "00111" when "011101010011001", -- t[15001] = 7
      "00111" when "011101010011010", -- t[15002] = 7
      "00111" when "011101010011011", -- t[15003] = 7
      "00111" when "011101010011100", -- t[15004] = 7
      "00111" when "011101010011101", -- t[15005] = 7
      "00111" when "011101010011110", -- t[15006] = 7
      "00111" when "011101010011111", -- t[15007] = 7
      "00111" when "011101010100000", -- t[15008] = 7
      "00111" when "011101010100001", -- t[15009] = 7
      "00111" when "011101010100010", -- t[15010] = 7
      "00111" when "011101010100011", -- t[15011] = 7
      "00111" when "011101010100100", -- t[15012] = 7
      "00111" when "011101010100101", -- t[15013] = 7
      "00111" when "011101010100110", -- t[15014] = 7
      "00111" when "011101010100111", -- t[15015] = 7
      "00111" when "011101010101000", -- t[15016] = 7
      "00111" when "011101010101001", -- t[15017] = 7
      "00111" when "011101010101010", -- t[15018] = 7
      "00111" when "011101010101011", -- t[15019] = 7
      "00111" when "011101010101100", -- t[15020] = 7
      "00111" when "011101010101101", -- t[15021] = 7
      "00111" when "011101010101110", -- t[15022] = 7
      "00111" when "011101010101111", -- t[15023] = 7
      "00111" when "011101010110000", -- t[15024] = 7
      "00111" when "011101010110001", -- t[15025] = 7
      "00111" when "011101010110010", -- t[15026] = 7
      "00111" when "011101010110011", -- t[15027] = 7
      "00111" when "011101010110100", -- t[15028] = 7
      "00111" when "011101010110101", -- t[15029] = 7
      "00111" when "011101010110110", -- t[15030] = 7
      "00111" when "011101010110111", -- t[15031] = 7
      "00111" when "011101010111000", -- t[15032] = 7
      "00111" when "011101010111001", -- t[15033] = 7
      "00111" when "011101010111010", -- t[15034] = 7
      "00111" when "011101010111011", -- t[15035] = 7
      "00111" when "011101010111100", -- t[15036] = 7
      "00111" when "011101010111101", -- t[15037] = 7
      "00111" when "011101010111110", -- t[15038] = 7
      "00111" when "011101010111111", -- t[15039] = 7
      "00111" when "011101011000000", -- t[15040] = 7
      "00111" when "011101011000001", -- t[15041] = 7
      "00111" when "011101011000010", -- t[15042] = 7
      "00111" when "011101011000011", -- t[15043] = 7
      "00111" when "011101011000100", -- t[15044] = 7
      "00111" when "011101011000101", -- t[15045] = 7
      "00111" when "011101011000110", -- t[15046] = 7
      "00111" when "011101011000111", -- t[15047] = 7
      "00111" when "011101011001000", -- t[15048] = 7
      "00111" when "011101011001001", -- t[15049] = 7
      "00111" when "011101011001010", -- t[15050] = 7
      "00111" when "011101011001011", -- t[15051] = 7
      "00111" when "011101011001100", -- t[15052] = 7
      "00111" when "011101011001101", -- t[15053] = 7
      "00111" when "011101011001110", -- t[15054] = 7
      "00111" when "011101011001111", -- t[15055] = 7
      "00111" when "011101011010000", -- t[15056] = 7
      "00111" when "011101011010001", -- t[15057] = 7
      "00111" when "011101011010010", -- t[15058] = 7
      "00111" when "011101011010011", -- t[15059] = 7
      "00111" when "011101011010100", -- t[15060] = 7
      "00111" when "011101011010101", -- t[15061] = 7
      "00111" when "011101011010110", -- t[15062] = 7
      "00111" when "011101011010111", -- t[15063] = 7
      "00111" when "011101011011000", -- t[15064] = 7
      "00111" when "011101011011001", -- t[15065] = 7
      "00111" when "011101011011010", -- t[15066] = 7
      "00111" when "011101011011011", -- t[15067] = 7
      "00111" when "011101011011100", -- t[15068] = 7
      "00111" when "011101011011101", -- t[15069] = 7
      "00111" when "011101011011110", -- t[15070] = 7
      "00111" when "011101011011111", -- t[15071] = 7
      "00111" when "011101011100000", -- t[15072] = 7
      "00111" when "011101011100001", -- t[15073] = 7
      "00111" when "011101011100010", -- t[15074] = 7
      "00111" when "011101011100011", -- t[15075] = 7
      "00111" when "011101011100100", -- t[15076] = 7
      "00111" when "011101011100101", -- t[15077] = 7
      "00111" when "011101011100110", -- t[15078] = 7
      "00111" when "011101011100111", -- t[15079] = 7
      "00111" when "011101011101000", -- t[15080] = 7
      "00111" when "011101011101001", -- t[15081] = 7
      "00111" when "011101011101010", -- t[15082] = 7
      "00111" when "011101011101011", -- t[15083] = 7
      "00111" when "011101011101100", -- t[15084] = 7
      "00111" when "011101011101101", -- t[15085] = 7
      "00111" when "011101011101110", -- t[15086] = 7
      "00111" when "011101011101111", -- t[15087] = 7
      "00111" when "011101011110000", -- t[15088] = 7
      "00111" when "011101011110001", -- t[15089] = 7
      "00111" when "011101011110010", -- t[15090] = 7
      "00111" when "011101011110011", -- t[15091] = 7
      "00111" when "011101011110100", -- t[15092] = 7
      "00111" when "011101011110101", -- t[15093] = 7
      "00111" when "011101011110110", -- t[15094] = 7
      "00111" when "011101011110111", -- t[15095] = 7
      "00111" when "011101011111000", -- t[15096] = 7
      "00111" when "011101011111001", -- t[15097] = 7
      "00111" when "011101011111010", -- t[15098] = 7
      "00111" when "011101011111011", -- t[15099] = 7
      "00111" when "011101011111100", -- t[15100] = 7
      "00111" when "011101011111101", -- t[15101] = 7
      "00111" when "011101011111110", -- t[15102] = 7
      "00111" when "011101011111111", -- t[15103] = 7
      "00111" when "011101100000000", -- t[15104] = 7
      "00111" when "011101100000001", -- t[15105] = 7
      "00111" when "011101100000010", -- t[15106] = 7
      "01000" when "011101100000011", -- t[15107] = 8
      "01000" when "011101100000100", -- t[15108] = 8
      "01000" when "011101100000101", -- t[15109] = 8
      "01000" when "011101100000110", -- t[15110] = 8
      "01000" when "011101100000111", -- t[15111] = 8
      "01000" when "011101100001000", -- t[15112] = 8
      "01000" when "011101100001001", -- t[15113] = 8
      "01000" when "011101100001010", -- t[15114] = 8
      "01000" when "011101100001011", -- t[15115] = 8
      "01000" when "011101100001100", -- t[15116] = 8
      "01000" when "011101100001101", -- t[15117] = 8
      "01000" when "011101100001110", -- t[15118] = 8
      "01000" when "011101100001111", -- t[15119] = 8
      "01000" when "011101100010000", -- t[15120] = 8
      "01000" when "011101100010001", -- t[15121] = 8
      "01000" when "011101100010010", -- t[15122] = 8
      "01000" when "011101100010011", -- t[15123] = 8
      "01000" when "011101100010100", -- t[15124] = 8
      "01000" when "011101100010101", -- t[15125] = 8
      "01000" when "011101100010110", -- t[15126] = 8
      "01000" when "011101100010111", -- t[15127] = 8
      "01000" when "011101100011000", -- t[15128] = 8
      "01000" when "011101100011001", -- t[15129] = 8
      "01000" when "011101100011010", -- t[15130] = 8
      "01000" when "011101100011011", -- t[15131] = 8
      "01000" when "011101100011100", -- t[15132] = 8
      "01000" when "011101100011101", -- t[15133] = 8
      "01000" when "011101100011110", -- t[15134] = 8
      "01000" when "011101100011111", -- t[15135] = 8
      "01000" when "011101100100000", -- t[15136] = 8
      "01000" when "011101100100001", -- t[15137] = 8
      "01000" when "011101100100010", -- t[15138] = 8
      "01000" when "011101100100011", -- t[15139] = 8
      "01000" when "011101100100100", -- t[15140] = 8
      "01000" when "011101100100101", -- t[15141] = 8
      "01000" when "011101100100110", -- t[15142] = 8
      "01000" when "011101100100111", -- t[15143] = 8
      "01000" when "011101100101000", -- t[15144] = 8
      "01000" when "011101100101001", -- t[15145] = 8
      "01000" when "011101100101010", -- t[15146] = 8
      "01000" when "011101100101011", -- t[15147] = 8
      "01000" when "011101100101100", -- t[15148] = 8
      "01000" when "011101100101101", -- t[15149] = 8
      "01000" when "011101100101110", -- t[15150] = 8
      "01000" when "011101100101111", -- t[15151] = 8
      "01000" when "011101100110000", -- t[15152] = 8
      "01000" when "011101100110001", -- t[15153] = 8
      "01000" when "011101100110010", -- t[15154] = 8
      "01000" when "011101100110011", -- t[15155] = 8
      "01000" when "011101100110100", -- t[15156] = 8
      "01000" when "011101100110101", -- t[15157] = 8
      "01000" when "011101100110110", -- t[15158] = 8
      "01000" when "011101100110111", -- t[15159] = 8
      "01000" when "011101100111000", -- t[15160] = 8
      "01000" when "011101100111001", -- t[15161] = 8
      "01000" when "011101100111010", -- t[15162] = 8
      "01000" when "011101100111011", -- t[15163] = 8
      "01000" when "011101100111100", -- t[15164] = 8
      "01000" when "011101100111101", -- t[15165] = 8
      "01000" when "011101100111110", -- t[15166] = 8
      "01000" when "011101100111111", -- t[15167] = 8
      "01000" when "011101101000000", -- t[15168] = 8
      "01000" when "011101101000001", -- t[15169] = 8
      "01000" when "011101101000010", -- t[15170] = 8
      "01000" when "011101101000011", -- t[15171] = 8
      "01000" when "011101101000100", -- t[15172] = 8
      "01000" when "011101101000101", -- t[15173] = 8
      "01000" when "011101101000110", -- t[15174] = 8
      "01000" when "011101101000111", -- t[15175] = 8
      "01000" when "011101101001000", -- t[15176] = 8
      "01000" when "011101101001001", -- t[15177] = 8
      "01000" when "011101101001010", -- t[15178] = 8
      "01000" when "011101101001011", -- t[15179] = 8
      "01000" when "011101101001100", -- t[15180] = 8
      "01000" when "011101101001101", -- t[15181] = 8
      "01000" when "011101101001110", -- t[15182] = 8
      "01000" when "011101101001111", -- t[15183] = 8
      "01000" when "011101101010000", -- t[15184] = 8
      "01000" when "011101101010001", -- t[15185] = 8
      "01000" when "011101101010010", -- t[15186] = 8
      "01000" when "011101101010011", -- t[15187] = 8
      "01000" when "011101101010100", -- t[15188] = 8
      "01000" when "011101101010101", -- t[15189] = 8
      "01000" when "011101101010110", -- t[15190] = 8
      "01000" when "011101101010111", -- t[15191] = 8
      "01000" when "011101101011000", -- t[15192] = 8
      "01000" when "011101101011001", -- t[15193] = 8
      "01000" when "011101101011010", -- t[15194] = 8
      "01000" when "011101101011011", -- t[15195] = 8
      "01000" when "011101101011100", -- t[15196] = 8
      "01000" when "011101101011101", -- t[15197] = 8
      "01000" when "011101101011110", -- t[15198] = 8
      "01000" when "011101101011111", -- t[15199] = 8
      "01000" when "011101101100000", -- t[15200] = 8
      "01000" when "011101101100001", -- t[15201] = 8
      "01000" when "011101101100010", -- t[15202] = 8
      "01000" when "011101101100011", -- t[15203] = 8
      "01000" when "011101101100100", -- t[15204] = 8
      "01000" when "011101101100101", -- t[15205] = 8
      "01000" when "011101101100110", -- t[15206] = 8
      "01000" when "011101101100111", -- t[15207] = 8
      "01000" when "011101101101000", -- t[15208] = 8
      "01000" when "011101101101001", -- t[15209] = 8
      "01000" when "011101101101010", -- t[15210] = 8
      "01000" when "011101101101011", -- t[15211] = 8
      "01000" when "011101101101100", -- t[15212] = 8
      "01000" when "011101101101101", -- t[15213] = 8
      "01000" when "011101101101110", -- t[15214] = 8
      "01000" when "011101101101111", -- t[15215] = 8
      "01000" when "011101101110000", -- t[15216] = 8
      "01000" when "011101101110001", -- t[15217] = 8
      "01000" when "011101101110010", -- t[15218] = 8
      "01000" when "011101101110011", -- t[15219] = 8
      "01000" when "011101101110100", -- t[15220] = 8
      "01000" when "011101101110101", -- t[15221] = 8
      "01000" when "011101101110110", -- t[15222] = 8
      "01000" when "011101101110111", -- t[15223] = 8
      "01000" when "011101101111000", -- t[15224] = 8
      "01000" when "011101101111001", -- t[15225] = 8
      "01000" when "011101101111010", -- t[15226] = 8
      "01000" when "011101101111011", -- t[15227] = 8
      "01000" when "011101101111100", -- t[15228] = 8
      "01000" when "011101101111101", -- t[15229] = 8
      "01000" when "011101101111110", -- t[15230] = 8
      "01000" when "011101101111111", -- t[15231] = 8
      "01000" when "011101110000000", -- t[15232] = 8
      "01000" when "011101110000001", -- t[15233] = 8
      "01000" when "011101110000010", -- t[15234] = 8
      "01000" when "011101110000011", -- t[15235] = 8
      "01000" when "011101110000100", -- t[15236] = 8
      "01000" when "011101110000101", -- t[15237] = 8
      "01000" when "011101110000110", -- t[15238] = 8
      "01000" when "011101110000111", -- t[15239] = 8
      "01000" when "011101110001000", -- t[15240] = 8
      "01000" when "011101110001001", -- t[15241] = 8
      "01000" when "011101110001010", -- t[15242] = 8
      "01000" when "011101110001011", -- t[15243] = 8
      "01000" when "011101110001100", -- t[15244] = 8
      "01000" when "011101110001101", -- t[15245] = 8
      "01000" when "011101110001110", -- t[15246] = 8
      "01000" when "011101110001111", -- t[15247] = 8
      "01000" when "011101110010000", -- t[15248] = 8
      "01000" when "011101110010001", -- t[15249] = 8
      "01000" when "011101110010010", -- t[15250] = 8
      "01000" when "011101110010011", -- t[15251] = 8
      "01000" when "011101110010100", -- t[15252] = 8
      "01000" when "011101110010101", -- t[15253] = 8
      "01000" when "011101110010110", -- t[15254] = 8
      "01000" when "011101110010111", -- t[15255] = 8
      "01000" when "011101110011000", -- t[15256] = 8
      "01000" when "011101110011001", -- t[15257] = 8
      "01000" when "011101110011010", -- t[15258] = 8
      "01000" when "011101110011011", -- t[15259] = 8
      "01000" when "011101110011100", -- t[15260] = 8
      "01000" when "011101110011101", -- t[15261] = 8
      "01000" when "011101110011110", -- t[15262] = 8
      "01000" when "011101110011111", -- t[15263] = 8
      "01000" when "011101110100000", -- t[15264] = 8
      "01000" when "011101110100001", -- t[15265] = 8
      "01000" when "011101110100010", -- t[15266] = 8
      "01000" when "011101110100011", -- t[15267] = 8
      "01000" when "011101110100100", -- t[15268] = 8
      "01000" when "011101110100101", -- t[15269] = 8
      "01000" when "011101110100110", -- t[15270] = 8
      "01000" when "011101110100111", -- t[15271] = 8
      "01000" when "011101110101000", -- t[15272] = 8
      "01000" when "011101110101001", -- t[15273] = 8
      "01000" when "011101110101010", -- t[15274] = 8
      "01000" when "011101110101011", -- t[15275] = 8
      "01000" when "011101110101100", -- t[15276] = 8
      "01000" when "011101110101101", -- t[15277] = 8
      "01000" when "011101110101110", -- t[15278] = 8
      "01000" when "011101110101111", -- t[15279] = 8
      "01000" when "011101110110000", -- t[15280] = 8
      "01000" when "011101110110001", -- t[15281] = 8
      "01000" when "011101110110010", -- t[15282] = 8
      "01000" when "011101110110011", -- t[15283] = 8
      "01000" when "011101110110100", -- t[15284] = 8
      "01000" when "011101110110101", -- t[15285] = 8
      "01000" when "011101110110110", -- t[15286] = 8
      "01000" when "011101110110111", -- t[15287] = 8
      "01000" when "011101110111000", -- t[15288] = 8
      "01000" when "011101110111001", -- t[15289] = 8
      "01000" when "011101110111010", -- t[15290] = 8
      "01000" when "011101110111011", -- t[15291] = 8
      "01000" when "011101110111100", -- t[15292] = 8
      "01000" when "011101110111101", -- t[15293] = 8
      "01000" when "011101110111110", -- t[15294] = 8
      "01000" when "011101110111111", -- t[15295] = 8
      "01000" when "011101111000000", -- t[15296] = 8
      "01000" when "011101111000001", -- t[15297] = 8
      "01000" when "011101111000010", -- t[15298] = 8
      "01000" when "011101111000011", -- t[15299] = 8
      "01000" when "011101111000100", -- t[15300] = 8
      "01000" when "011101111000101", -- t[15301] = 8
      "01000" when "011101111000110", -- t[15302] = 8
      "01000" when "011101111000111", -- t[15303] = 8
      "01000" when "011101111001000", -- t[15304] = 8
      "01000" when "011101111001001", -- t[15305] = 8
      "01000" when "011101111001010", -- t[15306] = 8
      "01000" when "011101111001011", -- t[15307] = 8
      "01000" when "011101111001100", -- t[15308] = 8
      "01000" when "011101111001101", -- t[15309] = 8
      "01000" when "011101111001110", -- t[15310] = 8
      "01000" when "011101111001111", -- t[15311] = 8
      "01000" when "011101111010000", -- t[15312] = 8
      "01000" when "011101111010001", -- t[15313] = 8
      "01000" when "011101111010010", -- t[15314] = 8
      "01000" when "011101111010011", -- t[15315] = 8
      "01000" when "011101111010100", -- t[15316] = 8
      "01000" when "011101111010101", -- t[15317] = 8
      "01000" when "011101111010110", -- t[15318] = 8
      "01000" when "011101111010111", -- t[15319] = 8
      "01000" when "011101111011000", -- t[15320] = 8
      "01000" when "011101111011001", -- t[15321] = 8
      "01000" when "011101111011010", -- t[15322] = 8
      "01000" when "011101111011011", -- t[15323] = 8
      "01000" when "011101111011100", -- t[15324] = 8
      "01000" when "011101111011101", -- t[15325] = 8
      "01000" when "011101111011110", -- t[15326] = 8
      "01000" when "011101111011111", -- t[15327] = 8
      "01000" when "011101111100000", -- t[15328] = 8
      "01000" when "011101111100001", -- t[15329] = 8
      "01000" when "011101111100010", -- t[15330] = 8
      "01000" when "011101111100011", -- t[15331] = 8
      "01000" when "011101111100100", -- t[15332] = 8
      "01000" when "011101111100101", -- t[15333] = 8
      "01000" when "011101111100110", -- t[15334] = 8
      "01000" when "011101111100111", -- t[15335] = 8
      "01000" when "011101111101000", -- t[15336] = 8
      "01000" when "011101111101001", -- t[15337] = 8
      "01000" when "011101111101010", -- t[15338] = 8
      "01000" when "011101111101011", -- t[15339] = 8
      "01000" when "011101111101100", -- t[15340] = 8
      "01000" when "011101111101101", -- t[15341] = 8
      "01000" when "011101111101110", -- t[15342] = 8
      "01000" when "011101111101111", -- t[15343] = 8
      "01000" when "011101111110000", -- t[15344] = 8
      "01000" when "011101111110001", -- t[15345] = 8
      "01000" when "011101111110010", -- t[15346] = 8
      "01000" when "011101111110011", -- t[15347] = 8
      "01000" when "011101111110100", -- t[15348] = 8
      "01000" when "011101111110101", -- t[15349] = 8
      "01000" when "011101111110110", -- t[15350] = 8
      "01000" when "011101111110111", -- t[15351] = 8
      "01000" when "011101111111000", -- t[15352] = 8
      "01000" when "011101111111001", -- t[15353] = 8
      "01000" when "011101111111010", -- t[15354] = 8
      "01000" when "011101111111011", -- t[15355] = 8
      "01000" when "011101111111100", -- t[15356] = 8
      "01000" when "011101111111101", -- t[15357] = 8
      "01000" when "011101111111110", -- t[15358] = 8
      "01000" when "011101111111111", -- t[15359] = 8
      "01000" when "011110000000000", -- t[15360] = 8
      "01000" when "011110000000001", -- t[15361] = 8
      "01000" when "011110000000010", -- t[15362] = 8
      "01000" when "011110000000011", -- t[15363] = 8
      "01000" when "011110000000100", -- t[15364] = 8
      "01000" when "011110000000101", -- t[15365] = 8
      "01000" when "011110000000110", -- t[15366] = 8
      "01000" when "011110000000111", -- t[15367] = 8
      "01000" when "011110000001000", -- t[15368] = 8
      "01000" when "011110000001001", -- t[15369] = 8
      "01000" when "011110000001010", -- t[15370] = 8
      "01000" when "011110000001011", -- t[15371] = 8
      "01000" when "011110000001100", -- t[15372] = 8
      "01000" when "011110000001101", -- t[15373] = 8
      "01000" when "011110000001110", -- t[15374] = 8
      "01000" when "011110000001111", -- t[15375] = 8
      "01000" when "011110000010000", -- t[15376] = 8
      "01000" when "011110000010001", -- t[15377] = 8
      "01000" when "011110000010010", -- t[15378] = 8
      "01000" when "011110000010011", -- t[15379] = 8
      "01000" when "011110000010100", -- t[15380] = 8
      "01000" when "011110000010101", -- t[15381] = 8
      "01000" when "011110000010110", -- t[15382] = 8
      "01000" when "011110000010111", -- t[15383] = 8
      "01000" when "011110000011000", -- t[15384] = 8
      "01000" when "011110000011001", -- t[15385] = 8
      "01000" when "011110000011010", -- t[15386] = 8
      "01000" when "011110000011011", -- t[15387] = 8
      "01000" when "011110000011100", -- t[15388] = 8
      "01000" when "011110000011101", -- t[15389] = 8
      "01000" when "011110000011110", -- t[15390] = 8
      "01000" when "011110000011111", -- t[15391] = 8
      "01000" when "011110000100000", -- t[15392] = 8
      "01000" when "011110000100001", -- t[15393] = 8
      "01000" when "011110000100010", -- t[15394] = 8
      "01000" when "011110000100011", -- t[15395] = 8
      "01000" when "011110000100100", -- t[15396] = 8
      "01000" when "011110000100101", -- t[15397] = 8
      "01000" when "011110000100110", -- t[15398] = 8
      "01000" when "011110000100111", -- t[15399] = 8
      "01000" when "011110000101000", -- t[15400] = 8
      "01000" when "011110000101001", -- t[15401] = 8
      "01000" when "011110000101010", -- t[15402] = 8
      "01000" when "011110000101011", -- t[15403] = 8
      "01000" when "011110000101100", -- t[15404] = 8
      "01000" when "011110000101101", -- t[15405] = 8
      "01000" when "011110000101110", -- t[15406] = 8
      "01000" when "011110000101111", -- t[15407] = 8
      "01000" when "011110000110000", -- t[15408] = 8
      "01000" when "011110000110001", -- t[15409] = 8
      "01000" when "011110000110010", -- t[15410] = 8
      "01000" when "011110000110011", -- t[15411] = 8
      "01000" when "011110000110100", -- t[15412] = 8
      "01000" when "011110000110101", -- t[15413] = 8
      "01000" when "011110000110110", -- t[15414] = 8
      "01000" when "011110000110111", -- t[15415] = 8
      "01000" when "011110000111000", -- t[15416] = 8
      "01000" when "011110000111001", -- t[15417] = 8
      "01000" when "011110000111010", -- t[15418] = 8
      "01000" when "011110000111011", -- t[15419] = 8
      "01000" when "011110000111100", -- t[15420] = 8
      "01000" when "011110000111101", -- t[15421] = 8
      "01000" when "011110000111110", -- t[15422] = 8
      "01000" when "011110000111111", -- t[15423] = 8
      "01000" when "011110001000000", -- t[15424] = 8
      "01000" when "011110001000001", -- t[15425] = 8
      "01000" when "011110001000010", -- t[15426] = 8
      "01000" when "011110001000011", -- t[15427] = 8
      "01000" when "011110001000100", -- t[15428] = 8
      "01000" when "011110001000101", -- t[15429] = 8
      "01000" when "011110001000110", -- t[15430] = 8
      "01000" when "011110001000111", -- t[15431] = 8
      "01000" when "011110001001000", -- t[15432] = 8
      "01000" when "011110001001001", -- t[15433] = 8
      "01000" when "011110001001010", -- t[15434] = 8
      "01000" when "011110001001011", -- t[15435] = 8
      "01000" when "011110001001100", -- t[15436] = 8
      "01000" when "011110001001101", -- t[15437] = 8
      "01000" when "011110001001110", -- t[15438] = 8
      "01000" when "011110001001111", -- t[15439] = 8
      "01000" when "011110001010000", -- t[15440] = 8
      "01000" when "011110001010001", -- t[15441] = 8
      "01000" when "011110001010010", -- t[15442] = 8
      "01000" when "011110001010011", -- t[15443] = 8
      "01000" when "011110001010100", -- t[15444] = 8
      "01000" when "011110001010101", -- t[15445] = 8
      "01000" when "011110001010110", -- t[15446] = 8
      "01000" when "011110001010111", -- t[15447] = 8
      "01000" when "011110001011000", -- t[15448] = 8
      "01000" when "011110001011001", -- t[15449] = 8
      "01000" when "011110001011010", -- t[15450] = 8
      "01000" when "011110001011011", -- t[15451] = 8
      "01000" when "011110001011100", -- t[15452] = 8
      "01000" when "011110001011101", -- t[15453] = 8
      "01000" when "011110001011110", -- t[15454] = 8
      "01000" when "011110001011111", -- t[15455] = 8
      "01000" when "011110001100000", -- t[15456] = 8
      "01000" when "011110001100001", -- t[15457] = 8
      "01000" when "011110001100010", -- t[15458] = 8
      "01000" when "011110001100011", -- t[15459] = 8
      "01000" when "011110001100100", -- t[15460] = 8
      "01000" when "011110001100101", -- t[15461] = 8
      "01000" when "011110001100110", -- t[15462] = 8
      "01000" when "011110001100111", -- t[15463] = 8
      "01000" when "011110001101000", -- t[15464] = 8
      "01000" when "011110001101001", -- t[15465] = 8
      "01000" when "011110001101010", -- t[15466] = 8
      "01000" when "011110001101011", -- t[15467] = 8
      "01000" when "011110001101100", -- t[15468] = 8
      "01000" when "011110001101101", -- t[15469] = 8
      "01000" when "011110001101110", -- t[15470] = 8
      "01000" when "011110001101111", -- t[15471] = 8
      "01000" when "011110001110000", -- t[15472] = 8
      "01000" when "011110001110001", -- t[15473] = 8
      "01000" when "011110001110010", -- t[15474] = 8
      "01000" when "011110001110011", -- t[15475] = 8
      "01001" when "011110001110100", -- t[15476] = 9
      "01001" when "011110001110101", -- t[15477] = 9
      "01001" when "011110001110110", -- t[15478] = 9
      "01001" when "011110001110111", -- t[15479] = 9
      "01001" when "011110001111000", -- t[15480] = 9
      "01001" when "011110001111001", -- t[15481] = 9
      "01001" when "011110001111010", -- t[15482] = 9
      "01001" when "011110001111011", -- t[15483] = 9
      "01001" when "011110001111100", -- t[15484] = 9
      "01001" when "011110001111101", -- t[15485] = 9
      "01001" when "011110001111110", -- t[15486] = 9
      "01001" when "011110001111111", -- t[15487] = 9
      "01001" when "011110010000000", -- t[15488] = 9
      "01001" when "011110010000001", -- t[15489] = 9
      "01001" when "011110010000010", -- t[15490] = 9
      "01001" when "011110010000011", -- t[15491] = 9
      "01001" when "011110010000100", -- t[15492] = 9
      "01001" when "011110010000101", -- t[15493] = 9
      "01001" when "011110010000110", -- t[15494] = 9
      "01001" when "011110010000111", -- t[15495] = 9
      "01001" when "011110010001000", -- t[15496] = 9
      "01001" when "011110010001001", -- t[15497] = 9
      "01001" when "011110010001010", -- t[15498] = 9
      "01001" when "011110010001011", -- t[15499] = 9
      "01001" when "011110010001100", -- t[15500] = 9
      "01001" when "011110010001101", -- t[15501] = 9
      "01001" when "011110010001110", -- t[15502] = 9
      "01001" when "011110010001111", -- t[15503] = 9
      "01001" when "011110010010000", -- t[15504] = 9
      "01001" when "011110010010001", -- t[15505] = 9
      "01001" when "011110010010010", -- t[15506] = 9
      "01001" when "011110010010011", -- t[15507] = 9
      "01001" when "011110010010100", -- t[15508] = 9
      "01001" when "011110010010101", -- t[15509] = 9
      "01001" when "011110010010110", -- t[15510] = 9
      "01001" when "011110010010111", -- t[15511] = 9
      "01001" when "011110010011000", -- t[15512] = 9
      "01001" when "011110010011001", -- t[15513] = 9
      "01001" when "011110010011010", -- t[15514] = 9
      "01001" when "011110010011011", -- t[15515] = 9
      "01001" when "011110010011100", -- t[15516] = 9
      "01001" when "011110010011101", -- t[15517] = 9
      "01001" when "011110010011110", -- t[15518] = 9
      "01001" when "011110010011111", -- t[15519] = 9
      "01001" when "011110010100000", -- t[15520] = 9
      "01001" when "011110010100001", -- t[15521] = 9
      "01001" when "011110010100010", -- t[15522] = 9
      "01001" when "011110010100011", -- t[15523] = 9
      "01001" when "011110010100100", -- t[15524] = 9
      "01001" when "011110010100101", -- t[15525] = 9
      "01001" when "011110010100110", -- t[15526] = 9
      "01001" when "011110010100111", -- t[15527] = 9
      "01001" when "011110010101000", -- t[15528] = 9
      "01001" when "011110010101001", -- t[15529] = 9
      "01001" when "011110010101010", -- t[15530] = 9
      "01001" when "011110010101011", -- t[15531] = 9
      "01001" when "011110010101100", -- t[15532] = 9
      "01001" when "011110010101101", -- t[15533] = 9
      "01001" when "011110010101110", -- t[15534] = 9
      "01001" when "011110010101111", -- t[15535] = 9
      "01001" when "011110010110000", -- t[15536] = 9
      "01001" when "011110010110001", -- t[15537] = 9
      "01001" when "011110010110010", -- t[15538] = 9
      "01001" when "011110010110011", -- t[15539] = 9
      "01001" when "011110010110100", -- t[15540] = 9
      "01001" when "011110010110101", -- t[15541] = 9
      "01001" when "011110010110110", -- t[15542] = 9
      "01001" when "011110010110111", -- t[15543] = 9
      "01001" when "011110010111000", -- t[15544] = 9
      "01001" when "011110010111001", -- t[15545] = 9
      "01001" when "011110010111010", -- t[15546] = 9
      "01001" when "011110010111011", -- t[15547] = 9
      "01001" when "011110010111100", -- t[15548] = 9
      "01001" when "011110010111101", -- t[15549] = 9
      "01001" when "011110010111110", -- t[15550] = 9
      "01001" when "011110010111111", -- t[15551] = 9
      "01001" when "011110011000000", -- t[15552] = 9
      "01001" when "011110011000001", -- t[15553] = 9
      "01001" when "011110011000010", -- t[15554] = 9
      "01001" when "011110011000011", -- t[15555] = 9
      "01001" when "011110011000100", -- t[15556] = 9
      "01001" when "011110011000101", -- t[15557] = 9
      "01001" when "011110011000110", -- t[15558] = 9
      "01001" when "011110011000111", -- t[15559] = 9
      "01001" when "011110011001000", -- t[15560] = 9
      "01001" when "011110011001001", -- t[15561] = 9
      "01001" when "011110011001010", -- t[15562] = 9
      "01001" when "011110011001011", -- t[15563] = 9
      "01001" when "011110011001100", -- t[15564] = 9
      "01001" when "011110011001101", -- t[15565] = 9
      "01001" when "011110011001110", -- t[15566] = 9
      "01001" when "011110011001111", -- t[15567] = 9
      "01001" when "011110011010000", -- t[15568] = 9
      "01001" when "011110011010001", -- t[15569] = 9
      "01001" when "011110011010010", -- t[15570] = 9
      "01001" when "011110011010011", -- t[15571] = 9
      "01001" when "011110011010100", -- t[15572] = 9
      "01001" when "011110011010101", -- t[15573] = 9
      "01001" when "011110011010110", -- t[15574] = 9
      "01001" when "011110011010111", -- t[15575] = 9
      "01001" when "011110011011000", -- t[15576] = 9
      "01001" when "011110011011001", -- t[15577] = 9
      "01001" when "011110011011010", -- t[15578] = 9
      "01001" when "011110011011011", -- t[15579] = 9
      "01001" when "011110011011100", -- t[15580] = 9
      "01001" when "011110011011101", -- t[15581] = 9
      "01001" when "011110011011110", -- t[15582] = 9
      "01001" when "011110011011111", -- t[15583] = 9
      "01001" when "011110011100000", -- t[15584] = 9
      "01001" when "011110011100001", -- t[15585] = 9
      "01001" when "011110011100010", -- t[15586] = 9
      "01001" when "011110011100011", -- t[15587] = 9
      "01001" when "011110011100100", -- t[15588] = 9
      "01001" when "011110011100101", -- t[15589] = 9
      "01001" when "011110011100110", -- t[15590] = 9
      "01001" when "011110011100111", -- t[15591] = 9
      "01001" when "011110011101000", -- t[15592] = 9
      "01001" when "011110011101001", -- t[15593] = 9
      "01001" when "011110011101010", -- t[15594] = 9
      "01001" when "011110011101011", -- t[15595] = 9
      "01001" when "011110011101100", -- t[15596] = 9
      "01001" when "011110011101101", -- t[15597] = 9
      "01001" when "011110011101110", -- t[15598] = 9
      "01001" when "011110011101111", -- t[15599] = 9
      "01001" when "011110011110000", -- t[15600] = 9
      "01001" when "011110011110001", -- t[15601] = 9
      "01001" when "011110011110010", -- t[15602] = 9
      "01001" when "011110011110011", -- t[15603] = 9
      "01001" when "011110011110100", -- t[15604] = 9
      "01001" when "011110011110101", -- t[15605] = 9
      "01001" when "011110011110110", -- t[15606] = 9
      "01001" when "011110011110111", -- t[15607] = 9
      "01001" when "011110011111000", -- t[15608] = 9
      "01001" when "011110011111001", -- t[15609] = 9
      "01001" when "011110011111010", -- t[15610] = 9
      "01001" when "011110011111011", -- t[15611] = 9
      "01001" when "011110011111100", -- t[15612] = 9
      "01001" when "011110011111101", -- t[15613] = 9
      "01001" when "011110011111110", -- t[15614] = 9
      "01001" when "011110011111111", -- t[15615] = 9
      "01001" when "011110100000000", -- t[15616] = 9
      "01001" when "011110100000001", -- t[15617] = 9
      "01001" when "011110100000010", -- t[15618] = 9
      "01001" when "011110100000011", -- t[15619] = 9
      "01001" when "011110100000100", -- t[15620] = 9
      "01001" when "011110100000101", -- t[15621] = 9
      "01001" when "011110100000110", -- t[15622] = 9
      "01001" when "011110100000111", -- t[15623] = 9
      "01001" when "011110100001000", -- t[15624] = 9
      "01001" when "011110100001001", -- t[15625] = 9
      "01001" when "011110100001010", -- t[15626] = 9
      "01001" when "011110100001011", -- t[15627] = 9
      "01001" when "011110100001100", -- t[15628] = 9
      "01001" when "011110100001101", -- t[15629] = 9
      "01001" when "011110100001110", -- t[15630] = 9
      "01001" when "011110100001111", -- t[15631] = 9
      "01001" when "011110100010000", -- t[15632] = 9
      "01001" when "011110100010001", -- t[15633] = 9
      "01001" when "011110100010010", -- t[15634] = 9
      "01001" when "011110100010011", -- t[15635] = 9
      "01001" when "011110100010100", -- t[15636] = 9
      "01001" when "011110100010101", -- t[15637] = 9
      "01001" when "011110100010110", -- t[15638] = 9
      "01001" when "011110100010111", -- t[15639] = 9
      "01001" when "011110100011000", -- t[15640] = 9
      "01001" when "011110100011001", -- t[15641] = 9
      "01001" when "011110100011010", -- t[15642] = 9
      "01001" when "011110100011011", -- t[15643] = 9
      "01001" when "011110100011100", -- t[15644] = 9
      "01001" when "011110100011101", -- t[15645] = 9
      "01001" when "011110100011110", -- t[15646] = 9
      "01001" when "011110100011111", -- t[15647] = 9
      "01001" when "011110100100000", -- t[15648] = 9
      "01001" when "011110100100001", -- t[15649] = 9
      "01001" when "011110100100010", -- t[15650] = 9
      "01001" when "011110100100011", -- t[15651] = 9
      "01001" when "011110100100100", -- t[15652] = 9
      "01001" when "011110100100101", -- t[15653] = 9
      "01001" when "011110100100110", -- t[15654] = 9
      "01001" when "011110100100111", -- t[15655] = 9
      "01001" when "011110100101000", -- t[15656] = 9
      "01001" when "011110100101001", -- t[15657] = 9
      "01001" when "011110100101010", -- t[15658] = 9
      "01001" when "011110100101011", -- t[15659] = 9
      "01001" when "011110100101100", -- t[15660] = 9
      "01001" when "011110100101101", -- t[15661] = 9
      "01001" when "011110100101110", -- t[15662] = 9
      "01001" when "011110100101111", -- t[15663] = 9
      "01001" when "011110100110000", -- t[15664] = 9
      "01001" when "011110100110001", -- t[15665] = 9
      "01001" when "011110100110010", -- t[15666] = 9
      "01001" when "011110100110011", -- t[15667] = 9
      "01001" when "011110100110100", -- t[15668] = 9
      "01001" when "011110100110101", -- t[15669] = 9
      "01001" when "011110100110110", -- t[15670] = 9
      "01001" when "011110100110111", -- t[15671] = 9
      "01001" when "011110100111000", -- t[15672] = 9
      "01001" when "011110100111001", -- t[15673] = 9
      "01001" when "011110100111010", -- t[15674] = 9
      "01001" when "011110100111011", -- t[15675] = 9
      "01001" when "011110100111100", -- t[15676] = 9
      "01001" when "011110100111101", -- t[15677] = 9
      "01001" when "011110100111110", -- t[15678] = 9
      "01001" when "011110100111111", -- t[15679] = 9
      "01001" when "011110101000000", -- t[15680] = 9
      "01001" when "011110101000001", -- t[15681] = 9
      "01001" when "011110101000010", -- t[15682] = 9
      "01001" when "011110101000011", -- t[15683] = 9
      "01001" when "011110101000100", -- t[15684] = 9
      "01001" when "011110101000101", -- t[15685] = 9
      "01001" when "011110101000110", -- t[15686] = 9
      "01001" when "011110101000111", -- t[15687] = 9
      "01001" when "011110101001000", -- t[15688] = 9
      "01001" when "011110101001001", -- t[15689] = 9
      "01001" when "011110101001010", -- t[15690] = 9
      "01001" when "011110101001011", -- t[15691] = 9
      "01001" when "011110101001100", -- t[15692] = 9
      "01001" when "011110101001101", -- t[15693] = 9
      "01001" when "011110101001110", -- t[15694] = 9
      "01001" when "011110101001111", -- t[15695] = 9
      "01001" when "011110101010000", -- t[15696] = 9
      "01001" when "011110101010001", -- t[15697] = 9
      "01001" when "011110101010010", -- t[15698] = 9
      "01001" when "011110101010011", -- t[15699] = 9
      "01001" when "011110101010100", -- t[15700] = 9
      "01001" when "011110101010101", -- t[15701] = 9
      "01001" when "011110101010110", -- t[15702] = 9
      "01001" when "011110101010111", -- t[15703] = 9
      "01001" when "011110101011000", -- t[15704] = 9
      "01001" when "011110101011001", -- t[15705] = 9
      "01001" when "011110101011010", -- t[15706] = 9
      "01001" when "011110101011011", -- t[15707] = 9
      "01001" when "011110101011100", -- t[15708] = 9
      "01001" when "011110101011101", -- t[15709] = 9
      "01001" when "011110101011110", -- t[15710] = 9
      "01001" when "011110101011111", -- t[15711] = 9
      "01001" when "011110101100000", -- t[15712] = 9
      "01001" when "011110101100001", -- t[15713] = 9
      "01001" when "011110101100010", -- t[15714] = 9
      "01001" when "011110101100011", -- t[15715] = 9
      "01001" when "011110101100100", -- t[15716] = 9
      "01001" when "011110101100101", -- t[15717] = 9
      "01001" when "011110101100110", -- t[15718] = 9
      "01001" when "011110101100111", -- t[15719] = 9
      "01001" when "011110101101000", -- t[15720] = 9
      "01001" when "011110101101001", -- t[15721] = 9
      "01001" when "011110101101010", -- t[15722] = 9
      "01001" when "011110101101011", -- t[15723] = 9
      "01001" when "011110101101100", -- t[15724] = 9
      "01001" when "011110101101101", -- t[15725] = 9
      "01001" when "011110101101110", -- t[15726] = 9
      "01001" when "011110101101111", -- t[15727] = 9
      "01001" when "011110101110000", -- t[15728] = 9
      "01001" when "011110101110001", -- t[15729] = 9
      "01001" when "011110101110010", -- t[15730] = 9
      "01001" when "011110101110011", -- t[15731] = 9
      "01001" when "011110101110100", -- t[15732] = 9
      "01001" when "011110101110101", -- t[15733] = 9
      "01001" when "011110101110110", -- t[15734] = 9
      "01001" when "011110101110111", -- t[15735] = 9
      "01001" when "011110101111000", -- t[15736] = 9
      "01001" when "011110101111001", -- t[15737] = 9
      "01001" when "011110101111010", -- t[15738] = 9
      "01001" when "011110101111011", -- t[15739] = 9
      "01001" when "011110101111100", -- t[15740] = 9
      "01001" when "011110101111101", -- t[15741] = 9
      "01001" when "011110101111110", -- t[15742] = 9
      "01001" when "011110101111111", -- t[15743] = 9
      "01001" when "011110110000000", -- t[15744] = 9
      "01001" when "011110110000001", -- t[15745] = 9
      "01001" when "011110110000010", -- t[15746] = 9
      "01001" when "011110110000011", -- t[15747] = 9
      "01001" when "011110110000100", -- t[15748] = 9
      "01001" when "011110110000101", -- t[15749] = 9
      "01001" when "011110110000110", -- t[15750] = 9
      "01001" when "011110110000111", -- t[15751] = 9
      "01001" when "011110110001000", -- t[15752] = 9
      "01001" when "011110110001001", -- t[15753] = 9
      "01001" when "011110110001010", -- t[15754] = 9
      "01001" when "011110110001011", -- t[15755] = 9
      "01001" when "011110110001100", -- t[15756] = 9
      "01001" when "011110110001101", -- t[15757] = 9
      "01001" when "011110110001110", -- t[15758] = 9
      "01001" when "011110110001111", -- t[15759] = 9
      "01001" when "011110110010000", -- t[15760] = 9
      "01001" when "011110110010001", -- t[15761] = 9
      "01001" when "011110110010010", -- t[15762] = 9
      "01001" when "011110110010011", -- t[15763] = 9
      "01001" when "011110110010100", -- t[15764] = 9
      "01001" when "011110110010101", -- t[15765] = 9
      "01001" when "011110110010110", -- t[15766] = 9
      "01001" when "011110110010111", -- t[15767] = 9
      "01001" when "011110110011000", -- t[15768] = 9
      "01001" when "011110110011001", -- t[15769] = 9
      "01001" when "011110110011010", -- t[15770] = 9
      "01001" when "011110110011011", -- t[15771] = 9
      "01001" when "011110110011100", -- t[15772] = 9
      "01001" when "011110110011101", -- t[15773] = 9
      "01001" when "011110110011110", -- t[15774] = 9
      "01001" when "011110110011111", -- t[15775] = 9
      "01001" when "011110110100000", -- t[15776] = 9
      "01001" when "011110110100001", -- t[15777] = 9
      "01001" when "011110110100010", -- t[15778] = 9
      "01001" when "011110110100011", -- t[15779] = 9
      "01001" when "011110110100100", -- t[15780] = 9
      "01001" when "011110110100101", -- t[15781] = 9
      "01001" when "011110110100110", -- t[15782] = 9
      "01001" when "011110110100111", -- t[15783] = 9
      "01001" when "011110110101000", -- t[15784] = 9
      "01001" when "011110110101001", -- t[15785] = 9
      "01001" when "011110110101010", -- t[15786] = 9
      "01001" when "011110110101011", -- t[15787] = 9
      "01001" when "011110110101100", -- t[15788] = 9
      "01001" when "011110110101101", -- t[15789] = 9
      "01001" when "011110110101110", -- t[15790] = 9
      "01001" when "011110110101111", -- t[15791] = 9
      "01001" when "011110110110000", -- t[15792] = 9
      "01001" when "011110110110001", -- t[15793] = 9
      "01001" when "011110110110010", -- t[15794] = 9
      "01001" when "011110110110011", -- t[15795] = 9
      "01001" when "011110110110100", -- t[15796] = 9
      "01001" when "011110110110101", -- t[15797] = 9
      "01001" when "011110110110110", -- t[15798] = 9
      "01001" when "011110110110111", -- t[15799] = 9
      "01001" when "011110110111000", -- t[15800] = 9
      "01001" when "011110110111001", -- t[15801] = 9
      "01001" when "011110110111010", -- t[15802] = 9
      "01001" when "011110110111011", -- t[15803] = 9
      "01001" when "011110110111100", -- t[15804] = 9
      "01010" when "011110110111101", -- t[15805] = 10
      "01010" when "011110110111110", -- t[15806] = 10
      "01010" when "011110110111111", -- t[15807] = 10
      "01010" when "011110111000000", -- t[15808] = 10
      "01010" when "011110111000001", -- t[15809] = 10
      "01010" when "011110111000010", -- t[15810] = 10
      "01010" when "011110111000011", -- t[15811] = 10
      "01010" when "011110111000100", -- t[15812] = 10
      "01010" when "011110111000101", -- t[15813] = 10
      "01010" when "011110111000110", -- t[15814] = 10
      "01010" when "011110111000111", -- t[15815] = 10
      "01010" when "011110111001000", -- t[15816] = 10
      "01010" when "011110111001001", -- t[15817] = 10
      "01010" when "011110111001010", -- t[15818] = 10
      "01010" when "011110111001011", -- t[15819] = 10
      "01010" when "011110111001100", -- t[15820] = 10
      "01010" when "011110111001101", -- t[15821] = 10
      "01010" when "011110111001110", -- t[15822] = 10
      "01010" when "011110111001111", -- t[15823] = 10
      "01010" when "011110111010000", -- t[15824] = 10
      "01010" when "011110111010001", -- t[15825] = 10
      "01010" when "011110111010010", -- t[15826] = 10
      "01010" when "011110111010011", -- t[15827] = 10
      "01010" when "011110111010100", -- t[15828] = 10
      "01010" when "011110111010101", -- t[15829] = 10
      "01010" when "011110111010110", -- t[15830] = 10
      "01010" when "011110111010111", -- t[15831] = 10
      "01010" when "011110111011000", -- t[15832] = 10
      "01010" when "011110111011001", -- t[15833] = 10
      "01010" when "011110111011010", -- t[15834] = 10
      "01010" when "011110111011011", -- t[15835] = 10
      "01010" when "011110111011100", -- t[15836] = 10
      "01010" when "011110111011101", -- t[15837] = 10
      "01010" when "011110111011110", -- t[15838] = 10
      "01010" when "011110111011111", -- t[15839] = 10
      "01010" when "011110111100000", -- t[15840] = 10
      "01010" when "011110111100001", -- t[15841] = 10
      "01010" when "011110111100010", -- t[15842] = 10
      "01010" when "011110111100011", -- t[15843] = 10
      "01010" when "011110111100100", -- t[15844] = 10
      "01010" when "011110111100101", -- t[15845] = 10
      "01010" when "011110111100110", -- t[15846] = 10
      "01010" when "011110111100111", -- t[15847] = 10
      "01010" when "011110111101000", -- t[15848] = 10
      "01010" when "011110111101001", -- t[15849] = 10
      "01010" when "011110111101010", -- t[15850] = 10
      "01010" when "011110111101011", -- t[15851] = 10
      "01010" when "011110111101100", -- t[15852] = 10
      "01010" when "011110111101101", -- t[15853] = 10
      "01010" when "011110111101110", -- t[15854] = 10
      "01010" when "011110111101111", -- t[15855] = 10
      "01010" when "011110111110000", -- t[15856] = 10
      "01010" when "011110111110001", -- t[15857] = 10
      "01010" when "011110111110010", -- t[15858] = 10
      "01010" when "011110111110011", -- t[15859] = 10
      "01010" when "011110111110100", -- t[15860] = 10
      "01010" when "011110111110101", -- t[15861] = 10
      "01010" when "011110111110110", -- t[15862] = 10
      "01010" when "011110111110111", -- t[15863] = 10
      "01010" when "011110111111000", -- t[15864] = 10
      "01010" when "011110111111001", -- t[15865] = 10
      "01010" when "011110111111010", -- t[15866] = 10
      "01010" when "011110111111011", -- t[15867] = 10
      "01010" when "011110111111100", -- t[15868] = 10
      "01010" when "011110111111101", -- t[15869] = 10
      "01010" when "011110111111110", -- t[15870] = 10
      "01010" when "011110111111111", -- t[15871] = 10
      "01010" when "011111000000000", -- t[15872] = 10
      "01010" when "011111000000001", -- t[15873] = 10
      "01010" when "011111000000010", -- t[15874] = 10
      "01010" when "011111000000011", -- t[15875] = 10
      "01010" when "011111000000100", -- t[15876] = 10
      "01010" when "011111000000101", -- t[15877] = 10
      "01010" when "011111000000110", -- t[15878] = 10
      "01010" when "011111000000111", -- t[15879] = 10
      "01010" when "011111000001000", -- t[15880] = 10
      "01010" when "011111000001001", -- t[15881] = 10
      "01010" when "011111000001010", -- t[15882] = 10
      "01010" when "011111000001011", -- t[15883] = 10
      "01010" when "011111000001100", -- t[15884] = 10
      "01010" when "011111000001101", -- t[15885] = 10
      "01010" when "011111000001110", -- t[15886] = 10
      "01010" when "011111000001111", -- t[15887] = 10
      "01010" when "011111000010000", -- t[15888] = 10
      "01010" when "011111000010001", -- t[15889] = 10
      "01010" when "011111000010010", -- t[15890] = 10
      "01010" when "011111000010011", -- t[15891] = 10
      "01010" when "011111000010100", -- t[15892] = 10
      "01010" when "011111000010101", -- t[15893] = 10
      "01010" when "011111000010110", -- t[15894] = 10
      "01010" when "011111000010111", -- t[15895] = 10
      "01010" when "011111000011000", -- t[15896] = 10
      "01010" when "011111000011001", -- t[15897] = 10
      "01010" when "011111000011010", -- t[15898] = 10
      "01010" when "011111000011011", -- t[15899] = 10
      "01010" when "011111000011100", -- t[15900] = 10
      "01010" when "011111000011101", -- t[15901] = 10
      "01010" when "011111000011110", -- t[15902] = 10
      "01010" when "011111000011111", -- t[15903] = 10
      "01010" when "011111000100000", -- t[15904] = 10
      "01010" when "011111000100001", -- t[15905] = 10
      "01010" when "011111000100010", -- t[15906] = 10
      "01010" when "011111000100011", -- t[15907] = 10
      "01010" when "011111000100100", -- t[15908] = 10
      "01010" when "011111000100101", -- t[15909] = 10
      "01010" when "011111000100110", -- t[15910] = 10
      "01010" when "011111000100111", -- t[15911] = 10
      "01010" when "011111000101000", -- t[15912] = 10
      "01010" when "011111000101001", -- t[15913] = 10
      "01010" when "011111000101010", -- t[15914] = 10
      "01010" when "011111000101011", -- t[15915] = 10
      "01010" when "011111000101100", -- t[15916] = 10
      "01010" when "011111000101101", -- t[15917] = 10
      "01010" when "011111000101110", -- t[15918] = 10
      "01010" when "011111000101111", -- t[15919] = 10
      "01010" when "011111000110000", -- t[15920] = 10
      "01010" when "011111000110001", -- t[15921] = 10
      "01010" when "011111000110010", -- t[15922] = 10
      "01010" when "011111000110011", -- t[15923] = 10
      "01010" when "011111000110100", -- t[15924] = 10
      "01010" when "011111000110101", -- t[15925] = 10
      "01010" when "011111000110110", -- t[15926] = 10
      "01010" when "011111000110111", -- t[15927] = 10
      "01010" when "011111000111000", -- t[15928] = 10
      "01010" when "011111000111001", -- t[15929] = 10
      "01010" when "011111000111010", -- t[15930] = 10
      "01010" when "011111000111011", -- t[15931] = 10
      "01010" when "011111000111100", -- t[15932] = 10
      "01010" when "011111000111101", -- t[15933] = 10
      "01010" when "011111000111110", -- t[15934] = 10
      "01010" when "011111000111111", -- t[15935] = 10
      "01010" when "011111001000000", -- t[15936] = 10
      "01010" when "011111001000001", -- t[15937] = 10
      "01010" when "011111001000010", -- t[15938] = 10
      "01010" when "011111001000011", -- t[15939] = 10
      "01010" when "011111001000100", -- t[15940] = 10
      "01010" when "011111001000101", -- t[15941] = 10
      "01010" when "011111001000110", -- t[15942] = 10
      "01010" when "011111001000111", -- t[15943] = 10
      "01010" when "011111001001000", -- t[15944] = 10
      "01010" when "011111001001001", -- t[15945] = 10
      "01010" when "011111001001010", -- t[15946] = 10
      "01010" when "011111001001011", -- t[15947] = 10
      "01010" when "011111001001100", -- t[15948] = 10
      "01010" when "011111001001101", -- t[15949] = 10
      "01010" when "011111001001110", -- t[15950] = 10
      "01010" when "011111001001111", -- t[15951] = 10
      "01010" when "011111001010000", -- t[15952] = 10
      "01010" when "011111001010001", -- t[15953] = 10
      "01010" when "011111001010010", -- t[15954] = 10
      "01010" when "011111001010011", -- t[15955] = 10
      "01010" when "011111001010100", -- t[15956] = 10
      "01010" when "011111001010101", -- t[15957] = 10
      "01010" when "011111001010110", -- t[15958] = 10
      "01010" when "011111001010111", -- t[15959] = 10
      "01010" when "011111001011000", -- t[15960] = 10
      "01010" when "011111001011001", -- t[15961] = 10
      "01010" when "011111001011010", -- t[15962] = 10
      "01010" when "011111001011011", -- t[15963] = 10
      "01010" when "011111001011100", -- t[15964] = 10
      "01010" when "011111001011101", -- t[15965] = 10
      "01010" when "011111001011110", -- t[15966] = 10
      "01010" when "011111001011111", -- t[15967] = 10
      "01010" when "011111001100000", -- t[15968] = 10
      "01010" when "011111001100001", -- t[15969] = 10
      "01010" when "011111001100010", -- t[15970] = 10
      "01010" when "011111001100011", -- t[15971] = 10
      "01010" when "011111001100100", -- t[15972] = 10
      "01010" when "011111001100101", -- t[15973] = 10
      "01010" when "011111001100110", -- t[15974] = 10
      "01010" when "011111001100111", -- t[15975] = 10
      "01010" when "011111001101000", -- t[15976] = 10
      "01010" when "011111001101001", -- t[15977] = 10
      "01010" when "011111001101010", -- t[15978] = 10
      "01010" when "011111001101011", -- t[15979] = 10
      "01010" when "011111001101100", -- t[15980] = 10
      "01010" when "011111001101101", -- t[15981] = 10
      "01010" when "011111001101110", -- t[15982] = 10
      "01010" when "011111001101111", -- t[15983] = 10
      "01010" when "011111001110000", -- t[15984] = 10
      "01010" when "011111001110001", -- t[15985] = 10
      "01010" when "011111001110010", -- t[15986] = 10
      "01010" when "011111001110011", -- t[15987] = 10
      "01010" when "011111001110100", -- t[15988] = 10
      "01010" when "011111001110101", -- t[15989] = 10
      "01010" when "011111001110110", -- t[15990] = 10
      "01010" when "011111001110111", -- t[15991] = 10
      "01010" when "011111001111000", -- t[15992] = 10
      "01010" when "011111001111001", -- t[15993] = 10
      "01010" when "011111001111010", -- t[15994] = 10
      "01010" when "011111001111011", -- t[15995] = 10
      "01010" when "011111001111100", -- t[15996] = 10
      "01010" when "011111001111101", -- t[15997] = 10
      "01010" when "011111001111110", -- t[15998] = 10
      "01010" when "011111001111111", -- t[15999] = 10
      "01010" when "011111010000000", -- t[16000] = 10
      "01010" when "011111010000001", -- t[16001] = 10
      "01010" when "011111010000010", -- t[16002] = 10
      "01010" when "011111010000011", -- t[16003] = 10
      "01010" when "011111010000100", -- t[16004] = 10
      "01010" when "011111010000101", -- t[16005] = 10
      "01010" when "011111010000110", -- t[16006] = 10
      "01010" when "011111010000111", -- t[16007] = 10
      "01010" when "011111010001000", -- t[16008] = 10
      "01010" when "011111010001001", -- t[16009] = 10
      "01010" when "011111010001010", -- t[16010] = 10
      "01010" when "011111010001011", -- t[16011] = 10
      "01010" when "011111010001100", -- t[16012] = 10
      "01010" when "011111010001101", -- t[16013] = 10
      "01010" when "011111010001110", -- t[16014] = 10
      "01010" when "011111010001111", -- t[16015] = 10
      "01010" when "011111010010000", -- t[16016] = 10
      "01010" when "011111010010001", -- t[16017] = 10
      "01010" when "011111010010010", -- t[16018] = 10
      "01010" when "011111010010011", -- t[16019] = 10
      "01010" when "011111010010100", -- t[16020] = 10
      "01010" when "011111010010101", -- t[16021] = 10
      "01010" when "011111010010110", -- t[16022] = 10
      "01010" when "011111010010111", -- t[16023] = 10
      "01010" when "011111010011000", -- t[16024] = 10
      "01010" when "011111010011001", -- t[16025] = 10
      "01010" when "011111010011010", -- t[16026] = 10
      "01010" when "011111010011011", -- t[16027] = 10
      "01010" when "011111010011100", -- t[16028] = 10
      "01010" when "011111010011101", -- t[16029] = 10
      "01010" when "011111010011110", -- t[16030] = 10
      "01010" when "011111010011111", -- t[16031] = 10
      "01010" when "011111010100000", -- t[16032] = 10
      "01010" when "011111010100001", -- t[16033] = 10
      "01010" when "011111010100010", -- t[16034] = 10
      "01010" when "011111010100011", -- t[16035] = 10
      "01010" when "011111010100100", -- t[16036] = 10
      "01010" when "011111010100101", -- t[16037] = 10
      "01010" when "011111010100110", -- t[16038] = 10
      "01010" when "011111010100111", -- t[16039] = 10
      "01010" when "011111010101000", -- t[16040] = 10
      "01010" when "011111010101001", -- t[16041] = 10
      "01010" when "011111010101010", -- t[16042] = 10
      "01010" when "011111010101011", -- t[16043] = 10
      "01010" when "011111010101100", -- t[16044] = 10
      "01010" when "011111010101101", -- t[16045] = 10
      "01010" when "011111010101110", -- t[16046] = 10
      "01010" when "011111010101111", -- t[16047] = 10
      "01010" when "011111010110000", -- t[16048] = 10
      "01010" when "011111010110001", -- t[16049] = 10
      "01010" when "011111010110010", -- t[16050] = 10
      "01010" when "011111010110011", -- t[16051] = 10
      "01010" when "011111010110100", -- t[16052] = 10
      "01010" when "011111010110101", -- t[16053] = 10
      "01010" when "011111010110110", -- t[16054] = 10
      "01010" when "011111010110111", -- t[16055] = 10
      "01010" when "011111010111000", -- t[16056] = 10
      "01010" when "011111010111001", -- t[16057] = 10
      "01010" when "011111010111010", -- t[16058] = 10
      "01010" when "011111010111011", -- t[16059] = 10
      "01010" when "011111010111100", -- t[16060] = 10
      "01010" when "011111010111101", -- t[16061] = 10
      "01010" when "011111010111110", -- t[16062] = 10
      "01010" when "011111010111111", -- t[16063] = 10
      "01010" when "011111011000000", -- t[16064] = 10
      "01010" when "011111011000001", -- t[16065] = 10
      "01010" when "011111011000010", -- t[16066] = 10
      "01010" when "011111011000011", -- t[16067] = 10
      "01010" when "011111011000100", -- t[16068] = 10
      "01010" when "011111011000101", -- t[16069] = 10
      "01010" when "011111011000110", -- t[16070] = 10
      "01010" when "011111011000111", -- t[16071] = 10
      "01010" when "011111011001000", -- t[16072] = 10
      "01010" when "011111011001001", -- t[16073] = 10
      "01010" when "011111011001010", -- t[16074] = 10
      "01010" when "011111011001011", -- t[16075] = 10
      "01010" when "011111011001100", -- t[16076] = 10
      "01010" when "011111011001101", -- t[16077] = 10
      "01010" when "011111011001110", -- t[16078] = 10
      "01010" when "011111011001111", -- t[16079] = 10
      "01010" when "011111011010000", -- t[16080] = 10
      "01010" when "011111011010001", -- t[16081] = 10
      "01010" when "011111011010010", -- t[16082] = 10
      "01010" when "011111011010011", -- t[16083] = 10
      "01010" when "011111011010100", -- t[16084] = 10
      "01010" when "011111011010101", -- t[16085] = 10
      "01010" when "011111011010110", -- t[16086] = 10
      "01010" when "011111011010111", -- t[16087] = 10
      "01010" when "011111011011000", -- t[16088] = 10
      "01010" when "011111011011001", -- t[16089] = 10
      "01010" when "011111011011010", -- t[16090] = 10
      "01010" when "011111011011011", -- t[16091] = 10
      "01010" when "011111011011100", -- t[16092] = 10
      "01010" when "011111011011101", -- t[16093] = 10
      "01010" when "011111011011110", -- t[16094] = 10
      "01010" when "011111011011111", -- t[16095] = 10
      "01010" when "011111011100000", -- t[16096] = 10
      "01010" when "011111011100001", -- t[16097] = 10
      "01010" when "011111011100010", -- t[16098] = 10
      "01010" when "011111011100011", -- t[16099] = 10
      "01011" when "011111011100100", -- t[16100] = 11
      "01011" when "011111011100101", -- t[16101] = 11
      "01011" when "011111011100110", -- t[16102] = 11
      "01011" when "011111011100111", -- t[16103] = 11
      "01011" when "011111011101000", -- t[16104] = 11
      "01011" when "011111011101001", -- t[16105] = 11
      "01011" when "011111011101010", -- t[16106] = 11
      "01011" when "011111011101011", -- t[16107] = 11
      "01011" when "011111011101100", -- t[16108] = 11
      "01011" when "011111011101101", -- t[16109] = 11
      "01011" when "011111011101110", -- t[16110] = 11
      "01011" when "011111011101111", -- t[16111] = 11
      "01011" when "011111011110000", -- t[16112] = 11
      "01011" when "011111011110001", -- t[16113] = 11
      "01011" when "011111011110010", -- t[16114] = 11
      "01011" when "011111011110011", -- t[16115] = 11
      "01011" when "011111011110100", -- t[16116] = 11
      "01011" when "011111011110101", -- t[16117] = 11
      "01011" when "011111011110110", -- t[16118] = 11
      "01011" when "011111011110111", -- t[16119] = 11
      "01011" when "011111011111000", -- t[16120] = 11
      "01011" when "011111011111001", -- t[16121] = 11
      "01011" when "011111011111010", -- t[16122] = 11
      "01011" when "011111011111011", -- t[16123] = 11
      "01011" when "011111011111100", -- t[16124] = 11
      "01011" when "011111011111101", -- t[16125] = 11
      "01011" when "011111011111110", -- t[16126] = 11
      "01011" when "011111011111111", -- t[16127] = 11
      "01011" when "011111100000000", -- t[16128] = 11
      "01011" when "011111100000001", -- t[16129] = 11
      "01011" when "011111100000010", -- t[16130] = 11
      "01011" when "011111100000011", -- t[16131] = 11
      "01011" when "011111100000100", -- t[16132] = 11
      "01011" when "011111100000101", -- t[16133] = 11
      "01011" when "011111100000110", -- t[16134] = 11
      "01011" when "011111100000111", -- t[16135] = 11
      "01011" when "011111100001000", -- t[16136] = 11
      "01011" when "011111100001001", -- t[16137] = 11
      "01011" when "011111100001010", -- t[16138] = 11
      "01011" when "011111100001011", -- t[16139] = 11
      "01011" when "011111100001100", -- t[16140] = 11
      "01011" when "011111100001101", -- t[16141] = 11
      "01011" when "011111100001110", -- t[16142] = 11
      "01011" when "011111100001111", -- t[16143] = 11
      "01011" when "011111100010000", -- t[16144] = 11
      "01011" when "011111100010001", -- t[16145] = 11
      "01011" when "011111100010010", -- t[16146] = 11
      "01011" when "011111100010011", -- t[16147] = 11
      "01011" when "011111100010100", -- t[16148] = 11
      "01011" when "011111100010101", -- t[16149] = 11
      "01011" when "011111100010110", -- t[16150] = 11
      "01011" when "011111100010111", -- t[16151] = 11
      "01011" when "011111100011000", -- t[16152] = 11
      "01011" when "011111100011001", -- t[16153] = 11
      "01011" when "011111100011010", -- t[16154] = 11
      "01011" when "011111100011011", -- t[16155] = 11
      "01011" when "011111100011100", -- t[16156] = 11
      "01011" when "011111100011101", -- t[16157] = 11
      "01011" when "011111100011110", -- t[16158] = 11
      "01011" when "011111100011111", -- t[16159] = 11
      "01011" when "011111100100000", -- t[16160] = 11
      "01011" when "011111100100001", -- t[16161] = 11
      "01011" when "011111100100010", -- t[16162] = 11
      "01011" when "011111100100011", -- t[16163] = 11
      "01011" when "011111100100100", -- t[16164] = 11
      "01011" when "011111100100101", -- t[16165] = 11
      "01011" when "011111100100110", -- t[16166] = 11
      "01011" when "011111100100111", -- t[16167] = 11
      "01011" when "011111100101000", -- t[16168] = 11
      "01011" when "011111100101001", -- t[16169] = 11
      "01011" when "011111100101010", -- t[16170] = 11
      "01011" when "011111100101011", -- t[16171] = 11
      "01011" when "011111100101100", -- t[16172] = 11
      "01011" when "011111100101101", -- t[16173] = 11
      "01011" when "011111100101110", -- t[16174] = 11
      "01011" when "011111100101111", -- t[16175] = 11
      "01011" when "011111100110000", -- t[16176] = 11
      "01011" when "011111100110001", -- t[16177] = 11
      "01011" when "011111100110010", -- t[16178] = 11
      "01011" when "011111100110011", -- t[16179] = 11
      "01011" when "011111100110100", -- t[16180] = 11
      "01011" when "011111100110101", -- t[16181] = 11
      "01011" when "011111100110110", -- t[16182] = 11
      "01011" when "011111100110111", -- t[16183] = 11
      "01011" when "011111100111000", -- t[16184] = 11
      "01011" when "011111100111001", -- t[16185] = 11
      "01011" when "011111100111010", -- t[16186] = 11
      "01011" when "011111100111011", -- t[16187] = 11
      "01011" when "011111100111100", -- t[16188] = 11
      "01011" when "011111100111101", -- t[16189] = 11
      "01011" when "011111100111110", -- t[16190] = 11
      "01011" when "011111100111111", -- t[16191] = 11
      "01011" when "011111101000000", -- t[16192] = 11
      "01011" when "011111101000001", -- t[16193] = 11
      "01011" when "011111101000010", -- t[16194] = 11
      "01011" when "011111101000011", -- t[16195] = 11
      "01011" when "011111101000100", -- t[16196] = 11
      "01011" when "011111101000101", -- t[16197] = 11
      "01011" when "011111101000110", -- t[16198] = 11
      "01011" when "011111101000111", -- t[16199] = 11
      "01011" when "011111101001000", -- t[16200] = 11
      "01011" when "011111101001001", -- t[16201] = 11
      "01011" when "011111101001010", -- t[16202] = 11
      "01011" when "011111101001011", -- t[16203] = 11
      "01011" when "011111101001100", -- t[16204] = 11
      "01011" when "011111101001101", -- t[16205] = 11
      "01011" when "011111101001110", -- t[16206] = 11
      "01011" when "011111101001111", -- t[16207] = 11
      "01011" when "011111101010000", -- t[16208] = 11
      "01011" when "011111101010001", -- t[16209] = 11
      "01011" when "011111101010010", -- t[16210] = 11
      "01011" when "011111101010011", -- t[16211] = 11
      "01011" when "011111101010100", -- t[16212] = 11
      "01011" when "011111101010101", -- t[16213] = 11
      "01011" when "011111101010110", -- t[16214] = 11
      "01011" when "011111101010111", -- t[16215] = 11
      "01011" when "011111101011000", -- t[16216] = 11
      "01011" when "011111101011001", -- t[16217] = 11
      "01011" when "011111101011010", -- t[16218] = 11
      "01011" when "011111101011011", -- t[16219] = 11
      "01011" when "011111101011100", -- t[16220] = 11
      "01011" when "011111101011101", -- t[16221] = 11
      "01011" when "011111101011110", -- t[16222] = 11
      "01011" when "011111101011111", -- t[16223] = 11
      "01011" when "011111101100000", -- t[16224] = 11
      "01011" when "011111101100001", -- t[16225] = 11
      "01011" when "011111101100010", -- t[16226] = 11
      "01011" when "011111101100011", -- t[16227] = 11
      "01011" when "011111101100100", -- t[16228] = 11
      "01011" when "011111101100101", -- t[16229] = 11
      "01011" when "011111101100110", -- t[16230] = 11
      "01011" when "011111101100111", -- t[16231] = 11
      "01011" when "011111101101000", -- t[16232] = 11
      "01011" when "011111101101001", -- t[16233] = 11
      "01011" when "011111101101010", -- t[16234] = 11
      "01011" when "011111101101011", -- t[16235] = 11
      "01011" when "011111101101100", -- t[16236] = 11
      "01011" when "011111101101101", -- t[16237] = 11
      "01011" when "011111101101110", -- t[16238] = 11
      "01011" when "011111101101111", -- t[16239] = 11
      "01011" when "011111101110000", -- t[16240] = 11
      "01011" when "011111101110001", -- t[16241] = 11
      "01011" when "011111101110010", -- t[16242] = 11
      "01011" when "011111101110011", -- t[16243] = 11
      "01011" when "011111101110100", -- t[16244] = 11
      "01011" when "011111101110101", -- t[16245] = 11
      "01011" when "011111101110110", -- t[16246] = 11
      "01011" when "011111101110111", -- t[16247] = 11
      "01011" when "011111101111000", -- t[16248] = 11
      "01011" when "011111101111001", -- t[16249] = 11
      "01011" when "011111101111010", -- t[16250] = 11
      "01011" when "011111101111011", -- t[16251] = 11
      "01011" when "011111101111100", -- t[16252] = 11
      "01011" when "011111101111101", -- t[16253] = 11
      "01011" when "011111101111110", -- t[16254] = 11
      "01011" when "011111101111111", -- t[16255] = 11
      "01011" when "011111110000000", -- t[16256] = 11
      "01011" when "011111110000001", -- t[16257] = 11
      "01011" when "011111110000010", -- t[16258] = 11
      "01011" when "011111110000011", -- t[16259] = 11
      "01011" when "011111110000100", -- t[16260] = 11
      "01011" when "011111110000101", -- t[16261] = 11
      "01011" when "011111110000110", -- t[16262] = 11
      "01011" when "011111110000111", -- t[16263] = 11
      "01011" when "011111110001000", -- t[16264] = 11
      "01011" when "011111110001001", -- t[16265] = 11
      "01011" when "011111110001010", -- t[16266] = 11
      "01011" when "011111110001011", -- t[16267] = 11
      "01011" when "011111110001100", -- t[16268] = 11
      "01011" when "011111110001101", -- t[16269] = 11
      "01011" when "011111110001110", -- t[16270] = 11
      "01011" when "011111110001111", -- t[16271] = 11
      "01011" when "011111110010000", -- t[16272] = 11
      "01011" when "011111110010001", -- t[16273] = 11
      "01011" when "011111110010010", -- t[16274] = 11
      "01011" when "011111110010011", -- t[16275] = 11
      "01011" when "011111110010100", -- t[16276] = 11
      "01011" when "011111110010101", -- t[16277] = 11
      "01011" when "011111110010110", -- t[16278] = 11
      "01011" when "011111110010111", -- t[16279] = 11
      "01011" when "011111110011000", -- t[16280] = 11
      "01011" when "011111110011001", -- t[16281] = 11
      "01011" when "011111110011010", -- t[16282] = 11
      "01011" when "011111110011011", -- t[16283] = 11
      "01011" when "011111110011100", -- t[16284] = 11
      "01011" when "011111110011101", -- t[16285] = 11
      "01011" when "011111110011110", -- t[16286] = 11
      "01011" when "011111110011111", -- t[16287] = 11
      "01011" when "011111110100000", -- t[16288] = 11
      "01011" when "011111110100001", -- t[16289] = 11
      "01011" when "011111110100010", -- t[16290] = 11
      "01011" when "011111110100011", -- t[16291] = 11
      "01011" when "011111110100100", -- t[16292] = 11
      "01011" when "011111110100101", -- t[16293] = 11
      "01011" when "011111110100110", -- t[16294] = 11
      "01011" when "011111110100111", -- t[16295] = 11
      "01011" when "011111110101000", -- t[16296] = 11
      "01011" when "011111110101001", -- t[16297] = 11
      "01011" when "011111110101010", -- t[16298] = 11
      "01011" when "011111110101011", -- t[16299] = 11
      "01011" when "011111110101100", -- t[16300] = 11
      "01011" when "011111110101101", -- t[16301] = 11
      "01011" when "011111110101110", -- t[16302] = 11
      "01011" when "011111110101111", -- t[16303] = 11
      "01011" when "011111110110000", -- t[16304] = 11
      "01011" when "011111110110001", -- t[16305] = 11
      "01011" when "011111110110010", -- t[16306] = 11
      "01011" when "011111110110011", -- t[16307] = 11
      "01011" when "011111110110100", -- t[16308] = 11
      "01011" when "011111110110101", -- t[16309] = 11
      "01011" when "011111110110110", -- t[16310] = 11
      "01011" when "011111110110111", -- t[16311] = 11
      "01011" when "011111110111000", -- t[16312] = 11
      "01011" when "011111110111001", -- t[16313] = 11
      "01011" when "011111110111010", -- t[16314] = 11
      "01011" when "011111110111011", -- t[16315] = 11
      "01011" when "011111110111100", -- t[16316] = 11
      "01011" when "011111110111101", -- t[16317] = 11
      "01011" when "011111110111110", -- t[16318] = 11
      "01011" when "011111110111111", -- t[16319] = 11
      "01011" when "011111111000000", -- t[16320] = 11
      "01011" when "011111111000001", -- t[16321] = 11
      "01011" when "011111111000010", -- t[16322] = 11
      "01011" when "011111111000011", -- t[16323] = 11
      "01011" when "011111111000100", -- t[16324] = 11
      "01011" when "011111111000101", -- t[16325] = 11
      "01011" when "011111111000110", -- t[16326] = 11
      "01011" when "011111111000111", -- t[16327] = 11
      "01011" when "011111111001000", -- t[16328] = 11
      "01011" when "011111111001001", -- t[16329] = 11
      "01011" when "011111111001010", -- t[16330] = 11
      "01011" when "011111111001011", -- t[16331] = 11
      "01011" when "011111111001100", -- t[16332] = 11
      "01011" when "011111111001101", -- t[16333] = 11
      "01011" when "011111111001110", -- t[16334] = 11
      "01011" when "011111111001111", -- t[16335] = 11
      "01011" when "011111111010000", -- t[16336] = 11
      "01011" when "011111111010001", -- t[16337] = 11
      "01011" when "011111111010010", -- t[16338] = 11
      "01011" when "011111111010011", -- t[16339] = 11
      "01011" when "011111111010100", -- t[16340] = 11
      "01011" when "011111111010101", -- t[16341] = 11
      "01011" when "011111111010110", -- t[16342] = 11
      "01011" when "011111111010111", -- t[16343] = 11
      "01011" when "011111111011000", -- t[16344] = 11
      "01011" when "011111111011001", -- t[16345] = 11
      "01011" when "011111111011010", -- t[16346] = 11
      "01011" when "011111111011011", -- t[16347] = 11
      "01011" when "011111111011100", -- t[16348] = 11
      "01011" when "011111111011101", -- t[16349] = 11
      "01011" when "011111111011110", -- t[16350] = 11
      "01011" when "011111111011111", -- t[16351] = 11
      "01011" when "011111111100000", -- t[16352] = 11
      "01011" when "011111111100001", -- t[16353] = 11
      "01011" when "011111111100010", -- t[16354] = 11
      "01011" when "011111111100011", -- t[16355] = 11
      "01011" when "011111111100100", -- t[16356] = 11
      "01011" when "011111111100101", -- t[16357] = 11
      "01011" when "011111111100110", -- t[16358] = 11
      "01011" when "011111111100111", -- t[16359] = 11
      "01011" when "011111111101000", -- t[16360] = 11
      "01011" when "011111111101001", -- t[16361] = 11
      "01011" when "011111111101010", -- t[16362] = 11
      "01011" when "011111111101011", -- t[16363] = 11
      "01011" when "011111111101100", -- t[16364] = 11
      "01011" when "011111111101101", -- t[16365] = 11
      "01011" when "011111111101110", -- t[16366] = 11
      "01011" when "011111111101111", -- t[16367] = 11
      "01100" when "011111111110000", -- t[16368] = 12
      "01100" when "011111111110001", -- t[16369] = 12
      "01100" when "011111111110010", -- t[16370] = 12
      "01100" when "011111111110011", -- t[16371] = 12
      "01100" when "011111111110100", -- t[16372] = 12
      "01100" when "011111111110101", -- t[16373] = 12
      "01100" when "011111111110110", -- t[16374] = 12
      "01100" when "011111111110111", -- t[16375] = 12
      "01100" when "011111111111000", -- t[16376] = 12
      "01100" when "011111111111001", -- t[16377] = 12
      "01100" when "011111111111010", -- t[16378] = 12
      "01100" when "011111111111011", -- t[16379] = 12
      "01100" when "011111111111100", -- t[16380] = 12
      "01100" when "011111111111101", -- t[16381] = 12
      "01100" when "011111111111110", -- t[16382] = 12
      "01100" when "011111111111111", -- t[16383] = 12
      "-----" when others;
end architecture;


-- Minimax-Defour: LNS subtraction function [ -8.000000, -4.000000 [ -> [ 0.000000, 0.125000 [
-- Input:  wE =   2, wF =  11, w =  13
-- Output: wE =  -3, wF =  11, w =   8
-- Decomposition: a  =  5, b  =  8
--                a0 =  5, b0 =  6, p0 =  5
--                a1 =  3, b1 =  2, p1 = 11
--                a2 =  3, b2 =  2, p2 =  5
--                g0 =  4, g1 =  -2
-- ROMs: 2^ 5 x 12  +  2^ 5 x  6  +  2^ 5 x  1  +  2^ 5 x  1  =     640 bits
-- Mult: 6 x 6 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T1_11 is
  component LNSSub_MNMX_T1_11_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_t2 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_t3 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T1_11_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_11_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_t0 is
begin
  with x select
    r <=
      "000011000010" when "00000", -- t[0] = 194
      "000011010011" when "00001", -- t[1] = 211
      "000011100101" when "00010", -- t[2] = 229
      "000011110111" when "00011", -- t[3] = 247
      "000100001110" when "00100", -- t[4] = 270
      "000100100111" when "00101", -- t[5] = 295
      "000100111110" when "00110", -- t[6] = 318
      "000101011011" when "00111", -- t[7] = 347
      "000101111100" when "01000", -- t[8] = 380
      "000110011011" when "01001", -- t[9] = 411
      "000111000010" when "01010", -- t[10] = 450
      "000111101011" when "01011", -- t[11] = 491
      "001000010101" when "01100", -- t[12] = 533
      "001001000100" when "01101", -- t[13] = 580
      "001001111010" when "01110", -- t[14] = 634
      "001010110010" when "01111", -- t[15] = 690
      "001011110010" when "10000", -- t[16] = 754
      "001100110110" when "10001", -- t[17] = 822
      "001110000000" when "10010", -- t[18] = 896
      "001111010000" when "10011", -- t[19] = 976
      "010000101001" when "10100", -- t[20] = 1065
      "010010001010" when "10101", -- t[21] = 1162
      "010011110101" when "10110", -- t[22] = 1269
      "010101100110" when "10111", -- t[23] = 1382
      "010111100110" when "11000", -- t[24] = 1510
      "011001101110" when "11001", -- t[25] = 1646
      "011100000101" when "11010", -- t[26] = 1797
      "011110101010" when "11011", -- t[27] = 1962
      "100001011111" when "11100", -- t[28] = 2143
      "100100100111" when "11101", -- t[29] = 2343
      "100111111111" when "11110", -- t[30] = 2559
      "101011101100" when "11111", -- t[31] = 2796
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_11_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_t1 is
begin
  with x select
    r <=
      "000010" when "00000", -- t[0] = 2
      "000010" when "00001", -- t[1] = 2
      "000010" when "00010", -- t[2] = 2
      "000011" when "00011", -- t[3] = 3
      "000011" when "00100", -- t[4] = 3
      "000011" when "00101", -- t[5] = 3
      "000100" when "00110", -- t[6] = 4
      "000100" when "00111", -- t[7] = 4
      "000100" when "01000", -- t[8] = 4
      "000101" when "01001", -- t[9] = 5
      "000101" when "01010", -- t[10] = 5
      "000101" when "01011", -- t[11] = 5
      "000110" when "01100", -- t[12] = 6
      "000111" when "01101", -- t[13] = 7
      "000111" when "01110", -- t[14] = 7
      "001000" when "01111", -- t[15] = 8
      "001000" when "10000", -- t[16] = 8
      "001001" when "10001", -- t[17] = 9
      "001010" when "10010", -- t[18] = 10
      "001011" when "10011", -- t[19] = 11
      "001100" when "10100", -- t[20] = 12
      "001101" when "10101", -- t[21] = 13
      "001110" when "10110", -- t[22] = 14
      "010000" when "10111", -- t[23] = 16
      "010001" when "11000", -- t[24] = 17
      "010011" when "11001", -- t[25] = 19
      "010101" when "11010", -- t[26] = 21
      "010111" when "11011", -- t[27] = 23
      "011001" when "11100", -- t[28] = 25
      "011011" when "11101", -- t[29] = 27
      "011110" when "11110", -- t[30] = 30
      "100001" when "11111", -- t[31] = 33
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_11_t2 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_t2 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "0" when "1101", -- t[13] = 0
      "0" when "1110", -- t[14] = 0
      "1" when "1111", -- t[15] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_11_t3 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_t3 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "1" when "1101", -- t[13] = 1
      "0" when "1110", -- t[14] = 0
      "1" when "1111", -- t[15] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_11.all;

entity LNSSub_MNMX_T1_11_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_mult is
  signal out_t : std_logic_vector(5 downto 0);
  signal r0    : std_logic_vector(11 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T1_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(11 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_11.all;

entity LNSSub_MNMX_T1_11_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T1_11_t2
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_11.all;

entity LNSSub_MNMX_T1_11_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T1_11_t3
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_11.all;

entity LNSSub_MNMX_T1_11 is
  port ( x : in  std_logic_vector(12 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_11 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(11 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(5 downto 0);
  signal r1  : std_logic_vector(11 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(11 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(11 downto 0);
  signal sum : std_logic_vector(11 downto 0);
begin
  a0 <= x(12 downto 8);
  inst_t0 : LNSSub_MNMX_T1_11_t0
    port map ( x => a0,
               r => r0(11 downto 0) );

  a1 <= x(12 downto 8);
  b1 <= x(7 downto 2);
  inst_mult : LNSSub_MNMX_T1_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(8 downto 0) );
  r1(11 downto 9) <= (11 downto 9 => '0');

  a2 <= x(12 downto 10);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T1_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(11 downto 0) );

  a3 <= x(12 downto 10);
  b3 <= x(7 downto 6);
  inst_xor3 : LNSSub_MNMX_T1_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(11 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(11 downto 4);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -4.000000, -2.000000 [ -> [ 0.000000, 0.500000 [
-- Input:  wE =   1, wF =  11, w =  12
-- Output: wE =  -1, wF =  11, w =  10
-- Decomposition: a  =  5, b  =  7
--                a0 =  5, b0 =  5, p0 =  5
--                a1 =  3, b1 =  2, p1 = 10
--                a2 =  3, b2 =  2, p2 =  5
--                g0 =  4, g1 =  -3
-- ROMs: 2^ 5 x 14  +  2^ 5 x  7  +  2^ 5 x  3  +  2^ 5 x  2  =     832 bits
-- Mult: 5 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T2_11 is
  component LNSSub_MNMX_T2_11_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_t2 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_t3 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MNMX_T2_11_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_11_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_t0 is
begin
  with x select
    r <=
      "00101111110111" when "00000", -- t[0] = 3063
      "00110010000001" when "00001", -- t[1] = 3201
      "00110100010100" when "00010", -- t[2] = 3348
      "00110110101100" when "00011", -- t[3] = 3500
      "00111001001101" when "00100", -- t[4] = 3661
      "00111011110101" when "00101", -- t[5] = 3829
      "00111110100110" when "00110", -- t[6] = 4006
      "01000001100000" when "00111", -- t[7] = 4192
      "01000100100010" when "01000", -- t[8] = 4386
      "01000111101011" when "01001", -- t[9] = 4587
      "01001011000001" when "01010", -- t[10] = 4801
      "01001110100011" when "01011", -- t[11] = 5027
      "01010010001100" when "01100", -- t[12] = 5260
      "01010110000101" when "01101", -- t[13] = 5509
      "01011010000110" when "01110", -- t[14] = 5766
      "01011110010100" when "01111", -- t[15] = 6036
      "01100010110101" when "10000", -- t[16] = 6325
      "01100111100001" when "10001", -- t[17] = 6625
      "01101100011101" when "10010", -- t[18] = 6941
      "01110001100100" when "10011", -- t[19] = 7268
      "01110111000010" when "10100", -- t[20] = 7618
      "01111100110010" when "10101", -- t[21] = 7986
      "10000010110011" when "10110", -- t[22] = 8371
      "10001001001001" when "10111", -- t[23] = 8777
      "10001111111001" when "11000", -- t[24] = 9209
      "10010110111001" when "11001", -- t[25] = 9657
      "10011110010111" when "11010", -- t[26] = 10135
      "10100110001111" when "11011", -- t[27] = 10639
      "10101110100000" when "11100", -- t[28] = 11168
      "10110111010001" when "11101", -- t[29] = 11729
      "11000000100100" when "11110", -- t[30] = 12324
      "11001010010101" when "11111", -- t[31] = 12949
      "--------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_11_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_t1 is
begin
  with x select
    r <=
      "0010001" when "00000", -- t[0] = 17
      "0010010" when "00001", -- t[1] = 18
      "0010011" when "00010", -- t[2] = 19
      "0010100" when "00011", -- t[3] = 20
      "0010101" when "00100", -- t[4] = 21
      "0010110" when "00101", -- t[5] = 22
      "0010111" when "00110", -- t[6] = 23
      "0011000" when "00111", -- t[7] = 24
      "0011001" when "01000", -- t[8] = 25
      "0011011" when "01001", -- t[9] = 27
      "0011100" when "01010", -- t[10] = 28
      "0011101" when "01011", -- t[11] = 29
      "0011111" when "01100", -- t[12] = 31
      "0100000" when "01101", -- t[13] = 32
      "0100010" when "01110", -- t[14] = 34
      "0100100" when "01111", -- t[15] = 36
      "0100101" when "10000", -- t[16] = 37
      "0100111" when "10001", -- t[17] = 39
      "0101001" when "10010", -- t[18] = 41
      "0101100" when "10011", -- t[19] = 44
      "0101110" when "10100", -- t[20] = 46
      "0110000" when "10101", -- t[21] = 48
      "0110011" when "10110", -- t[22] = 51
      "0110110" when "10111", -- t[23] = 54
      "0111000" when "11000", -- t[24] = 56
      "0111100" when "11001", -- t[25] = 60
      "0111111" when "11010", -- t[26] = 63
      "1000010" when "11011", -- t[27] = 66
      "1000110" when "11100", -- t[28] = 70
      "1001010" when "11101", -- t[29] = 74
      "1001110" when "11110", -- t[30] = 78
      "1010011" when "11111", -- t[31] = 83
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_11_t2 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_t2 is
begin
  with x select
    r <=
      "000" when "0000", -- t[0] = 0
      "001" when "0001", -- t[1] = 1
      "000" when "0010", -- t[2] = 0
      "010" when "0011", -- t[3] = 2
      "000" when "0100", -- t[4] = 0
      "010" when "0101", -- t[5] = 2
      "001" when "0110", -- t[6] = 1
      "011" when "0111", -- t[7] = 3
      "001" when "1000", -- t[8] = 1
      "011" when "1001", -- t[9] = 3
      "001" when "1010", -- t[10] = 1
      "100" when "1011", -- t[11] = 4
      "001" when "1100", -- t[12] = 1
      "101" when "1101", -- t[13] = 5
      "010" when "1110", -- t[14] = 2
      "111" when "1111", -- t[15] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_11_t3 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_t3 is
begin
  with x select
    r <=
      "00" when "0000", -- t[0] = 0
      "00" when "0001", -- t[1] = 0
      "00" when "0010", -- t[2] = 0
      "00" when "0011", -- t[3] = 0
      "00" when "0100", -- t[4] = 0
      "00" when "0101", -- t[5] = 0
      "00" when "0110", -- t[6] = 0
      "00" when "0111", -- t[7] = 0
      "00" when "1000", -- t[8] = 0
      "01" when "1001", -- t[9] = 1
      "00" when "1010", -- t[10] = 0
      "01" when "1011", -- t[11] = 1
      "00" when "1100", -- t[12] = 0
      "01" when "1101", -- t[13] = 1
      "00" when "1110", -- t[14] = 0
      "10" when "1111", -- t[15] = 2
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_11.all;

entity LNSSub_MNMX_T2_11_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(11 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T2_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(11 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_11.all;

entity LNSSub_MNMX_T2_11_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T2_11_t2
    port map ( x => in_t,
               r => out_t );

  r(13 downto 3) <= (13 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_11.all;

entity LNSSub_MNMX_T2_11_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T2_11_t3
    port map ( x => in_t,
               r => out_t );

  r(13 downto 2) <= (13 downto 2 => '0');
  r(0) <= out_t(0);
  r(1) <= out_t(1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_11.all;

entity LNSSub_MNMX_T2_11 is
  port ( x : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_11 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(13 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(4 downto 0);
  signal r1  : std_logic_vector(13 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(13 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(13 downto 0);
  signal sum : std_logic_vector(13 downto 0);
begin
  a0 <= x(11 downto 7);
  inst_t0 : LNSSub_MNMX_T2_11_t0
    port map ( x => a0,
               r => r0(13 downto 0) );

  a1 <= x(11 downto 7);
  b1 <= x(6 downto 2);
  inst_mult : LNSSub_MNMX_T2_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(9 downto 0) );
  r1(13 downto 10) <= (13 downto 10 => '0');

  a2 <= x(11 downto 9);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T2_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(13 downto 0) );

  a3 <= x(11 downto 9);
  b3 <= x(6 downto 5);
  inst_xor3 : LNSSub_MNMX_T2_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(13 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(13 downto 4);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -2.000000, -1.000000 [ -> [ 0.000000, 1.000000 [
-- Input:  wE =   0, wF =  11, w =  11
-- Output: wE =   0, wF =  11, w =  11
-- Decomposition: a  =  5, b  =  6
--                a0 =  5, b0 =  4, p0 =  5
--                a1 =  3, b1 =  2, p1 =  9
--                a2 =  3, b2 =  2, p2 =  5
--                g0 =  3, g1 =  -4
-- ROMs: 2^ 5 x 14  +  2^ 5 x  7  +  2^ 5 x  4  +  2^ 5 x  1  =     832 bits
-- Mult: 4 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T3_11 is
  component LNSSub_MNMX_T3_11_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_t2 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_t3 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;

  component LNSSub_MNMX_T3_11_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(13 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_11_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_t0 is
begin
  with x select
    r <=
      "01101010011000" when "00000", -- t[0] = 6808
      "01101101000100" when "00001", -- t[1] = 6980
      "01101111110111" when "00010", -- t[2] = 7159
      "01110010110000" when "00011", -- t[3] = 7344
      "01110101101100" when "00100", -- t[4] = 7532
      "01111000110000" when "00101", -- t[5] = 7728
      "01111011110111" when "00110", -- t[6] = 7927
      "01111111001000" when "00111", -- t[7] = 8136
      "10000010011101" when "01000", -- t[8] = 8349
      "10000101111001" when "01001", -- t[9] = 8569
      "10001001011100" when "01010", -- t[10] = 8796
      "10001101000111" when "01011", -- t[11] = 9031
      "10010000111001" when "01100", -- t[12] = 9273
      "10010100110011" when "01101", -- t[13] = 9523
      "10011000110011" when "01110", -- t[14] = 9779
      "10011100111110" when "01111", -- t[15] = 10046
      "10100001010011" when "10000", -- t[16] = 10323
      "10100101101111" when "10001", -- t[17] = 10607
      "10101010010110" when "10010", -- t[18] = 10902
      "10101111000111" when "10011", -- t[19] = 11207
      "10110100000011" when "10100", -- t[20] = 11523
      "10111001001010" when "10101", -- t[21] = 11850
      "10111110011101" when "10110", -- t[22] = 12189
      "11000011111110" when "10111", -- t[23] = 12542
      "11001001101001" when "11000", -- t[24] = 12905
      "11001111100101" when "11001", -- t[25] = 13285
      "11010101101110" when "11010", -- t[26] = 13678
      "11011100000111" when "11011", -- t[27] = 14087
      "11100010110000" when "11100", -- t[28] = 14512
      "11101001101011" when "11101", -- t[29] = 14955
      "11110000111000" when "11110", -- t[30] = 15416
      "11111000011001" when "11111", -- t[31] = 15897
      "--------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_11_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_t1 is
begin
  with x select
    r <=
      "0101011" when "00000", -- t[0] = 43
      "0101101" when "00001", -- t[1] = 45
      "0101110" when "00010", -- t[2] = 46
      "0101111" when "00011", -- t[3] = 47
      "0110001" when "00100", -- t[4] = 49
      "0110010" when "00101", -- t[5] = 50
      "0110100" when "00110", -- t[6] = 52
      "0110101" when "00111", -- t[7] = 53
      "0110111" when "01000", -- t[8] = 55
      "0111001" when "01001", -- t[9] = 57
      "0111011" when "01010", -- t[10] = 59
      "0111100" when "01011", -- t[11] = 60
      "0111110" when "01100", -- t[12] = 62
      "1000000" when "01101", -- t[13] = 64
      "1000011" when "01110", -- t[14] = 67
      "1000101" when "01111", -- t[15] = 69
      "1000111" when "10000", -- t[16] = 71
      "1001010" when "10001", -- t[17] = 74
      "1001100" when "10010", -- t[18] = 76
      "1001111" when "10011", -- t[19] = 79
      "1010010" when "10100", -- t[20] = 82
      "1010101" when "10101", -- t[21] = 85
      "1011000" when "10110", -- t[22] = 88
      "1011011" when "10111", -- t[23] = 91
      "1011111" when "11000", -- t[24] = 95
      "1100010" when "11001", -- t[25] = 98
      "1100110" when "11010", -- t[26] = 102
      "1101010" when "11011", -- t[27] = 106
      "1101111" when "11100", -- t[28] = 111
      "1110011" when "11101", -- t[29] = 115
      "1111000" when "11110", -- t[30] = 120
      "1111101" when "11111", -- t[31] = 125
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_11_t2 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_t2 is
begin
  with x select
    r <=
      "0001" when "0000", -- t[0] = 1
      "0100" when "0001", -- t[1] = 4
      "0001" when "0010", -- t[2] = 1
      "0100" when "0011", -- t[3] = 4
      "0001" when "0100", -- t[4] = 1
      "0101" when "0101", -- t[5] = 5
      "0010" when "0110", -- t[6] = 2
      "0110" when "0111", -- t[7] = 6
      "0010" when "1000", -- t[8] = 2
      "0111" when "1001", -- t[9] = 7
      "0010" when "1010", -- t[10] = 2
      "1000" when "1011", -- t[11] = 8
      "0011" when "1100", -- t[12] = 3
      "1001" when "1101", -- t[13] = 9
      "0011" when "1110", -- t[14] = 3
      "1011" when "1111", -- t[15] = 11
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_11_t3 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_t3 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "1" when "1101", -- t[13] = 1
      "0" when "1110", -- t[14] = 0
      "1" when "1111", -- t[15] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_11.all;

entity LNSSub_MNMX_T3_11_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(10 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T3_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(10 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_11.all;

entity LNSSub_MNMX_T3_11_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T3_11_t2
    port map ( x => in_t,
               r => out_t );

  r(13 downto 4) <= (13 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_11.all;

entity LNSSub_MNMX_T3_11_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T3_11_t3
    port map ( x => in_t,
               r => out_t );

  r(13 downto 1) <= (13 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_11.all;

entity LNSSub_MNMX_T3_11 is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_11 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(13 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(13 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(13 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(13 downto 0);
  signal sum : std_logic_vector(13 downto 0);
begin
  a0 <= x(10 downto 6);
  inst_t0 : LNSSub_MNMX_T3_11_t0
    port map ( x => a0,
               r => r0(13 downto 0) );

  a1 <= x(10 downto 6);
  b1 <= x(5 downto 2);
  inst_mult : LNSSub_MNMX_T3_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(8 downto 0) );
  r1(13 downto 9) <= (13 downto 9 => '0');

  a2 <= x(10 downto 8);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T3_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(13 downto 0) );

  a3 <= x(10 downto 8);
  b3 <= x(5 downto 4);
  inst_xor3 : LNSSub_MNMX_T3_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(13 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(13 downto 3);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -1.000000, -0.500000 [ -> [ 0.000000, 2.000000 [
-- Input:  wE =  -1, wF =  11, w =  10
-- Output: wE =   1, wF =  11, w =  12
-- Decomposition: a  =  4, b  =  6
--                a0 =  4, b0 =  4, p0 =  4
--                a1 =  2, b1 =  2, p1 =  8
--                a2 =  2, b2 =  2, p2 =  4
--                g0 =  0, g1 =  -4
-- ROMs: 2^ 4 x 12  +  2^ 4 x  9  +  2^ 4 x  2  +  2^ 4 x  0  =     368 bits
-- Mult: 4 x 9 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T4_11 is
  component LNSSub_MNMX_T4_11_t0 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_t1 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_t2 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_t3 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_mult is
    port ( a : in  std_logic_vector(3 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T4_11_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_11_t0 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_t0 is
begin
  with x select
    r <=
      "100000000010" when "0000", -- t[0] = 2050
      "100001000100" when "0001", -- t[1] = 2116
      "100010001000" when "0010", -- t[2] = 2184
      "100011010000" when "0011", -- t[3] = 2256
      "100100011011" when "0100", -- t[4] = 2331
      "100101101001" when "0101", -- t[5] = 2409
      "100110111100" when "0110", -- t[6] = 2492
      "101000010011" when "0111", -- t[7] = 2579
      "101001101110" when "1000", -- t[8] = 2670
      "101011001111" when "1001", -- t[9] = 2767
      "101100110101" when "1010", -- t[10] = 2869
      "101110100001" when "1011", -- t[11] = 2977
      "110000010100" when "1100", -- t[12] = 3092
      "110010001110" when "1101", -- t[13] = 3214
      "110100010000" when "1110", -- t[14] = 3344
      "110110011011" when "1111", -- t[15] = 3483
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_11_t1 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_t1 is
begin
  with x select
    r <=
      "010000011" when "0000", -- t[0] = 131
      "010001001" when "0001", -- t[1] = 137
      "010001111" when "0010", -- t[2] = 143
      "010010110" when "0011", -- t[3] = 150
      "010011101" when "0100", -- t[4] = 157
      "010100101" when "0101", -- t[5] = 165
      "010101110" when "0110", -- t[6] = 174
      "010110111" when "0111", -- t[7] = 183
      "011000001" when "1000", -- t[8] = 193
      "011001100" when "1001", -- t[9] = 204
      "011011000" when "1010", -- t[10] = 216
      "011100101" when "1011", -- t[11] = 229
      "011110011" when "1100", -- t[12] = 243
      "100000100" when "1101", -- t[13] = 260
      "100010110" when "1110", -- t[14] = 278
      "100101010" when "1111", -- t[15] = 298
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_11_t2 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_t2 is
begin
  with x select
    r <=
      "00" when "000", -- t[0] = 0
      "01" when "001", -- t[1] = 1
      "00" when "010", -- t[2] = 0
      "01" when "011", -- t[3] = 1
      "00" when "100", -- t[4] = 0
      "10" when "101", -- t[5] = 2
      "01" when "110", -- t[6] = 1
      "11" when "111", -- t[7] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_11_t3 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_t3 is
begin
  with x select
    r <=
      "0" when "000", -- t[0] = 0
      "0" when "001", -- t[1] = 0
      "0" when "010", -- t[2] = 0
      "0" when "011", -- t[3] = 0
      "0" when "100", -- t[4] = 0
      "0" when "101", -- t[5] = 0
      "0" when "110", -- t[6] = 0
      "0" when "111", -- t[7] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_11.all;

entity LNSSub_MNMX_T4_11_mult is
  port ( a : in  std_logic_vector(3 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_mult is
  signal out_t : std_logic_vector(8 downto 0);
  signal r0    : std_logic_vector(12 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T4_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(12 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_11.all;

entity LNSSub_MNMX_T4_11_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T4_11_t2
    port map ( x => in_t,
               r => out_t );

  r(11 downto 2) <= (11 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_11.all;

entity LNSSub_MNMX_T4_11_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T4_11_t3
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_11.all;

entity LNSSub_MNMX_T4_11 is
  port ( x : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_11 is
  signal a0  : std_logic_vector(3 downto 0);
  signal r0  : std_logic_vector(11 downto 0);
  signal a1  : std_logic_vector(3 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(11 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(11 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(11 downto 0);
  signal sum : std_logic_vector(11 downto 0);
begin
  a0 <= x(9 downto 6);
  inst_t0 : LNSSub_MNMX_T4_11_t0
    port map ( x => a0,
               r => r0(11 downto 0) );

  a1 <= x(9 downto 6);
  b1 <= x(5 downto 2);
  inst_mult : LNSSub_MNMX_T4_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(11 downto 8) <= (11 downto 8 => '0');

  a2 <= x(9 downto 8);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T4_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(11 downto 0) );

  a3 <= x(9 downto 8);
  b3 <= x(5 downto 4);
  inst_xor3 : LNSSub_MNMX_T4_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(11 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(11 downto 0);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.500000, -0.250000 [ -> [ 0.000000, 4.000000 [
-- Input:  wE =  -2, wF =  11, w =   9
-- Output: wE =   2, wF =   9, w =  11
-- Decomposition: a  =  3, b  =  6
--                a0 =  3, b0 =  4, p0 =  3
--                a1 =  2, b1 =  2, p1 =  7
--                a2 =  2, b2 =  2, p2 =  3
--                g0 =  2, g1 =  -5
-- ROMs: 2^ 3 x 13  +  2^ 3 x  7  +  2^ 4 x  3  +  2^ 4 x  2  =     240 bits
-- Mult: 4 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T5_11 is
  component LNSSub_MNMX_T5_11_t0 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_t1 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_t2 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_t3 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_mult is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MNMX_T5_11_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_11_t0 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_t0 is
begin
  with x select
    r <=
      "0111000110001" when "000", -- t[0] = 3633
      "0111011010011" when "001", -- t[1] = 3795
      "0111101111111" when "010", -- t[2] = 3967
      "1000000111101" when "011", -- t[3] = 4157
      "1000100001010" when "100", -- t[4] = 4362
      "1000111101100" when "101", -- t[5] = 4588
      "1001011101000" when "110", -- t[6] = 4840
      "1010000000000" when "111", -- t[7] = 5120
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_11_t1 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_t1 is
begin
  with x select
    r <=
      "0101000" when "000", -- t[0] = 40
      "0101011" when "001", -- t[1] = 43
      "0101111" when "010", -- t[2] = 47
      "0110011" when "011", -- t[3] = 51
      "0111001" when "100", -- t[4] = 57
      "0111111" when "101", -- t[5] = 63
      "1000110" when "110", -- t[6] = 70
      "1001111" when "111", -- t[7] = 79
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_11_t2 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_t2 is
begin
  with x select
    r <=
      "001" when "000", -- t[0] = 1
      "011" when "001", -- t[1] = 3
      "001" when "010", -- t[2] = 1
      "100" when "011", -- t[3] = 4
      "001" when "100", -- t[4] = 1
      "101" when "101", -- t[5] = 5
      "010" when "110", -- t[6] = 2
      "110" when "111", -- t[7] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_11_t3 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_t3 is
begin
  with x select
    r <=
      "00" when "000", -- t[0] = 0
      "00" when "001", -- t[1] = 0
      "00" when "010", -- t[2] = 0
      "01" when "011", -- t[3] = 1
      "00" when "100", -- t[4] = 0
      "01" when "101", -- t[5] = 1
      "00" when "110", -- t[6] = 0
      "10" when "111", -- t[7] = 2
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_11.all;

entity LNSSub_MNMX_T5_11_mult is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(10 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T5_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(10 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_11.all;

entity LNSSub_MNMX_T5_11_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T5_11_t2
    port map ( x => in_t,
               r => out_t );

  r(12 downto 3) <= (12 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_11.all;

entity LNSSub_MNMX_T5_11_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T5_11_t3
    port map ( x => in_t,
               r => out_t );

  r(12 downto 2) <= (12 downto 2 => '0');
  r(0) <= out_t(0);
  r(1) <= out_t(1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_11.all;

entity LNSSub_MNMX_T5_11 is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_11 is
  signal a0  : std_logic_vector(2 downto 0);
  signal r0  : std_logic_vector(12 downto 0);
  signal a1  : std_logic_vector(2 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(12 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(12 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(12 downto 0);
  signal sum : std_logic_vector(12 downto 0);
begin
  a0 <= x(8 downto 6);
  inst_t0 : LNSSub_MNMX_T5_11_t0
    port map ( x => a0,
               r => r0(12 downto 0) );

  a1 <= x(8 downto 6);
  b1 <= x(5 downto 2);
  inst_mult : LNSSub_MNMX_T5_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(8 downto 0) );
  r1(12 downto 9) <= (12 downto 9 => '0');

  a2 <= x(8 downto 7);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T5_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(12 downto 0) );

  a3 <= x(8 downto 7);
  b3 <= x(5 downto 4);
  inst_xor3 : LNSSub_MNMX_T5_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(12 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(12 downto 2);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.250000, -0.125000 [ -> [ 0.000000, 4.000000 [
-- Input:  wE =  -3, wF =  11, w =   8
-- Output: wE =   2, wF =   8, w =  10
-- Decomposition: a  =  3, b  =  5
--                a0 =  3, b0 =  4, p0 =  3
--                a1 =  2, b1 =  1, p1 =  7
--                a2 =  2, b2 =  1, p2 =  3
--                g0 =  2, g1 =  -7
-- ROMs: 2^ 3 x 12  +  2^ 3 x  5  +  2^ 3 x  2  +  2^ 3 x  0  =     152 bits
-- Mult: 4 x 5 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T6_11 is
  component LNSSub_MNMX_T6_11_t0 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_t1 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_t2 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_t3 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_mult is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T6_11_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_11_t0 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_t0 is
begin
  with x select
    r <=
      "101010011111" when "000", -- t[0] = 2719
      "101011110110" when "001", -- t[1] = 2806
      "101101010100" when "010", -- t[2] = 2900
      "101110111001" when "011", -- t[3] = 3001
      "110000101001" when "100", -- t[4] = 3113
      "110010011111" when "101", -- t[5] = 3231
      "110100101000" when "110", -- t[6] = 3368
      "110110111010" when "111", -- t[7] = 3514
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_11_t1 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_t1 is
begin
  with x select
    r <=
      "01011" when "000", -- t[0] = 11
      "01100" when "001", -- t[1] = 12
      "01101" when "010", -- t[2] = 13
      "01110" when "011", -- t[3] = 14
      "01111" when "100", -- t[4] = 15
      "10001" when "101", -- t[5] = 17
      "10010" when "110", -- t[6] = 18
      "10101" when "111", -- t[7] = 21
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_11_t2 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_t2 is
begin
  with x select
    r <=
      "01" when "00", -- t[0] = 1
      "01" when "01", -- t[1] = 1
      "01" when "10", -- t[2] = 1
      "10" when "11", -- t[3] = 2
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_11_t3 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_t3 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "0" when "01", -- t[1] = 0
      "0" when "10", -- t[2] = 0
      "0" when "11", -- t[3] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_11.all;

entity LNSSub_MNMX_T6_11_mult is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_mult is
  signal out_t : std_logic_vector(4 downto 0);
  signal r0    : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T6_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(8 downto 1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_11.all;

entity LNSSub_MNMX_T6_11_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T6_11_t2
    port map ( x => in_t,
               r => out_t );

  r(11 downto 2) <= (11 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_11.all;

entity LNSSub_MNMX_T6_11_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T6_11_t3
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_11.all;

entity LNSSub_MNMX_T6_11 is
  port ( x : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_11 is
  signal a0  : std_logic_vector(2 downto 0);
  signal r0  : std_logic_vector(11 downto 0);
  signal a1  : std_logic_vector(2 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(11 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(11 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(11 downto 0);
  signal sum : std_logic_vector(11 downto 0);
begin
  a0 <= x(7 downto 5);
  inst_t0 : LNSSub_MNMX_T6_11_t0
    port map ( x => a0,
               r => r0(11 downto 0) );

  a1 <= x(7 downto 5);
  b1 <= x(4 downto 1);
  inst_mult : LNSSub_MNMX_T6_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(11 downto 8) <= (11 downto 8 => '0');

  a2 <= x(7 downto 6);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T6_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(11 downto 0) );

  a3 <= x(7 downto 6);
  b3 <= x(4 downto 4);
  inst_xor3 : LNSSub_MNMX_T6_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(11 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(11 downto 2);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.125000, -0.062500 [ -> [ 0.000000, 8.000000 [
-- Input:  wE =  -4, wF =  11, w =   7
-- Output: wE =   3, wF =   7, w =  10
-- Decomposition: a  =  2, b  =  5
--                a0 =  2, b0 =  2, p0 =  2
--                a1 =  1, b1 =  3, p1 =  4
--                a2 =  1, b2 =  1, p2 =  2
--                g0 =  2, g1 =  -5
-- ROMs: 2^ 2 x 12  +  2^ 2 x  7  +  2^ 4 x  4  +  2^ 2 x  0  =     140 bits
-- Mult: 2 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T7_11 is
  component LNSSub_MNMX_T7_11_t0 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_t1 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_t2 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_t3 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_mult is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_xor2 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T7_11_xor3 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_11_t0 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_t0 is
begin
  with x select
    r <=
      "011100111010" when "00", -- t[0] = 1850
      "011110011010" when "01", -- t[1] = 1946
      "100000001001" when "10", -- t[2] = 2057
      "100010001111" when "11", -- t[3] = 2191
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_11_t1 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_t1 is
begin
  with x select
    r <=
      "0101111" when "00", -- t[0] = 47
      "0110111" when "01", -- t[1] = 55
      "1000001" when "10", -- t[2] = 65
      "1010000" when "11", -- t[3] = 80
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_11_t2 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_t2 is
begin
  with x select
    r <=
      "0001" when "000", -- t[0] = 1
      "0100" when "001", -- t[1] = 4
      "0111" when "010", -- t[2] = 7
      "1011" when "011", -- t[3] = 11
      "0010" when "100", -- t[4] = 2
      "0110" when "101", -- t[5] = 6
      "1011" when "110", -- t[6] = 11
      "1111" when "111", -- t[7] = 15
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_11_t3 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_t3 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_11.all;

entity LNSSub_MNMX_T7_11_mult is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T7_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(8 downto 1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_11.all;

entity LNSSub_MNMX_T7_11_xor2 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(2);
  in_t(2 downto 2) <= a;
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_t2 : LNSSub_MNMX_T7_11_t2
    port map ( x => in_t,
               r => out_t );

  r(11 downto 4) <= (11 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_11.all;

entity LNSSub_MNMX_T7_11_xor3 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T7_11_t3
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_11.all;

entity LNSSub_MNMX_T7_11 is
  port ( x : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_11 is
  signal a0  : std_logic_vector(1 downto 0);
  signal r0  : std_logic_vector(11 downto 0);
  signal a1  : std_logic_vector(1 downto 0);
  signal b1  : std_logic_vector(1 downto 0);
  signal r1  : std_logic_vector(11 downto 0);
  signal a2  : std_logic_vector(0 downto 0);
  signal b2  : std_logic_vector(2 downto 0);
  signal r2  : std_logic_vector(11 downto 0);
  signal a3  : std_logic_vector(0 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(11 downto 0);
  signal sum : std_logic_vector(11 downto 0);
begin
  a0 <= x(6 downto 5);
  inst_t0 : LNSSub_MNMX_T7_11_t0
    port map ( x => a0,
               r => r0(11 downto 0) );

  a1 <= x(6 downto 5);
  b1 <= x(4 downto 3);
  inst_mult : LNSSub_MNMX_T7_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(11 downto 8) <= (11 downto 8 => '0');

  a2 <= x(6 downto 6);
  b2 <= x(2 downto 0);
  inst_xor2 : LNSSub_MNMX_T7_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(11 downto 0) );

  a3 <= x(6 downto 6);
  b3 <= x(4 downto 4);
  inst_xor3 : LNSSub_MNMX_T7_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(11 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(11 downto 2);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.062500, -0.031250 [ -> [ 0.000000, 8.000000 [
-- Input:  wE =  -5, wF =  11, w =   6
-- Output: wE =   3, wF =   6, w =   9
-- Decomposition: a  =  2, b  =  4
--                a0 =  2, b0 =  2, p0 =  2
--                a1 =  1, b1 =  2, p1 =  4
--                a2 =  1, b2 =  1, p2 =  2
--                g0 =  1, g1 =  -5
-- ROMs: 2^ 2 x 10  +  2^ 2 x  7  +  2^ 3 x  2  +  2^ 2 x  0  =      84 bits
-- Mult: 2 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T8_11 is
  component LNSSub_MNMX_T8_11_t0 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_t1 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_t2 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_t3 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_mult is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_xor2 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T8_11_xor3 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_11_t0 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_t0 is
begin
  with x select
    r <=
      "1001001011" when "00", -- t[0] = 587
      "1001100011" when "01", -- t[1] = 611
      "1010000000" when "10", -- t[2] = 640
      "1010100001" when "11", -- t[3] = 673
      "----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_11_t1 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_t1 is
begin
  with x select
    r <=
      "0110000" when "00", -- t[0] = 48
      "0111000" when "01", -- t[1] = 56
      "1000010" when "10", -- t[2] = 66
      "1010001" when "11", -- t[3] = 81
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_11_t2 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_t2 is
begin
  with x select
    r <=
      "00" when "00", -- t[0] = 0
      "10" when "01", -- t[1] = 2
      "01" when "10", -- t[2] = 1
      "11" when "11", -- t[3] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_11_t3 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_t3 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_11.all;

entity LNSSub_MNMX_T8_11_mult is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T8_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(8 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_11.all;

entity LNSSub_MNMX_T8_11_xor2 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T8_11_t2
    port map ( x => in_t,
               r => out_t );

  r(9 downto 2) <= (9 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_11.all;

entity LNSSub_MNMX_T8_11_xor3 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T8_11_t3
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_11.all;

entity LNSSub_MNMX_T8_11 is
  port ( x : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_11 is
  signal a0  : std_logic_vector(1 downto 0);
  signal r0  : std_logic_vector(9 downto 0);
  signal a1  : std_logic_vector(1 downto 0);
  signal b1  : std_logic_vector(1 downto 0);
  signal r1  : std_logic_vector(9 downto 0);
  signal a2  : std_logic_vector(0 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(9 downto 0);
  signal a3  : std_logic_vector(0 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(9 downto 0);
  signal sum : std_logic_vector(9 downto 0);
begin
  a0 <= x(5 downto 4);
  inst_t0 : LNSSub_MNMX_T8_11_t0
    port map ( x => a0,
               r => r0(9 downto 0) );

  a1 <= x(5 downto 4);
  b1 <= x(3 downto 2);
  inst_mult : LNSSub_MNMX_T8_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(5 downto 0) );
  r1(9 downto 6) <= (9 downto 6 => '0');

  a2 <= x(5 downto 5);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T8_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(9 downto 0) );

  a3 <= x(5 downto 5);
  b3 <= x(3 downto 3);
  inst_xor3 : LNSSub_MNMX_T8_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(9 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(9 downto 1);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.031250, -0.015625 [ -> [ 0.000000, 8.000000 [
-- Input:  wE =  -6, wF =  11, w =   5
-- Output: wE =   3, wF =   5, w =   8
-- Decomposition: a  =  2, b  =  3
--                a0 =  2, b0 =  2, p0 =  2
--                a1 =  1, b1 =  1, p1 =  4
--                a2 =  1, b2 =  1, p2 =  2
--                g0 =  1, g1 =  -4
-- ROMs: 2^ 2 x  9  +  2^ 2 x  8  +  2^ 2 x  1  +  2^ 2 x  0  =      72 bits
-- Mult: 2 x 8 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T9_11 is
  component LNSSub_MNMX_T9_11_t0 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_t1 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_t2 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_t3 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_mult is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_xor2 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T9_11_xor3 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T9_11_t0 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_t0 is
begin
  with x select
    r <=
      "101100101" when "00", -- t[0] = 357
      "101110001" when "01", -- t[1] = 369
      "101111111" when "10", -- t[2] = 383
      "110010000" when "11", -- t[3] = 400
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T9_11_t1 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_t1 is
begin
  with x select
    r <=
      "01100001" when "00", -- t[0] = 97
      "01110000" when "01", -- t[1] = 112
      "10000100" when "10", -- t[2] = 132
      "10100001" when "11", -- t[3] = 161
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T9_11_t2 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_t2 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "1" when "1", -- t[1] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T9_11_t3 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_t3 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T9_11.all;

entity LNSSub_MNMX_T9_11_mult is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_mult is
  signal out_t : std_logic_vector(7 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T9_11_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T9_11.all;

entity LNSSub_MNMX_T9_11_xor2 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T9_11_t2
    port map ( x => in_t,
               r => out_t );

  r(8 downto 1) <= (8 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T9_11.all;

entity LNSSub_MNMX_T9_11_xor3 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T9_11_t3
    port map ( x => in_t,
               r => out_t );

  r(8 downto 1) <= (8 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T9_11.all;

entity LNSSub_MNMX_T9_11 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_11 is
  signal a0  : std_logic_vector(1 downto 0);
  signal r0  : std_logic_vector(8 downto 0);
  signal a1  : std_logic_vector(1 downto 0);
  signal b1  : std_logic_vector(1 downto 0);
  signal r1  : std_logic_vector(8 downto 0);
  signal a2  : std_logic_vector(0 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(8 downto 0);
  signal a3  : std_logic_vector(0 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(8 downto 0);
  signal sum : std_logic_vector(8 downto 0);
begin
  a0 <= x(4 downto 3);
  inst_t0 : LNSSub_MNMX_T9_11_t0
    port map ( x => a0,
               r => r0(8 downto 0) );

  a1 <= x(4 downto 3);
  b1 <= x(2 downto 1);
  inst_mult : LNSSub_MNMX_T9_11_mult
    port map ( a => a1,
               b => b1,
               r => r1(4 downto 0) );
  r1(8 downto 5) <= (8 downto 5 => '0');

  a2 <= x(4 downto 4);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T9_11_xor2
    port map ( a => a2,
               b => b2,
               r => r2(8 downto 0) );

  a3 <= x(4 downto 4);
  b3 <= x(2 downto 2);
  inst_xor3 : LNSSub_MNMX_T9_11_xor3
    port map ( a => a3,
               b => b3,
               r => r3(8 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(8 downto 1);
end architecture;


-- Simple table: LNS subtraction function [ -0.015625, 0.000000 [ -> [ 0.000000, 16.000000 [
-- Input:  wE =  -6, wF =  11, w =   5
-- Output: wE =   4, wF =   4, w =   8

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T10_11 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T10_11 is
begin
  with x select
    r <=
      "01101001" when "00000", -- t[0] = 105
      "01101001" when "00001", -- t[1] = 105
      "01101010" when "00010", -- t[2] = 106
      "01101011" when "00011", -- t[3] = 107
      "01101100" when "00100", -- t[4] = 108
      "01101100" when "00101", -- t[5] = 108
      "01101101" when "00110", -- t[6] = 109
      "01101110" when "00111", -- t[7] = 110
      "01101111" when "01000", -- t[8] = 111
      "01110000" when "01001", -- t[9] = 112
      "01110001" when "01010", -- t[10] = 113
      "01110010" when "01011", -- t[11] = 114
      "01110011" when "01100", -- t[12] = 115
      "01110101" when "01101", -- t[13] = 117
      "01110110" when "01110", -- t[14] = 118
      "01110111" when "01111", -- t[15] = 119
      "01111001" when "10000", -- t[16] = 121
      "01111010" when "10001", -- t[17] = 122
      "01111100" when "10010", -- t[18] = 124
      "01111101" when "10011", -- t[19] = 125
      "01111111" when "10100", -- t[20] = 127
      "10000001" when "10101", -- t[21] = 129
      "10000011" when "10110", -- t[22] = 131
      "10000110" when "10111", -- t[23] = 134
      "10001000" when "11000", -- t[24] = 136
      "10001100" when "11001", -- t[25] = 140
      "10001111" when "11010", -- t[26] = 143
      "10010011" when "11011", -- t[27] = 147
      "10011000" when "11100", -- t[28] = 152
      "10011111" when "11101", -- t[29] = 159
      "10101000" when "11110", -- t[30] = 168
      "10111000" when "11111", -- t[31] = 184
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_lnssub_mnmx_11.all;

entity LNSSub_MNMX_11 is
  port ( x : in  std_logic_vector(14 downto 0);
         r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_11 is
  signal out_t0 : std_logic_vector(4 downto 0);
  signal out_t1 : std_logic_vector(7 downto 0);
  signal out_t2 : std_logic_vector(9 downto 0);
  signal out_t3 : std_logic_vector(10 downto 0);
  signal out_t4 : std_logic_vector(11 downto 0);
  signal out_t5 : std_logic_vector(10 downto 0);
  signal out_t6 : std_logic_vector(9 downto 0);
  signal out_t7 : std_logic_vector(9 downto 0);
  signal out_t8 : std_logic_vector(8 downto 0);
  signal out_t9 : std_logic_vector(7 downto 0);
  signal out_t10 : std_logic_vector(7 downto 0);
begin
  inst_t0 : LNSSub_MNMX_T0_11
    port map ( x => x(14 downto 0),
               r => out_t0 );

  inst_t1 : LNSSub_MNMX_T1_11
    port map ( x => x(12 downto 0),
               r => out_t1 );

  inst_t2 : LNSSub_MNMX_T2_11
    port map ( x => x(11 downto 0),
               r => out_t2 );

  inst_t3 : LNSSub_MNMX_T3_11
    port map ( x => x(10 downto 0),
               r => out_t3 );

  inst_t4 : LNSSub_MNMX_T4_11
    port map ( x => x(9 downto 0),
               r => out_t4 );

  inst_t5 : LNSSub_MNMX_T5_11
    port map ( x => x(8 downto 0),
               r => out_t5 );

  inst_t6 : LNSSub_MNMX_T6_11
    port map ( x => x(7 downto 0),
               r => out_t6 );

  inst_t7 : LNSSub_MNMX_T7_11
    port map ( x => x(6 downto 0),
               r => out_t7 );

  inst_t8 : LNSSub_MNMX_T8_11
    port map ( x => x(5 downto 0),
               r => out_t8 );

  inst_t9 : LNSSub_MNMX_T9_11
    port map ( x => x(4 downto 0),
               r => out_t9 );

  inst_t10 : LNSSub_MNMX_T10_11
    port map ( x => x(4 downto 0),
               r => out_t10 );

  r <= (14 downto 5 => '0') & out_t0
         when x(14 downto 14) /= (14 downto 14 => '1') else
       (14 downto 8 => '0') & out_t1
         when x(13) /= '1' else
       (14 downto 10 => '0') & out_t2
         when x(12) /= '1' else
       (14 downto 11 => '0') & out_t3
         when x(11) /= '1' else
       (14 downto 12 => '0') & out_t4
         when x(10) /= '1' else
       (14 downto 13 => '0') & out_t5 & (1 downto 0 => '0')
         when x(9) /= '1' else
       (14 downto 13 => '0') & out_t6 & (2 downto 0 => '0')
         when x(8) /= '1' else
       (14 downto 14 => '0') & out_t7 & (3 downto 0 => '0')
         when x(7) /= '1' else
       (14 downto 14 => '0') & out_t8 & (4 downto 0 => '0')
         when x(6) /= '1' else
       (14 downto 14 => '0') & out_t9 & (5 downto 0 => '0')
         when x(5) /= '1' else
       out_t10 & (6 downto 0 => '0');
end architecture;
