-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of LNS sub function with 8-bit integer part and 10-bit fractional part
-- wI = 14 bits
-- wO = 14 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnssub_mnmx_10 is
  component LNSSub_MNMX_T0_10 is
    port ( x : in  std_logic_vector(13 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10 is
    port ( x : in  std_logic_vector(11 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10 is
    port ( x : in  std_logic_vector(10 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10 is
    port ( x : in  std_logic_vector(9 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10 is
    port ( x : in  std_logic_vector(8 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10 is
    port ( x : in  std_logic_vector(7 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10 is
    port ( x : in  std_logic_vector(6 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10 is
    port ( x : in  std_logic_vector(5 downto 0);
           r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T9_10 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
end package;


-- Simple table: LNS subtraction function [ -16.000000, 0.000000 [ -> [ 0.000000, 0.015625 [
-- (restricted to [ -16.000000, -8.000000 [ )
-- Input:  wE =   4, wF =  10, w =  14
-- Output: wE =  -6, wF =  10, w =   4

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T0_10 is
  port ( x : in  std_logic_vector(13 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T0_10 is
  signal r0 : std_logic_vector(3 downto 0);
begin
--  r <= "0000";

  with x select
    r <=
      "0000" when "00000000000000", -- t[0] = 0
      "0000" when "00000000000001", -- t[1] = 0
      "0000" when "00000000000010", -- t[2] = 0
      "0000" when "00000000000011", -- t[3] = 0
      "0000" when "00000000000100", -- t[4] = 0
      "0000" when "00000000000101", -- t[5] = 0
      "0000" when "00000000000110", -- t[6] = 0
      "0000" when "00000000000111", -- t[7] = 0
      "0000" when "00000000001000", -- t[8] = 0
      "0000" when "00000000001001", -- t[9] = 0
      "0000" when "00000000001010", -- t[10] = 0
      "0000" when "00000000001011", -- t[11] = 0
      "0000" when "00000000001100", -- t[12] = 0
      "0000" when "00000000001101", -- t[13] = 0
      "0000" when "00000000001110", -- t[14] = 0
      "0000" when "00000000001111", -- t[15] = 0
      "0000" when "00000000010000", -- t[16] = 0
      "0000" when "00000000010001", -- t[17] = 0
      "0000" when "00000000010010", -- t[18] = 0
      "0000" when "00000000010011", -- t[19] = 0
      "0000" when "00000000010100", -- t[20] = 0
      "0000" when "00000000010101", -- t[21] = 0
      "0000" when "00000000010110", -- t[22] = 0
      "0000" when "00000000010111", -- t[23] = 0
      "0000" when "00000000011000", -- t[24] = 0
      "0000" when "00000000011001", -- t[25] = 0
      "0000" when "00000000011010", -- t[26] = 0
      "0000" when "00000000011011", -- t[27] = 0
      "0000" when "00000000011100", -- t[28] = 0
      "0000" when "00000000011101", -- t[29] = 0
      "0000" when "00000000011110", -- t[30] = 0
      "0000" when "00000000011111", -- t[31] = 0
      "0000" when "00000000100000", -- t[32] = 0
      "0000" when "00000000100001", -- t[33] = 0
      "0000" when "00000000100010", -- t[34] = 0
      "0000" when "00000000100011", -- t[35] = 0
      "0000" when "00000000100100", -- t[36] = 0
      "0000" when "00000000100101", -- t[37] = 0
      "0000" when "00000000100110", -- t[38] = 0
      "0000" when "00000000100111", -- t[39] = 0
      "0000" when "00000000101000", -- t[40] = 0
      "0000" when "00000000101001", -- t[41] = 0
      "0000" when "00000000101010", -- t[42] = 0
      "0000" when "00000000101011", -- t[43] = 0
      "0000" when "00000000101100", -- t[44] = 0
      "0000" when "00000000101101", -- t[45] = 0
      "0000" when "00000000101110", -- t[46] = 0
      "0000" when "00000000101111", -- t[47] = 0
      "0000" when "00000000110000", -- t[48] = 0
      "0000" when "00000000110001", -- t[49] = 0
      "0000" when "00000000110010", -- t[50] = 0
      "0000" when "00000000110011", -- t[51] = 0
      "0000" when "00000000110100", -- t[52] = 0
      "0000" when "00000000110101", -- t[53] = 0
      "0000" when "00000000110110", -- t[54] = 0
      "0000" when "00000000110111", -- t[55] = 0
      "0000" when "00000000111000", -- t[56] = 0
      "0000" when "00000000111001", -- t[57] = 0
      "0000" when "00000000111010", -- t[58] = 0
      "0000" when "00000000111011", -- t[59] = 0
      "0000" when "00000000111100", -- t[60] = 0
      "0000" when "00000000111101", -- t[61] = 0
      "0000" when "00000000111110", -- t[62] = 0
      "0000" when "00000000111111", -- t[63] = 0
      "0000" when "00000001000000", -- t[64] = 0
      "0000" when "00000001000001", -- t[65] = 0
      "0000" when "00000001000010", -- t[66] = 0
      "0000" when "00000001000011", -- t[67] = 0
      "0000" when "00000001000100", -- t[68] = 0
      "0000" when "00000001000101", -- t[69] = 0
      "0000" when "00000001000110", -- t[70] = 0
      "0000" when "00000001000111", -- t[71] = 0
      "0000" when "00000001001000", -- t[72] = 0
      "0000" when "00000001001001", -- t[73] = 0
      "0000" when "00000001001010", -- t[74] = 0
      "0000" when "00000001001011", -- t[75] = 0
      "0000" when "00000001001100", -- t[76] = 0
      "0000" when "00000001001101", -- t[77] = 0
      "0000" when "00000001001110", -- t[78] = 0
      "0000" when "00000001001111", -- t[79] = 0
      "0000" when "00000001010000", -- t[80] = 0
      "0000" when "00000001010001", -- t[81] = 0
      "0000" when "00000001010010", -- t[82] = 0
      "0000" when "00000001010011", -- t[83] = 0
      "0000" when "00000001010100", -- t[84] = 0
      "0000" when "00000001010101", -- t[85] = 0
      "0000" when "00000001010110", -- t[86] = 0
      "0000" when "00000001010111", -- t[87] = 0
      "0000" when "00000001011000", -- t[88] = 0
      "0000" when "00000001011001", -- t[89] = 0
      "0000" when "00000001011010", -- t[90] = 0
      "0000" when "00000001011011", -- t[91] = 0
      "0000" when "00000001011100", -- t[92] = 0
      "0000" when "00000001011101", -- t[93] = 0
      "0000" when "00000001011110", -- t[94] = 0
      "0000" when "00000001011111", -- t[95] = 0
      "0000" when "00000001100000", -- t[96] = 0
      "0000" when "00000001100001", -- t[97] = 0
      "0000" when "00000001100010", -- t[98] = 0
      "0000" when "00000001100011", -- t[99] = 0
      "0000" when "00000001100100", -- t[100] = 0
      "0000" when "00000001100101", -- t[101] = 0
      "0000" when "00000001100110", -- t[102] = 0
      "0000" when "00000001100111", -- t[103] = 0
      "0000" when "00000001101000", -- t[104] = 0
      "0000" when "00000001101001", -- t[105] = 0
      "0000" when "00000001101010", -- t[106] = 0
      "0000" when "00000001101011", -- t[107] = 0
      "0000" when "00000001101100", -- t[108] = 0
      "0000" when "00000001101101", -- t[109] = 0
      "0000" when "00000001101110", -- t[110] = 0
      "0000" when "00000001101111", -- t[111] = 0
      "0000" when "00000001110000", -- t[112] = 0
      "0000" when "00000001110001", -- t[113] = 0
      "0000" when "00000001110010", -- t[114] = 0
      "0000" when "00000001110011", -- t[115] = 0
      "0000" when "00000001110100", -- t[116] = 0
      "0000" when "00000001110101", -- t[117] = 0
      "0000" when "00000001110110", -- t[118] = 0
      "0000" when "00000001110111", -- t[119] = 0
      "0000" when "00000001111000", -- t[120] = 0
      "0000" when "00000001111001", -- t[121] = 0
      "0000" when "00000001111010", -- t[122] = 0
      "0000" when "00000001111011", -- t[123] = 0
      "0000" when "00000001111100", -- t[124] = 0
      "0000" when "00000001111101", -- t[125] = 0
      "0000" when "00000001111110", -- t[126] = 0
      "0000" when "00000001111111", -- t[127] = 0
      "0000" when "00000010000000", -- t[128] = 0
      "0000" when "00000010000001", -- t[129] = 0
      "0000" when "00000010000010", -- t[130] = 0
      "0000" when "00000010000011", -- t[131] = 0
      "0000" when "00000010000100", -- t[132] = 0
      "0000" when "00000010000101", -- t[133] = 0
      "0000" when "00000010000110", -- t[134] = 0
      "0000" when "00000010000111", -- t[135] = 0
      "0000" when "00000010001000", -- t[136] = 0
      "0000" when "00000010001001", -- t[137] = 0
      "0000" when "00000010001010", -- t[138] = 0
      "0000" when "00000010001011", -- t[139] = 0
      "0000" when "00000010001100", -- t[140] = 0
      "0000" when "00000010001101", -- t[141] = 0
      "0000" when "00000010001110", -- t[142] = 0
      "0000" when "00000010001111", -- t[143] = 0
      "0000" when "00000010010000", -- t[144] = 0
      "0000" when "00000010010001", -- t[145] = 0
      "0000" when "00000010010010", -- t[146] = 0
      "0000" when "00000010010011", -- t[147] = 0
      "0000" when "00000010010100", -- t[148] = 0
      "0000" when "00000010010101", -- t[149] = 0
      "0000" when "00000010010110", -- t[150] = 0
      "0000" when "00000010010111", -- t[151] = 0
      "0000" when "00000010011000", -- t[152] = 0
      "0000" when "00000010011001", -- t[153] = 0
      "0000" when "00000010011010", -- t[154] = 0
      "0000" when "00000010011011", -- t[155] = 0
      "0000" when "00000010011100", -- t[156] = 0
      "0000" when "00000010011101", -- t[157] = 0
      "0000" when "00000010011110", -- t[158] = 0
      "0000" when "00000010011111", -- t[159] = 0
      "0000" when "00000010100000", -- t[160] = 0
      "0000" when "00000010100001", -- t[161] = 0
      "0000" when "00000010100010", -- t[162] = 0
      "0000" when "00000010100011", -- t[163] = 0
      "0000" when "00000010100100", -- t[164] = 0
      "0000" when "00000010100101", -- t[165] = 0
      "0000" when "00000010100110", -- t[166] = 0
      "0000" when "00000010100111", -- t[167] = 0
      "0000" when "00000010101000", -- t[168] = 0
      "0000" when "00000010101001", -- t[169] = 0
      "0000" when "00000010101010", -- t[170] = 0
      "0000" when "00000010101011", -- t[171] = 0
      "0000" when "00000010101100", -- t[172] = 0
      "0000" when "00000010101101", -- t[173] = 0
      "0000" when "00000010101110", -- t[174] = 0
      "0000" when "00000010101111", -- t[175] = 0
      "0000" when "00000010110000", -- t[176] = 0
      "0000" when "00000010110001", -- t[177] = 0
      "0000" when "00000010110010", -- t[178] = 0
      "0000" when "00000010110011", -- t[179] = 0
      "0000" when "00000010110100", -- t[180] = 0
      "0000" when "00000010110101", -- t[181] = 0
      "0000" when "00000010110110", -- t[182] = 0
      "0000" when "00000010110111", -- t[183] = 0
      "0000" when "00000010111000", -- t[184] = 0
      "0000" when "00000010111001", -- t[185] = 0
      "0000" when "00000010111010", -- t[186] = 0
      "0000" when "00000010111011", -- t[187] = 0
      "0000" when "00000010111100", -- t[188] = 0
      "0000" when "00000010111101", -- t[189] = 0
      "0000" when "00000010111110", -- t[190] = 0
      "0000" when "00000010111111", -- t[191] = 0
      "0000" when "00000011000000", -- t[192] = 0
      "0000" when "00000011000001", -- t[193] = 0
      "0000" when "00000011000010", -- t[194] = 0
      "0000" when "00000011000011", -- t[195] = 0
      "0000" when "00000011000100", -- t[196] = 0
      "0000" when "00000011000101", -- t[197] = 0
      "0000" when "00000011000110", -- t[198] = 0
      "0000" when "00000011000111", -- t[199] = 0
      "0000" when "00000011001000", -- t[200] = 0
      "0000" when "00000011001001", -- t[201] = 0
      "0000" when "00000011001010", -- t[202] = 0
      "0000" when "00000011001011", -- t[203] = 0
      "0000" when "00000011001100", -- t[204] = 0
      "0000" when "00000011001101", -- t[205] = 0
      "0000" when "00000011001110", -- t[206] = 0
      "0000" when "00000011001111", -- t[207] = 0
      "0000" when "00000011010000", -- t[208] = 0
      "0000" when "00000011010001", -- t[209] = 0
      "0000" when "00000011010010", -- t[210] = 0
      "0000" when "00000011010011", -- t[211] = 0
      "0000" when "00000011010100", -- t[212] = 0
      "0000" when "00000011010101", -- t[213] = 0
      "0000" when "00000011010110", -- t[214] = 0
      "0000" when "00000011010111", -- t[215] = 0
      "0000" when "00000011011000", -- t[216] = 0
      "0000" when "00000011011001", -- t[217] = 0
      "0000" when "00000011011010", -- t[218] = 0
      "0000" when "00000011011011", -- t[219] = 0
      "0000" when "00000011011100", -- t[220] = 0
      "0000" when "00000011011101", -- t[221] = 0
      "0000" when "00000011011110", -- t[222] = 0
      "0000" when "00000011011111", -- t[223] = 0
      "0000" when "00000011100000", -- t[224] = 0
      "0000" when "00000011100001", -- t[225] = 0
      "0000" when "00000011100010", -- t[226] = 0
      "0000" when "00000011100011", -- t[227] = 0
      "0000" when "00000011100100", -- t[228] = 0
      "0000" when "00000011100101", -- t[229] = 0
      "0000" when "00000011100110", -- t[230] = 0
      "0000" when "00000011100111", -- t[231] = 0
      "0000" when "00000011101000", -- t[232] = 0
      "0000" when "00000011101001", -- t[233] = 0
      "0000" when "00000011101010", -- t[234] = 0
      "0000" when "00000011101011", -- t[235] = 0
      "0000" when "00000011101100", -- t[236] = 0
      "0000" when "00000011101101", -- t[237] = 0
      "0000" when "00000011101110", -- t[238] = 0
      "0000" when "00000011101111", -- t[239] = 0
      "0000" when "00000011110000", -- t[240] = 0
      "0000" when "00000011110001", -- t[241] = 0
      "0000" when "00000011110010", -- t[242] = 0
      "0000" when "00000011110011", -- t[243] = 0
      "0000" when "00000011110100", -- t[244] = 0
      "0000" when "00000011110101", -- t[245] = 0
      "0000" when "00000011110110", -- t[246] = 0
      "0000" when "00000011110111", -- t[247] = 0
      "0000" when "00000011111000", -- t[248] = 0
      "0000" when "00000011111001", -- t[249] = 0
      "0000" when "00000011111010", -- t[250] = 0
      "0000" when "00000011111011", -- t[251] = 0
      "0000" when "00000011111100", -- t[252] = 0
      "0000" when "00000011111101", -- t[253] = 0
      "0000" when "00000011111110", -- t[254] = 0
      "0000" when "00000011111111", -- t[255] = 0
      "0000" when "00000100000000", -- t[256] = 0
      "0000" when "00000100000001", -- t[257] = 0
      "0000" when "00000100000010", -- t[258] = 0
      "0000" when "00000100000011", -- t[259] = 0
      "0000" when "00000100000100", -- t[260] = 0
      "0000" when "00000100000101", -- t[261] = 0
      "0000" when "00000100000110", -- t[262] = 0
      "0000" when "00000100000111", -- t[263] = 0
      "0000" when "00000100001000", -- t[264] = 0
      "0000" when "00000100001001", -- t[265] = 0
      "0000" when "00000100001010", -- t[266] = 0
      "0000" when "00000100001011", -- t[267] = 0
      "0000" when "00000100001100", -- t[268] = 0
      "0000" when "00000100001101", -- t[269] = 0
      "0000" when "00000100001110", -- t[270] = 0
      "0000" when "00000100001111", -- t[271] = 0
      "0000" when "00000100010000", -- t[272] = 0
      "0000" when "00000100010001", -- t[273] = 0
      "0000" when "00000100010010", -- t[274] = 0
      "0000" when "00000100010011", -- t[275] = 0
      "0000" when "00000100010100", -- t[276] = 0
      "0000" when "00000100010101", -- t[277] = 0
      "0000" when "00000100010110", -- t[278] = 0
      "0000" when "00000100010111", -- t[279] = 0
      "0000" when "00000100011000", -- t[280] = 0
      "0000" when "00000100011001", -- t[281] = 0
      "0000" when "00000100011010", -- t[282] = 0
      "0000" when "00000100011011", -- t[283] = 0
      "0000" when "00000100011100", -- t[284] = 0
      "0000" when "00000100011101", -- t[285] = 0
      "0000" when "00000100011110", -- t[286] = 0
      "0000" when "00000100011111", -- t[287] = 0
      "0000" when "00000100100000", -- t[288] = 0
      "0000" when "00000100100001", -- t[289] = 0
      "0000" when "00000100100010", -- t[290] = 0
      "0000" when "00000100100011", -- t[291] = 0
      "0000" when "00000100100100", -- t[292] = 0
      "0000" when "00000100100101", -- t[293] = 0
      "0000" when "00000100100110", -- t[294] = 0
      "0000" when "00000100100111", -- t[295] = 0
      "0000" when "00000100101000", -- t[296] = 0
      "0000" when "00000100101001", -- t[297] = 0
      "0000" when "00000100101010", -- t[298] = 0
      "0000" when "00000100101011", -- t[299] = 0
      "0000" when "00000100101100", -- t[300] = 0
      "0000" when "00000100101101", -- t[301] = 0
      "0000" when "00000100101110", -- t[302] = 0
      "0000" when "00000100101111", -- t[303] = 0
      "0000" when "00000100110000", -- t[304] = 0
      "0000" when "00000100110001", -- t[305] = 0
      "0000" when "00000100110010", -- t[306] = 0
      "0000" when "00000100110011", -- t[307] = 0
      "0000" when "00000100110100", -- t[308] = 0
      "0000" when "00000100110101", -- t[309] = 0
      "0000" when "00000100110110", -- t[310] = 0
      "0000" when "00000100110111", -- t[311] = 0
      "0000" when "00000100111000", -- t[312] = 0
      "0000" when "00000100111001", -- t[313] = 0
      "0000" when "00000100111010", -- t[314] = 0
      "0000" when "00000100111011", -- t[315] = 0
      "0000" when "00000100111100", -- t[316] = 0
      "0000" when "00000100111101", -- t[317] = 0
      "0000" when "00000100111110", -- t[318] = 0
      "0000" when "00000100111111", -- t[319] = 0
      "0000" when "00000101000000", -- t[320] = 0
      "0000" when "00000101000001", -- t[321] = 0
      "0000" when "00000101000010", -- t[322] = 0
      "0000" when "00000101000011", -- t[323] = 0
      "0000" when "00000101000100", -- t[324] = 0
      "0000" when "00000101000101", -- t[325] = 0
      "0000" when "00000101000110", -- t[326] = 0
      "0000" when "00000101000111", -- t[327] = 0
      "0000" when "00000101001000", -- t[328] = 0
      "0000" when "00000101001001", -- t[329] = 0
      "0000" when "00000101001010", -- t[330] = 0
      "0000" when "00000101001011", -- t[331] = 0
      "0000" when "00000101001100", -- t[332] = 0
      "0000" when "00000101001101", -- t[333] = 0
      "0000" when "00000101001110", -- t[334] = 0
      "0000" when "00000101001111", -- t[335] = 0
      "0000" when "00000101010000", -- t[336] = 0
      "0000" when "00000101010001", -- t[337] = 0
      "0000" when "00000101010010", -- t[338] = 0
      "0000" when "00000101010011", -- t[339] = 0
      "0000" when "00000101010100", -- t[340] = 0
      "0000" when "00000101010101", -- t[341] = 0
      "0000" when "00000101010110", -- t[342] = 0
      "0000" when "00000101010111", -- t[343] = 0
      "0000" when "00000101011000", -- t[344] = 0
      "0000" when "00000101011001", -- t[345] = 0
      "0000" when "00000101011010", -- t[346] = 0
      "0000" when "00000101011011", -- t[347] = 0
      "0000" when "00000101011100", -- t[348] = 0
      "0000" when "00000101011101", -- t[349] = 0
      "0000" when "00000101011110", -- t[350] = 0
      "0000" when "00000101011111", -- t[351] = 0
      "0000" when "00000101100000", -- t[352] = 0
      "0000" when "00000101100001", -- t[353] = 0
      "0000" when "00000101100010", -- t[354] = 0
      "0000" when "00000101100011", -- t[355] = 0
      "0000" when "00000101100100", -- t[356] = 0
      "0000" when "00000101100101", -- t[357] = 0
      "0000" when "00000101100110", -- t[358] = 0
      "0000" when "00000101100111", -- t[359] = 0
      "0000" when "00000101101000", -- t[360] = 0
      "0000" when "00000101101001", -- t[361] = 0
      "0000" when "00000101101010", -- t[362] = 0
      "0000" when "00000101101011", -- t[363] = 0
      "0000" when "00000101101100", -- t[364] = 0
      "0000" when "00000101101101", -- t[365] = 0
      "0000" when "00000101101110", -- t[366] = 0
      "0000" when "00000101101111", -- t[367] = 0
      "0000" when "00000101110000", -- t[368] = 0
      "0000" when "00000101110001", -- t[369] = 0
      "0000" when "00000101110010", -- t[370] = 0
      "0000" when "00000101110011", -- t[371] = 0
      "0000" when "00000101110100", -- t[372] = 0
      "0000" when "00000101110101", -- t[373] = 0
      "0000" when "00000101110110", -- t[374] = 0
      "0000" when "00000101110111", -- t[375] = 0
      "0000" when "00000101111000", -- t[376] = 0
      "0000" when "00000101111001", -- t[377] = 0
      "0000" when "00000101111010", -- t[378] = 0
      "0000" when "00000101111011", -- t[379] = 0
      "0000" when "00000101111100", -- t[380] = 0
      "0000" when "00000101111101", -- t[381] = 0
      "0000" when "00000101111110", -- t[382] = 0
      "0000" when "00000101111111", -- t[383] = 0
      "0000" when "00000110000000", -- t[384] = 0
      "0000" when "00000110000001", -- t[385] = 0
      "0000" when "00000110000010", -- t[386] = 0
      "0000" when "00000110000011", -- t[387] = 0
      "0000" when "00000110000100", -- t[388] = 0
      "0000" when "00000110000101", -- t[389] = 0
      "0000" when "00000110000110", -- t[390] = 0
      "0000" when "00000110000111", -- t[391] = 0
      "0000" when "00000110001000", -- t[392] = 0
      "0000" when "00000110001001", -- t[393] = 0
      "0000" when "00000110001010", -- t[394] = 0
      "0000" when "00000110001011", -- t[395] = 0
      "0000" when "00000110001100", -- t[396] = 0
      "0000" when "00000110001101", -- t[397] = 0
      "0000" when "00000110001110", -- t[398] = 0
      "0000" when "00000110001111", -- t[399] = 0
      "0000" when "00000110010000", -- t[400] = 0
      "0000" when "00000110010001", -- t[401] = 0
      "0000" when "00000110010010", -- t[402] = 0
      "0000" when "00000110010011", -- t[403] = 0
      "0000" when "00000110010100", -- t[404] = 0
      "0000" when "00000110010101", -- t[405] = 0
      "0000" when "00000110010110", -- t[406] = 0
      "0000" when "00000110010111", -- t[407] = 0
      "0000" when "00000110011000", -- t[408] = 0
      "0000" when "00000110011001", -- t[409] = 0
      "0000" when "00000110011010", -- t[410] = 0
      "0000" when "00000110011011", -- t[411] = 0
      "0000" when "00000110011100", -- t[412] = 0
      "0000" when "00000110011101", -- t[413] = 0
      "0000" when "00000110011110", -- t[414] = 0
      "0000" when "00000110011111", -- t[415] = 0
      "0000" when "00000110100000", -- t[416] = 0
      "0000" when "00000110100001", -- t[417] = 0
      "0000" when "00000110100010", -- t[418] = 0
      "0000" when "00000110100011", -- t[419] = 0
      "0000" when "00000110100100", -- t[420] = 0
      "0000" when "00000110100101", -- t[421] = 0
      "0000" when "00000110100110", -- t[422] = 0
      "0000" when "00000110100111", -- t[423] = 0
      "0000" when "00000110101000", -- t[424] = 0
      "0000" when "00000110101001", -- t[425] = 0
      "0000" when "00000110101010", -- t[426] = 0
      "0000" when "00000110101011", -- t[427] = 0
      "0000" when "00000110101100", -- t[428] = 0
      "0000" when "00000110101101", -- t[429] = 0
      "0000" when "00000110101110", -- t[430] = 0
      "0000" when "00000110101111", -- t[431] = 0
      "0000" when "00000110110000", -- t[432] = 0
      "0000" when "00000110110001", -- t[433] = 0
      "0000" when "00000110110010", -- t[434] = 0
      "0000" when "00000110110011", -- t[435] = 0
      "0000" when "00000110110100", -- t[436] = 0
      "0000" when "00000110110101", -- t[437] = 0
      "0000" when "00000110110110", -- t[438] = 0
      "0000" when "00000110110111", -- t[439] = 0
      "0000" when "00000110111000", -- t[440] = 0
      "0000" when "00000110111001", -- t[441] = 0
      "0000" when "00000110111010", -- t[442] = 0
      "0000" when "00000110111011", -- t[443] = 0
      "0000" when "00000110111100", -- t[444] = 0
      "0000" when "00000110111101", -- t[445] = 0
      "0000" when "00000110111110", -- t[446] = 0
      "0000" when "00000110111111", -- t[447] = 0
      "0000" when "00000111000000", -- t[448] = 0
      "0000" when "00000111000001", -- t[449] = 0
      "0000" when "00000111000010", -- t[450] = 0
      "0000" when "00000111000011", -- t[451] = 0
      "0000" when "00000111000100", -- t[452] = 0
      "0000" when "00000111000101", -- t[453] = 0
      "0000" when "00000111000110", -- t[454] = 0
      "0000" when "00000111000111", -- t[455] = 0
      "0000" when "00000111001000", -- t[456] = 0
      "0000" when "00000111001001", -- t[457] = 0
      "0000" when "00000111001010", -- t[458] = 0
      "0000" when "00000111001011", -- t[459] = 0
      "0000" when "00000111001100", -- t[460] = 0
      "0000" when "00000111001101", -- t[461] = 0
      "0000" when "00000111001110", -- t[462] = 0
      "0000" when "00000111001111", -- t[463] = 0
      "0000" when "00000111010000", -- t[464] = 0
      "0000" when "00000111010001", -- t[465] = 0
      "0000" when "00000111010010", -- t[466] = 0
      "0000" when "00000111010011", -- t[467] = 0
      "0000" when "00000111010100", -- t[468] = 0
      "0000" when "00000111010101", -- t[469] = 0
      "0000" when "00000111010110", -- t[470] = 0
      "0000" when "00000111010111", -- t[471] = 0
      "0000" when "00000111011000", -- t[472] = 0
      "0000" when "00000111011001", -- t[473] = 0
      "0000" when "00000111011010", -- t[474] = 0
      "0000" when "00000111011011", -- t[475] = 0
      "0000" when "00000111011100", -- t[476] = 0
      "0000" when "00000111011101", -- t[477] = 0
      "0000" when "00000111011110", -- t[478] = 0
      "0000" when "00000111011111", -- t[479] = 0
      "0000" when "00000111100000", -- t[480] = 0
      "0000" when "00000111100001", -- t[481] = 0
      "0000" when "00000111100010", -- t[482] = 0
      "0000" when "00000111100011", -- t[483] = 0
      "0000" when "00000111100100", -- t[484] = 0
      "0000" when "00000111100101", -- t[485] = 0
      "0000" when "00000111100110", -- t[486] = 0
      "0000" when "00000111100111", -- t[487] = 0
      "0000" when "00000111101000", -- t[488] = 0
      "0000" when "00000111101001", -- t[489] = 0
      "0000" when "00000111101010", -- t[490] = 0
      "0000" when "00000111101011", -- t[491] = 0
      "0000" when "00000111101100", -- t[492] = 0
      "0000" when "00000111101101", -- t[493] = 0
      "0000" when "00000111101110", -- t[494] = 0
      "0000" when "00000111101111", -- t[495] = 0
      "0000" when "00000111110000", -- t[496] = 0
      "0000" when "00000111110001", -- t[497] = 0
      "0000" when "00000111110010", -- t[498] = 0
      "0000" when "00000111110011", -- t[499] = 0
      "0000" when "00000111110100", -- t[500] = 0
      "0000" when "00000111110101", -- t[501] = 0
      "0000" when "00000111110110", -- t[502] = 0
      "0000" when "00000111110111", -- t[503] = 0
      "0000" when "00000111111000", -- t[504] = 0
      "0000" when "00000111111001", -- t[505] = 0
      "0000" when "00000111111010", -- t[506] = 0
      "0000" when "00000111111011", -- t[507] = 0
      "0000" when "00000111111100", -- t[508] = 0
      "0000" when "00000111111101", -- t[509] = 0
      "0000" when "00000111111110", -- t[510] = 0
      "0000" when "00000111111111", -- t[511] = 0
      "0000" when "00001000000000", -- t[512] = 0
      "0000" when "00001000000001", -- t[513] = 0
      "0000" when "00001000000010", -- t[514] = 0
      "0000" when "00001000000011", -- t[515] = 0
      "0000" when "00001000000100", -- t[516] = 0
      "0000" when "00001000000101", -- t[517] = 0
      "0000" when "00001000000110", -- t[518] = 0
      "0000" when "00001000000111", -- t[519] = 0
      "0000" when "00001000001000", -- t[520] = 0
      "0000" when "00001000001001", -- t[521] = 0
      "0000" when "00001000001010", -- t[522] = 0
      "0000" when "00001000001011", -- t[523] = 0
      "0000" when "00001000001100", -- t[524] = 0
      "0000" when "00001000001101", -- t[525] = 0
      "0000" when "00001000001110", -- t[526] = 0
      "0000" when "00001000001111", -- t[527] = 0
      "0000" when "00001000010000", -- t[528] = 0
      "0000" when "00001000010001", -- t[529] = 0
      "0000" when "00001000010010", -- t[530] = 0
      "0000" when "00001000010011", -- t[531] = 0
      "0000" when "00001000010100", -- t[532] = 0
      "0000" when "00001000010101", -- t[533] = 0
      "0000" when "00001000010110", -- t[534] = 0
      "0000" when "00001000010111", -- t[535] = 0
      "0000" when "00001000011000", -- t[536] = 0
      "0000" when "00001000011001", -- t[537] = 0
      "0000" when "00001000011010", -- t[538] = 0
      "0000" when "00001000011011", -- t[539] = 0
      "0000" when "00001000011100", -- t[540] = 0
      "0000" when "00001000011101", -- t[541] = 0
      "0000" when "00001000011110", -- t[542] = 0
      "0000" when "00001000011111", -- t[543] = 0
      "0000" when "00001000100000", -- t[544] = 0
      "0000" when "00001000100001", -- t[545] = 0
      "0000" when "00001000100010", -- t[546] = 0
      "0000" when "00001000100011", -- t[547] = 0
      "0000" when "00001000100100", -- t[548] = 0
      "0000" when "00001000100101", -- t[549] = 0
      "0000" when "00001000100110", -- t[550] = 0
      "0000" when "00001000100111", -- t[551] = 0
      "0000" when "00001000101000", -- t[552] = 0
      "0000" when "00001000101001", -- t[553] = 0
      "0000" when "00001000101010", -- t[554] = 0
      "0000" when "00001000101011", -- t[555] = 0
      "0000" when "00001000101100", -- t[556] = 0
      "0000" when "00001000101101", -- t[557] = 0
      "0000" when "00001000101110", -- t[558] = 0
      "0000" when "00001000101111", -- t[559] = 0
      "0000" when "00001000110000", -- t[560] = 0
      "0000" when "00001000110001", -- t[561] = 0
      "0000" when "00001000110010", -- t[562] = 0
      "0000" when "00001000110011", -- t[563] = 0
      "0000" when "00001000110100", -- t[564] = 0
      "0000" when "00001000110101", -- t[565] = 0
      "0000" when "00001000110110", -- t[566] = 0
      "0000" when "00001000110111", -- t[567] = 0
      "0000" when "00001000111000", -- t[568] = 0
      "0000" when "00001000111001", -- t[569] = 0
      "0000" when "00001000111010", -- t[570] = 0
      "0000" when "00001000111011", -- t[571] = 0
      "0000" when "00001000111100", -- t[572] = 0
      "0000" when "00001000111101", -- t[573] = 0
      "0000" when "00001000111110", -- t[574] = 0
      "0000" when "00001000111111", -- t[575] = 0
      "0000" when "00001001000000", -- t[576] = 0
      "0000" when "00001001000001", -- t[577] = 0
      "0000" when "00001001000010", -- t[578] = 0
      "0000" when "00001001000011", -- t[579] = 0
      "0000" when "00001001000100", -- t[580] = 0
      "0000" when "00001001000101", -- t[581] = 0
      "0000" when "00001001000110", -- t[582] = 0
      "0000" when "00001001000111", -- t[583] = 0
      "0000" when "00001001001000", -- t[584] = 0
      "0000" when "00001001001001", -- t[585] = 0
      "0000" when "00001001001010", -- t[586] = 0
      "0000" when "00001001001011", -- t[587] = 0
      "0000" when "00001001001100", -- t[588] = 0
      "0000" when "00001001001101", -- t[589] = 0
      "0000" when "00001001001110", -- t[590] = 0
      "0000" when "00001001001111", -- t[591] = 0
      "0000" when "00001001010000", -- t[592] = 0
      "0000" when "00001001010001", -- t[593] = 0
      "0000" when "00001001010010", -- t[594] = 0
      "0000" when "00001001010011", -- t[595] = 0
      "0000" when "00001001010100", -- t[596] = 0
      "0000" when "00001001010101", -- t[597] = 0
      "0000" when "00001001010110", -- t[598] = 0
      "0000" when "00001001010111", -- t[599] = 0
      "0000" when "00001001011000", -- t[600] = 0
      "0000" when "00001001011001", -- t[601] = 0
      "0000" when "00001001011010", -- t[602] = 0
      "0000" when "00001001011011", -- t[603] = 0
      "0000" when "00001001011100", -- t[604] = 0
      "0000" when "00001001011101", -- t[605] = 0
      "0000" when "00001001011110", -- t[606] = 0
      "0000" when "00001001011111", -- t[607] = 0
      "0000" when "00001001100000", -- t[608] = 0
      "0000" when "00001001100001", -- t[609] = 0
      "0000" when "00001001100010", -- t[610] = 0
      "0000" when "00001001100011", -- t[611] = 0
      "0000" when "00001001100100", -- t[612] = 0
      "0000" when "00001001100101", -- t[613] = 0
      "0000" when "00001001100110", -- t[614] = 0
      "0000" when "00001001100111", -- t[615] = 0
      "0000" when "00001001101000", -- t[616] = 0
      "0000" when "00001001101001", -- t[617] = 0
      "0000" when "00001001101010", -- t[618] = 0
      "0000" when "00001001101011", -- t[619] = 0
      "0000" when "00001001101100", -- t[620] = 0
      "0000" when "00001001101101", -- t[621] = 0
      "0000" when "00001001101110", -- t[622] = 0
      "0000" when "00001001101111", -- t[623] = 0
      "0000" when "00001001110000", -- t[624] = 0
      "0000" when "00001001110001", -- t[625] = 0
      "0000" when "00001001110010", -- t[626] = 0
      "0000" when "00001001110011", -- t[627] = 0
      "0000" when "00001001110100", -- t[628] = 0
      "0000" when "00001001110101", -- t[629] = 0
      "0000" when "00001001110110", -- t[630] = 0
      "0000" when "00001001110111", -- t[631] = 0
      "0000" when "00001001111000", -- t[632] = 0
      "0000" when "00001001111001", -- t[633] = 0
      "0000" when "00001001111010", -- t[634] = 0
      "0000" when "00001001111011", -- t[635] = 0
      "0000" when "00001001111100", -- t[636] = 0
      "0000" when "00001001111101", -- t[637] = 0
      "0000" when "00001001111110", -- t[638] = 0
      "0000" when "00001001111111", -- t[639] = 0
      "0000" when "00001010000000", -- t[640] = 0
      "0000" when "00001010000001", -- t[641] = 0
      "0000" when "00001010000010", -- t[642] = 0
      "0000" when "00001010000011", -- t[643] = 0
      "0000" when "00001010000100", -- t[644] = 0
      "0000" when "00001010000101", -- t[645] = 0
      "0000" when "00001010000110", -- t[646] = 0
      "0000" when "00001010000111", -- t[647] = 0
      "0000" when "00001010001000", -- t[648] = 0
      "0000" when "00001010001001", -- t[649] = 0
      "0000" when "00001010001010", -- t[650] = 0
      "0000" when "00001010001011", -- t[651] = 0
      "0000" when "00001010001100", -- t[652] = 0
      "0000" when "00001010001101", -- t[653] = 0
      "0000" when "00001010001110", -- t[654] = 0
      "0000" when "00001010001111", -- t[655] = 0
      "0000" when "00001010010000", -- t[656] = 0
      "0000" when "00001010010001", -- t[657] = 0
      "0000" when "00001010010010", -- t[658] = 0
      "0000" when "00001010010011", -- t[659] = 0
      "0000" when "00001010010100", -- t[660] = 0
      "0000" when "00001010010101", -- t[661] = 0
      "0000" when "00001010010110", -- t[662] = 0
      "0000" when "00001010010111", -- t[663] = 0
      "0000" when "00001010011000", -- t[664] = 0
      "0000" when "00001010011001", -- t[665] = 0
      "0000" when "00001010011010", -- t[666] = 0
      "0000" when "00001010011011", -- t[667] = 0
      "0000" when "00001010011100", -- t[668] = 0
      "0000" when "00001010011101", -- t[669] = 0
      "0000" when "00001010011110", -- t[670] = 0
      "0000" when "00001010011111", -- t[671] = 0
      "0000" when "00001010100000", -- t[672] = 0
      "0000" when "00001010100001", -- t[673] = 0
      "0000" when "00001010100010", -- t[674] = 0
      "0000" when "00001010100011", -- t[675] = 0
      "0000" when "00001010100100", -- t[676] = 0
      "0000" when "00001010100101", -- t[677] = 0
      "0000" when "00001010100110", -- t[678] = 0
      "0000" when "00001010100111", -- t[679] = 0
      "0000" when "00001010101000", -- t[680] = 0
      "0000" when "00001010101001", -- t[681] = 0
      "0000" when "00001010101010", -- t[682] = 0
      "0000" when "00001010101011", -- t[683] = 0
      "0000" when "00001010101100", -- t[684] = 0
      "0000" when "00001010101101", -- t[685] = 0
      "0000" when "00001010101110", -- t[686] = 0
      "0000" when "00001010101111", -- t[687] = 0
      "0000" when "00001010110000", -- t[688] = 0
      "0000" when "00001010110001", -- t[689] = 0
      "0000" when "00001010110010", -- t[690] = 0
      "0000" when "00001010110011", -- t[691] = 0
      "0000" when "00001010110100", -- t[692] = 0
      "0000" when "00001010110101", -- t[693] = 0
      "0000" when "00001010110110", -- t[694] = 0
      "0000" when "00001010110111", -- t[695] = 0
      "0000" when "00001010111000", -- t[696] = 0
      "0000" when "00001010111001", -- t[697] = 0
      "0000" when "00001010111010", -- t[698] = 0
      "0000" when "00001010111011", -- t[699] = 0
      "0000" when "00001010111100", -- t[700] = 0
      "0000" when "00001010111101", -- t[701] = 0
      "0000" when "00001010111110", -- t[702] = 0
      "0000" when "00001010111111", -- t[703] = 0
      "0000" when "00001011000000", -- t[704] = 0
      "0000" when "00001011000001", -- t[705] = 0
      "0000" when "00001011000010", -- t[706] = 0
      "0000" when "00001011000011", -- t[707] = 0
      "0000" when "00001011000100", -- t[708] = 0
      "0000" when "00001011000101", -- t[709] = 0
      "0000" when "00001011000110", -- t[710] = 0
      "0000" when "00001011000111", -- t[711] = 0
      "0000" when "00001011001000", -- t[712] = 0
      "0000" when "00001011001001", -- t[713] = 0
      "0000" when "00001011001010", -- t[714] = 0
      "0000" when "00001011001011", -- t[715] = 0
      "0000" when "00001011001100", -- t[716] = 0
      "0000" when "00001011001101", -- t[717] = 0
      "0000" when "00001011001110", -- t[718] = 0
      "0000" when "00001011001111", -- t[719] = 0
      "0000" when "00001011010000", -- t[720] = 0
      "0000" when "00001011010001", -- t[721] = 0
      "0000" when "00001011010010", -- t[722] = 0
      "0000" when "00001011010011", -- t[723] = 0
      "0000" when "00001011010100", -- t[724] = 0
      "0000" when "00001011010101", -- t[725] = 0
      "0000" when "00001011010110", -- t[726] = 0
      "0000" when "00001011010111", -- t[727] = 0
      "0000" when "00001011011000", -- t[728] = 0
      "0000" when "00001011011001", -- t[729] = 0
      "0000" when "00001011011010", -- t[730] = 0
      "0000" when "00001011011011", -- t[731] = 0
      "0000" when "00001011011100", -- t[732] = 0
      "0000" when "00001011011101", -- t[733] = 0
      "0000" when "00001011011110", -- t[734] = 0
      "0000" when "00001011011111", -- t[735] = 0
      "0000" when "00001011100000", -- t[736] = 0
      "0000" when "00001011100001", -- t[737] = 0
      "0000" when "00001011100010", -- t[738] = 0
      "0000" when "00001011100011", -- t[739] = 0
      "0000" when "00001011100100", -- t[740] = 0
      "0000" when "00001011100101", -- t[741] = 0
      "0000" when "00001011100110", -- t[742] = 0
      "0000" when "00001011100111", -- t[743] = 0
      "0000" when "00001011101000", -- t[744] = 0
      "0000" when "00001011101001", -- t[745] = 0
      "0000" when "00001011101010", -- t[746] = 0
      "0000" when "00001011101011", -- t[747] = 0
      "0000" when "00001011101100", -- t[748] = 0
      "0000" when "00001011101101", -- t[749] = 0
      "0000" when "00001011101110", -- t[750] = 0
      "0000" when "00001011101111", -- t[751] = 0
      "0000" when "00001011110000", -- t[752] = 0
      "0000" when "00001011110001", -- t[753] = 0
      "0000" when "00001011110010", -- t[754] = 0
      "0000" when "00001011110011", -- t[755] = 0
      "0000" when "00001011110100", -- t[756] = 0
      "0000" when "00001011110101", -- t[757] = 0
      "0000" when "00001011110110", -- t[758] = 0
      "0000" when "00001011110111", -- t[759] = 0
      "0000" when "00001011111000", -- t[760] = 0
      "0000" when "00001011111001", -- t[761] = 0
      "0000" when "00001011111010", -- t[762] = 0
      "0000" when "00001011111011", -- t[763] = 0
      "0000" when "00001011111100", -- t[764] = 0
      "0000" when "00001011111101", -- t[765] = 0
      "0000" when "00001011111110", -- t[766] = 0
      "0000" when "00001011111111", -- t[767] = 0
      "0000" when "00001100000000", -- t[768] = 0
      "0000" when "00001100000001", -- t[769] = 0
      "0000" when "00001100000010", -- t[770] = 0
      "0000" when "00001100000011", -- t[771] = 0
      "0000" when "00001100000100", -- t[772] = 0
      "0000" when "00001100000101", -- t[773] = 0
      "0000" when "00001100000110", -- t[774] = 0
      "0000" when "00001100000111", -- t[775] = 0
      "0000" when "00001100001000", -- t[776] = 0
      "0000" when "00001100001001", -- t[777] = 0
      "0000" when "00001100001010", -- t[778] = 0
      "0000" when "00001100001011", -- t[779] = 0
      "0000" when "00001100001100", -- t[780] = 0
      "0000" when "00001100001101", -- t[781] = 0
      "0000" when "00001100001110", -- t[782] = 0
      "0000" when "00001100001111", -- t[783] = 0
      "0000" when "00001100010000", -- t[784] = 0
      "0000" when "00001100010001", -- t[785] = 0
      "0000" when "00001100010010", -- t[786] = 0
      "0000" when "00001100010011", -- t[787] = 0
      "0000" when "00001100010100", -- t[788] = 0
      "0000" when "00001100010101", -- t[789] = 0
      "0000" when "00001100010110", -- t[790] = 0
      "0000" when "00001100010111", -- t[791] = 0
      "0000" when "00001100011000", -- t[792] = 0
      "0000" when "00001100011001", -- t[793] = 0
      "0000" when "00001100011010", -- t[794] = 0
      "0000" when "00001100011011", -- t[795] = 0
      "0000" when "00001100011100", -- t[796] = 0
      "0000" when "00001100011101", -- t[797] = 0
      "0000" when "00001100011110", -- t[798] = 0
      "0000" when "00001100011111", -- t[799] = 0
      "0000" when "00001100100000", -- t[800] = 0
      "0000" when "00001100100001", -- t[801] = 0
      "0000" when "00001100100010", -- t[802] = 0
      "0000" when "00001100100011", -- t[803] = 0
      "0000" when "00001100100100", -- t[804] = 0
      "0000" when "00001100100101", -- t[805] = 0
      "0000" when "00001100100110", -- t[806] = 0
      "0000" when "00001100100111", -- t[807] = 0
      "0000" when "00001100101000", -- t[808] = 0
      "0000" when "00001100101001", -- t[809] = 0
      "0000" when "00001100101010", -- t[810] = 0
      "0000" when "00001100101011", -- t[811] = 0
      "0000" when "00001100101100", -- t[812] = 0
      "0000" when "00001100101101", -- t[813] = 0
      "0000" when "00001100101110", -- t[814] = 0
      "0000" when "00001100101111", -- t[815] = 0
      "0000" when "00001100110000", -- t[816] = 0
      "0000" when "00001100110001", -- t[817] = 0
      "0000" when "00001100110010", -- t[818] = 0
      "0000" when "00001100110011", -- t[819] = 0
      "0000" when "00001100110100", -- t[820] = 0
      "0000" when "00001100110101", -- t[821] = 0
      "0000" when "00001100110110", -- t[822] = 0
      "0000" when "00001100110111", -- t[823] = 0
      "0000" when "00001100111000", -- t[824] = 0
      "0000" when "00001100111001", -- t[825] = 0
      "0000" when "00001100111010", -- t[826] = 0
      "0000" when "00001100111011", -- t[827] = 0
      "0000" when "00001100111100", -- t[828] = 0
      "0000" when "00001100111101", -- t[829] = 0
      "0000" when "00001100111110", -- t[830] = 0
      "0000" when "00001100111111", -- t[831] = 0
      "0000" when "00001101000000", -- t[832] = 0
      "0000" when "00001101000001", -- t[833] = 0
      "0000" when "00001101000010", -- t[834] = 0
      "0000" when "00001101000011", -- t[835] = 0
      "0000" when "00001101000100", -- t[836] = 0
      "0000" when "00001101000101", -- t[837] = 0
      "0000" when "00001101000110", -- t[838] = 0
      "0000" when "00001101000111", -- t[839] = 0
      "0000" when "00001101001000", -- t[840] = 0
      "0000" when "00001101001001", -- t[841] = 0
      "0000" when "00001101001010", -- t[842] = 0
      "0000" when "00001101001011", -- t[843] = 0
      "0000" when "00001101001100", -- t[844] = 0
      "0000" when "00001101001101", -- t[845] = 0
      "0000" when "00001101001110", -- t[846] = 0
      "0000" when "00001101001111", -- t[847] = 0
      "0000" when "00001101010000", -- t[848] = 0
      "0000" when "00001101010001", -- t[849] = 0
      "0000" when "00001101010010", -- t[850] = 0
      "0000" when "00001101010011", -- t[851] = 0
      "0000" when "00001101010100", -- t[852] = 0
      "0000" when "00001101010101", -- t[853] = 0
      "0000" when "00001101010110", -- t[854] = 0
      "0000" when "00001101010111", -- t[855] = 0
      "0000" when "00001101011000", -- t[856] = 0
      "0000" when "00001101011001", -- t[857] = 0
      "0000" when "00001101011010", -- t[858] = 0
      "0000" when "00001101011011", -- t[859] = 0
      "0000" when "00001101011100", -- t[860] = 0
      "0000" when "00001101011101", -- t[861] = 0
      "0000" when "00001101011110", -- t[862] = 0
      "0000" when "00001101011111", -- t[863] = 0
      "0000" when "00001101100000", -- t[864] = 0
      "0000" when "00001101100001", -- t[865] = 0
      "0000" when "00001101100010", -- t[866] = 0
      "0000" when "00001101100011", -- t[867] = 0
      "0000" when "00001101100100", -- t[868] = 0
      "0000" when "00001101100101", -- t[869] = 0
      "0000" when "00001101100110", -- t[870] = 0
      "0000" when "00001101100111", -- t[871] = 0
      "0000" when "00001101101000", -- t[872] = 0
      "0000" when "00001101101001", -- t[873] = 0
      "0000" when "00001101101010", -- t[874] = 0
      "0000" when "00001101101011", -- t[875] = 0
      "0000" when "00001101101100", -- t[876] = 0
      "0000" when "00001101101101", -- t[877] = 0
      "0000" when "00001101101110", -- t[878] = 0
      "0000" when "00001101101111", -- t[879] = 0
      "0000" when "00001101110000", -- t[880] = 0
      "0000" when "00001101110001", -- t[881] = 0
      "0000" when "00001101110010", -- t[882] = 0
      "0000" when "00001101110011", -- t[883] = 0
      "0000" when "00001101110100", -- t[884] = 0
      "0000" when "00001101110101", -- t[885] = 0
      "0000" when "00001101110110", -- t[886] = 0
      "0000" when "00001101110111", -- t[887] = 0
      "0000" when "00001101111000", -- t[888] = 0
      "0000" when "00001101111001", -- t[889] = 0
      "0000" when "00001101111010", -- t[890] = 0
      "0000" when "00001101111011", -- t[891] = 0
      "0000" when "00001101111100", -- t[892] = 0
      "0000" when "00001101111101", -- t[893] = 0
      "0000" when "00001101111110", -- t[894] = 0
      "0000" when "00001101111111", -- t[895] = 0
      "0000" when "00001110000000", -- t[896] = 0
      "0000" when "00001110000001", -- t[897] = 0
      "0000" when "00001110000010", -- t[898] = 0
      "0000" when "00001110000011", -- t[899] = 0
      "0000" when "00001110000100", -- t[900] = 0
      "0000" when "00001110000101", -- t[901] = 0
      "0000" when "00001110000110", -- t[902] = 0
      "0000" when "00001110000111", -- t[903] = 0
      "0000" when "00001110001000", -- t[904] = 0
      "0000" when "00001110001001", -- t[905] = 0
      "0000" when "00001110001010", -- t[906] = 0
      "0000" when "00001110001011", -- t[907] = 0
      "0000" when "00001110001100", -- t[908] = 0
      "0000" when "00001110001101", -- t[909] = 0
      "0000" when "00001110001110", -- t[910] = 0
      "0000" when "00001110001111", -- t[911] = 0
      "0000" when "00001110010000", -- t[912] = 0
      "0000" when "00001110010001", -- t[913] = 0
      "0000" when "00001110010010", -- t[914] = 0
      "0000" when "00001110010011", -- t[915] = 0
      "0000" when "00001110010100", -- t[916] = 0
      "0000" when "00001110010101", -- t[917] = 0
      "0000" when "00001110010110", -- t[918] = 0
      "0000" when "00001110010111", -- t[919] = 0
      "0000" when "00001110011000", -- t[920] = 0
      "0000" when "00001110011001", -- t[921] = 0
      "0000" when "00001110011010", -- t[922] = 0
      "0000" when "00001110011011", -- t[923] = 0
      "0000" when "00001110011100", -- t[924] = 0
      "0000" when "00001110011101", -- t[925] = 0
      "0000" when "00001110011110", -- t[926] = 0
      "0000" when "00001110011111", -- t[927] = 0
      "0000" when "00001110100000", -- t[928] = 0
      "0000" when "00001110100001", -- t[929] = 0
      "0000" when "00001110100010", -- t[930] = 0
      "0000" when "00001110100011", -- t[931] = 0
      "0000" when "00001110100100", -- t[932] = 0
      "0000" when "00001110100101", -- t[933] = 0
      "0000" when "00001110100110", -- t[934] = 0
      "0000" when "00001110100111", -- t[935] = 0
      "0000" when "00001110101000", -- t[936] = 0
      "0000" when "00001110101001", -- t[937] = 0
      "0000" when "00001110101010", -- t[938] = 0
      "0000" when "00001110101011", -- t[939] = 0
      "0000" when "00001110101100", -- t[940] = 0
      "0000" when "00001110101101", -- t[941] = 0
      "0000" when "00001110101110", -- t[942] = 0
      "0000" when "00001110101111", -- t[943] = 0
      "0000" when "00001110110000", -- t[944] = 0
      "0000" when "00001110110001", -- t[945] = 0
      "0000" when "00001110110010", -- t[946] = 0
      "0000" when "00001110110011", -- t[947] = 0
      "0000" when "00001110110100", -- t[948] = 0
      "0000" when "00001110110101", -- t[949] = 0
      "0000" when "00001110110110", -- t[950] = 0
      "0000" when "00001110110111", -- t[951] = 0
      "0000" when "00001110111000", -- t[952] = 0
      "0000" when "00001110111001", -- t[953] = 0
      "0000" when "00001110111010", -- t[954] = 0
      "0000" when "00001110111011", -- t[955] = 0
      "0000" when "00001110111100", -- t[956] = 0
      "0000" when "00001110111101", -- t[957] = 0
      "0000" when "00001110111110", -- t[958] = 0
      "0000" when "00001110111111", -- t[959] = 0
      "0000" when "00001111000000", -- t[960] = 0
      "0000" when "00001111000001", -- t[961] = 0
      "0000" when "00001111000010", -- t[962] = 0
      "0000" when "00001111000011", -- t[963] = 0
      "0000" when "00001111000100", -- t[964] = 0
      "0000" when "00001111000101", -- t[965] = 0
      "0000" when "00001111000110", -- t[966] = 0
      "0000" when "00001111000111", -- t[967] = 0
      "0000" when "00001111001000", -- t[968] = 0
      "0000" when "00001111001001", -- t[969] = 0
      "0000" when "00001111001010", -- t[970] = 0
      "0000" when "00001111001011", -- t[971] = 0
      "0000" when "00001111001100", -- t[972] = 0
      "0000" when "00001111001101", -- t[973] = 0
      "0000" when "00001111001110", -- t[974] = 0
      "0000" when "00001111001111", -- t[975] = 0
      "0000" when "00001111010000", -- t[976] = 0
      "0000" when "00001111010001", -- t[977] = 0
      "0000" when "00001111010010", -- t[978] = 0
      "0000" when "00001111010011", -- t[979] = 0
      "0000" when "00001111010100", -- t[980] = 0
      "0000" when "00001111010101", -- t[981] = 0
      "0000" when "00001111010110", -- t[982] = 0
      "0000" when "00001111010111", -- t[983] = 0
      "0000" when "00001111011000", -- t[984] = 0
      "0000" when "00001111011001", -- t[985] = 0
      "0000" when "00001111011010", -- t[986] = 0
      "0000" when "00001111011011", -- t[987] = 0
      "0000" when "00001111011100", -- t[988] = 0
      "0000" when "00001111011101", -- t[989] = 0
      "0000" when "00001111011110", -- t[990] = 0
      "0000" when "00001111011111", -- t[991] = 0
      "0000" when "00001111100000", -- t[992] = 0
      "0000" when "00001111100001", -- t[993] = 0
      "0000" when "00001111100010", -- t[994] = 0
      "0000" when "00001111100011", -- t[995] = 0
      "0000" when "00001111100100", -- t[996] = 0
      "0000" when "00001111100101", -- t[997] = 0
      "0000" when "00001111100110", -- t[998] = 0
      "0000" when "00001111100111", -- t[999] = 0
      "0000" when "00001111101000", -- t[1000] = 0
      "0000" when "00001111101001", -- t[1001] = 0
      "0000" when "00001111101010", -- t[1002] = 0
      "0000" when "00001111101011", -- t[1003] = 0
      "0000" when "00001111101100", -- t[1004] = 0
      "0000" when "00001111101101", -- t[1005] = 0
      "0000" when "00001111101110", -- t[1006] = 0
      "0000" when "00001111101111", -- t[1007] = 0
      "0000" when "00001111110000", -- t[1008] = 0
      "0000" when "00001111110001", -- t[1009] = 0
      "0000" when "00001111110010", -- t[1010] = 0
      "0000" when "00001111110011", -- t[1011] = 0
      "0000" when "00001111110100", -- t[1012] = 0
      "0000" when "00001111110101", -- t[1013] = 0
      "0000" when "00001111110110", -- t[1014] = 0
      "0000" when "00001111110111", -- t[1015] = 0
      "0000" when "00001111111000", -- t[1016] = 0
      "0000" when "00001111111001", -- t[1017] = 0
      "0000" when "00001111111010", -- t[1018] = 0
      "0000" when "00001111111011", -- t[1019] = 0
      "0000" when "00001111111100", -- t[1020] = 0
      "0000" when "00001111111101", -- t[1021] = 0
      "0000" when "00001111111110", -- t[1022] = 0
      "0000" when "00001111111111", -- t[1023] = 0
      "0000" when "00010000000000", -- t[1024] = 0
      "0000" when "00010000000001", -- t[1025] = 0
      "0000" when "00010000000010", -- t[1026] = 0
      "0000" when "00010000000011", -- t[1027] = 0
      "0000" when "00010000000100", -- t[1028] = 0
      "0000" when "00010000000101", -- t[1029] = 0
      "0000" when "00010000000110", -- t[1030] = 0
      "0000" when "00010000000111", -- t[1031] = 0
      "0000" when "00010000001000", -- t[1032] = 0
      "0000" when "00010000001001", -- t[1033] = 0
      "0000" when "00010000001010", -- t[1034] = 0
      "0000" when "00010000001011", -- t[1035] = 0
      "0000" when "00010000001100", -- t[1036] = 0
      "0000" when "00010000001101", -- t[1037] = 0
      "0000" when "00010000001110", -- t[1038] = 0
      "0000" when "00010000001111", -- t[1039] = 0
      "0000" when "00010000010000", -- t[1040] = 0
      "0000" when "00010000010001", -- t[1041] = 0
      "0000" when "00010000010010", -- t[1042] = 0
      "0000" when "00010000010011", -- t[1043] = 0
      "0000" when "00010000010100", -- t[1044] = 0
      "0000" when "00010000010101", -- t[1045] = 0
      "0000" when "00010000010110", -- t[1046] = 0
      "0000" when "00010000010111", -- t[1047] = 0
      "0000" when "00010000011000", -- t[1048] = 0
      "0000" when "00010000011001", -- t[1049] = 0
      "0000" when "00010000011010", -- t[1050] = 0
      "0000" when "00010000011011", -- t[1051] = 0
      "0000" when "00010000011100", -- t[1052] = 0
      "0000" when "00010000011101", -- t[1053] = 0
      "0000" when "00010000011110", -- t[1054] = 0
      "0000" when "00010000011111", -- t[1055] = 0
      "0000" when "00010000100000", -- t[1056] = 0
      "0000" when "00010000100001", -- t[1057] = 0
      "0000" when "00010000100010", -- t[1058] = 0
      "0000" when "00010000100011", -- t[1059] = 0
      "0000" when "00010000100100", -- t[1060] = 0
      "0000" when "00010000100101", -- t[1061] = 0
      "0000" when "00010000100110", -- t[1062] = 0
      "0000" when "00010000100111", -- t[1063] = 0
      "0000" when "00010000101000", -- t[1064] = 0
      "0000" when "00010000101001", -- t[1065] = 0
      "0000" when "00010000101010", -- t[1066] = 0
      "0000" when "00010000101011", -- t[1067] = 0
      "0000" when "00010000101100", -- t[1068] = 0
      "0000" when "00010000101101", -- t[1069] = 0
      "0000" when "00010000101110", -- t[1070] = 0
      "0000" when "00010000101111", -- t[1071] = 0
      "0000" when "00010000110000", -- t[1072] = 0
      "0000" when "00010000110001", -- t[1073] = 0
      "0000" when "00010000110010", -- t[1074] = 0
      "0000" when "00010000110011", -- t[1075] = 0
      "0000" when "00010000110100", -- t[1076] = 0
      "0000" when "00010000110101", -- t[1077] = 0
      "0000" when "00010000110110", -- t[1078] = 0
      "0000" when "00010000110111", -- t[1079] = 0
      "0000" when "00010000111000", -- t[1080] = 0
      "0000" when "00010000111001", -- t[1081] = 0
      "0000" when "00010000111010", -- t[1082] = 0
      "0000" when "00010000111011", -- t[1083] = 0
      "0000" when "00010000111100", -- t[1084] = 0
      "0000" when "00010000111101", -- t[1085] = 0
      "0000" when "00010000111110", -- t[1086] = 0
      "0000" when "00010000111111", -- t[1087] = 0
      "0000" when "00010001000000", -- t[1088] = 0
      "0000" when "00010001000001", -- t[1089] = 0
      "0000" when "00010001000010", -- t[1090] = 0
      "0000" when "00010001000011", -- t[1091] = 0
      "0000" when "00010001000100", -- t[1092] = 0
      "0000" when "00010001000101", -- t[1093] = 0
      "0000" when "00010001000110", -- t[1094] = 0
      "0000" when "00010001000111", -- t[1095] = 0
      "0000" when "00010001001000", -- t[1096] = 0
      "0000" when "00010001001001", -- t[1097] = 0
      "0000" when "00010001001010", -- t[1098] = 0
      "0000" when "00010001001011", -- t[1099] = 0
      "0000" when "00010001001100", -- t[1100] = 0
      "0000" when "00010001001101", -- t[1101] = 0
      "0000" when "00010001001110", -- t[1102] = 0
      "0000" when "00010001001111", -- t[1103] = 0
      "0000" when "00010001010000", -- t[1104] = 0
      "0000" when "00010001010001", -- t[1105] = 0
      "0000" when "00010001010010", -- t[1106] = 0
      "0000" when "00010001010011", -- t[1107] = 0
      "0000" when "00010001010100", -- t[1108] = 0
      "0000" when "00010001010101", -- t[1109] = 0
      "0000" when "00010001010110", -- t[1110] = 0
      "0000" when "00010001010111", -- t[1111] = 0
      "0000" when "00010001011000", -- t[1112] = 0
      "0000" when "00010001011001", -- t[1113] = 0
      "0000" when "00010001011010", -- t[1114] = 0
      "0000" when "00010001011011", -- t[1115] = 0
      "0000" when "00010001011100", -- t[1116] = 0
      "0000" when "00010001011101", -- t[1117] = 0
      "0000" when "00010001011110", -- t[1118] = 0
      "0000" when "00010001011111", -- t[1119] = 0
      "0000" when "00010001100000", -- t[1120] = 0
      "0000" when "00010001100001", -- t[1121] = 0
      "0000" when "00010001100010", -- t[1122] = 0
      "0000" when "00010001100011", -- t[1123] = 0
      "0000" when "00010001100100", -- t[1124] = 0
      "0000" when "00010001100101", -- t[1125] = 0
      "0000" when "00010001100110", -- t[1126] = 0
      "0000" when "00010001100111", -- t[1127] = 0
      "0000" when "00010001101000", -- t[1128] = 0
      "0000" when "00010001101001", -- t[1129] = 0
      "0000" when "00010001101010", -- t[1130] = 0
      "0000" when "00010001101011", -- t[1131] = 0
      "0000" when "00010001101100", -- t[1132] = 0
      "0000" when "00010001101101", -- t[1133] = 0
      "0000" when "00010001101110", -- t[1134] = 0
      "0000" when "00010001101111", -- t[1135] = 0
      "0000" when "00010001110000", -- t[1136] = 0
      "0000" when "00010001110001", -- t[1137] = 0
      "0000" when "00010001110010", -- t[1138] = 0
      "0000" when "00010001110011", -- t[1139] = 0
      "0000" when "00010001110100", -- t[1140] = 0
      "0000" when "00010001110101", -- t[1141] = 0
      "0000" when "00010001110110", -- t[1142] = 0
      "0000" when "00010001110111", -- t[1143] = 0
      "0000" when "00010001111000", -- t[1144] = 0
      "0000" when "00010001111001", -- t[1145] = 0
      "0000" when "00010001111010", -- t[1146] = 0
      "0000" when "00010001111011", -- t[1147] = 0
      "0000" when "00010001111100", -- t[1148] = 0
      "0000" when "00010001111101", -- t[1149] = 0
      "0000" when "00010001111110", -- t[1150] = 0
      "0000" when "00010001111111", -- t[1151] = 0
      "0000" when "00010010000000", -- t[1152] = 0
      "0000" when "00010010000001", -- t[1153] = 0
      "0000" when "00010010000010", -- t[1154] = 0
      "0000" when "00010010000011", -- t[1155] = 0
      "0000" when "00010010000100", -- t[1156] = 0
      "0000" when "00010010000101", -- t[1157] = 0
      "0000" when "00010010000110", -- t[1158] = 0
      "0000" when "00010010000111", -- t[1159] = 0
      "0000" when "00010010001000", -- t[1160] = 0
      "0000" when "00010010001001", -- t[1161] = 0
      "0000" when "00010010001010", -- t[1162] = 0
      "0000" when "00010010001011", -- t[1163] = 0
      "0000" when "00010010001100", -- t[1164] = 0
      "0000" when "00010010001101", -- t[1165] = 0
      "0000" when "00010010001110", -- t[1166] = 0
      "0000" when "00010010001111", -- t[1167] = 0
      "0000" when "00010010010000", -- t[1168] = 0
      "0000" when "00010010010001", -- t[1169] = 0
      "0000" when "00010010010010", -- t[1170] = 0
      "0000" when "00010010010011", -- t[1171] = 0
      "0000" when "00010010010100", -- t[1172] = 0
      "0000" when "00010010010101", -- t[1173] = 0
      "0000" when "00010010010110", -- t[1174] = 0
      "0000" when "00010010010111", -- t[1175] = 0
      "0000" when "00010010011000", -- t[1176] = 0
      "0000" when "00010010011001", -- t[1177] = 0
      "0000" when "00010010011010", -- t[1178] = 0
      "0000" when "00010010011011", -- t[1179] = 0
      "0000" when "00010010011100", -- t[1180] = 0
      "0000" when "00010010011101", -- t[1181] = 0
      "0000" when "00010010011110", -- t[1182] = 0
      "0000" when "00010010011111", -- t[1183] = 0
      "0000" when "00010010100000", -- t[1184] = 0
      "0000" when "00010010100001", -- t[1185] = 0
      "0000" when "00010010100010", -- t[1186] = 0
      "0000" when "00010010100011", -- t[1187] = 0
      "0000" when "00010010100100", -- t[1188] = 0
      "0000" when "00010010100101", -- t[1189] = 0
      "0000" when "00010010100110", -- t[1190] = 0
      "0000" when "00010010100111", -- t[1191] = 0
      "0000" when "00010010101000", -- t[1192] = 0
      "0000" when "00010010101001", -- t[1193] = 0
      "0000" when "00010010101010", -- t[1194] = 0
      "0000" when "00010010101011", -- t[1195] = 0
      "0000" when "00010010101100", -- t[1196] = 0
      "0000" when "00010010101101", -- t[1197] = 0
      "0000" when "00010010101110", -- t[1198] = 0
      "0000" when "00010010101111", -- t[1199] = 0
      "0000" when "00010010110000", -- t[1200] = 0
      "0000" when "00010010110001", -- t[1201] = 0
      "0000" when "00010010110010", -- t[1202] = 0
      "0000" when "00010010110011", -- t[1203] = 0
      "0000" when "00010010110100", -- t[1204] = 0
      "0000" when "00010010110101", -- t[1205] = 0
      "0000" when "00010010110110", -- t[1206] = 0
      "0000" when "00010010110111", -- t[1207] = 0
      "0000" when "00010010111000", -- t[1208] = 0
      "0000" when "00010010111001", -- t[1209] = 0
      "0000" when "00010010111010", -- t[1210] = 0
      "0000" when "00010010111011", -- t[1211] = 0
      "0000" when "00010010111100", -- t[1212] = 0
      "0000" when "00010010111101", -- t[1213] = 0
      "0000" when "00010010111110", -- t[1214] = 0
      "0000" when "00010010111111", -- t[1215] = 0
      "0000" when "00010011000000", -- t[1216] = 0
      "0000" when "00010011000001", -- t[1217] = 0
      "0000" when "00010011000010", -- t[1218] = 0
      "0000" when "00010011000011", -- t[1219] = 0
      "0000" when "00010011000100", -- t[1220] = 0
      "0000" when "00010011000101", -- t[1221] = 0
      "0000" when "00010011000110", -- t[1222] = 0
      "0000" when "00010011000111", -- t[1223] = 0
      "0000" when "00010011001000", -- t[1224] = 0
      "0000" when "00010011001001", -- t[1225] = 0
      "0000" when "00010011001010", -- t[1226] = 0
      "0000" when "00010011001011", -- t[1227] = 0
      "0000" when "00010011001100", -- t[1228] = 0
      "0000" when "00010011001101", -- t[1229] = 0
      "0000" when "00010011001110", -- t[1230] = 0
      "0000" when "00010011001111", -- t[1231] = 0
      "0000" when "00010011010000", -- t[1232] = 0
      "0000" when "00010011010001", -- t[1233] = 0
      "0000" when "00010011010010", -- t[1234] = 0
      "0000" when "00010011010011", -- t[1235] = 0
      "0000" when "00010011010100", -- t[1236] = 0
      "0000" when "00010011010101", -- t[1237] = 0
      "0000" when "00010011010110", -- t[1238] = 0
      "0000" when "00010011010111", -- t[1239] = 0
      "0000" when "00010011011000", -- t[1240] = 0
      "0000" when "00010011011001", -- t[1241] = 0
      "0000" when "00010011011010", -- t[1242] = 0
      "0000" when "00010011011011", -- t[1243] = 0
      "0000" when "00010011011100", -- t[1244] = 0
      "0000" when "00010011011101", -- t[1245] = 0
      "0000" when "00010011011110", -- t[1246] = 0
      "0000" when "00010011011111", -- t[1247] = 0
      "0000" when "00010011100000", -- t[1248] = 0
      "0000" when "00010011100001", -- t[1249] = 0
      "0000" when "00010011100010", -- t[1250] = 0
      "0000" when "00010011100011", -- t[1251] = 0
      "0000" when "00010011100100", -- t[1252] = 0
      "0000" when "00010011100101", -- t[1253] = 0
      "0000" when "00010011100110", -- t[1254] = 0
      "0000" when "00010011100111", -- t[1255] = 0
      "0000" when "00010011101000", -- t[1256] = 0
      "0000" when "00010011101001", -- t[1257] = 0
      "0000" when "00010011101010", -- t[1258] = 0
      "0000" when "00010011101011", -- t[1259] = 0
      "0000" when "00010011101100", -- t[1260] = 0
      "0000" when "00010011101101", -- t[1261] = 0
      "0000" when "00010011101110", -- t[1262] = 0
      "0000" when "00010011101111", -- t[1263] = 0
      "0000" when "00010011110000", -- t[1264] = 0
      "0000" when "00010011110001", -- t[1265] = 0
      "0000" when "00010011110010", -- t[1266] = 0
      "0000" when "00010011110011", -- t[1267] = 0
      "0000" when "00010011110100", -- t[1268] = 0
      "0000" when "00010011110101", -- t[1269] = 0
      "0000" when "00010011110110", -- t[1270] = 0
      "0000" when "00010011110111", -- t[1271] = 0
      "0000" when "00010011111000", -- t[1272] = 0
      "0000" when "00010011111001", -- t[1273] = 0
      "0000" when "00010011111010", -- t[1274] = 0
      "0000" when "00010011111011", -- t[1275] = 0
      "0000" when "00010011111100", -- t[1276] = 0
      "0000" when "00010011111101", -- t[1277] = 0
      "0000" when "00010011111110", -- t[1278] = 0
      "0000" when "00010011111111", -- t[1279] = 0
      "0000" when "00010100000000", -- t[1280] = 0
      "0000" when "00010100000001", -- t[1281] = 0
      "0000" when "00010100000010", -- t[1282] = 0
      "0000" when "00010100000011", -- t[1283] = 0
      "0000" when "00010100000100", -- t[1284] = 0
      "0000" when "00010100000101", -- t[1285] = 0
      "0000" when "00010100000110", -- t[1286] = 0
      "0000" when "00010100000111", -- t[1287] = 0
      "0000" when "00010100001000", -- t[1288] = 0
      "0000" when "00010100001001", -- t[1289] = 0
      "0000" when "00010100001010", -- t[1290] = 0
      "0000" when "00010100001011", -- t[1291] = 0
      "0000" when "00010100001100", -- t[1292] = 0
      "0000" when "00010100001101", -- t[1293] = 0
      "0000" when "00010100001110", -- t[1294] = 0
      "0000" when "00010100001111", -- t[1295] = 0
      "0000" when "00010100010000", -- t[1296] = 0
      "0000" when "00010100010001", -- t[1297] = 0
      "0000" when "00010100010010", -- t[1298] = 0
      "0000" when "00010100010011", -- t[1299] = 0
      "0000" when "00010100010100", -- t[1300] = 0
      "0000" when "00010100010101", -- t[1301] = 0
      "0000" when "00010100010110", -- t[1302] = 0
      "0000" when "00010100010111", -- t[1303] = 0
      "0000" when "00010100011000", -- t[1304] = 0
      "0000" when "00010100011001", -- t[1305] = 0
      "0000" when "00010100011010", -- t[1306] = 0
      "0000" when "00010100011011", -- t[1307] = 0
      "0000" when "00010100011100", -- t[1308] = 0
      "0000" when "00010100011101", -- t[1309] = 0
      "0000" when "00010100011110", -- t[1310] = 0
      "0000" when "00010100011111", -- t[1311] = 0
      "0000" when "00010100100000", -- t[1312] = 0
      "0000" when "00010100100001", -- t[1313] = 0
      "0000" when "00010100100010", -- t[1314] = 0
      "0000" when "00010100100011", -- t[1315] = 0
      "0000" when "00010100100100", -- t[1316] = 0
      "0000" when "00010100100101", -- t[1317] = 0
      "0000" when "00010100100110", -- t[1318] = 0
      "0000" when "00010100100111", -- t[1319] = 0
      "0000" when "00010100101000", -- t[1320] = 0
      "0000" when "00010100101001", -- t[1321] = 0
      "0000" when "00010100101010", -- t[1322] = 0
      "0000" when "00010100101011", -- t[1323] = 0
      "0000" when "00010100101100", -- t[1324] = 0
      "0000" when "00010100101101", -- t[1325] = 0
      "0000" when "00010100101110", -- t[1326] = 0
      "0000" when "00010100101111", -- t[1327] = 0
      "0000" when "00010100110000", -- t[1328] = 0
      "0000" when "00010100110001", -- t[1329] = 0
      "0000" when "00010100110010", -- t[1330] = 0
      "0000" when "00010100110011", -- t[1331] = 0
      "0000" when "00010100110100", -- t[1332] = 0
      "0000" when "00010100110101", -- t[1333] = 0
      "0000" when "00010100110110", -- t[1334] = 0
      "0000" when "00010100110111", -- t[1335] = 0
      "0000" when "00010100111000", -- t[1336] = 0
      "0000" when "00010100111001", -- t[1337] = 0
      "0000" when "00010100111010", -- t[1338] = 0
      "0000" when "00010100111011", -- t[1339] = 0
      "0000" when "00010100111100", -- t[1340] = 0
      "0000" when "00010100111101", -- t[1341] = 0
      "0000" when "00010100111110", -- t[1342] = 0
      "0000" when "00010100111111", -- t[1343] = 0
      "0000" when "00010101000000", -- t[1344] = 0
      "0000" when "00010101000001", -- t[1345] = 0
      "0000" when "00010101000010", -- t[1346] = 0
      "0000" when "00010101000011", -- t[1347] = 0
      "0000" when "00010101000100", -- t[1348] = 0
      "0000" when "00010101000101", -- t[1349] = 0
      "0000" when "00010101000110", -- t[1350] = 0
      "0000" when "00010101000111", -- t[1351] = 0
      "0000" when "00010101001000", -- t[1352] = 0
      "0000" when "00010101001001", -- t[1353] = 0
      "0000" when "00010101001010", -- t[1354] = 0
      "0000" when "00010101001011", -- t[1355] = 0
      "0000" when "00010101001100", -- t[1356] = 0
      "0000" when "00010101001101", -- t[1357] = 0
      "0000" when "00010101001110", -- t[1358] = 0
      "0000" when "00010101001111", -- t[1359] = 0
      "0000" when "00010101010000", -- t[1360] = 0
      "0000" when "00010101010001", -- t[1361] = 0
      "0000" when "00010101010010", -- t[1362] = 0
      "0000" when "00010101010011", -- t[1363] = 0
      "0000" when "00010101010100", -- t[1364] = 0
      "0000" when "00010101010101", -- t[1365] = 0
      "0000" when "00010101010110", -- t[1366] = 0
      "0000" when "00010101010111", -- t[1367] = 0
      "0000" when "00010101011000", -- t[1368] = 0
      "0000" when "00010101011001", -- t[1369] = 0
      "0000" when "00010101011010", -- t[1370] = 0
      "0000" when "00010101011011", -- t[1371] = 0
      "0000" when "00010101011100", -- t[1372] = 0
      "0000" when "00010101011101", -- t[1373] = 0
      "0000" when "00010101011110", -- t[1374] = 0
      "0000" when "00010101011111", -- t[1375] = 0
      "0000" when "00010101100000", -- t[1376] = 0
      "0000" when "00010101100001", -- t[1377] = 0
      "0000" when "00010101100010", -- t[1378] = 0
      "0000" when "00010101100011", -- t[1379] = 0
      "0000" when "00010101100100", -- t[1380] = 0
      "0000" when "00010101100101", -- t[1381] = 0
      "0000" when "00010101100110", -- t[1382] = 0
      "0000" when "00010101100111", -- t[1383] = 0
      "0000" when "00010101101000", -- t[1384] = 0
      "0000" when "00010101101001", -- t[1385] = 0
      "0000" when "00010101101010", -- t[1386] = 0
      "0000" when "00010101101011", -- t[1387] = 0
      "0000" when "00010101101100", -- t[1388] = 0
      "0000" when "00010101101101", -- t[1389] = 0
      "0000" when "00010101101110", -- t[1390] = 0
      "0000" when "00010101101111", -- t[1391] = 0
      "0000" when "00010101110000", -- t[1392] = 0
      "0000" when "00010101110001", -- t[1393] = 0
      "0000" when "00010101110010", -- t[1394] = 0
      "0000" when "00010101110011", -- t[1395] = 0
      "0000" when "00010101110100", -- t[1396] = 0
      "0000" when "00010101110101", -- t[1397] = 0
      "0000" when "00010101110110", -- t[1398] = 0
      "0000" when "00010101110111", -- t[1399] = 0
      "0000" when "00010101111000", -- t[1400] = 0
      "0000" when "00010101111001", -- t[1401] = 0
      "0000" when "00010101111010", -- t[1402] = 0
      "0000" when "00010101111011", -- t[1403] = 0
      "0000" when "00010101111100", -- t[1404] = 0
      "0000" when "00010101111101", -- t[1405] = 0
      "0000" when "00010101111110", -- t[1406] = 0
      "0000" when "00010101111111", -- t[1407] = 0
      "0000" when "00010110000000", -- t[1408] = 0
      "0000" when "00010110000001", -- t[1409] = 0
      "0000" when "00010110000010", -- t[1410] = 0
      "0000" when "00010110000011", -- t[1411] = 0
      "0000" when "00010110000100", -- t[1412] = 0
      "0000" when "00010110000101", -- t[1413] = 0
      "0000" when "00010110000110", -- t[1414] = 0
      "0000" when "00010110000111", -- t[1415] = 0
      "0000" when "00010110001000", -- t[1416] = 0
      "0000" when "00010110001001", -- t[1417] = 0
      "0000" when "00010110001010", -- t[1418] = 0
      "0000" when "00010110001011", -- t[1419] = 0
      "0000" when "00010110001100", -- t[1420] = 0
      "0000" when "00010110001101", -- t[1421] = 0
      "0000" when "00010110001110", -- t[1422] = 0
      "0000" when "00010110001111", -- t[1423] = 0
      "0000" when "00010110010000", -- t[1424] = 0
      "0000" when "00010110010001", -- t[1425] = 0
      "0000" when "00010110010010", -- t[1426] = 0
      "0000" when "00010110010011", -- t[1427] = 0
      "0000" when "00010110010100", -- t[1428] = 0
      "0000" when "00010110010101", -- t[1429] = 0
      "0000" when "00010110010110", -- t[1430] = 0
      "0000" when "00010110010111", -- t[1431] = 0
      "0000" when "00010110011000", -- t[1432] = 0
      "0000" when "00010110011001", -- t[1433] = 0
      "0000" when "00010110011010", -- t[1434] = 0
      "0000" when "00010110011011", -- t[1435] = 0
      "0000" when "00010110011100", -- t[1436] = 0
      "0000" when "00010110011101", -- t[1437] = 0
      "0000" when "00010110011110", -- t[1438] = 0
      "0000" when "00010110011111", -- t[1439] = 0
      "0000" when "00010110100000", -- t[1440] = 0
      "0000" when "00010110100001", -- t[1441] = 0
      "0000" when "00010110100010", -- t[1442] = 0
      "0000" when "00010110100011", -- t[1443] = 0
      "0000" when "00010110100100", -- t[1444] = 0
      "0000" when "00010110100101", -- t[1445] = 0
      "0000" when "00010110100110", -- t[1446] = 0
      "0000" when "00010110100111", -- t[1447] = 0
      "0000" when "00010110101000", -- t[1448] = 0
      "0000" when "00010110101001", -- t[1449] = 0
      "0000" when "00010110101010", -- t[1450] = 0
      "0000" when "00010110101011", -- t[1451] = 0
      "0000" when "00010110101100", -- t[1452] = 0
      "0000" when "00010110101101", -- t[1453] = 0
      "0000" when "00010110101110", -- t[1454] = 0
      "0000" when "00010110101111", -- t[1455] = 0
      "0000" when "00010110110000", -- t[1456] = 0
      "0000" when "00010110110001", -- t[1457] = 0
      "0000" when "00010110110010", -- t[1458] = 0
      "0000" when "00010110110011", -- t[1459] = 0
      "0000" when "00010110110100", -- t[1460] = 0
      "0000" when "00010110110101", -- t[1461] = 0
      "0000" when "00010110110110", -- t[1462] = 0
      "0000" when "00010110110111", -- t[1463] = 0
      "0000" when "00010110111000", -- t[1464] = 0
      "0000" when "00010110111001", -- t[1465] = 0
      "0000" when "00010110111010", -- t[1466] = 0
      "0000" when "00010110111011", -- t[1467] = 0
      "0000" when "00010110111100", -- t[1468] = 0
      "0000" when "00010110111101", -- t[1469] = 0
      "0000" when "00010110111110", -- t[1470] = 0
      "0000" when "00010110111111", -- t[1471] = 0
      "0000" when "00010111000000", -- t[1472] = 0
      "0000" when "00010111000001", -- t[1473] = 0
      "0000" when "00010111000010", -- t[1474] = 0
      "0000" when "00010111000011", -- t[1475] = 0
      "0000" when "00010111000100", -- t[1476] = 0
      "0000" when "00010111000101", -- t[1477] = 0
      "0000" when "00010111000110", -- t[1478] = 0
      "0000" when "00010111000111", -- t[1479] = 0
      "0000" when "00010111001000", -- t[1480] = 0
      "0000" when "00010111001001", -- t[1481] = 0
      "0000" when "00010111001010", -- t[1482] = 0
      "0000" when "00010111001011", -- t[1483] = 0
      "0000" when "00010111001100", -- t[1484] = 0
      "0000" when "00010111001101", -- t[1485] = 0
      "0000" when "00010111001110", -- t[1486] = 0
      "0000" when "00010111001111", -- t[1487] = 0
      "0000" when "00010111010000", -- t[1488] = 0
      "0000" when "00010111010001", -- t[1489] = 0
      "0000" when "00010111010010", -- t[1490] = 0
      "0000" when "00010111010011", -- t[1491] = 0
      "0000" when "00010111010100", -- t[1492] = 0
      "0000" when "00010111010101", -- t[1493] = 0
      "0000" when "00010111010110", -- t[1494] = 0
      "0000" when "00010111010111", -- t[1495] = 0
      "0000" when "00010111011000", -- t[1496] = 0
      "0000" when "00010111011001", -- t[1497] = 0
      "0000" when "00010111011010", -- t[1498] = 0
      "0000" when "00010111011011", -- t[1499] = 0
      "0000" when "00010111011100", -- t[1500] = 0
      "0000" when "00010111011101", -- t[1501] = 0
      "0000" when "00010111011110", -- t[1502] = 0
      "0000" when "00010111011111", -- t[1503] = 0
      "0000" when "00010111100000", -- t[1504] = 0
      "0000" when "00010111100001", -- t[1505] = 0
      "0000" when "00010111100010", -- t[1506] = 0
      "0000" when "00010111100011", -- t[1507] = 0
      "0000" when "00010111100100", -- t[1508] = 0
      "0000" when "00010111100101", -- t[1509] = 0
      "0000" when "00010111100110", -- t[1510] = 0
      "0000" when "00010111100111", -- t[1511] = 0
      "0000" when "00010111101000", -- t[1512] = 0
      "0000" when "00010111101001", -- t[1513] = 0
      "0000" when "00010111101010", -- t[1514] = 0
      "0000" when "00010111101011", -- t[1515] = 0
      "0000" when "00010111101100", -- t[1516] = 0
      "0000" when "00010111101101", -- t[1517] = 0
      "0000" when "00010111101110", -- t[1518] = 0
      "0000" when "00010111101111", -- t[1519] = 0
      "0000" when "00010111110000", -- t[1520] = 0
      "0000" when "00010111110001", -- t[1521] = 0
      "0000" when "00010111110010", -- t[1522] = 0
      "0000" when "00010111110011", -- t[1523] = 0
      "0000" when "00010111110100", -- t[1524] = 0
      "0000" when "00010111110101", -- t[1525] = 0
      "0000" when "00010111110110", -- t[1526] = 0
      "0000" when "00010111110111", -- t[1527] = 0
      "0000" when "00010111111000", -- t[1528] = 0
      "0000" when "00010111111001", -- t[1529] = 0
      "0000" when "00010111111010", -- t[1530] = 0
      "0000" when "00010111111011", -- t[1531] = 0
      "0000" when "00010111111100", -- t[1532] = 0
      "0000" when "00010111111101", -- t[1533] = 0
      "0000" when "00010111111110", -- t[1534] = 0
      "0000" when "00010111111111", -- t[1535] = 0
      "0000" when "00011000000000", -- t[1536] = 0
      "0000" when "00011000000001", -- t[1537] = 0
      "0000" when "00011000000010", -- t[1538] = 0
      "0000" when "00011000000011", -- t[1539] = 0
      "0000" when "00011000000100", -- t[1540] = 0
      "0000" when "00011000000101", -- t[1541] = 0
      "0000" when "00011000000110", -- t[1542] = 0
      "0000" when "00011000000111", -- t[1543] = 0
      "0000" when "00011000001000", -- t[1544] = 0
      "0000" when "00011000001001", -- t[1545] = 0
      "0000" when "00011000001010", -- t[1546] = 0
      "0000" when "00011000001011", -- t[1547] = 0
      "0000" when "00011000001100", -- t[1548] = 0
      "0000" when "00011000001101", -- t[1549] = 0
      "0000" when "00011000001110", -- t[1550] = 0
      "0000" when "00011000001111", -- t[1551] = 0
      "0000" when "00011000010000", -- t[1552] = 0
      "0000" when "00011000010001", -- t[1553] = 0
      "0000" when "00011000010010", -- t[1554] = 0
      "0000" when "00011000010011", -- t[1555] = 0
      "0000" when "00011000010100", -- t[1556] = 0
      "0000" when "00011000010101", -- t[1557] = 0
      "0000" when "00011000010110", -- t[1558] = 0
      "0000" when "00011000010111", -- t[1559] = 0
      "0000" when "00011000011000", -- t[1560] = 0
      "0000" when "00011000011001", -- t[1561] = 0
      "0000" when "00011000011010", -- t[1562] = 0
      "0000" when "00011000011011", -- t[1563] = 0
      "0000" when "00011000011100", -- t[1564] = 0
      "0000" when "00011000011101", -- t[1565] = 0
      "0000" when "00011000011110", -- t[1566] = 0
      "0000" when "00011000011111", -- t[1567] = 0
      "0000" when "00011000100000", -- t[1568] = 0
      "0000" when "00011000100001", -- t[1569] = 0
      "0000" when "00011000100010", -- t[1570] = 0
      "0000" when "00011000100011", -- t[1571] = 0
      "0000" when "00011000100100", -- t[1572] = 0
      "0000" when "00011000100101", -- t[1573] = 0
      "0000" when "00011000100110", -- t[1574] = 0
      "0000" when "00011000100111", -- t[1575] = 0
      "0000" when "00011000101000", -- t[1576] = 0
      "0000" when "00011000101001", -- t[1577] = 0
      "0000" when "00011000101010", -- t[1578] = 0
      "0000" when "00011000101011", -- t[1579] = 0
      "0000" when "00011000101100", -- t[1580] = 0
      "0000" when "00011000101101", -- t[1581] = 0
      "0000" when "00011000101110", -- t[1582] = 0
      "0000" when "00011000101111", -- t[1583] = 0
      "0000" when "00011000110000", -- t[1584] = 0
      "0000" when "00011000110001", -- t[1585] = 0
      "0000" when "00011000110010", -- t[1586] = 0
      "0000" when "00011000110011", -- t[1587] = 0
      "0000" when "00011000110100", -- t[1588] = 0
      "0000" when "00011000110101", -- t[1589] = 0
      "0000" when "00011000110110", -- t[1590] = 0
      "0000" when "00011000110111", -- t[1591] = 0
      "0000" when "00011000111000", -- t[1592] = 0
      "0000" when "00011000111001", -- t[1593] = 0
      "0000" when "00011000111010", -- t[1594] = 0
      "0000" when "00011000111011", -- t[1595] = 0
      "0000" when "00011000111100", -- t[1596] = 0
      "0000" when "00011000111101", -- t[1597] = 0
      "0000" when "00011000111110", -- t[1598] = 0
      "0000" when "00011000111111", -- t[1599] = 0
      "0000" when "00011001000000", -- t[1600] = 0
      "0000" when "00011001000001", -- t[1601] = 0
      "0000" when "00011001000010", -- t[1602] = 0
      "0000" when "00011001000011", -- t[1603] = 0
      "0000" when "00011001000100", -- t[1604] = 0
      "0000" when "00011001000101", -- t[1605] = 0
      "0000" when "00011001000110", -- t[1606] = 0
      "0000" when "00011001000111", -- t[1607] = 0
      "0000" when "00011001001000", -- t[1608] = 0
      "0000" when "00011001001001", -- t[1609] = 0
      "0000" when "00011001001010", -- t[1610] = 0
      "0000" when "00011001001011", -- t[1611] = 0
      "0000" when "00011001001100", -- t[1612] = 0
      "0000" when "00011001001101", -- t[1613] = 0
      "0000" when "00011001001110", -- t[1614] = 0
      "0000" when "00011001001111", -- t[1615] = 0
      "0000" when "00011001010000", -- t[1616] = 0
      "0000" when "00011001010001", -- t[1617] = 0
      "0000" when "00011001010010", -- t[1618] = 0
      "0000" when "00011001010011", -- t[1619] = 0
      "0000" when "00011001010100", -- t[1620] = 0
      "0000" when "00011001010101", -- t[1621] = 0
      "0000" when "00011001010110", -- t[1622] = 0
      "0000" when "00011001010111", -- t[1623] = 0
      "0000" when "00011001011000", -- t[1624] = 0
      "0000" when "00011001011001", -- t[1625] = 0
      "0000" when "00011001011010", -- t[1626] = 0
      "0000" when "00011001011011", -- t[1627] = 0
      "0000" when "00011001011100", -- t[1628] = 0
      "0000" when "00011001011101", -- t[1629] = 0
      "0000" when "00011001011110", -- t[1630] = 0
      "0000" when "00011001011111", -- t[1631] = 0
      "0000" when "00011001100000", -- t[1632] = 0
      "0000" when "00011001100001", -- t[1633] = 0
      "0000" when "00011001100010", -- t[1634] = 0
      "0000" when "00011001100011", -- t[1635] = 0
      "0000" when "00011001100100", -- t[1636] = 0
      "0000" when "00011001100101", -- t[1637] = 0
      "0000" when "00011001100110", -- t[1638] = 0
      "0000" when "00011001100111", -- t[1639] = 0
      "0000" when "00011001101000", -- t[1640] = 0
      "0000" when "00011001101001", -- t[1641] = 0
      "0000" when "00011001101010", -- t[1642] = 0
      "0000" when "00011001101011", -- t[1643] = 0
      "0000" when "00011001101100", -- t[1644] = 0
      "0000" when "00011001101101", -- t[1645] = 0
      "0000" when "00011001101110", -- t[1646] = 0
      "0000" when "00011001101111", -- t[1647] = 0
      "0000" when "00011001110000", -- t[1648] = 0
      "0000" when "00011001110001", -- t[1649] = 0
      "0000" when "00011001110010", -- t[1650] = 0
      "0000" when "00011001110011", -- t[1651] = 0
      "0000" when "00011001110100", -- t[1652] = 0
      "0000" when "00011001110101", -- t[1653] = 0
      "0000" when "00011001110110", -- t[1654] = 0
      "0000" when "00011001110111", -- t[1655] = 0
      "0000" when "00011001111000", -- t[1656] = 0
      "0000" when "00011001111001", -- t[1657] = 0
      "0000" when "00011001111010", -- t[1658] = 0
      "0000" when "00011001111011", -- t[1659] = 0
      "0000" when "00011001111100", -- t[1660] = 0
      "0000" when "00011001111101", -- t[1661] = 0
      "0000" when "00011001111110", -- t[1662] = 0
      "0000" when "00011001111111", -- t[1663] = 0
      "0000" when "00011010000000", -- t[1664] = 0
      "0000" when "00011010000001", -- t[1665] = 0
      "0000" when "00011010000010", -- t[1666] = 0
      "0000" when "00011010000011", -- t[1667] = 0
      "0000" when "00011010000100", -- t[1668] = 0
      "0000" when "00011010000101", -- t[1669] = 0
      "0000" when "00011010000110", -- t[1670] = 0
      "0000" when "00011010000111", -- t[1671] = 0
      "0000" when "00011010001000", -- t[1672] = 0
      "0000" when "00011010001001", -- t[1673] = 0
      "0000" when "00011010001010", -- t[1674] = 0
      "0000" when "00011010001011", -- t[1675] = 0
      "0000" when "00011010001100", -- t[1676] = 0
      "0000" when "00011010001101", -- t[1677] = 0
      "0000" when "00011010001110", -- t[1678] = 0
      "0000" when "00011010001111", -- t[1679] = 0
      "0000" when "00011010010000", -- t[1680] = 0
      "0000" when "00011010010001", -- t[1681] = 0
      "0000" when "00011010010010", -- t[1682] = 0
      "0000" when "00011010010011", -- t[1683] = 0
      "0000" when "00011010010100", -- t[1684] = 0
      "0000" when "00011010010101", -- t[1685] = 0
      "0000" when "00011010010110", -- t[1686] = 0
      "0000" when "00011010010111", -- t[1687] = 0
      "0000" when "00011010011000", -- t[1688] = 0
      "0000" when "00011010011001", -- t[1689] = 0
      "0000" when "00011010011010", -- t[1690] = 0
      "0000" when "00011010011011", -- t[1691] = 0
      "0000" when "00011010011100", -- t[1692] = 0
      "0000" when "00011010011101", -- t[1693] = 0
      "0000" when "00011010011110", -- t[1694] = 0
      "0000" when "00011010011111", -- t[1695] = 0
      "0000" when "00011010100000", -- t[1696] = 0
      "0000" when "00011010100001", -- t[1697] = 0
      "0000" when "00011010100010", -- t[1698] = 0
      "0000" when "00011010100011", -- t[1699] = 0
      "0000" when "00011010100100", -- t[1700] = 0
      "0000" when "00011010100101", -- t[1701] = 0
      "0000" when "00011010100110", -- t[1702] = 0
      "0000" when "00011010100111", -- t[1703] = 0
      "0000" when "00011010101000", -- t[1704] = 0
      "0000" when "00011010101001", -- t[1705] = 0
      "0000" when "00011010101010", -- t[1706] = 0
      "0000" when "00011010101011", -- t[1707] = 0
      "0000" when "00011010101100", -- t[1708] = 0
      "0000" when "00011010101101", -- t[1709] = 0
      "0000" when "00011010101110", -- t[1710] = 0
      "0000" when "00011010101111", -- t[1711] = 0
      "0000" when "00011010110000", -- t[1712] = 0
      "0000" when "00011010110001", -- t[1713] = 0
      "0000" when "00011010110010", -- t[1714] = 0
      "0000" when "00011010110011", -- t[1715] = 0
      "0000" when "00011010110100", -- t[1716] = 0
      "0000" when "00011010110101", -- t[1717] = 0
      "0000" when "00011010110110", -- t[1718] = 0
      "0000" when "00011010110111", -- t[1719] = 0
      "0000" when "00011010111000", -- t[1720] = 0
      "0000" when "00011010111001", -- t[1721] = 0
      "0000" when "00011010111010", -- t[1722] = 0
      "0000" when "00011010111011", -- t[1723] = 0
      "0000" when "00011010111100", -- t[1724] = 0
      "0000" when "00011010111101", -- t[1725] = 0
      "0000" when "00011010111110", -- t[1726] = 0
      "0000" when "00011010111111", -- t[1727] = 0
      "0000" when "00011011000000", -- t[1728] = 0
      "0000" when "00011011000001", -- t[1729] = 0
      "0000" when "00011011000010", -- t[1730] = 0
      "0000" when "00011011000011", -- t[1731] = 0
      "0000" when "00011011000100", -- t[1732] = 0
      "0000" when "00011011000101", -- t[1733] = 0
      "0000" when "00011011000110", -- t[1734] = 0
      "0000" when "00011011000111", -- t[1735] = 0
      "0000" when "00011011001000", -- t[1736] = 0
      "0000" when "00011011001001", -- t[1737] = 0
      "0000" when "00011011001010", -- t[1738] = 0
      "0000" when "00011011001011", -- t[1739] = 0
      "0000" when "00011011001100", -- t[1740] = 0
      "0000" when "00011011001101", -- t[1741] = 0
      "0000" when "00011011001110", -- t[1742] = 0
      "0000" when "00011011001111", -- t[1743] = 0
      "0000" when "00011011010000", -- t[1744] = 0
      "0000" when "00011011010001", -- t[1745] = 0
      "0000" when "00011011010010", -- t[1746] = 0
      "0000" when "00011011010011", -- t[1747] = 0
      "0000" when "00011011010100", -- t[1748] = 0
      "0000" when "00011011010101", -- t[1749] = 0
      "0000" when "00011011010110", -- t[1750] = 0
      "0000" when "00011011010111", -- t[1751] = 0
      "0000" when "00011011011000", -- t[1752] = 0
      "0000" when "00011011011001", -- t[1753] = 0
      "0000" when "00011011011010", -- t[1754] = 0
      "0000" when "00011011011011", -- t[1755] = 0
      "0000" when "00011011011100", -- t[1756] = 0
      "0000" when "00011011011101", -- t[1757] = 0
      "0000" when "00011011011110", -- t[1758] = 0
      "0000" when "00011011011111", -- t[1759] = 0
      "0000" when "00011011100000", -- t[1760] = 0
      "0000" when "00011011100001", -- t[1761] = 0
      "0000" when "00011011100010", -- t[1762] = 0
      "0000" when "00011011100011", -- t[1763] = 0
      "0000" when "00011011100100", -- t[1764] = 0
      "0000" when "00011011100101", -- t[1765] = 0
      "0000" when "00011011100110", -- t[1766] = 0
      "0000" when "00011011100111", -- t[1767] = 0
      "0000" when "00011011101000", -- t[1768] = 0
      "0000" when "00011011101001", -- t[1769] = 0
      "0000" when "00011011101010", -- t[1770] = 0
      "0000" when "00011011101011", -- t[1771] = 0
      "0000" when "00011011101100", -- t[1772] = 0
      "0000" when "00011011101101", -- t[1773] = 0
      "0000" when "00011011101110", -- t[1774] = 0
      "0000" when "00011011101111", -- t[1775] = 0
      "0000" when "00011011110000", -- t[1776] = 0
      "0000" when "00011011110001", -- t[1777] = 0
      "0000" when "00011011110010", -- t[1778] = 0
      "0000" when "00011011110011", -- t[1779] = 0
      "0000" when "00011011110100", -- t[1780] = 0
      "0000" when "00011011110101", -- t[1781] = 0
      "0000" when "00011011110110", -- t[1782] = 0
      "0000" when "00011011110111", -- t[1783] = 0
      "0000" when "00011011111000", -- t[1784] = 0
      "0000" when "00011011111001", -- t[1785] = 0
      "0000" when "00011011111010", -- t[1786] = 0
      "0000" when "00011011111011", -- t[1787] = 0
      "0000" when "00011011111100", -- t[1788] = 0
      "0000" when "00011011111101", -- t[1789] = 0
      "0000" when "00011011111110", -- t[1790] = 0
      "0000" when "00011011111111", -- t[1791] = 0
      "0000" when "00011100000000", -- t[1792] = 0
      "0000" when "00011100000001", -- t[1793] = 0
      "0000" when "00011100000010", -- t[1794] = 0
      "0000" when "00011100000011", -- t[1795] = 0
      "0000" when "00011100000100", -- t[1796] = 0
      "0000" when "00011100000101", -- t[1797] = 0
      "0000" when "00011100000110", -- t[1798] = 0
      "0000" when "00011100000111", -- t[1799] = 0
      "0000" when "00011100001000", -- t[1800] = 0
      "0000" when "00011100001001", -- t[1801] = 0
      "0000" when "00011100001010", -- t[1802] = 0
      "0000" when "00011100001011", -- t[1803] = 0
      "0000" when "00011100001100", -- t[1804] = 0
      "0000" when "00011100001101", -- t[1805] = 0
      "0000" when "00011100001110", -- t[1806] = 0
      "0000" when "00011100001111", -- t[1807] = 0
      "0000" when "00011100010000", -- t[1808] = 0
      "0000" when "00011100010001", -- t[1809] = 0
      "0000" when "00011100010010", -- t[1810] = 0
      "0000" when "00011100010011", -- t[1811] = 0
      "0000" when "00011100010100", -- t[1812] = 0
      "0000" when "00011100010101", -- t[1813] = 0
      "0000" when "00011100010110", -- t[1814] = 0
      "0000" when "00011100010111", -- t[1815] = 0
      "0000" when "00011100011000", -- t[1816] = 0
      "0000" when "00011100011001", -- t[1817] = 0
      "0000" when "00011100011010", -- t[1818] = 0
      "0000" when "00011100011011", -- t[1819] = 0
      "0000" when "00011100011100", -- t[1820] = 0
      "0000" when "00011100011101", -- t[1821] = 0
      "0000" when "00011100011110", -- t[1822] = 0
      "0000" when "00011100011111", -- t[1823] = 0
      "0000" when "00011100100000", -- t[1824] = 0
      "0000" when "00011100100001", -- t[1825] = 0
      "0000" when "00011100100010", -- t[1826] = 0
      "0000" when "00011100100011", -- t[1827] = 0
      "0000" when "00011100100100", -- t[1828] = 0
      "0000" when "00011100100101", -- t[1829] = 0
      "0000" when "00011100100110", -- t[1830] = 0
      "0000" when "00011100100111", -- t[1831] = 0
      "0000" when "00011100101000", -- t[1832] = 0
      "0000" when "00011100101001", -- t[1833] = 0
      "0000" when "00011100101010", -- t[1834] = 0
      "0000" when "00011100101011", -- t[1835] = 0
      "0000" when "00011100101100", -- t[1836] = 0
      "0000" when "00011100101101", -- t[1837] = 0
      "0000" when "00011100101110", -- t[1838] = 0
      "0000" when "00011100101111", -- t[1839] = 0
      "0000" when "00011100110000", -- t[1840] = 0
      "0000" when "00011100110001", -- t[1841] = 0
      "0000" when "00011100110010", -- t[1842] = 0
      "0000" when "00011100110011", -- t[1843] = 0
      "0000" when "00011100110100", -- t[1844] = 0
      "0000" when "00011100110101", -- t[1845] = 0
      "0000" when "00011100110110", -- t[1846] = 0
      "0000" when "00011100110111", -- t[1847] = 0
      "0000" when "00011100111000", -- t[1848] = 0
      "0000" when "00011100111001", -- t[1849] = 0
      "0000" when "00011100111010", -- t[1850] = 0
      "0000" when "00011100111011", -- t[1851] = 0
      "0000" when "00011100111100", -- t[1852] = 0
      "0000" when "00011100111101", -- t[1853] = 0
      "0000" when "00011100111110", -- t[1854] = 0
      "0000" when "00011100111111", -- t[1855] = 0
      "0000" when "00011101000000", -- t[1856] = 0
      "0000" when "00011101000001", -- t[1857] = 0
      "0000" when "00011101000010", -- t[1858] = 0
      "0000" when "00011101000011", -- t[1859] = 0
      "0000" when "00011101000100", -- t[1860] = 0
      "0000" when "00011101000101", -- t[1861] = 0
      "0000" when "00011101000110", -- t[1862] = 0
      "0000" when "00011101000111", -- t[1863] = 0
      "0000" when "00011101001000", -- t[1864] = 0
      "0000" when "00011101001001", -- t[1865] = 0
      "0000" when "00011101001010", -- t[1866] = 0
      "0000" when "00011101001011", -- t[1867] = 0
      "0000" when "00011101001100", -- t[1868] = 0
      "0000" when "00011101001101", -- t[1869] = 0
      "0000" when "00011101001110", -- t[1870] = 0
      "0000" when "00011101001111", -- t[1871] = 0
      "0000" when "00011101010000", -- t[1872] = 0
      "0000" when "00011101010001", -- t[1873] = 0
      "0000" when "00011101010010", -- t[1874] = 0
      "0000" when "00011101010011", -- t[1875] = 0
      "0000" when "00011101010100", -- t[1876] = 0
      "0000" when "00011101010101", -- t[1877] = 0
      "0000" when "00011101010110", -- t[1878] = 0
      "0000" when "00011101010111", -- t[1879] = 0
      "0000" when "00011101011000", -- t[1880] = 0
      "0000" when "00011101011001", -- t[1881] = 0
      "0000" when "00011101011010", -- t[1882] = 0
      "0000" when "00011101011011", -- t[1883] = 0
      "0000" when "00011101011100", -- t[1884] = 0
      "0000" when "00011101011101", -- t[1885] = 0
      "0000" when "00011101011110", -- t[1886] = 0
      "0000" when "00011101011111", -- t[1887] = 0
      "0000" when "00011101100000", -- t[1888] = 0
      "0000" when "00011101100001", -- t[1889] = 0
      "0000" when "00011101100010", -- t[1890] = 0
      "0000" when "00011101100011", -- t[1891] = 0
      "0000" when "00011101100100", -- t[1892] = 0
      "0000" when "00011101100101", -- t[1893] = 0
      "0000" when "00011101100110", -- t[1894] = 0
      "0000" when "00011101100111", -- t[1895] = 0
      "0000" when "00011101101000", -- t[1896] = 0
      "0000" when "00011101101001", -- t[1897] = 0
      "0000" when "00011101101010", -- t[1898] = 0
      "0000" when "00011101101011", -- t[1899] = 0
      "0000" when "00011101101100", -- t[1900] = 0
      "0000" when "00011101101101", -- t[1901] = 0
      "0000" when "00011101101110", -- t[1902] = 0
      "0000" when "00011101101111", -- t[1903] = 0
      "0000" when "00011101110000", -- t[1904] = 0
      "0000" when "00011101110001", -- t[1905] = 0
      "0000" when "00011101110010", -- t[1906] = 0
      "0000" when "00011101110011", -- t[1907] = 0
      "0000" when "00011101110100", -- t[1908] = 0
      "0000" when "00011101110101", -- t[1909] = 0
      "0000" when "00011101110110", -- t[1910] = 0
      "0000" when "00011101110111", -- t[1911] = 0
      "0000" when "00011101111000", -- t[1912] = 0
      "0000" when "00011101111001", -- t[1913] = 0
      "0000" when "00011101111010", -- t[1914] = 0
      "0000" when "00011101111011", -- t[1915] = 0
      "0000" when "00011101111100", -- t[1916] = 0
      "0000" when "00011101111101", -- t[1917] = 0
      "0000" when "00011101111110", -- t[1918] = 0
      "0000" when "00011101111111", -- t[1919] = 0
      "0000" when "00011110000000", -- t[1920] = 0
      "0000" when "00011110000001", -- t[1921] = 0
      "0000" when "00011110000010", -- t[1922] = 0
      "0000" when "00011110000011", -- t[1923] = 0
      "0000" when "00011110000100", -- t[1924] = 0
      "0000" when "00011110000101", -- t[1925] = 0
      "0000" when "00011110000110", -- t[1926] = 0
      "0000" when "00011110000111", -- t[1927] = 0
      "0000" when "00011110001000", -- t[1928] = 0
      "0000" when "00011110001001", -- t[1929] = 0
      "0000" when "00011110001010", -- t[1930] = 0
      "0000" when "00011110001011", -- t[1931] = 0
      "0000" when "00011110001100", -- t[1932] = 0
      "0000" when "00011110001101", -- t[1933] = 0
      "0000" when "00011110001110", -- t[1934] = 0
      "0000" when "00011110001111", -- t[1935] = 0
      "0000" when "00011110010000", -- t[1936] = 0
      "0000" when "00011110010001", -- t[1937] = 0
      "0000" when "00011110010010", -- t[1938] = 0
      "0000" when "00011110010011", -- t[1939] = 0
      "0000" when "00011110010100", -- t[1940] = 0
      "0000" when "00011110010101", -- t[1941] = 0
      "0000" when "00011110010110", -- t[1942] = 0
      "0000" when "00011110010111", -- t[1943] = 0
      "0000" when "00011110011000", -- t[1944] = 0
      "0000" when "00011110011001", -- t[1945] = 0
      "0000" when "00011110011010", -- t[1946] = 0
      "0000" when "00011110011011", -- t[1947] = 0
      "0000" when "00011110011100", -- t[1948] = 0
      "0000" when "00011110011101", -- t[1949] = 0
      "0000" when "00011110011110", -- t[1950] = 0
      "0000" when "00011110011111", -- t[1951] = 0
      "0000" when "00011110100000", -- t[1952] = 0
      "0000" when "00011110100001", -- t[1953] = 0
      "0000" when "00011110100010", -- t[1954] = 0
      "0000" when "00011110100011", -- t[1955] = 0
      "0000" when "00011110100100", -- t[1956] = 0
      "0000" when "00011110100101", -- t[1957] = 0
      "0000" when "00011110100110", -- t[1958] = 0
      "0000" when "00011110100111", -- t[1959] = 0
      "0000" when "00011110101000", -- t[1960] = 0
      "0000" when "00011110101001", -- t[1961] = 0
      "0000" when "00011110101010", -- t[1962] = 0
      "0000" when "00011110101011", -- t[1963] = 0
      "0000" when "00011110101100", -- t[1964] = 0
      "0000" when "00011110101101", -- t[1965] = 0
      "0000" when "00011110101110", -- t[1966] = 0
      "0000" when "00011110101111", -- t[1967] = 0
      "0000" when "00011110110000", -- t[1968] = 0
      "0000" when "00011110110001", -- t[1969] = 0
      "0000" when "00011110110010", -- t[1970] = 0
      "0000" when "00011110110011", -- t[1971] = 0
      "0000" when "00011110110100", -- t[1972] = 0
      "0000" when "00011110110101", -- t[1973] = 0
      "0000" when "00011110110110", -- t[1974] = 0
      "0000" when "00011110110111", -- t[1975] = 0
      "0000" when "00011110111000", -- t[1976] = 0
      "0000" when "00011110111001", -- t[1977] = 0
      "0000" when "00011110111010", -- t[1978] = 0
      "0000" when "00011110111011", -- t[1979] = 0
      "0000" when "00011110111100", -- t[1980] = 0
      "0000" when "00011110111101", -- t[1981] = 0
      "0000" when "00011110111110", -- t[1982] = 0
      "0000" when "00011110111111", -- t[1983] = 0
      "0000" when "00011111000000", -- t[1984] = 0
      "0000" when "00011111000001", -- t[1985] = 0
      "0000" when "00011111000010", -- t[1986] = 0
      "0000" when "00011111000011", -- t[1987] = 0
      "0000" when "00011111000100", -- t[1988] = 0
      "0000" when "00011111000101", -- t[1989] = 0
      "0000" when "00011111000110", -- t[1990] = 0
      "0000" when "00011111000111", -- t[1991] = 0
      "0000" when "00011111001000", -- t[1992] = 0
      "0000" when "00011111001001", -- t[1993] = 0
      "0000" when "00011111001010", -- t[1994] = 0
      "0000" when "00011111001011", -- t[1995] = 0
      "0000" when "00011111001100", -- t[1996] = 0
      "0000" when "00011111001101", -- t[1997] = 0
      "0000" when "00011111001110", -- t[1998] = 0
      "0000" when "00011111001111", -- t[1999] = 0
      "0000" when "00011111010000", -- t[2000] = 0
      "0000" when "00011111010001", -- t[2001] = 0
      "0000" when "00011111010010", -- t[2002] = 0
      "0000" when "00011111010011", -- t[2003] = 0
      "0000" when "00011111010100", -- t[2004] = 0
      "0000" when "00011111010101", -- t[2005] = 0
      "0000" when "00011111010110", -- t[2006] = 0
      "0000" when "00011111010111", -- t[2007] = 0
      "0000" when "00011111011000", -- t[2008] = 0
      "0000" when "00011111011001", -- t[2009] = 0
      "0000" when "00011111011010", -- t[2010] = 0
      "0000" when "00011111011011", -- t[2011] = 0
      "0000" when "00011111011100", -- t[2012] = 0
      "0000" when "00011111011101", -- t[2013] = 0
      "0000" when "00011111011110", -- t[2014] = 0
      "0000" when "00011111011111", -- t[2015] = 0
      "0000" when "00011111100000", -- t[2016] = 0
      "0000" when "00011111100001", -- t[2017] = 0
      "0000" when "00011111100010", -- t[2018] = 0
      "0000" when "00011111100011", -- t[2019] = 0
      "0000" when "00011111100100", -- t[2020] = 0
      "0000" when "00011111100101", -- t[2021] = 0
      "0000" when "00011111100110", -- t[2022] = 0
      "0000" when "00011111100111", -- t[2023] = 0
      "0000" when "00011111101000", -- t[2024] = 0
      "0000" when "00011111101001", -- t[2025] = 0
      "0000" when "00011111101010", -- t[2026] = 0
      "0000" when "00011111101011", -- t[2027] = 0
      "0000" when "00011111101100", -- t[2028] = 0
      "0000" when "00011111101101", -- t[2029] = 0
      "0000" when "00011111101110", -- t[2030] = 0
      "0000" when "00011111101111", -- t[2031] = 0
      "0000" when "00011111110000", -- t[2032] = 0
      "0000" when "00011111110001", -- t[2033] = 0
      "0000" when "00011111110010", -- t[2034] = 0
      "0000" when "00011111110011", -- t[2035] = 0
      "0000" when "00011111110100", -- t[2036] = 0
      "0000" when "00011111110101", -- t[2037] = 0
      "0000" when "00011111110110", -- t[2038] = 0
      "0000" when "00011111110111", -- t[2039] = 0
      "0000" when "00011111111000", -- t[2040] = 0
      "0000" when "00011111111001", -- t[2041] = 0
      "0000" when "00011111111010", -- t[2042] = 0
      "0000" when "00011111111011", -- t[2043] = 0
      "0000" when "00011111111100", -- t[2044] = 0
      "0000" when "00011111111101", -- t[2045] = 0
      "0000" when "00011111111110", -- t[2046] = 0
      "0000" when "00011111111111", -- t[2047] = 0
      "0000" when "00100000000000", -- t[2048] = 0
      "0000" when "00100000000001", -- t[2049] = 0
      "0000" when "00100000000010", -- t[2050] = 0
      "0000" when "00100000000011", -- t[2051] = 0
      "0000" when "00100000000100", -- t[2052] = 0
      "0000" when "00100000000101", -- t[2053] = 0
      "0000" when "00100000000110", -- t[2054] = 0
      "0000" when "00100000000111", -- t[2055] = 0
      "0000" when "00100000001000", -- t[2056] = 0
      "0000" when "00100000001001", -- t[2057] = 0
      "0000" when "00100000001010", -- t[2058] = 0
      "0000" when "00100000001011", -- t[2059] = 0
      "0000" when "00100000001100", -- t[2060] = 0
      "0000" when "00100000001101", -- t[2061] = 0
      "0000" when "00100000001110", -- t[2062] = 0
      "0000" when "00100000001111", -- t[2063] = 0
      "0000" when "00100000010000", -- t[2064] = 0
      "0000" when "00100000010001", -- t[2065] = 0
      "0000" when "00100000010010", -- t[2066] = 0
      "0000" when "00100000010011", -- t[2067] = 0
      "0000" when "00100000010100", -- t[2068] = 0
      "0000" when "00100000010101", -- t[2069] = 0
      "0000" when "00100000010110", -- t[2070] = 0
      "0000" when "00100000010111", -- t[2071] = 0
      "0000" when "00100000011000", -- t[2072] = 0
      "0000" when "00100000011001", -- t[2073] = 0
      "0000" when "00100000011010", -- t[2074] = 0
      "0000" when "00100000011011", -- t[2075] = 0
      "0000" when "00100000011100", -- t[2076] = 0
      "0000" when "00100000011101", -- t[2077] = 0
      "0000" when "00100000011110", -- t[2078] = 0
      "0000" when "00100000011111", -- t[2079] = 0
      "0000" when "00100000100000", -- t[2080] = 0
      "0000" when "00100000100001", -- t[2081] = 0
      "0000" when "00100000100010", -- t[2082] = 0
      "0000" when "00100000100011", -- t[2083] = 0
      "0000" when "00100000100100", -- t[2084] = 0
      "0000" when "00100000100101", -- t[2085] = 0
      "0000" when "00100000100110", -- t[2086] = 0
      "0000" when "00100000100111", -- t[2087] = 0
      "0000" when "00100000101000", -- t[2088] = 0
      "0000" when "00100000101001", -- t[2089] = 0
      "0000" when "00100000101010", -- t[2090] = 0
      "0000" when "00100000101011", -- t[2091] = 0
      "0000" when "00100000101100", -- t[2092] = 0
      "0000" when "00100000101101", -- t[2093] = 0
      "0000" when "00100000101110", -- t[2094] = 0
      "0000" when "00100000101111", -- t[2095] = 0
      "0000" when "00100000110000", -- t[2096] = 0
      "0000" when "00100000110001", -- t[2097] = 0
      "0000" when "00100000110010", -- t[2098] = 0
      "0000" when "00100000110011", -- t[2099] = 0
      "0000" when "00100000110100", -- t[2100] = 0
      "0000" when "00100000110101", -- t[2101] = 0
      "0000" when "00100000110110", -- t[2102] = 0
      "0000" when "00100000110111", -- t[2103] = 0
      "0000" when "00100000111000", -- t[2104] = 0
      "0000" when "00100000111001", -- t[2105] = 0
      "0000" when "00100000111010", -- t[2106] = 0
      "0000" when "00100000111011", -- t[2107] = 0
      "0000" when "00100000111100", -- t[2108] = 0
      "0000" when "00100000111101", -- t[2109] = 0
      "0000" when "00100000111110", -- t[2110] = 0
      "0000" when "00100000111111", -- t[2111] = 0
      "0000" when "00100001000000", -- t[2112] = 0
      "0000" when "00100001000001", -- t[2113] = 0
      "0000" when "00100001000010", -- t[2114] = 0
      "0000" when "00100001000011", -- t[2115] = 0
      "0000" when "00100001000100", -- t[2116] = 0
      "0000" when "00100001000101", -- t[2117] = 0
      "0000" when "00100001000110", -- t[2118] = 0
      "0000" when "00100001000111", -- t[2119] = 0
      "0000" when "00100001001000", -- t[2120] = 0
      "0000" when "00100001001001", -- t[2121] = 0
      "0000" when "00100001001010", -- t[2122] = 0
      "0000" when "00100001001011", -- t[2123] = 0
      "0000" when "00100001001100", -- t[2124] = 0
      "0000" when "00100001001101", -- t[2125] = 0
      "0000" when "00100001001110", -- t[2126] = 0
      "0000" when "00100001001111", -- t[2127] = 0
      "0000" when "00100001010000", -- t[2128] = 0
      "0000" when "00100001010001", -- t[2129] = 0
      "0000" when "00100001010010", -- t[2130] = 0
      "0000" when "00100001010011", -- t[2131] = 0
      "0000" when "00100001010100", -- t[2132] = 0
      "0000" when "00100001010101", -- t[2133] = 0
      "0000" when "00100001010110", -- t[2134] = 0
      "0000" when "00100001010111", -- t[2135] = 0
      "0000" when "00100001011000", -- t[2136] = 0
      "0000" when "00100001011001", -- t[2137] = 0
      "0000" when "00100001011010", -- t[2138] = 0
      "0000" when "00100001011011", -- t[2139] = 0
      "0000" when "00100001011100", -- t[2140] = 0
      "0000" when "00100001011101", -- t[2141] = 0
      "0000" when "00100001011110", -- t[2142] = 0
      "0000" when "00100001011111", -- t[2143] = 0
      "0000" when "00100001100000", -- t[2144] = 0
      "0000" when "00100001100001", -- t[2145] = 0
      "0000" when "00100001100010", -- t[2146] = 0
      "0000" when "00100001100011", -- t[2147] = 0
      "0000" when "00100001100100", -- t[2148] = 0
      "0000" when "00100001100101", -- t[2149] = 0
      "0000" when "00100001100110", -- t[2150] = 0
      "0000" when "00100001100111", -- t[2151] = 0
      "0000" when "00100001101000", -- t[2152] = 0
      "0000" when "00100001101001", -- t[2153] = 0
      "0000" when "00100001101010", -- t[2154] = 0
      "0000" when "00100001101011", -- t[2155] = 0
      "0000" when "00100001101100", -- t[2156] = 0
      "0000" when "00100001101101", -- t[2157] = 0
      "0000" when "00100001101110", -- t[2158] = 0
      "0000" when "00100001101111", -- t[2159] = 0
      "0000" when "00100001110000", -- t[2160] = 0
      "0000" when "00100001110001", -- t[2161] = 0
      "0000" when "00100001110010", -- t[2162] = 0
      "0000" when "00100001110011", -- t[2163] = 0
      "0000" when "00100001110100", -- t[2164] = 0
      "0000" when "00100001110101", -- t[2165] = 0
      "0000" when "00100001110110", -- t[2166] = 0
      "0000" when "00100001110111", -- t[2167] = 0
      "0000" when "00100001111000", -- t[2168] = 0
      "0000" when "00100001111001", -- t[2169] = 0
      "0000" when "00100001111010", -- t[2170] = 0
      "0000" when "00100001111011", -- t[2171] = 0
      "0000" when "00100001111100", -- t[2172] = 0
      "0000" when "00100001111101", -- t[2173] = 0
      "0000" when "00100001111110", -- t[2174] = 0
      "0000" when "00100001111111", -- t[2175] = 0
      "0000" when "00100010000000", -- t[2176] = 0
      "0000" when "00100010000001", -- t[2177] = 0
      "0000" when "00100010000010", -- t[2178] = 0
      "0000" when "00100010000011", -- t[2179] = 0
      "0000" when "00100010000100", -- t[2180] = 0
      "0000" when "00100010000101", -- t[2181] = 0
      "0000" when "00100010000110", -- t[2182] = 0
      "0000" when "00100010000111", -- t[2183] = 0
      "0000" when "00100010001000", -- t[2184] = 0
      "0000" when "00100010001001", -- t[2185] = 0
      "0000" when "00100010001010", -- t[2186] = 0
      "0000" when "00100010001011", -- t[2187] = 0
      "0000" when "00100010001100", -- t[2188] = 0
      "0000" when "00100010001101", -- t[2189] = 0
      "0000" when "00100010001110", -- t[2190] = 0
      "0000" when "00100010001111", -- t[2191] = 0
      "0000" when "00100010010000", -- t[2192] = 0
      "0000" when "00100010010001", -- t[2193] = 0
      "0000" when "00100010010010", -- t[2194] = 0
      "0000" when "00100010010011", -- t[2195] = 0
      "0000" when "00100010010100", -- t[2196] = 0
      "0000" when "00100010010101", -- t[2197] = 0
      "0000" when "00100010010110", -- t[2198] = 0
      "0000" when "00100010010111", -- t[2199] = 0
      "0000" when "00100010011000", -- t[2200] = 0
      "0000" when "00100010011001", -- t[2201] = 0
      "0000" when "00100010011010", -- t[2202] = 0
      "0000" when "00100010011011", -- t[2203] = 0
      "0000" when "00100010011100", -- t[2204] = 0
      "0000" when "00100010011101", -- t[2205] = 0
      "0000" when "00100010011110", -- t[2206] = 0
      "0000" when "00100010011111", -- t[2207] = 0
      "0000" when "00100010100000", -- t[2208] = 0
      "0000" when "00100010100001", -- t[2209] = 0
      "0000" when "00100010100010", -- t[2210] = 0
      "0000" when "00100010100011", -- t[2211] = 0
      "0000" when "00100010100100", -- t[2212] = 0
      "0000" when "00100010100101", -- t[2213] = 0
      "0000" when "00100010100110", -- t[2214] = 0
      "0000" when "00100010100111", -- t[2215] = 0
      "0000" when "00100010101000", -- t[2216] = 0
      "0000" when "00100010101001", -- t[2217] = 0
      "0000" when "00100010101010", -- t[2218] = 0
      "0000" when "00100010101011", -- t[2219] = 0
      "0000" when "00100010101100", -- t[2220] = 0
      "0000" when "00100010101101", -- t[2221] = 0
      "0000" when "00100010101110", -- t[2222] = 0
      "0000" when "00100010101111", -- t[2223] = 0
      "0000" when "00100010110000", -- t[2224] = 0
      "0000" when "00100010110001", -- t[2225] = 0
      "0000" when "00100010110010", -- t[2226] = 0
      "0000" when "00100010110011", -- t[2227] = 0
      "0000" when "00100010110100", -- t[2228] = 0
      "0000" when "00100010110101", -- t[2229] = 0
      "0000" when "00100010110110", -- t[2230] = 0
      "0000" when "00100010110111", -- t[2231] = 0
      "0000" when "00100010111000", -- t[2232] = 0
      "0000" when "00100010111001", -- t[2233] = 0
      "0000" when "00100010111010", -- t[2234] = 0
      "0000" when "00100010111011", -- t[2235] = 0
      "0000" when "00100010111100", -- t[2236] = 0
      "0000" when "00100010111101", -- t[2237] = 0
      "0000" when "00100010111110", -- t[2238] = 0
      "0000" when "00100010111111", -- t[2239] = 0
      "0000" when "00100011000000", -- t[2240] = 0
      "0000" when "00100011000001", -- t[2241] = 0
      "0000" when "00100011000010", -- t[2242] = 0
      "0000" when "00100011000011", -- t[2243] = 0
      "0000" when "00100011000100", -- t[2244] = 0
      "0000" when "00100011000101", -- t[2245] = 0
      "0000" when "00100011000110", -- t[2246] = 0
      "0000" when "00100011000111", -- t[2247] = 0
      "0000" when "00100011001000", -- t[2248] = 0
      "0000" when "00100011001001", -- t[2249] = 0
      "0000" when "00100011001010", -- t[2250] = 0
      "0000" when "00100011001011", -- t[2251] = 0
      "0000" when "00100011001100", -- t[2252] = 0
      "0000" when "00100011001101", -- t[2253] = 0
      "0000" when "00100011001110", -- t[2254] = 0
      "0000" when "00100011001111", -- t[2255] = 0
      "0000" when "00100011010000", -- t[2256] = 0
      "0000" when "00100011010001", -- t[2257] = 0
      "0000" when "00100011010010", -- t[2258] = 0
      "0000" when "00100011010011", -- t[2259] = 0
      "0000" when "00100011010100", -- t[2260] = 0
      "0000" when "00100011010101", -- t[2261] = 0
      "0000" when "00100011010110", -- t[2262] = 0
      "0000" when "00100011010111", -- t[2263] = 0
      "0000" when "00100011011000", -- t[2264] = 0
      "0000" when "00100011011001", -- t[2265] = 0
      "0000" when "00100011011010", -- t[2266] = 0
      "0000" when "00100011011011", -- t[2267] = 0
      "0000" when "00100011011100", -- t[2268] = 0
      "0000" when "00100011011101", -- t[2269] = 0
      "0000" when "00100011011110", -- t[2270] = 0
      "0000" when "00100011011111", -- t[2271] = 0
      "0000" when "00100011100000", -- t[2272] = 0
      "0000" when "00100011100001", -- t[2273] = 0
      "0000" when "00100011100010", -- t[2274] = 0
      "0000" when "00100011100011", -- t[2275] = 0
      "0000" when "00100011100100", -- t[2276] = 0
      "0000" when "00100011100101", -- t[2277] = 0
      "0000" when "00100011100110", -- t[2278] = 0
      "0000" when "00100011100111", -- t[2279] = 0
      "0000" when "00100011101000", -- t[2280] = 0
      "0000" when "00100011101001", -- t[2281] = 0
      "0000" when "00100011101010", -- t[2282] = 0
      "0000" when "00100011101011", -- t[2283] = 0
      "0000" when "00100011101100", -- t[2284] = 0
      "0000" when "00100011101101", -- t[2285] = 0
      "0000" when "00100011101110", -- t[2286] = 0
      "0000" when "00100011101111", -- t[2287] = 0
      "0000" when "00100011110000", -- t[2288] = 0
      "0000" when "00100011110001", -- t[2289] = 0
      "0000" when "00100011110010", -- t[2290] = 0
      "0000" when "00100011110011", -- t[2291] = 0
      "0000" when "00100011110100", -- t[2292] = 0
      "0000" when "00100011110101", -- t[2293] = 0
      "0000" when "00100011110110", -- t[2294] = 0
      "0000" when "00100011110111", -- t[2295] = 0
      "0000" when "00100011111000", -- t[2296] = 0
      "0000" when "00100011111001", -- t[2297] = 0
      "0000" when "00100011111010", -- t[2298] = 0
      "0000" when "00100011111011", -- t[2299] = 0
      "0000" when "00100011111100", -- t[2300] = 0
      "0000" when "00100011111101", -- t[2301] = 0
      "0000" when "00100011111110", -- t[2302] = 0
      "0000" when "00100011111111", -- t[2303] = 0
      "0000" when "00100100000000", -- t[2304] = 0
      "0000" when "00100100000001", -- t[2305] = 0
      "0000" when "00100100000010", -- t[2306] = 0
      "0000" when "00100100000011", -- t[2307] = 0
      "0000" when "00100100000100", -- t[2308] = 0
      "0000" when "00100100000101", -- t[2309] = 0
      "0000" when "00100100000110", -- t[2310] = 0
      "0000" when "00100100000111", -- t[2311] = 0
      "0000" when "00100100001000", -- t[2312] = 0
      "0000" when "00100100001001", -- t[2313] = 0
      "0000" when "00100100001010", -- t[2314] = 0
      "0000" when "00100100001011", -- t[2315] = 0
      "0000" when "00100100001100", -- t[2316] = 0
      "0000" when "00100100001101", -- t[2317] = 0
      "0000" when "00100100001110", -- t[2318] = 0
      "0000" when "00100100001111", -- t[2319] = 0
      "0000" when "00100100010000", -- t[2320] = 0
      "0000" when "00100100010001", -- t[2321] = 0
      "0000" when "00100100010010", -- t[2322] = 0
      "0000" when "00100100010011", -- t[2323] = 0
      "0000" when "00100100010100", -- t[2324] = 0
      "0000" when "00100100010101", -- t[2325] = 0
      "0000" when "00100100010110", -- t[2326] = 0
      "0000" when "00100100010111", -- t[2327] = 0
      "0000" when "00100100011000", -- t[2328] = 0
      "0000" when "00100100011001", -- t[2329] = 0
      "0000" when "00100100011010", -- t[2330] = 0
      "0000" when "00100100011011", -- t[2331] = 0
      "0000" when "00100100011100", -- t[2332] = 0
      "0000" when "00100100011101", -- t[2333] = 0
      "0000" when "00100100011110", -- t[2334] = 0
      "0000" when "00100100011111", -- t[2335] = 0
      "0000" when "00100100100000", -- t[2336] = 0
      "0000" when "00100100100001", -- t[2337] = 0
      "0000" when "00100100100010", -- t[2338] = 0
      "0000" when "00100100100011", -- t[2339] = 0
      "0000" when "00100100100100", -- t[2340] = 0
      "0000" when "00100100100101", -- t[2341] = 0
      "0000" when "00100100100110", -- t[2342] = 0
      "0000" when "00100100100111", -- t[2343] = 0
      "0000" when "00100100101000", -- t[2344] = 0
      "0000" when "00100100101001", -- t[2345] = 0
      "0000" when "00100100101010", -- t[2346] = 0
      "0000" when "00100100101011", -- t[2347] = 0
      "0000" when "00100100101100", -- t[2348] = 0
      "0000" when "00100100101101", -- t[2349] = 0
      "0000" when "00100100101110", -- t[2350] = 0
      "0000" when "00100100101111", -- t[2351] = 0
      "0000" when "00100100110000", -- t[2352] = 0
      "0000" when "00100100110001", -- t[2353] = 0
      "0000" when "00100100110010", -- t[2354] = 0
      "0000" when "00100100110011", -- t[2355] = 0
      "0000" when "00100100110100", -- t[2356] = 0
      "0000" when "00100100110101", -- t[2357] = 0
      "0000" when "00100100110110", -- t[2358] = 0
      "0000" when "00100100110111", -- t[2359] = 0
      "0000" when "00100100111000", -- t[2360] = 0
      "0000" when "00100100111001", -- t[2361] = 0
      "0000" when "00100100111010", -- t[2362] = 0
      "0000" when "00100100111011", -- t[2363] = 0
      "0000" when "00100100111100", -- t[2364] = 0
      "0000" when "00100100111101", -- t[2365] = 0
      "0000" when "00100100111110", -- t[2366] = 0
      "0000" when "00100100111111", -- t[2367] = 0
      "0000" when "00100101000000", -- t[2368] = 0
      "0000" when "00100101000001", -- t[2369] = 0
      "0000" when "00100101000010", -- t[2370] = 0
      "0000" when "00100101000011", -- t[2371] = 0
      "0000" when "00100101000100", -- t[2372] = 0
      "0000" when "00100101000101", -- t[2373] = 0
      "0000" when "00100101000110", -- t[2374] = 0
      "0000" when "00100101000111", -- t[2375] = 0
      "0000" when "00100101001000", -- t[2376] = 0
      "0000" when "00100101001001", -- t[2377] = 0
      "0000" when "00100101001010", -- t[2378] = 0
      "0000" when "00100101001011", -- t[2379] = 0
      "0000" when "00100101001100", -- t[2380] = 0
      "0000" when "00100101001101", -- t[2381] = 0
      "0000" when "00100101001110", -- t[2382] = 0
      "0000" when "00100101001111", -- t[2383] = 0
      "0000" when "00100101010000", -- t[2384] = 0
      "0000" when "00100101010001", -- t[2385] = 0
      "0000" when "00100101010010", -- t[2386] = 0
      "0000" when "00100101010011", -- t[2387] = 0
      "0000" when "00100101010100", -- t[2388] = 0
      "0000" when "00100101010101", -- t[2389] = 0
      "0000" when "00100101010110", -- t[2390] = 0
      "0000" when "00100101010111", -- t[2391] = 0
      "0000" when "00100101011000", -- t[2392] = 0
      "0000" when "00100101011001", -- t[2393] = 0
      "0000" when "00100101011010", -- t[2394] = 0
      "0000" when "00100101011011", -- t[2395] = 0
      "0000" when "00100101011100", -- t[2396] = 0
      "0000" when "00100101011101", -- t[2397] = 0
      "0000" when "00100101011110", -- t[2398] = 0
      "0000" when "00100101011111", -- t[2399] = 0
      "0000" when "00100101100000", -- t[2400] = 0
      "0000" when "00100101100001", -- t[2401] = 0
      "0000" when "00100101100010", -- t[2402] = 0
      "0000" when "00100101100011", -- t[2403] = 0
      "0000" when "00100101100100", -- t[2404] = 0
      "0000" when "00100101100101", -- t[2405] = 0
      "0000" when "00100101100110", -- t[2406] = 0
      "0000" when "00100101100111", -- t[2407] = 0
      "0000" when "00100101101000", -- t[2408] = 0
      "0000" when "00100101101001", -- t[2409] = 0
      "0000" when "00100101101010", -- t[2410] = 0
      "0000" when "00100101101011", -- t[2411] = 0
      "0000" when "00100101101100", -- t[2412] = 0
      "0000" when "00100101101101", -- t[2413] = 0
      "0000" when "00100101101110", -- t[2414] = 0
      "0000" when "00100101101111", -- t[2415] = 0
      "0000" when "00100101110000", -- t[2416] = 0
      "0000" when "00100101110001", -- t[2417] = 0
      "0000" when "00100101110010", -- t[2418] = 0
      "0000" when "00100101110011", -- t[2419] = 0
      "0000" when "00100101110100", -- t[2420] = 0
      "0000" when "00100101110101", -- t[2421] = 0
      "0000" when "00100101110110", -- t[2422] = 0
      "0000" when "00100101110111", -- t[2423] = 0
      "0000" when "00100101111000", -- t[2424] = 0
      "0000" when "00100101111001", -- t[2425] = 0
      "0000" when "00100101111010", -- t[2426] = 0
      "0000" when "00100101111011", -- t[2427] = 0
      "0000" when "00100101111100", -- t[2428] = 0
      "0000" when "00100101111101", -- t[2429] = 0
      "0000" when "00100101111110", -- t[2430] = 0
      "0000" when "00100101111111", -- t[2431] = 0
      "0000" when "00100110000000", -- t[2432] = 0
      "0000" when "00100110000001", -- t[2433] = 0
      "0000" when "00100110000010", -- t[2434] = 0
      "0000" when "00100110000011", -- t[2435] = 0
      "0000" when "00100110000100", -- t[2436] = 0
      "0000" when "00100110000101", -- t[2437] = 0
      "0000" when "00100110000110", -- t[2438] = 0
      "0000" when "00100110000111", -- t[2439] = 0
      "0000" when "00100110001000", -- t[2440] = 0
      "0000" when "00100110001001", -- t[2441] = 0
      "0000" when "00100110001010", -- t[2442] = 0
      "0000" when "00100110001011", -- t[2443] = 0
      "0000" when "00100110001100", -- t[2444] = 0
      "0000" when "00100110001101", -- t[2445] = 0
      "0000" when "00100110001110", -- t[2446] = 0
      "0000" when "00100110001111", -- t[2447] = 0
      "0000" when "00100110010000", -- t[2448] = 0
      "0000" when "00100110010001", -- t[2449] = 0
      "0000" when "00100110010010", -- t[2450] = 0
      "0000" when "00100110010011", -- t[2451] = 0
      "0000" when "00100110010100", -- t[2452] = 0
      "0000" when "00100110010101", -- t[2453] = 0
      "0000" when "00100110010110", -- t[2454] = 0
      "0000" when "00100110010111", -- t[2455] = 0
      "0000" when "00100110011000", -- t[2456] = 0
      "0000" when "00100110011001", -- t[2457] = 0
      "0000" when "00100110011010", -- t[2458] = 0
      "0000" when "00100110011011", -- t[2459] = 0
      "0000" when "00100110011100", -- t[2460] = 0
      "0000" when "00100110011101", -- t[2461] = 0
      "0000" when "00100110011110", -- t[2462] = 0
      "0000" when "00100110011111", -- t[2463] = 0
      "0000" when "00100110100000", -- t[2464] = 0
      "0000" when "00100110100001", -- t[2465] = 0
      "0000" when "00100110100010", -- t[2466] = 0
      "0000" when "00100110100011", -- t[2467] = 0
      "0000" when "00100110100100", -- t[2468] = 0
      "0000" when "00100110100101", -- t[2469] = 0
      "0000" when "00100110100110", -- t[2470] = 0
      "0000" when "00100110100111", -- t[2471] = 0
      "0000" when "00100110101000", -- t[2472] = 0
      "0000" when "00100110101001", -- t[2473] = 0
      "0000" when "00100110101010", -- t[2474] = 0
      "0000" when "00100110101011", -- t[2475] = 0
      "0000" when "00100110101100", -- t[2476] = 0
      "0000" when "00100110101101", -- t[2477] = 0
      "0000" when "00100110101110", -- t[2478] = 0
      "0000" when "00100110101111", -- t[2479] = 0
      "0000" when "00100110110000", -- t[2480] = 0
      "0000" when "00100110110001", -- t[2481] = 0
      "0000" when "00100110110010", -- t[2482] = 0
      "0000" when "00100110110011", -- t[2483] = 0
      "0000" when "00100110110100", -- t[2484] = 0
      "0000" when "00100110110101", -- t[2485] = 0
      "0000" when "00100110110110", -- t[2486] = 0
      "0000" when "00100110110111", -- t[2487] = 0
      "0000" when "00100110111000", -- t[2488] = 0
      "0000" when "00100110111001", -- t[2489] = 0
      "0000" when "00100110111010", -- t[2490] = 0
      "0000" when "00100110111011", -- t[2491] = 0
      "0000" when "00100110111100", -- t[2492] = 0
      "0000" when "00100110111101", -- t[2493] = 0
      "0000" when "00100110111110", -- t[2494] = 0
      "0000" when "00100110111111", -- t[2495] = 0
      "0000" when "00100111000000", -- t[2496] = 0
      "0000" when "00100111000001", -- t[2497] = 0
      "0000" when "00100111000010", -- t[2498] = 0
      "0000" when "00100111000011", -- t[2499] = 0
      "0000" when "00100111000100", -- t[2500] = 0
      "0000" when "00100111000101", -- t[2501] = 0
      "0000" when "00100111000110", -- t[2502] = 0
      "0000" when "00100111000111", -- t[2503] = 0
      "0000" when "00100111001000", -- t[2504] = 0
      "0000" when "00100111001001", -- t[2505] = 0
      "0000" when "00100111001010", -- t[2506] = 0
      "0000" when "00100111001011", -- t[2507] = 0
      "0000" when "00100111001100", -- t[2508] = 0
      "0000" when "00100111001101", -- t[2509] = 0
      "0000" when "00100111001110", -- t[2510] = 0
      "0000" when "00100111001111", -- t[2511] = 0
      "0000" when "00100111010000", -- t[2512] = 0
      "0000" when "00100111010001", -- t[2513] = 0
      "0000" when "00100111010010", -- t[2514] = 0
      "0000" when "00100111010011", -- t[2515] = 0
      "0000" when "00100111010100", -- t[2516] = 0
      "0000" when "00100111010101", -- t[2517] = 0
      "0000" when "00100111010110", -- t[2518] = 0
      "0000" when "00100111010111", -- t[2519] = 0
      "0000" when "00100111011000", -- t[2520] = 0
      "0000" when "00100111011001", -- t[2521] = 0
      "0000" when "00100111011010", -- t[2522] = 0
      "0000" when "00100111011011", -- t[2523] = 0
      "0000" when "00100111011100", -- t[2524] = 0
      "0000" when "00100111011101", -- t[2525] = 0
      "0000" when "00100111011110", -- t[2526] = 0
      "0000" when "00100111011111", -- t[2527] = 0
      "0000" when "00100111100000", -- t[2528] = 0
      "0000" when "00100111100001", -- t[2529] = 0
      "0000" when "00100111100010", -- t[2530] = 0
      "0000" when "00100111100011", -- t[2531] = 0
      "0000" when "00100111100100", -- t[2532] = 0
      "0000" when "00100111100101", -- t[2533] = 0
      "0000" when "00100111100110", -- t[2534] = 0
      "0000" when "00100111100111", -- t[2535] = 0
      "0000" when "00100111101000", -- t[2536] = 0
      "0000" when "00100111101001", -- t[2537] = 0
      "0000" when "00100111101010", -- t[2538] = 0
      "0000" when "00100111101011", -- t[2539] = 0
      "0000" when "00100111101100", -- t[2540] = 0
      "0000" when "00100111101101", -- t[2541] = 0
      "0000" when "00100111101110", -- t[2542] = 0
      "0000" when "00100111101111", -- t[2543] = 0
      "0000" when "00100111110000", -- t[2544] = 0
      "0000" when "00100111110001", -- t[2545] = 0
      "0000" when "00100111110010", -- t[2546] = 0
      "0000" when "00100111110011", -- t[2547] = 0
      "0000" when "00100111110100", -- t[2548] = 0
      "0000" when "00100111110101", -- t[2549] = 0
      "0000" when "00100111110110", -- t[2550] = 0
      "0000" when "00100111110111", -- t[2551] = 0
      "0000" when "00100111111000", -- t[2552] = 0
      "0000" when "00100111111001", -- t[2553] = 0
      "0000" when "00100111111010", -- t[2554] = 0
      "0000" when "00100111111011", -- t[2555] = 0
      "0000" when "00100111111100", -- t[2556] = 0
      "0000" when "00100111111101", -- t[2557] = 0
      "0000" when "00100111111110", -- t[2558] = 0
      "0000" when "00100111111111", -- t[2559] = 0
      "0000" when "00101000000000", -- t[2560] = 0
      "0000" when "00101000000001", -- t[2561] = 0
      "0000" when "00101000000010", -- t[2562] = 0
      "0000" when "00101000000011", -- t[2563] = 0
      "0000" when "00101000000100", -- t[2564] = 0
      "0000" when "00101000000101", -- t[2565] = 0
      "0000" when "00101000000110", -- t[2566] = 0
      "0000" when "00101000000111", -- t[2567] = 0
      "0000" when "00101000001000", -- t[2568] = 0
      "0000" when "00101000001001", -- t[2569] = 0
      "0000" when "00101000001010", -- t[2570] = 0
      "0000" when "00101000001011", -- t[2571] = 0
      "0000" when "00101000001100", -- t[2572] = 0
      "0000" when "00101000001101", -- t[2573] = 0
      "0000" when "00101000001110", -- t[2574] = 0
      "0000" when "00101000001111", -- t[2575] = 0
      "0000" when "00101000010000", -- t[2576] = 0
      "0000" when "00101000010001", -- t[2577] = 0
      "0000" when "00101000010010", -- t[2578] = 0
      "0000" when "00101000010011", -- t[2579] = 0
      "0000" when "00101000010100", -- t[2580] = 0
      "0000" when "00101000010101", -- t[2581] = 0
      "0000" when "00101000010110", -- t[2582] = 0
      "0000" when "00101000010111", -- t[2583] = 0
      "0000" when "00101000011000", -- t[2584] = 0
      "0000" when "00101000011001", -- t[2585] = 0
      "0000" when "00101000011010", -- t[2586] = 0
      "0000" when "00101000011011", -- t[2587] = 0
      "0000" when "00101000011100", -- t[2588] = 0
      "0000" when "00101000011101", -- t[2589] = 0
      "0000" when "00101000011110", -- t[2590] = 0
      "0000" when "00101000011111", -- t[2591] = 0
      "0000" when "00101000100000", -- t[2592] = 0
      "0000" when "00101000100001", -- t[2593] = 0
      "0000" when "00101000100010", -- t[2594] = 0
      "0000" when "00101000100011", -- t[2595] = 0
      "0000" when "00101000100100", -- t[2596] = 0
      "0000" when "00101000100101", -- t[2597] = 0
      "0000" when "00101000100110", -- t[2598] = 0
      "0000" when "00101000100111", -- t[2599] = 0
      "0000" when "00101000101000", -- t[2600] = 0
      "0000" when "00101000101001", -- t[2601] = 0
      "0000" when "00101000101010", -- t[2602] = 0
      "0000" when "00101000101011", -- t[2603] = 0
      "0000" when "00101000101100", -- t[2604] = 0
      "0000" when "00101000101101", -- t[2605] = 0
      "0000" when "00101000101110", -- t[2606] = 0
      "0000" when "00101000101111", -- t[2607] = 0
      "0000" when "00101000110000", -- t[2608] = 0
      "0000" when "00101000110001", -- t[2609] = 0
      "0000" when "00101000110010", -- t[2610] = 0
      "0000" when "00101000110011", -- t[2611] = 0
      "0000" when "00101000110100", -- t[2612] = 0
      "0000" when "00101000110101", -- t[2613] = 0
      "0000" when "00101000110110", -- t[2614] = 0
      "0000" when "00101000110111", -- t[2615] = 0
      "0000" when "00101000111000", -- t[2616] = 0
      "0000" when "00101000111001", -- t[2617] = 0
      "0000" when "00101000111010", -- t[2618] = 0
      "0000" when "00101000111011", -- t[2619] = 0
      "0000" when "00101000111100", -- t[2620] = 0
      "0000" when "00101000111101", -- t[2621] = 0
      "0000" when "00101000111110", -- t[2622] = 0
      "0000" when "00101000111111", -- t[2623] = 0
      "0000" when "00101001000000", -- t[2624] = 0
      "0000" when "00101001000001", -- t[2625] = 0
      "0000" when "00101001000010", -- t[2626] = 0
      "0000" when "00101001000011", -- t[2627] = 0
      "0000" when "00101001000100", -- t[2628] = 0
      "0000" when "00101001000101", -- t[2629] = 0
      "0000" when "00101001000110", -- t[2630] = 0
      "0000" when "00101001000111", -- t[2631] = 0
      "0000" when "00101001001000", -- t[2632] = 0
      "0000" when "00101001001001", -- t[2633] = 0
      "0000" when "00101001001010", -- t[2634] = 0
      "0000" when "00101001001011", -- t[2635] = 0
      "0000" when "00101001001100", -- t[2636] = 0
      "0000" when "00101001001101", -- t[2637] = 0
      "0000" when "00101001001110", -- t[2638] = 0
      "0000" when "00101001001111", -- t[2639] = 0
      "0000" when "00101001010000", -- t[2640] = 0
      "0000" when "00101001010001", -- t[2641] = 0
      "0000" when "00101001010010", -- t[2642] = 0
      "0000" when "00101001010011", -- t[2643] = 0
      "0000" when "00101001010100", -- t[2644] = 0
      "0000" when "00101001010101", -- t[2645] = 0
      "0000" when "00101001010110", -- t[2646] = 0
      "0000" when "00101001010111", -- t[2647] = 0
      "0000" when "00101001011000", -- t[2648] = 0
      "0000" when "00101001011001", -- t[2649] = 0
      "0000" when "00101001011010", -- t[2650] = 0
      "0000" when "00101001011011", -- t[2651] = 0
      "0000" when "00101001011100", -- t[2652] = 0
      "0000" when "00101001011101", -- t[2653] = 0
      "0000" when "00101001011110", -- t[2654] = 0
      "0000" when "00101001011111", -- t[2655] = 0
      "0000" when "00101001100000", -- t[2656] = 0
      "0000" when "00101001100001", -- t[2657] = 0
      "0000" when "00101001100010", -- t[2658] = 0
      "0000" when "00101001100011", -- t[2659] = 0
      "0000" when "00101001100100", -- t[2660] = 0
      "0000" when "00101001100101", -- t[2661] = 0
      "0000" when "00101001100110", -- t[2662] = 0
      "0000" when "00101001100111", -- t[2663] = 0
      "0000" when "00101001101000", -- t[2664] = 0
      "0000" when "00101001101001", -- t[2665] = 0
      "0000" when "00101001101010", -- t[2666] = 0
      "0000" when "00101001101011", -- t[2667] = 0
      "0000" when "00101001101100", -- t[2668] = 0
      "0000" when "00101001101101", -- t[2669] = 0
      "0000" when "00101001101110", -- t[2670] = 0
      "0000" when "00101001101111", -- t[2671] = 0
      "0000" when "00101001110000", -- t[2672] = 0
      "0000" when "00101001110001", -- t[2673] = 0
      "0000" when "00101001110010", -- t[2674] = 0
      "0000" when "00101001110011", -- t[2675] = 0
      "0000" when "00101001110100", -- t[2676] = 0
      "0000" when "00101001110101", -- t[2677] = 0
      "0000" when "00101001110110", -- t[2678] = 0
      "0000" when "00101001110111", -- t[2679] = 0
      "0000" when "00101001111000", -- t[2680] = 0
      "0000" when "00101001111001", -- t[2681] = 0
      "0000" when "00101001111010", -- t[2682] = 0
      "0000" when "00101001111011", -- t[2683] = 0
      "0000" when "00101001111100", -- t[2684] = 0
      "0000" when "00101001111101", -- t[2685] = 0
      "0000" when "00101001111110", -- t[2686] = 0
      "0000" when "00101001111111", -- t[2687] = 0
      "0000" when "00101010000000", -- t[2688] = 0
      "0000" when "00101010000001", -- t[2689] = 0
      "0000" when "00101010000010", -- t[2690] = 0
      "0000" when "00101010000011", -- t[2691] = 0
      "0000" when "00101010000100", -- t[2692] = 0
      "0000" when "00101010000101", -- t[2693] = 0
      "0000" when "00101010000110", -- t[2694] = 0
      "0000" when "00101010000111", -- t[2695] = 0
      "0000" when "00101010001000", -- t[2696] = 0
      "0000" when "00101010001001", -- t[2697] = 0
      "0000" when "00101010001010", -- t[2698] = 0
      "0000" when "00101010001011", -- t[2699] = 0
      "0000" when "00101010001100", -- t[2700] = 0
      "0000" when "00101010001101", -- t[2701] = 0
      "0000" when "00101010001110", -- t[2702] = 0
      "0000" when "00101010001111", -- t[2703] = 0
      "0000" when "00101010010000", -- t[2704] = 0
      "0000" when "00101010010001", -- t[2705] = 0
      "0000" when "00101010010010", -- t[2706] = 0
      "0000" when "00101010010011", -- t[2707] = 0
      "0000" when "00101010010100", -- t[2708] = 0
      "0000" when "00101010010101", -- t[2709] = 0
      "0000" when "00101010010110", -- t[2710] = 0
      "0000" when "00101010010111", -- t[2711] = 0
      "0000" when "00101010011000", -- t[2712] = 0
      "0000" when "00101010011001", -- t[2713] = 0
      "0000" when "00101010011010", -- t[2714] = 0
      "0000" when "00101010011011", -- t[2715] = 0
      "0000" when "00101010011100", -- t[2716] = 0
      "0000" when "00101010011101", -- t[2717] = 0
      "0000" when "00101010011110", -- t[2718] = 0
      "0000" when "00101010011111", -- t[2719] = 0
      "0000" when "00101010100000", -- t[2720] = 0
      "0000" when "00101010100001", -- t[2721] = 0
      "0000" when "00101010100010", -- t[2722] = 0
      "0000" when "00101010100011", -- t[2723] = 0
      "0000" when "00101010100100", -- t[2724] = 0
      "0000" when "00101010100101", -- t[2725] = 0
      "0000" when "00101010100110", -- t[2726] = 0
      "0000" when "00101010100111", -- t[2727] = 0
      "0000" when "00101010101000", -- t[2728] = 0
      "0000" when "00101010101001", -- t[2729] = 0
      "0000" when "00101010101010", -- t[2730] = 0
      "0000" when "00101010101011", -- t[2731] = 0
      "0000" when "00101010101100", -- t[2732] = 0
      "0000" when "00101010101101", -- t[2733] = 0
      "0000" when "00101010101110", -- t[2734] = 0
      "0000" when "00101010101111", -- t[2735] = 0
      "0000" when "00101010110000", -- t[2736] = 0
      "0000" when "00101010110001", -- t[2737] = 0
      "0000" when "00101010110010", -- t[2738] = 0
      "0000" when "00101010110011", -- t[2739] = 0
      "0000" when "00101010110100", -- t[2740] = 0
      "0000" when "00101010110101", -- t[2741] = 0
      "0000" when "00101010110110", -- t[2742] = 0
      "0000" when "00101010110111", -- t[2743] = 0
      "0000" when "00101010111000", -- t[2744] = 0
      "0000" when "00101010111001", -- t[2745] = 0
      "0000" when "00101010111010", -- t[2746] = 0
      "0000" when "00101010111011", -- t[2747] = 0
      "0000" when "00101010111100", -- t[2748] = 0
      "0000" when "00101010111101", -- t[2749] = 0
      "0000" when "00101010111110", -- t[2750] = 0
      "0000" when "00101010111111", -- t[2751] = 0
      "0000" when "00101011000000", -- t[2752] = 0
      "0000" when "00101011000001", -- t[2753] = 0
      "0000" when "00101011000010", -- t[2754] = 0
      "0000" when "00101011000011", -- t[2755] = 0
      "0000" when "00101011000100", -- t[2756] = 0
      "0000" when "00101011000101", -- t[2757] = 0
      "0000" when "00101011000110", -- t[2758] = 0
      "0000" when "00101011000111", -- t[2759] = 0
      "0000" when "00101011001000", -- t[2760] = 0
      "0000" when "00101011001001", -- t[2761] = 0
      "0000" when "00101011001010", -- t[2762] = 0
      "0000" when "00101011001011", -- t[2763] = 0
      "0000" when "00101011001100", -- t[2764] = 0
      "0000" when "00101011001101", -- t[2765] = 0
      "0000" when "00101011001110", -- t[2766] = 0
      "0000" when "00101011001111", -- t[2767] = 0
      "0000" when "00101011010000", -- t[2768] = 0
      "0000" when "00101011010001", -- t[2769] = 0
      "0000" when "00101011010010", -- t[2770] = 0
      "0000" when "00101011010011", -- t[2771] = 0
      "0000" when "00101011010100", -- t[2772] = 0
      "0000" when "00101011010101", -- t[2773] = 0
      "0000" when "00101011010110", -- t[2774] = 0
      "0000" when "00101011010111", -- t[2775] = 0
      "0000" when "00101011011000", -- t[2776] = 0
      "0000" when "00101011011001", -- t[2777] = 0
      "0000" when "00101011011010", -- t[2778] = 0
      "0000" when "00101011011011", -- t[2779] = 0
      "0000" when "00101011011100", -- t[2780] = 0
      "0000" when "00101011011101", -- t[2781] = 0
      "0000" when "00101011011110", -- t[2782] = 0
      "0000" when "00101011011111", -- t[2783] = 0
      "0000" when "00101011100000", -- t[2784] = 0
      "0000" when "00101011100001", -- t[2785] = 0
      "0000" when "00101011100010", -- t[2786] = 0
      "0000" when "00101011100011", -- t[2787] = 0
      "0000" when "00101011100100", -- t[2788] = 0
      "0000" when "00101011100101", -- t[2789] = 0
      "0000" when "00101011100110", -- t[2790] = 0
      "0000" when "00101011100111", -- t[2791] = 0
      "0000" when "00101011101000", -- t[2792] = 0
      "0000" when "00101011101001", -- t[2793] = 0
      "0000" when "00101011101010", -- t[2794] = 0
      "0000" when "00101011101011", -- t[2795] = 0
      "0000" when "00101011101100", -- t[2796] = 0
      "0000" when "00101011101101", -- t[2797] = 0
      "0000" when "00101011101110", -- t[2798] = 0
      "0000" when "00101011101111", -- t[2799] = 0
      "0000" when "00101011110000", -- t[2800] = 0
      "0000" when "00101011110001", -- t[2801] = 0
      "0000" when "00101011110010", -- t[2802] = 0
      "0000" when "00101011110011", -- t[2803] = 0
      "0000" when "00101011110100", -- t[2804] = 0
      "0000" when "00101011110101", -- t[2805] = 0
      "0000" when "00101011110110", -- t[2806] = 0
      "0000" when "00101011110111", -- t[2807] = 0
      "0000" when "00101011111000", -- t[2808] = 0
      "0000" when "00101011111001", -- t[2809] = 0
      "0000" when "00101011111010", -- t[2810] = 0
      "0000" when "00101011111011", -- t[2811] = 0
      "0000" when "00101011111100", -- t[2812] = 0
      "0000" when "00101011111101", -- t[2813] = 0
      "0000" when "00101011111110", -- t[2814] = 0
      "0000" when "00101011111111", -- t[2815] = 0
      "0000" when "00101100000000", -- t[2816] = 0
      "0000" when "00101100000001", -- t[2817] = 0
      "0000" when "00101100000010", -- t[2818] = 0
      "0000" when "00101100000011", -- t[2819] = 0
      "0000" when "00101100000100", -- t[2820] = 0
      "0000" when "00101100000101", -- t[2821] = 0
      "0000" when "00101100000110", -- t[2822] = 0
      "0000" when "00101100000111", -- t[2823] = 0
      "0000" when "00101100001000", -- t[2824] = 0
      "0000" when "00101100001001", -- t[2825] = 0
      "0000" when "00101100001010", -- t[2826] = 0
      "0000" when "00101100001011", -- t[2827] = 0
      "0000" when "00101100001100", -- t[2828] = 0
      "0000" when "00101100001101", -- t[2829] = 0
      "0000" when "00101100001110", -- t[2830] = 0
      "0000" when "00101100001111", -- t[2831] = 0
      "0000" when "00101100010000", -- t[2832] = 0
      "0000" when "00101100010001", -- t[2833] = 0
      "0000" when "00101100010010", -- t[2834] = 0
      "0000" when "00101100010011", -- t[2835] = 0
      "0000" when "00101100010100", -- t[2836] = 0
      "0000" when "00101100010101", -- t[2837] = 0
      "0000" when "00101100010110", -- t[2838] = 0
      "0000" when "00101100010111", -- t[2839] = 0
      "0000" when "00101100011000", -- t[2840] = 0
      "0000" when "00101100011001", -- t[2841] = 0
      "0000" when "00101100011010", -- t[2842] = 0
      "0000" when "00101100011011", -- t[2843] = 0
      "0000" when "00101100011100", -- t[2844] = 0
      "0000" when "00101100011101", -- t[2845] = 0
      "0000" when "00101100011110", -- t[2846] = 0
      "0000" when "00101100011111", -- t[2847] = 0
      "0000" when "00101100100000", -- t[2848] = 0
      "0000" when "00101100100001", -- t[2849] = 0
      "0000" when "00101100100010", -- t[2850] = 0
      "0000" when "00101100100011", -- t[2851] = 0
      "0000" when "00101100100100", -- t[2852] = 0
      "0000" when "00101100100101", -- t[2853] = 0
      "0000" when "00101100100110", -- t[2854] = 0
      "0000" when "00101100100111", -- t[2855] = 0
      "0000" when "00101100101000", -- t[2856] = 0
      "0000" when "00101100101001", -- t[2857] = 0
      "0000" when "00101100101010", -- t[2858] = 0
      "0000" when "00101100101011", -- t[2859] = 0
      "0000" when "00101100101100", -- t[2860] = 0
      "0000" when "00101100101101", -- t[2861] = 0
      "0000" when "00101100101110", -- t[2862] = 0
      "0000" when "00101100101111", -- t[2863] = 0
      "0000" when "00101100110000", -- t[2864] = 0
      "0000" when "00101100110001", -- t[2865] = 0
      "0000" when "00101100110010", -- t[2866] = 0
      "0000" when "00101100110011", -- t[2867] = 0
      "0000" when "00101100110100", -- t[2868] = 0
      "0000" when "00101100110101", -- t[2869] = 0
      "0000" when "00101100110110", -- t[2870] = 0
      "0000" when "00101100110111", -- t[2871] = 0
      "0000" when "00101100111000", -- t[2872] = 0
      "0000" when "00101100111001", -- t[2873] = 0
      "0000" when "00101100111010", -- t[2874] = 0
      "0000" when "00101100111011", -- t[2875] = 0
      "0000" when "00101100111100", -- t[2876] = 0
      "0000" when "00101100111101", -- t[2877] = 0
      "0000" when "00101100111110", -- t[2878] = 0
      "0000" when "00101100111111", -- t[2879] = 0
      "0000" when "00101101000000", -- t[2880] = 0
      "0000" when "00101101000001", -- t[2881] = 0
      "0000" when "00101101000010", -- t[2882] = 0
      "0000" when "00101101000011", -- t[2883] = 0
      "0000" when "00101101000100", -- t[2884] = 0
      "0000" when "00101101000101", -- t[2885] = 0
      "0000" when "00101101000110", -- t[2886] = 0
      "0000" when "00101101000111", -- t[2887] = 0
      "0000" when "00101101001000", -- t[2888] = 0
      "0000" when "00101101001001", -- t[2889] = 0
      "0000" when "00101101001010", -- t[2890] = 0
      "0000" when "00101101001011", -- t[2891] = 0
      "0000" when "00101101001100", -- t[2892] = 0
      "0000" when "00101101001101", -- t[2893] = 0
      "0000" when "00101101001110", -- t[2894] = 0
      "0000" when "00101101001111", -- t[2895] = 0
      "0000" when "00101101010000", -- t[2896] = 0
      "0000" when "00101101010001", -- t[2897] = 0
      "0000" when "00101101010010", -- t[2898] = 0
      "0000" when "00101101010011", -- t[2899] = 0
      "0000" when "00101101010100", -- t[2900] = 0
      "0000" when "00101101010101", -- t[2901] = 0
      "0000" when "00101101010110", -- t[2902] = 0
      "0000" when "00101101010111", -- t[2903] = 0
      "0000" when "00101101011000", -- t[2904] = 0
      "0000" when "00101101011001", -- t[2905] = 0
      "0000" when "00101101011010", -- t[2906] = 0
      "0000" when "00101101011011", -- t[2907] = 0
      "0000" when "00101101011100", -- t[2908] = 0
      "0000" when "00101101011101", -- t[2909] = 0
      "0000" when "00101101011110", -- t[2910] = 0
      "0000" when "00101101011111", -- t[2911] = 0
      "0000" when "00101101100000", -- t[2912] = 0
      "0000" when "00101101100001", -- t[2913] = 0
      "0000" when "00101101100010", -- t[2914] = 0
      "0000" when "00101101100011", -- t[2915] = 0
      "0000" when "00101101100100", -- t[2916] = 0
      "0000" when "00101101100101", -- t[2917] = 0
      "0000" when "00101101100110", -- t[2918] = 0
      "0000" when "00101101100111", -- t[2919] = 0
      "0000" when "00101101101000", -- t[2920] = 0
      "0000" when "00101101101001", -- t[2921] = 0
      "0000" when "00101101101010", -- t[2922] = 0
      "0000" when "00101101101011", -- t[2923] = 0
      "0000" when "00101101101100", -- t[2924] = 0
      "0000" when "00101101101101", -- t[2925] = 0
      "0000" when "00101101101110", -- t[2926] = 0
      "0000" when "00101101101111", -- t[2927] = 0
      "0000" when "00101101110000", -- t[2928] = 0
      "0000" when "00101101110001", -- t[2929] = 0
      "0000" when "00101101110010", -- t[2930] = 0
      "0000" when "00101101110011", -- t[2931] = 0
      "0000" when "00101101110100", -- t[2932] = 0
      "0000" when "00101101110101", -- t[2933] = 0
      "0000" when "00101101110110", -- t[2934] = 0
      "0000" when "00101101110111", -- t[2935] = 0
      "0000" when "00101101111000", -- t[2936] = 0
      "0000" when "00101101111001", -- t[2937] = 0
      "0000" when "00101101111010", -- t[2938] = 0
      "0000" when "00101101111011", -- t[2939] = 0
      "0000" when "00101101111100", -- t[2940] = 0
      "0000" when "00101101111101", -- t[2941] = 0
      "0000" when "00101101111110", -- t[2942] = 0
      "0000" when "00101101111111", -- t[2943] = 0
      "0000" when "00101110000000", -- t[2944] = 0
      "0000" when "00101110000001", -- t[2945] = 0
      "0000" when "00101110000010", -- t[2946] = 0
      "0000" when "00101110000011", -- t[2947] = 0
      "0000" when "00101110000100", -- t[2948] = 0
      "0000" when "00101110000101", -- t[2949] = 0
      "0000" when "00101110000110", -- t[2950] = 0
      "0000" when "00101110000111", -- t[2951] = 0
      "0000" when "00101110001000", -- t[2952] = 0
      "0000" when "00101110001001", -- t[2953] = 0
      "0000" when "00101110001010", -- t[2954] = 0
      "0000" when "00101110001011", -- t[2955] = 0
      "0000" when "00101110001100", -- t[2956] = 0
      "0000" when "00101110001101", -- t[2957] = 0
      "0000" when "00101110001110", -- t[2958] = 0
      "0000" when "00101110001111", -- t[2959] = 0
      "0000" when "00101110010000", -- t[2960] = 0
      "0000" when "00101110010001", -- t[2961] = 0
      "0000" when "00101110010010", -- t[2962] = 0
      "0000" when "00101110010011", -- t[2963] = 0
      "0000" when "00101110010100", -- t[2964] = 0
      "0000" when "00101110010101", -- t[2965] = 0
      "0000" when "00101110010110", -- t[2966] = 0
      "0000" when "00101110010111", -- t[2967] = 0
      "0000" when "00101110011000", -- t[2968] = 0
      "0000" when "00101110011001", -- t[2969] = 0
      "0000" when "00101110011010", -- t[2970] = 0
      "0000" when "00101110011011", -- t[2971] = 0
      "0000" when "00101110011100", -- t[2972] = 0
      "0000" when "00101110011101", -- t[2973] = 0
      "0000" when "00101110011110", -- t[2974] = 0
      "0000" when "00101110011111", -- t[2975] = 0
      "0000" when "00101110100000", -- t[2976] = 0
      "0000" when "00101110100001", -- t[2977] = 0
      "0000" when "00101110100010", -- t[2978] = 0
      "0000" when "00101110100011", -- t[2979] = 0
      "0000" when "00101110100100", -- t[2980] = 0
      "0000" when "00101110100101", -- t[2981] = 0
      "0000" when "00101110100110", -- t[2982] = 0
      "0000" when "00101110100111", -- t[2983] = 0
      "0000" when "00101110101000", -- t[2984] = 0
      "0000" when "00101110101001", -- t[2985] = 0
      "0000" when "00101110101010", -- t[2986] = 0
      "0000" when "00101110101011", -- t[2987] = 0
      "0000" when "00101110101100", -- t[2988] = 0
      "0000" when "00101110101101", -- t[2989] = 0
      "0000" when "00101110101110", -- t[2990] = 0
      "0000" when "00101110101111", -- t[2991] = 0
      "0000" when "00101110110000", -- t[2992] = 0
      "0000" when "00101110110001", -- t[2993] = 0
      "0000" when "00101110110010", -- t[2994] = 0
      "0000" when "00101110110011", -- t[2995] = 0
      "0000" when "00101110110100", -- t[2996] = 0
      "0000" when "00101110110101", -- t[2997] = 0
      "0000" when "00101110110110", -- t[2998] = 0
      "0000" when "00101110110111", -- t[2999] = 0
      "0000" when "00101110111000", -- t[3000] = 0
      "0000" when "00101110111001", -- t[3001] = 0
      "0000" when "00101110111010", -- t[3002] = 0
      "0000" when "00101110111011", -- t[3003] = 0
      "0000" when "00101110111100", -- t[3004] = 0
      "0000" when "00101110111101", -- t[3005] = 0
      "0000" when "00101110111110", -- t[3006] = 0
      "0000" when "00101110111111", -- t[3007] = 0
      "0000" when "00101111000000", -- t[3008] = 0
      "0000" when "00101111000001", -- t[3009] = 0
      "0000" when "00101111000010", -- t[3010] = 0
      "0000" when "00101111000011", -- t[3011] = 0
      "0000" when "00101111000100", -- t[3012] = 0
      "0000" when "00101111000101", -- t[3013] = 0
      "0000" when "00101111000110", -- t[3014] = 0
      "0000" when "00101111000111", -- t[3015] = 0
      "0000" when "00101111001000", -- t[3016] = 0
      "0000" when "00101111001001", -- t[3017] = 0
      "0000" when "00101111001010", -- t[3018] = 0
      "0000" when "00101111001011", -- t[3019] = 0
      "0000" when "00101111001100", -- t[3020] = 0
      "0000" when "00101111001101", -- t[3021] = 0
      "0000" when "00101111001110", -- t[3022] = 0
      "0000" when "00101111001111", -- t[3023] = 0
      "0000" when "00101111010000", -- t[3024] = 0
      "0000" when "00101111010001", -- t[3025] = 0
      "0000" when "00101111010010", -- t[3026] = 0
      "0000" when "00101111010011", -- t[3027] = 0
      "0000" when "00101111010100", -- t[3028] = 0
      "0000" when "00101111010101", -- t[3029] = 0
      "0000" when "00101111010110", -- t[3030] = 0
      "0000" when "00101111010111", -- t[3031] = 0
      "0000" when "00101111011000", -- t[3032] = 0
      "0000" when "00101111011001", -- t[3033] = 0
      "0000" when "00101111011010", -- t[3034] = 0
      "0000" when "00101111011011", -- t[3035] = 0
      "0000" when "00101111011100", -- t[3036] = 0
      "0000" when "00101111011101", -- t[3037] = 0
      "0000" when "00101111011110", -- t[3038] = 0
      "0000" when "00101111011111", -- t[3039] = 0
      "0000" when "00101111100000", -- t[3040] = 0
      "0000" when "00101111100001", -- t[3041] = 0
      "0000" when "00101111100010", -- t[3042] = 0
      "0000" when "00101111100011", -- t[3043] = 0
      "0000" when "00101111100100", -- t[3044] = 0
      "0000" when "00101111100101", -- t[3045] = 0
      "0000" when "00101111100110", -- t[3046] = 0
      "0000" when "00101111100111", -- t[3047] = 0
      "0000" when "00101111101000", -- t[3048] = 0
      "0000" when "00101111101001", -- t[3049] = 0
      "0000" when "00101111101010", -- t[3050] = 0
      "0000" when "00101111101011", -- t[3051] = 0
      "0000" when "00101111101100", -- t[3052] = 0
      "0000" when "00101111101101", -- t[3053] = 0
      "0000" when "00101111101110", -- t[3054] = 0
      "0000" when "00101111101111", -- t[3055] = 0
      "0000" when "00101111110000", -- t[3056] = 0
      "0000" when "00101111110001", -- t[3057] = 0
      "0000" when "00101111110010", -- t[3058] = 0
      "0000" when "00101111110011", -- t[3059] = 0
      "0000" when "00101111110100", -- t[3060] = 0
      "0000" when "00101111110101", -- t[3061] = 0
      "0000" when "00101111110110", -- t[3062] = 0
      "0000" when "00101111110111", -- t[3063] = 0
      "0000" when "00101111111000", -- t[3064] = 0
      "0000" when "00101111111001", -- t[3065] = 0
      "0000" when "00101111111010", -- t[3066] = 0
      "0000" when "00101111111011", -- t[3067] = 0
      "0000" when "00101111111100", -- t[3068] = 0
      "0000" when "00101111111101", -- t[3069] = 0
      "0000" when "00101111111110", -- t[3070] = 0
      "0000" when "00101111111111", -- t[3071] = 0
      "0000" when "00110000000000", -- t[3072] = 0
      "0000" when "00110000000001", -- t[3073] = 0
      "0000" when "00110000000010", -- t[3074] = 0
      "0000" when "00110000000011", -- t[3075] = 0
      "0000" when "00110000000100", -- t[3076] = 0
      "0000" when "00110000000101", -- t[3077] = 0
      "0000" when "00110000000110", -- t[3078] = 0
      "0000" when "00110000000111", -- t[3079] = 0
      "0000" when "00110000001000", -- t[3080] = 0
      "0000" when "00110000001001", -- t[3081] = 0
      "0000" when "00110000001010", -- t[3082] = 0
      "0000" when "00110000001011", -- t[3083] = 0
      "0000" when "00110000001100", -- t[3084] = 0
      "0000" when "00110000001101", -- t[3085] = 0
      "0000" when "00110000001110", -- t[3086] = 0
      "0000" when "00110000001111", -- t[3087] = 0
      "0000" when "00110000010000", -- t[3088] = 0
      "0000" when "00110000010001", -- t[3089] = 0
      "0000" when "00110000010010", -- t[3090] = 0
      "0000" when "00110000010011", -- t[3091] = 0
      "0000" when "00110000010100", -- t[3092] = 0
      "0000" when "00110000010101", -- t[3093] = 0
      "0000" when "00110000010110", -- t[3094] = 0
      "0000" when "00110000010111", -- t[3095] = 0
      "0000" when "00110000011000", -- t[3096] = 0
      "0000" when "00110000011001", -- t[3097] = 0
      "0000" when "00110000011010", -- t[3098] = 0
      "0000" when "00110000011011", -- t[3099] = 0
      "0000" when "00110000011100", -- t[3100] = 0
      "0000" when "00110000011101", -- t[3101] = 0
      "0000" when "00110000011110", -- t[3102] = 0
      "0000" when "00110000011111", -- t[3103] = 0
      "0000" when "00110000100000", -- t[3104] = 0
      "0000" when "00110000100001", -- t[3105] = 0
      "0000" when "00110000100010", -- t[3106] = 0
      "0000" when "00110000100011", -- t[3107] = 0
      "0000" when "00110000100100", -- t[3108] = 0
      "0000" when "00110000100101", -- t[3109] = 0
      "0000" when "00110000100110", -- t[3110] = 0
      "0000" when "00110000100111", -- t[3111] = 0
      "0000" when "00110000101000", -- t[3112] = 0
      "0000" when "00110000101001", -- t[3113] = 0
      "0000" when "00110000101010", -- t[3114] = 0
      "0000" when "00110000101011", -- t[3115] = 0
      "0000" when "00110000101100", -- t[3116] = 0
      "0000" when "00110000101101", -- t[3117] = 0
      "0000" when "00110000101110", -- t[3118] = 0
      "0000" when "00110000101111", -- t[3119] = 0
      "0000" when "00110000110000", -- t[3120] = 0
      "0000" when "00110000110001", -- t[3121] = 0
      "0000" when "00110000110010", -- t[3122] = 0
      "0000" when "00110000110011", -- t[3123] = 0
      "0000" when "00110000110100", -- t[3124] = 0
      "0000" when "00110000110101", -- t[3125] = 0
      "0000" when "00110000110110", -- t[3126] = 0
      "0000" when "00110000110111", -- t[3127] = 0
      "0000" when "00110000111000", -- t[3128] = 0
      "0000" when "00110000111001", -- t[3129] = 0
      "0000" when "00110000111010", -- t[3130] = 0
      "0000" when "00110000111011", -- t[3131] = 0
      "0000" when "00110000111100", -- t[3132] = 0
      "0000" when "00110000111101", -- t[3133] = 0
      "0000" when "00110000111110", -- t[3134] = 0
      "0000" when "00110000111111", -- t[3135] = 0
      "0000" when "00110001000000", -- t[3136] = 0
      "0000" when "00110001000001", -- t[3137] = 0
      "0000" when "00110001000010", -- t[3138] = 0
      "0000" when "00110001000011", -- t[3139] = 0
      "0000" when "00110001000100", -- t[3140] = 0
      "0000" when "00110001000101", -- t[3141] = 0
      "0000" when "00110001000110", -- t[3142] = 0
      "0000" when "00110001000111", -- t[3143] = 0
      "0000" when "00110001001000", -- t[3144] = 0
      "0000" when "00110001001001", -- t[3145] = 0
      "0000" when "00110001001010", -- t[3146] = 0
      "0000" when "00110001001011", -- t[3147] = 0
      "0000" when "00110001001100", -- t[3148] = 0
      "0000" when "00110001001101", -- t[3149] = 0
      "0000" when "00110001001110", -- t[3150] = 0
      "0000" when "00110001001111", -- t[3151] = 0
      "0000" when "00110001010000", -- t[3152] = 0
      "0000" when "00110001010001", -- t[3153] = 0
      "0000" when "00110001010010", -- t[3154] = 0
      "0000" when "00110001010011", -- t[3155] = 0
      "0000" when "00110001010100", -- t[3156] = 0
      "0000" when "00110001010101", -- t[3157] = 0
      "0000" when "00110001010110", -- t[3158] = 0
      "0000" when "00110001010111", -- t[3159] = 0
      "0000" when "00110001011000", -- t[3160] = 0
      "0000" when "00110001011001", -- t[3161] = 0
      "0000" when "00110001011010", -- t[3162] = 0
      "0000" when "00110001011011", -- t[3163] = 0
      "0000" when "00110001011100", -- t[3164] = 0
      "0000" when "00110001011101", -- t[3165] = 0
      "0000" when "00110001011110", -- t[3166] = 0
      "0000" when "00110001011111", -- t[3167] = 0
      "0000" when "00110001100000", -- t[3168] = 0
      "0000" when "00110001100001", -- t[3169] = 0
      "0000" when "00110001100010", -- t[3170] = 0
      "0000" when "00110001100011", -- t[3171] = 0
      "0000" when "00110001100100", -- t[3172] = 0
      "0000" when "00110001100101", -- t[3173] = 0
      "0000" when "00110001100110", -- t[3174] = 0
      "0000" when "00110001100111", -- t[3175] = 0
      "0000" when "00110001101000", -- t[3176] = 0
      "0000" when "00110001101001", -- t[3177] = 0
      "0000" when "00110001101010", -- t[3178] = 0
      "0000" when "00110001101011", -- t[3179] = 0
      "0000" when "00110001101100", -- t[3180] = 0
      "0000" when "00110001101101", -- t[3181] = 0
      "0000" when "00110001101110", -- t[3182] = 0
      "0000" when "00110001101111", -- t[3183] = 0
      "0000" when "00110001110000", -- t[3184] = 0
      "0000" when "00110001110001", -- t[3185] = 0
      "0000" when "00110001110010", -- t[3186] = 0
      "0000" when "00110001110011", -- t[3187] = 0
      "0000" when "00110001110100", -- t[3188] = 0
      "0000" when "00110001110101", -- t[3189] = 0
      "0000" when "00110001110110", -- t[3190] = 0
      "0000" when "00110001110111", -- t[3191] = 0
      "0000" when "00110001111000", -- t[3192] = 0
      "0000" when "00110001111001", -- t[3193] = 0
      "0000" when "00110001111010", -- t[3194] = 0
      "0000" when "00110001111011", -- t[3195] = 0
      "0000" when "00110001111100", -- t[3196] = 0
      "0000" when "00110001111101", -- t[3197] = 0
      "0000" when "00110001111110", -- t[3198] = 0
      "0000" when "00110001111111", -- t[3199] = 0
      "0000" when "00110010000000", -- t[3200] = 0
      "0000" when "00110010000001", -- t[3201] = 0
      "0000" when "00110010000010", -- t[3202] = 0
      "0000" when "00110010000011", -- t[3203] = 0
      "0000" when "00110010000100", -- t[3204] = 0
      "0000" when "00110010000101", -- t[3205] = 0
      "0000" when "00110010000110", -- t[3206] = 0
      "0000" when "00110010000111", -- t[3207] = 0
      "0000" when "00110010001000", -- t[3208] = 0
      "0000" when "00110010001001", -- t[3209] = 0
      "0000" when "00110010001010", -- t[3210] = 0
      "0000" when "00110010001011", -- t[3211] = 0
      "0000" when "00110010001100", -- t[3212] = 0
      "0000" when "00110010001101", -- t[3213] = 0
      "0000" when "00110010001110", -- t[3214] = 0
      "0000" when "00110010001111", -- t[3215] = 0
      "0000" when "00110010010000", -- t[3216] = 0
      "0000" when "00110010010001", -- t[3217] = 0
      "0000" when "00110010010010", -- t[3218] = 0
      "0000" when "00110010010011", -- t[3219] = 0
      "0000" when "00110010010100", -- t[3220] = 0
      "0000" when "00110010010101", -- t[3221] = 0
      "0000" when "00110010010110", -- t[3222] = 0
      "0000" when "00110010010111", -- t[3223] = 0
      "0000" when "00110010011000", -- t[3224] = 0
      "0000" when "00110010011001", -- t[3225] = 0
      "0000" when "00110010011010", -- t[3226] = 0
      "0000" when "00110010011011", -- t[3227] = 0
      "0000" when "00110010011100", -- t[3228] = 0
      "0000" when "00110010011101", -- t[3229] = 0
      "0000" when "00110010011110", -- t[3230] = 0
      "0000" when "00110010011111", -- t[3231] = 0
      "0000" when "00110010100000", -- t[3232] = 0
      "0000" when "00110010100001", -- t[3233] = 0
      "0000" when "00110010100010", -- t[3234] = 0
      "0000" when "00110010100011", -- t[3235] = 0
      "0000" when "00110010100100", -- t[3236] = 0
      "0000" when "00110010100101", -- t[3237] = 0
      "0000" when "00110010100110", -- t[3238] = 0
      "0000" when "00110010100111", -- t[3239] = 0
      "0000" when "00110010101000", -- t[3240] = 0
      "0000" when "00110010101001", -- t[3241] = 0
      "0000" when "00110010101010", -- t[3242] = 0
      "0000" when "00110010101011", -- t[3243] = 0
      "0000" when "00110010101100", -- t[3244] = 0
      "0000" when "00110010101101", -- t[3245] = 0
      "0000" when "00110010101110", -- t[3246] = 0
      "0000" when "00110010101111", -- t[3247] = 0
      "0000" when "00110010110000", -- t[3248] = 0
      "0000" when "00110010110001", -- t[3249] = 0
      "0000" when "00110010110010", -- t[3250] = 0
      "0000" when "00110010110011", -- t[3251] = 0
      "0000" when "00110010110100", -- t[3252] = 0
      "0000" when "00110010110101", -- t[3253] = 0
      "0000" when "00110010110110", -- t[3254] = 0
      "0000" when "00110010110111", -- t[3255] = 0
      "0000" when "00110010111000", -- t[3256] = 0
      "0000" when "00110010111001", -- t[3257] = 0
      "0000" when "00110010111010", -- t[3258] = 0
      "0000" when "00110010111011", -- t[3259] = 0
      "0000" when "00110010111100", -- t[3260] = 0
      "0000" when "00110010111101", -- t[3261] = 0
      "0000" when "00110010111110", -- t[3262] = 0
      "0000" when "00110010111111", -- t[3263] = 0
      "0000" when "00110011000000", -- t[3264] = 0
      "0000" when "00110011000001", -- t[3265] = 0
      "0000" when "00110011000010", -- t[3266] = 0
      "0000" when "00110011000011", -- t[3267] = 0
      "0000" when "00110011000100", -- t[3268] = 0
      "0000" when "00110011000101", -- t[3269] = 0
      "0000" when "00110011000110", -- t[3270] = 0
      "0000" when "00110011000111", -- t[3271] = 0
      "0000" when "00110011001000", -- t[3272] = 0
      "0000" when "00110011001001", -- t[3273] = 0
      "0000" when "00110011001010", -- t[3274] = 0
      "0000" when "00110011001011", -- t[3275] = 0
      "0000" when "00110011001100", -- t[3276] = 0
      "0000" when "00110011001101", -- t[3277] = 0
      "0000" when "00110011001110", -- t[3278] = 0
      "0000" when "00110011001111", -- t[3279] = 0
      "0000" when "00110011010000", -- t[3280] = 0
      "0000" when "00110011010001", -- t[3281] = 0
      "0000" when "00110011010010", -- t[3282] = 0
      "0000" when "00110011010011", -- t[3283] = 0
      "0000" when "00110011010100", -- t[3284] = 0
      "0000" when "00110011010101", -- t[3285] = 0
      "0000" when "00110011010110", -- t[3286] = 0
      "0000" when "00110011010111", -- t[3287] = 0
      "0000" when "00110011011000", -- t[3288] = 0
      "0000" when "00110011011001", -- t[3289] = 0
      "0000" when "00110011011010", -- t[3290] = 0
      "0000" when "00110011011011", -- t[3291] = 0
      "0000" when "00110011011100", -- t[3292] = 0
      "0000" when "00110011011101", -- t[3293] = 0
      "0000" when "00110011011110", -- t[3294] = 0
      "0000" when "00110011011111", -- t[3295] = 0
      "0000" when "00110011100000", -- t[3296] = 0
      "0000" when "00110011100001", -- t[3297] = 0
      "0000" when "00110011100010", -- t[3298] = 0
      "0000" when "00110011100011", -- t[3299] = 0
      "0000" when "00110011100100", -- t[3300] = 0
      "0000" when "00110011100101", -- t[3301] = 0
      "0000" when "00110011100110", -- t[3302] = 0
      "0000" when "00110011100111", -- t[3303] = 0
      "0000" when "00110011101000", -- t[3304] = 0
      "0000" when "00110011101001", -- t[3305] = 0
      "0000" when "00110011101010", -- t[3306] = 0
      "0000" when "00110011101011", -- t[3307] = 0
      "0000" when "00110011101100", -- t[3308] = 0
      "0000" when "00110011101101", -- t[3309] = 0
      "0000" when "00110011101110", -- t[3310] = 0
      "0000" when "00110011101111", -- t[3311] = 0
      "0000" when "00110011110000", -- t[3312] = 0
      "0000" when "00110011110001", -- t[3313] = 0
      "0000" when "00110011110010", -- t[3314] = 0
      "0000" when "00110011110011", -- t[3315] = 0
      "0000" when "00110011110100", -- t[3316] = 0
      "0000" when "00110011110101", -- t[3317] = 0
      "0000" when "00110011110110", -- t[3318] = 0
      "0000" when "00110011110111", -- t[3319] = 0
      "0000" when "00110011111000", -- t[3320] = 0
      "0000" when "00110011111001", -- t[3321] = 0
      "0000" when "00110011111010", -- t[3322] = 0
      "0000" when "00110011111011", -- t[3323] = 0
      "0000" when "00110011111100", -- t[3324] = 0
      "0000" when "00110011111101", -- t[3325] = 0
      "0000" when "00110011111110", -- t[3326] = 0
      "0000" when "00110011111111", -- t[3327] = 0
      "0000" when "00110100000000", -- t[3328] = 0
      "0000" when "00110100000001", -- t[3329] = 0
      "0000" when "00110100000010", -- t[3330] = 0
      "0000" when "00110100000011", -- t[3331] = 0
      "0000" when "00110100000100", -- t[3332] = 0
      "0000" when "00110100000101", -- t[3333] = 0
      "0000" when "00110100000110", -- t[3334] = 0
      "0000" when "00110100000111", -- t[3335] = 0
      "0000" when "00110100001000", -- t[3336] = 0
      "0000" when "00110100001001", -- t[3337] = 0
      "0000" when "00110100001010", -- t[3338] = 0
      "0000" when "00110100001011", -- t[3339] = 0
      "0000" when "00110100001100", -- t[3340] = 0
      "0000" when "00110100001101", -- t[3341] = 0
      "0000" when "00110100001110", -- t[3342] = 0
      "0000" when "00110100001111", -- t[3343] = 0
      "0000" when "00110100010000", -- t[3344] = 0
      "0000" when "00110100010001", -- t[3345] = 0
      "0000" when "00110100010010", -- t[3346] = 0
      "0000" when "00110100010011", -- t[3347] = 0
      "0000" when "00110100010100", -- t[3348] = 0
      "0000" when "00110100010101", -- t[3349] = 0
      "0000" when "00110100010110", -- t[3350] = 0
      "0000" when "00110100010111", -- t[3351] = 0
      "0000" when "00110100011000", -- t[3352] = 0
      "0000" when "00110100011001", -- t[3353] = 0
      "0000" when "00110100011010", -- t[3354] = 0
      "0000" when "00110100011011", -- t[3355] = 0
      "0000" when "00110100011100", -- t[3356] = 0
      "0000" when "00110100011101", -- t[3357] = 0
      "0000" when "00110100011110", -- t[3358] = 0
      "0000" when "00110100011111", -- t[3359] = 0
      "0000" when "00110100100000", -- t[3360] = 0
      "0000" when "00110100100001", -- t[3361] = 0
      "0000" when "00110100100010", -- t[3362] = 0
      "0000" when "00110100100011", -- t[3363] = 0
      "0000" when "00110100100100", -- t[3364] = 0
      "0000" when "00110100100101", -- t[3365] = 0
      "0000" when "00110100100110", -- t[3366] = 0
      "0000" when "00110100100111", -- t[3367] = 0
      "0000" when "00110100101000", -- t[3368] = 0
      "0000" when "00110100101001", -- t[3369] = 0
      "0000" when "00110100101010", -- t[3370] = 0
      "0000" when "00110100101011", -- t[3371] = 0
      "0000" when "00110100101100", -- t[3372] = 0
      "0000" when "00110100101101", -- t[3373] = 0
      "0000" when "00110100101110", -- t[3374] = 0
      "0000" when "00110100101111", -- t[3375] = 0
      "0000" when "00110100110000", -- t[3376] = 0
      "0000" when "00110100110001", -- t[3377] = 0
      "0000" when "00110100110010", -- t[3378] = 0
      "0000" when "00110100110011", -- t[3379] = 0
      "0000" when "00110100110100", -- t[3380] = 0
      "0000" when "00110100110101", -- t[3381] = 0
      "0000" when "00110100110110", -- t[3382] = 0
      "0000" when "00110100110111", -- t[3383] = 0
      "0000" when "00110100111000", -- t[3384] = 0
      "0000" when "00110100111001", -- t[3385] = 0
      "0000" when "00110100111010", -- t[3386] = 0
      "0000" when "00110100111011", -- t[3387] = 0
      "0000" when "00110100111100", -- t[3388] = 0
      "0000" when "00110100111101", -- t[3389] = 0
      "0000" when "00110100111110", -- t[3390] = 0
      "0000" when "00110100111111", -- t[3391] = 0
      "0000" when "00110101000000", -- t[3392] = 0
      "0000" when "00110101000001", -- t[3393] = 0
      "0000" when "00110101000010", -- t[3394] = 0
      "0000" when "00110101000011", -- t[3395] = 0
      "0000" when "00110101000100", -- t[3396] = 0
      "0000" when "00110101000101", -- t[3397] = 0
      "0000" when "00110101000110", -- t[3398] = 0
      "0000" when "00110101000111", -- t[3399] = 0
      "0000" when "00110101001000", -- t[3400] = 0
      "0000" when "00110101001001", -- t[3401] = 0
      "0000" when "00110101001010", -- t[3402] = 0
      "0000" when "00110101001011", -- t[3403] = 0
      "0000" when "00110101001100", -- t[3404] = 0
      "0000" when "00110101001101", -- t[3405] = 0
      "0000" when "00110101001110", -- t[3406] = 0
      "0000" when "00110101001111", -- t[3407] = 0
      "0000" when "00110101010000", -- t[3408] = 0
      "0000" when "00110101010001", -- t[3409] = 0
      "0000" when "00110101010010", -- t[3410] = 0
      "0000" when "00110101010011", -- t[3411] = 0
      "0000" when "00110101010100", -- t[3412] = 0
      "0000" when "00110101010101", -- t[3413] = 0
      "0000" when "00110101010110", -- t[3414] = 0
      "0000" when "00110101010111", -- t[3415] = 0
      "0000" when "00110101011000", -- t[3416] = 0
      "0000" when "00110101011001", -- t[3417] = 0
      "0000" when "00110101011010", -- t[3418] = 0
      "0000" when "00110101011011", -- t[3419] = 0
      "0000" when "00110101011100", -- t[3420] = 0
      "0000" when "00110101011101", -- t[3421] = 0
      "0000" when "00110101011110", -- t[3422] = 0
      "0000" when "00110101011111", -- t[3423] = 0
      "0000" when "00110101100000", -- t[3424] = 0
      "0000" when "00110101100001", -- t[3425] = 0
      "0000" when "00110101100010", -- t[3426] = 0
      "0000" when "00110101100011", -- t[3427] = 0
      "0000" when "00110101100100", -- t[3428] = 0
      "0000" when "00110101100101", -- t[3429] = 0
      "0000" when "00110101100110", -- t[3430] = 0
      "0000" when "00110101100111", -- t[3431] = 0
      "0000" when "00110101101000", -- t[3432] = 0
      "0000" when "00110101101001", -- t[3433] = 0
      "0000" when "00110101101010", -- t[3434] = 0
      "0000" when "00110101101011", -- t[3435] = 0
      "0000" when "00110101101100", -- t[3436] = 0
      "0000" when "00110101101101", -- t[3437] = 0
      "0000" when "00110101101110", -- t[3438] = 0
      "0000" when "00110101101111", -- t[3439] = 0
      "0000" when "00110101110000", -- t[3440] = 0
      "0000" when "00110101110001", -- t[3441] = 0
      "0000" when "00110101110010", -- t[3442] = 0
      "0000" when "00110101110011", -- t[3443] = 0
      "0000" when "00110101110100", -- t[3444] = 0
      "0000" when "00110101110101", -- t[3445] = 0
      "0000" when "00110101110110", -- t[3446] = 0
      "0000" when "00110101110111", -- t[3447] = 0
      "0000" when "00110101111000", -- t[3448] = 0
      "0000" when "00110101111001", -- t[3449] = 0
      "0000" when "00110101111010", -- t[3450] = 0
      "0000" when "00110101111011", -- t[3451] = 0
      "0000" when "00110101111100", -- t[3452] = 0
      "0000" when "00110101111101", -- t[3453] = 0
      "0000" when "00110101111110", -- t[3454] = 0
      "0000" when "00110101111111", -- t[3455] = 0
      "0000" when "00110110000000", -- t[3456] = 0
      "0000" when "00110110000001", -- t[3457] = 0
      "0000" when "00110110000010", -- t[3458] = 0
      "0000" when "00110110000011", -- t[3459] = 0
      "0000" when "00110110000100", -- t[3460] = 0
      "0000" when "00110110000101", -- t[3461] = 0
      "0000" when "00110110000110", -- t[3462] = 0
      "0000" when "00110110000111", -- t[3463] = 0
      "0000" when "00110110001000", -- t[3464] = 0
      "0000" when "00110110001001", -- t[3465] = 0
      "0000" when "00110110001010", -- t[3466] = 0
      "0000" when "00110110001011", -- t[3467] = 0
      "0000" when "00110110001100", -- t[3468] = 0
      "0000" when "00110110001101", -- t[3469] = 0
      "0000" when "00110110001110", -- t[3470] = 0
      "0000" when "00110110001111", -- t[3471] = 0
      "0000" when "00110110010000", -- t[3472] = 0
      "0000" when "00110110010001", -- t[3473] = 0
      "0000" when "00110110010010", -- t[3474] = 0
      "0000" when "00110110010011", -- t[3475] = 0
      "0000" when "00110110010100", -- t[3476] = 0
      "0000" when "00110110010101", -- t[3477] = 0
      "0000" when "00110110010110", -- t[3478] = 0
      "0000" when "00110110010111", -- t[3479] = 0
      "0000" when "00110110011000", -- t[3480] = 0
      "0000" when "00110110011001", -- t[3481] = 0
      "0000" when "00110110011010", -- t[3482] = 0
      "0000" when "00110110011011", -- t[3483] = 0
      "0000" when "00110110011100", -- t[3484] = 0
      "0000" when "00110110011101", -- t[3485] = 0
      "0000" when "00110110011110", -- t[3486] = 0
      "0000" when "00110110011111", -- t[3487] = 0
      "0000" when "00110110100000", -- t[3488] = 0
      "0000" when "00110110100001", -- t[3489] = 0
      "0000" when "00110110100010", -- t[3490] = 0
      "0000" when "00110110100011", -- t[3491] = 0
      "0000" when "00110110100100", -- t[3492] = 0
      "0000" when "00110110100101", -- t[3493] = 0
      "0000" when "00110110100110", -- t[3494] = 0
      "0000" when "00110110100111", -- t[3495] = 0
      "0000" when "00110110101000", -- t[3496] = 0
      "0000" when "00110110101001", -- t[3497] = 0
      "0000" when "00110110101010", -- t[3498] = 0
      "0000" when "00110110101011", -- t[3499] = 0
      "0000" when "00110110101100", -- t[3500] = 0
      "0000" when "00110110101101", -- t[3501] = 0
      "0000" when "00110110101110", -- t[3502] = 0
      "0000" when "00110110101111", -- t[3503] = 0
      "0000" when "00110110110000", -- t[3504] = 0
      "0000" when "00110110110001", -- t[3505] = 0
      "0000" when "00110110110010", -- t[3506] = 0
      "0000" when "00110110110011", -- t[3507] = 0
      "0000" when "00110110110100", -- t[3508] = 0
      "0000" when "00110110110101", -- t[3509] = 0
      "0000" when "00110110110110", -- t[3510] = 0
      "0000" when "00110110110111", -- t[3511] = 0
      "0000" when "00110110111000", -- t[3512] = 0
      "0000" when "00110110111001", -- t[3513] = 0
      "0000" when "00110110111010", -- t[3514] = 0
      "0000" when "00110110111011", -- t[3515] = 0
      "0000" when "00110110111100", -- t[3516] = 0
      "0000" when "00110110111101", -- t[3517] = 0
      "0000" when "00110110111110", -- t[3518] = 0
      "0000" when "00110110111111", -- t[3519] = 0
      "0000" when "00110111000000", -- t[3520] = 0
      "0000" when "00110111000001", -- t[3521] = 0
      "0000" when "00110111000010", -- t[3522] = 0
      "0000" when "00110111000011", -- t[3523] = 0
      "0000" when "00110111000100", -- t[3524] = 0
      "0000" when "00110111000101", -- t[3525] = 0
      "0000" when "00110111000110", -- t[3526] = 0
      "0000" when "00110111000111", -- t[3527] = 0
      "0000" when "00110111001000", -- t[3528] = 0
      "0000" when "00110111001001", -- t[3529] = 0
      "0000" when "00110111001010", -- t[3530] = 0
      "0000" when "00110111001011", -- t[3531] = 0
      "0000" when "00110111001100", -- t[3532] = 0
      "0000" when "00110111001101", -- t[3533] = 0
      "0000" when "00110111001110", -- t[3534] = 0
      "0000" when "00110111001111", -- t[3535] = 0
      "0000" when "00110111010000", -- t[3536] = 0
      "0000" when "00110111010001", -- t[3537] = 0
      "0000" when "00110111010010", -- t[3538] = 0
      "0000" when "00110111010011", -- t[3539] = 0
      "0000" when "00110111010100", -- t[3540] = 0
      "0000" when "00110111010101", -- t[3541] = 0
      "0000" when "00110111010110", -- t[3542] = 0
      "0000" when "00110111010111", -- t[3543] = 0
      "0000" when "00110111011000", -- t[3544] = 0
      "0000" when "00110111011001", -- t[3545] = 0
      "0000" when "00110111011010", -- t[3546] = 0
      "0000" when "00110111011011", -- t[3547] = 0
      "0000" when "00110111011100", -- t[3548] = 0
      "0000" when "00110111011101", -- t[3549] = 0
      "0000" when "00110111011110", -- t[3550] = 0
      "0000" when "00110111011111", -- t[3551] = 0
      "0000" when "00110111100000", -- t[3552] = 0
      "0000" when "00110111100001", -- t[3553] = 0
      "0000" when "00110111100010", -- t[3554] = 0
      "0000" when "00110111100011", -- t[3555] = 0
      "0000" when "00110111100100", -- t[3556] = 0
      "0000" when "00110111100101", -- t[3557] = 0
      "0000" when "00110111100110", -- t[3558] = 0
      "0000" when "00110111100111", -- t[3559] = 0
      "0000" when "00110111101000", -- t[3560] = 0
      "0000" when "00110111101001", -- t[3561] = 0
      "0000" when "00110111101010", -- t[3562] = 0
      "0000" when "00110111101011", -- t[3563] = 0
      "0000" when "00110111101100", -- t[3564] = 0
      "0000" when "00110111101101", -- t[3565] = 0
      "0000" when "00110111101110", -- t[3566] = 0
      "0000" when "00110111101111", -- t[3567] = 0
      "0000" when "00110111110000", -- t[3568] = 0
      "0000" when "00110111110001", -- t[3569] = 0
      "0000" when "00110111110010", -- t[3570] = 0
      "0000" when "00110111110011", -- t[3571] = 0
      "0000" when "00110111110100", -- t[3572] = 0
      "0000" when "00110111110101", -- t[3573] = 0
      "0000" when "00110111110110", -- t[3574] = 0
      "0000" when "00110111110111", -- t[3575] = 0
      "0000" when "00110111111000", -- t[3576] = 0
      "0000" when "00110111111001", -- t[3577] = 0
      "0000" when "00110111111010", -- t[3578] = 0
      "0000" when "00110111111011", -- t[3579] = 0
      "0000" when "00110111111100", -- t[3580] = 0
      "0000" when "00110111111101", -- t[3581] = 0
      "0000" when "00110111111110", -- t[3582] = 0
      "0000" when "00110111111111", -- t[3583] = 0
      "0000" when "00111000000000", -- t[3584] = 0
      "0000" when "00111000000001", -- t[3585] = 0
      "0000" when "00111000000010", -- t[3586] = 0
      "0000" when "00111000000011", -- t[3587] = 0
      "0000" when "00111000000100", -- t[3588] = 0
      "0000" when "00111000000101", -- t[3589] = 0
      "0000" when "00111000000110", -- t[3590] = 0
      "0000" when "00111000000111", -- t[3591] = 0
      "0000" when "00111000001000", -- t[3592] = 0
      "0000" when "00111000001001", -- t[3593] = 0
      "0000" when "00111000001010", -- t[3594] = 0
      "0000" when "00111000001011", -- t[3595] = 0
      "0000" when "00111000001100", -- t[3596] = 0
      "0000" when "00111000001101", -- t[3597] = 0
      "0000" when "00111000001110", -- t[3598] = 0
      "0000" when "00111000001111", -- t[3599] = 0
      "0000" when "00111000010000", -- t[3600] = 0
      "0000" when "00111000010001", -- t[3601] = 0
      "0000" when "00111000010010", -- t[3602] = 0
      "0000" when "00111000010011", -- t[3603] = 0
      "0000" when "00111000010100", -- t[3604] = 0
      "0000" when "00111000010101", -- t[3605] = 0
      "0000" when "00111000010110", -- t[3606] = 0
      "0000" when "00111000010111", -- t[3607] = 0
      "0000" when "00111000011000", -- t[3608] = 0
      "0000" when "00111000011001", -- t[3609] = 0
      "0000" when "00111000011010", -- t[3610] = 0
      "0000" when "00111000011011", -- t[3611] = 0
      "0000" when "00111000011100", -- t[3612] = 0
      "0000" when "00111000011101", -- t[3613] = 0
      "0000" when "00111000011110", -- t[3614] = 0
      "0000" when "00111000011111", -- t[3615] = 0
      "0000" when "00111000100000", -- t[3616] = 0
      "0000" when "00111000100001", -- t[3617] = 0
      "0000" when "00111000100010", -- t[3618] = 0
      "0000" when "00111000100011", -- t[3619] = 0
      "0000" when "00111000100100", -- t[3620] = 0
      "0000" when "00111000100101", -- t[3621] = 0
      "0000" when "00111000100110", -- t[3622] = 0
      "0000" when "00111000100111", -- t[3623] = 0
      "0000" when "00111000101000", -- t[3624] = 0
      "0000" when "00111000101001", -- t[3625] = 0
      "0000" when "00111000101010", -- t[3626] = 0
      "0000" when "00111000101011", -- t[3627] = 0
      "0000" when "00111000101100", -- t[3628] = 0
      "0000" when "00111000101101", -- t[3629] = 0
      "0000" when "00111000101110", -- t[3630] = 0
      "0000" when "00111000101111", -- t[3631] = 0
      "0000" when "00111000110000", -- t[3632] = 0
      "0000" when "00111000110001", -- t[3633] = 0
      "0000" when "00111000110010", -- t[3634] = 0
      "0000" when "00111000110011", -- t[3635] = 0
      "0000" when "00111000110100", -- t[3636] = 0
      "0000" when "00111000110101", -- t[3637] = 0
      "0000" when "00111000110110", -- t[3638] = 0
      "0000" when "00111000110111", -- t[3639] = 0
      "0000" when "00111000111000", -- t[3640] = 0
      "0000" when "00111000111001", -- t[3641] = 0
      "0000" when "00111000111010", -- t[3642] = 0
      "0000" when "00111000111011", -- t[3643] = 0
      "0000" when "00111000111100", -- t[3644] = 0
      "0000" when "00111000111101", -- t[3645] = 0
      "0000" when "00111000111110", -- t[3646] = 0
      "0000" when "00111000111111", -- t[3647] = 0
      "0000" when "00111001000000", -- t[3648] = 0
      "0000" when "00111001000001", -- t[3649] = 0
      "0000" when "00111001000010", -- t[3650] = 0
      "0000" when "00111001000011", -- t[3651] = 0
      "0000" when "00111001000100", -- t[3652] = 0
      "0000" when "00111001000101", -- t[3653] = 0
      "0000" when "00111001000110", -- t[3654] = 0
      "0000" when "00111001000111", -- t[3655] = 0
      "0000" when "00111001001000", -- t[3656] = 0
      "0000" when "00111001001001", -- t[3657] = 0
      "0000" when "00111001001010", -- t[3658] = 0
      "0000" when "00111001001011", -- t[3659] = 0
      "0000" when "00111001001100", -- t[3660] = 0
      "0000" when "00111001001101", -- t[3661] = 0
      "0000" when "00111001001110", -- t[3662] = 0
      "0000" when "00111001001111", -- t[3663] = 0
      "0000" when "00111001010000", -- t[3664] = 0
      "0000" when "00111001010001", -- t[3665] = 0
      "0000" when "00111001010010", -- t[3666] = 0
      "0000" when "00111001010011", -- t[3667] = 0
      "0000" when "00111001010100", -- t[3668] = 0
      "0000" when "00111001010101", -- t[3669] = 0
      "0000" when "00111001010110", -- t[3670] = 0
      "0000" when "00111001010111", -- t[3671] = 0
      "0000" when "00111001011000", -- t[3672] = 0
      "0000" when "00111001011001", -- t[3673] = 0
      "0000" when "00111001011010", -- t[3674] = 0
      "0000" when "00111001011011", -- t[3675] = 0
      "0000" when "00111001011100", -- t[3676] = 0
      "0000" when "00111001011101", -- t[3677] = 0
      "0000" when "00111001011110", -- t[3678] = 0
      "0000" when "00111001011111", -- t[3679] = 0
      "0000" when "00111001100000", -- t[3680] = 0
      "0000" when "00111001100001", -- t[3681] = 0
      "0000" when "00111001100010", -- t[3682] = 0
      "0000" when "00111001100011", -- t[3683] = 0
      "0000" when "00111001100100", -- t[3684] = 0
      "0000" when "00111001100101", -- t[3685] = 0
      "0000" when "00111001100110", -- t[3686] = 0
      "0000" when "00111001100111", -- t[3687] = 0
      "0000" when "00111001101000", -- t[3688] = 0
      "0000" when "00111001101001", -- t[3689] = 0
      "0000" when "00111001101010", -- t[3690] = 0
      "0000" when "00111001101011", -- t[3691] = 0
      "0000" when "00111001101100", -- t[3692] = 0
      "0000" when "00111001101101", -- t[3693] = 0
      "0000" when "00111001101110", -- t[3694] = 0
      "0000" when "00111001101111", -- t[3695] = 0
      "0000" when "00111001110000", -- t[3696] = 0
      "0000" when "00111001110001", -- t[3697] = 0
      "0000" when "00111001110010", -- t[3698] = 0
      "0000" when "00111001110011", -- t[3699] = 0
      "0000" when "00111001110100", -- t[3700] = 0
      "0000" when "00111001110101", -- t[3701] = 0
      "0000" when "00111001110110", -- t[3702] = 0
      "0000" when "00111001110111", -- t[3703] = 0
      "0000" when "00111001111000", -- t[3704] = 0
      "0000" when "00111001111001", -- t[3705] = 0
      "0000" when "00111001111010", -- t[3706] = 0
      "0000" when "00111001111011", -- t[3707] = 0
      "0000" when "00111001111100", -- t[3708] = 0
      "0000" when "00111001111101", -- t[3709] = 0
      "0000" when "00111001111110", -- t[3710] = 0
      "0000" when "00111001111111", -- t[3711] = 0
      "0000" when "00111010000000", -- t[3712] = 0
      "0000" when "00111010000001", -- t[3713] = 0
      "0000" when "00111010000010", -- t[3714] = 0
      "0000" when "00111010000011", -- t[3715] = 0
      "0000" when "00111010000100", -- t[3716] = 0
      "0000" when "00111010000101", -- t[3717] = 0
      "0000" when "00111010000110", -- t[3718] = 0
      "0000" when "00111010000111", -- t[3719] = 0
      "0000" when "00111010001000", -- t[3720] = 0
      "0000" when "00111010001001", -- t[3721] = 0
      "0000" when "00111010001010", -- t[3722] = 0
      "0000" when "00111010001011", -- t[3723] = 0
      "0000" when "00111010001100", -- t[3724] = 0
      "0000" when "00111010001101", -- t[3725] = 0
      "0000" when "00111010001110", -- t[3726] = 0
      "0000" when "00111010001111", -- t[3727] = 0
      "0000" when "00111010010000", -- t[3728] = 0
      "0000" when "00111010010001", -- t[3729] = 0
      "0000" when "00111010010010", -- t[3730] = 0
      "0000" when "00111010010011", -- t[3731] = 0
      "0000" when "00111010010100", -- t[3732] = 0
      "0000" when "00111010010101", -- t[3733] = 0
      "0000" when "00111010010110", -- t[3734] = 0
      "0000" when "00111010010111", -- t[3735] = 0
      "0000" when "00111010011000", -- t[3736] = 0
      "0000" when "00111010011001", -- t[3737] = 0
      "0000" when "00111010011010", -- t[3738] = 0
      "0000" when "00111010011011", -- t[3739] = 0
      "0000" when "00111010011100", -- t[3740] = 0
      "0000" when "00111010011101", -- t[3741] = 0
      "0000" when "00111010011110", -- t[3742] = 0
      "0000" when "00111010011111", -- t[3743] = 0
      "0000" when "00111010100000", -- t[3744] = 0
      "0000" when "00111010100001", -- t[3745] = 0
      "0000" when "00111010100010", -- t[3746] = 0
      "0000" when "00111010100011", -- t[3747] = 0
      "0000" when "00111010100100", -- t[3748] = 0
      "0000" when "00111010100101", -- t[3749] = 0
      "0000" when "00111010100110", -- t[3750] = 0
      "0000" when "00111010100111", -- t[3751] = 0
      "0000" when "00111010101000", -- t[3752] = 0
      "0000" when "00111010101001", -- t[3753] = 0
      "0000" when "00111010101010", -- t[3754] = 0
      "0000" when "00111010101011", -- t[3755] = 0
      "0000" when "00111010101100", -- t[3756] = 0
      "0000" when "00111010101101", -- t[3757] = 0
      "0000" when "00111010101110", -- t[3758] = 0
      "0000" when "00111010101111", -- t[3759] = 0
      "0000" when "00111010110000", -- t[3760] = 0
      "0000" when "00111010110001", -- t[3761] = 0
      "0000" when "00111010110010", -- t[3762] = 0
      "0000" when "00111010110011", -- t[3763] = 0
      "0000" when "00111010110100", -- t[3764] = 0
      "0000" when "00111010110101", -- t[3765] = 0
      "0000" when "00111010110110", -- t[3766] = 0
      "0000" when "00111010110111", -- t[3767] = 0
      "0000" when "00111010111000", -- t[3768] = 0
      "0000" when "00111010111001", -- t[3769] = 0
      "0000" when "00111010111010", -- t[3770] = 0
      "0000" when "00111010111011", -- t[3771] = 0
      "0000" when "00111010111100", -- t[3772] = 0
      "0000" when "00111010111101", -- t[3773] = 0
      "0000" when "00111010111110", -- t[3774] = 0
      "0000" when "00111010111111", -- t[3775] = 0
      "0000" when "00111011000000", -- t[3776] = 0
      "0000" when "00111011000001", -- t[3777] = 0
      "0000" when "00111011000010", -- t[3778] = 0
      "0000" when "00111011000011", -- t[3779] = 0
      "0000" when "00111011000100", -- t[3780] = 0
      "0000" when "00111011000101", -- t[3781] = 0
      "0000" when "00111011000110", -- t[3782] = 0
      "0000" when "00111011000111", -- t[3783] = 0
      "0000" when "00111011001000", -- t[3784] = 0
      "0000" when "00111011001001", -- t[3785] = 0
      "0000" when "00111011001010", -- t[3786] = 0
      "0000" when "00111011001011", -- t[3787] = 0
      "0000" when "00111011001100", -- t[3788] = 0
      "0000" when "00111011001101", -- t[3789] = 0
      "0000" when "00111011001110", -- t[3790] = 0
      "0000" when "00111011001111", -- t[3791] = 0
      "0000" when "00111011010000", -- t[3792] = 0
      "0000" when "00111011010001", -- t[3793] = 0
      "0000" when "00111011010010", -- t[3794] = 0
      "0000" when "00111011010011", -- t[3795] = 0
      "0000" when "00111011010100", -- t[3796] = 0
      "0000" when "00111011010101", -- t[3797] = 0
      "0000" when "00111011010110", -- t[3798] = 0
      "0000" when "00111011010111", -- t[3799] = 0
      "0000" when "00111011011000", -- t[3800] = 0
      "0000" when "00111011011001", -- t[3801] = 0
      "0000" when "00111011011010", -- t[3802] = 0
      "0000" when "00111011011011", -- t[3803] = 0
      "0000" when "00111011011100", -- t[3804] = 0
      "0000" when "00111011011101", -- t[3805] = 0
      "0000" when "00111011011110", -- t[3806] = 0
      "0000" when "00111011011111", -- t[3807] = 0
      "0000" when "00111011100000", -- t[3808] = 0
      "0000" when "00111011100001", -- t[3809] = 0
      "0000" when "00111011100010", -- t[3810] = 0
      "0000" when "00111011100011", -- t[3811] = 0
      "0000" when "00111011100100", -- t[3812] = 0
      "0000" when "00111011100101", -- t[3813] = 0
      "0000" when "00111011100110", -- t[3814] = 0
      "0000" when "00111011100111", -- t[3815] = 0
      "0000" when "00111011101000", -- t[3816] = 0
      "0000" when "00111011101001", -- t[3817] = 0
      "0000" when "00111011101010", -- t[3818] = 0
      "0000" when "00111011101011", -- t[3819] = 0
      "0000" when "00111011101100", -- t[3820] = 0
      "0000" when "00111011101101", -- t[3821] = 0
      "0000" when "00111011101110", -- t[3822] = 0
      "0000" when "00111011101111", -- t[3823] = 0
      "0000" when "00111011110000", -- t[3824] = 0
      "0000" when "00111011110001", -- t[3825] = 0
      "0000" when "00111011110010", -- t[3826] = 0
      "0000" when "00111011110011", -- t[3827] = 0
      "0000" when "00111011110100", -- t[3828] = 0
      "0000" when "00111011110101", -- t[3829] = 0
      "0000" when "00111011110110", -- t[3830] = 0
      "0000" when "00111011110111", -- t[3831] = 0
      "0000" when "00111011111000", -- t[3832] = 0
      "0000" when "00111011111001", -- t[3833] = 0
      "0000" when "00111011111010", -- t[3834] = 0
      "0000" when "00111011111011", -- t[3835] = 0
      "0000" when "00111011111100", -- t[3836] = 0
      "0000" when "00111011111101", -- t[3837] = 0
      "0000" when "00111011111110", -- t[3838] = 0
      "0000" when "00111011111111", -- t[3839] = 0
      "0000" when "00111100000000", -- t[3840] = 0
      "0000" when "00111100000001", -- t[3841] = 0
      "0000" when "00111100000010", -- t[3842] = 0
      "0000" when "00111100000011", -- t[3843] = 0
      "0000" when "00111100000100", -- t[3844] = 0
      "0000" when "00111100000101", -- t[3845] = 0
      "0000" when "00111100000110", -- t[3846] = 0
      "0000" when "00111100000111", -- t[3847] = 0
      "0000" when "00111100001000", -- t[3848] = 0
      "0000" when "00111100001001", -- t[3849] = 0
      "0000" when "00111100001010", -- t[3850] = 0
      "0000" when "00111100001011", -- t[3851] = 0
      "0000" when "00111100001100", -- t[3852] = 0
      "0000" when "00111100001101", -- t[3853] = 0
      "0000" when "00111100001110", -- t[3854] = 0
      "0000" when "00111100001111", -- t[3855] = 0
      "0000" when "00111100010000", -- t[3856] = 0
      "0000" when "00111100010001", -- t[3857] = 0
      "0000" when "00111100010010", -- t[3858] = 0
      "0000" when "00111100010011", -- t[3859] = 0
      "0000" when "00111100010100", -- t[3860] = 0
      "0000" when "00111100010101", -- t[3861] = 0
      "0000" when "00111100010110", -- t[3862] = 0
      "0000" when "00111100010111", -- t[3863] = 0
      "0000" when "00111100011000", -- t[3864] = 0
      "0000" when "00111100011001", -- t[3865] = 0
      "0000" when "00111100011010", -- t[3866] = 0
      "0000" when "00111100011011", -- t[3867] = 0
      "0000" when "00111100011100", -- t[3868] = 0
      "0000" when "00111100011101", -- t[3869] = 0
      "0000" when "00111100011110", -- t[3870] = 0
      "0000" when "00111100011111", -- t[3871] = 0
      "0000" when "00111100100000", -- t[3872] = 0
      "0000" when "00111100100001", -- t[3873] = 0
      "0000" when "00111100100010", -- t[3874] = 0
      "0000" when "00111100100011", -- t[3875] = 0
      "0000" when "00111100100100", -- t[3876] = 0
      "0000" when "00111100100101", -- t[3877] = 0
      "0000" when "00111100100110", -- t[3878] = 0
      "0000" when "00111100100111", -- t[3879] = 0
      "0000" when "00111100101000", -- t[3880] = 0
      "0000" when "00111100101001", -- t[3881] = 0
      "0000" when "00111100101010", -- t[3882] = 0
      "0000" when "00111100101011", -- t[3883] = 0
      "0000" when "00111100101100", -- t[3884] = 0
      "0000" when "00111100101101", -- t[3885] = 0
      "0000" when "00111100101110", -- t[3886] = 0
      "0000" when "00111100101111", -- t[3887] = 0
      "0000" when "00111100110000", -- t[3888] = 0
      "0000" when "00111100110001", -- t[3889] = 0
      "0000" when "00111100110010", -- t[3890] = 0
      "0000" when "00111100110011", -- t[3891] = 0
      "0000" when "00111100110100", -- t[3892] = 0
      "0000" when "00111100110101", -- t[3893] = 0
      "0000" when "00111100110110", -- t[3894] = 0
      "0000" when "00111100110111", -- t[3895] = 0
      "0000" when "00111100111000", -- t[3896] = 0
      "0000" when "00111100111001", -- t[3897] = 0
      "0000" when "00111100111010", -- t[3898] = 0
      "0000" when "00111100111011", -- t[3899] = 0
      "0000" when "00111100111100", -- t[3900] = 0
      "0000" when "00111100111101", -- t[3901] = 0
      "0000" when "00111100111110", -- t[3902] = 0
      "0000" when "00111100111111", -- t[3903] = 0
      "0000" when "00111101000000", -- t[3904] = 0
      "0000" when "00111101000001", -- t[3905] = 0
      "0000" when "00111101000010", -- t[3906] = 0
      "0000" when "00111101000011", -- t[3907] = 0
      "0000" when "00111101000100", -- t[3908] = 0
      "0000" when "00111101000101", -- t[3909] = 0
      "0000" when "00111101000110", -- t[3910] = 0
      "0000" when "00111101000111", -- t[3911] = 0
      "0000" when "00111101001000", -- t[3912] = 0
      "0000" when "00111101001001", -- t[3913] = 0
      "0000" when "00111101001010", -- t[3914] = 0
      "0000" when "00111101001011", -- t[3915] = 0
      "0000" when "00111101001100", -- t[3916] = 0
      "0000" when "00111101001101", -- t[3917] = 0
      "0000" when "00111101001110", -- t[3918] = 0
      "0000" when "00111101001111", -- t[3919] = 0
      "0000" when "00111101010000", -- t[3920] = 0
      "0000" when "00111101010001", -- t[3921] = 0
      "0000" when "00111101010010", -- t[3922] = 0
      "0000" when "00111101010011", -- t[3923] = 0
      "0000" when "00111101010100", -- t[3924] = 0
      "0000" when "00111101010101", -- t[3925] = 0
      "0000" when "00111101010110", -- t[3926] = 0
      "0000" when "00111101010111", -- t[3927] = 0
      "0000" when "00111101011000", -- t[3928] = 0
      "0000" when "00111101011001", -- t[3929] = 0
      "0000" when "00111101011010", -- t[3930] = 0
      "0000" when "00111101011011", -- t[3931] = 0
      "0000" when "00111101011100", -- t[3932] = 0
      "0000" when "00111101011101", -- t[3933] = 0
      "0000" when "00111101011110", -- t[3934] = 0
      "0000" when "00111101011111", -- t[3935] = 0
      "0000" when "00111101100000", -- t[3936] = 0
      "0000" when "00111101100001", -- t[3937] = 0
      "0000" when "00111101100010", -- t[3938] = 0
      "0000" when "00111101100011", -- t[3939] = 0
      "0000" when "00111101100100", -- t[3940] = 0
      "0000" when "00111101100101", -- t[3941] = 0
      "0000" when "00111101100110", -- t[3942] = 0
      "0000" when "00111101100111", -- t[3943] = 0
      "0000" when "00111101101000", -- t[3944] = 0
      "0000" when "00111101101001", -- t[3945] = 0
      "0000" when "00111101101010", -- t[3946] = 0
      "0000" when "00111101101011", -- t[3947] = 0
      "0000" when "00111101101100", -- t[3948] = 0
      "0000" when "00111101101101", -- t[3949] = 0
      "0000" when "00111101101110", -- t[3950] = 0
      "0000" when "00111101101111", -- t[3951] = 0
      "0000" when "00111101110000", -- t[3952] = 0
      "0000" when "00111101110001", -- t[3953] = 0
      "0000" when "00111101110010", -- t[3954] = 0
      "0000" when "00111101110011", -- t[3955] = 0
      "0000" when "00111101110100", -- t[3956] = 0
      "0000" when "00111101110101", -- t[3957] = 0
      "0000" when "00111101110110", -- t[3958] = 0
      "0000" when "00111101110111", -- t[3959] = 0
      "0000" when "00111101111000", -- t[3960] = 0
      "0000" when "00111101111001", -- t[3961] = 0
      "0000" when "00111101111010", -- t[3962] = 0
      "0000" when "00111101111011", -- t[3963] = 0
      "0000" when "00111101111100", -- t[3964] = 0
      "0000" when "00111101111101", -- t[3965] = 0
      "0000" when "00111101111110", -- t[3966] = 0
      "0000" when "00111101111111", -- t[3967] = 0
      "0000" when "00111110000000", -- t[3968] = 0
      "0000" when "00111110000001", -- t[3969] = 0
      "0000" when "00111110000010", -- t[3970] = 0
      "0000" when "00111110000011", -- t[3971] = 0
      "0000" when "00111110000100", -- t[3972] = 0
      "0000" when "00111110000101", -- t[3973] = 0
      "0000" when "00111110000110", -- t[3974] = 0
      "0000" when "00111110000111", -- t[3975] = 0
      "0000" when "00111110001000", -- t[3976] = 0
      "0000" when "00111110001001", -- t[3977] = 0
      "0000" when "00111110001010", -- t[3978] = 0
      "0000" when "00111110001011", -- t[3979] = 0
      "0000" when "00111110001100", -- t[3980] = 0
      "0000" when "00111110001101", -- t[3981] = 0
      "0000" when "00111110001110", -- t[3982] = 0
      "0000" when "00111110001111", -- t[3983] = 0
      "0000" when "00111110010000", -- t[3984] = 0
      "0000" when "00111110010001", -- t[3985] = 0
      "0000" when "00111110010010", -- t[3986] = 0
      "0000" when "00111110010011", -- t[3987] = 0
      "0000" when "00111110010100", -- t[3988] = 0
      "0000" when "00111110010101", -- t[3989] = 0
      "0000" when "00111110010110", -- t[3990] = 0
      "0000" when "00111110010111", -- t[3991] = 0
      "0000" when "00111110011000", -- t[3992] = 0
      "0000" when "00111110011001", -- t[3993] = 0
      "0000" when "00111110011010", -- t[3994] = 0
      "0000" when "00111110011011", -- t[3995] = 0
      "0000" when "00111110011100", -- t[3996] = 0
      "0000" when "00111110011101", -- t[3997] = 0
      "0000" when "00111110011110", -- t[3998] = 0
      "0000" when "00111110011111", -- t[3999] = 0
      "0000" when "00111110100000", -- t[4000] = 0
      "0000" when "00111110100001", -- t[4001] = 0
      "0000" when "00111110100010", -- t[4002] = 0
      "0000" when "00111110100011", -- t[4003] = 0
      "0000" when "00111110100100", -- t[4004] = 0
      "0000" when "00111110100101", -- t[4005] = 0
      "0000" when "00111110100110", -- t[4006] = 0
      "0000" when "00111110100111", -- t[4007] = 0
      "0000" when "00111110101000", -- t[4008] = 0
      "0000" when "00111110101001", -- t[4009] = 0
      "0000" when "00111110101010", -- t[4010] = 0
      "0000" when "00111110101011", -- t[4011] = 0
      "0000" when "00111110101100", -- t[4012] = 0
      "0000" when "00111110101101", -- t[4013] = 0
      "0000" when "00111110101110", -- t[4014] = 0
      "0000" when "00111110101111", -- t[4015] = 0
      "0000" when "00111110110000", -- t[4016] = 0
      "0000" when "00111110110001", -- t[4017] = 0
      "0000" when "00111110110010", -- t[4018] = 0
      "0000" when "00111110110011", -- t[4019] = 0
      "0000" when "00111110110100", -- t[4020] = 0
      "0000" when "00111110110101", -- t[4021] = 0
      "0000" when "00111110110110", -- t[4022] = 0
      "0000" when "00111110110111", -- t[4023] = 0
      "0000" when "00111110111000", -- t[4024] = 0
      "0000" when "00111110111001", -- t[4025] = 0
      "0000" when "00111110111010", -- t[4026] = 0
      "0000" when "00111110111011", -- t[4027] = 0
      "0000" when "00111110111100", -- t[4028] = 0
      "0000" when "00111110111101", -- t[4029] = 0
      "0000" when "00111110111110", -- t[4030] = 0
      "0000" when "00111110111111", -- t[4031] = 0
      "0000" when "00111111000000", -- t[4032] = 0
      "0000" when "00111111000001", -- t[4033] = 0
      "0000" when "00111111000010", -- t[4034] = 0
      "0000" when "00111111000011", -- t[4035] = 0
      "0000" when "00111111000100", -- t[4036] = 0
      "0000" when "00111111000101", -- t[4037] = 0
      "0000" when "00111111000110", -- t[4038] = 0
      "0000" when "00111111000111", -- t[4039] = 0
      "0000" when "00111111001000", -- t[4040] = 0
      "0000" when "00111111001001", -- t[4041] = 0
      "0000" when "00111111001010", -- t[4042] = 0
      "0000" when "00111111001011", -- t[4043] = 0
      "0000" when "00111111001100", -- t[4044] = 0
      "0000" when "00111111001101", -- t[4045] = 0
      "0000" when "00111111001110", -- t[4046] = 0
      "0000" when "00111111001111", -- t[4047] = 0
      "0000" when "00111111010000", -- t[4048] = 0
      "0000" when "00111111010001", -- t[4049] = 0
      "0000" when "00111111010010", -- t[4050] = 0
      "0000" when "00111111010011", -- t[4051] = 0
      "0000" when "00111111010100", -- t[4052] = 0
      "0000" when "00111111010101", -- t[4053] = 0
      "0000" when "00111111010110", -- t[4054] = 0
      "0000" when "00111111010111", -- t[4055] = 0
      "0000" when "00111111011000", -- t[4056] = 0
      "0000" when "00111111011001", -- t[4057] = 0
      "0000" when "00111111011010", -- t[4058] = 0
      "0000" when "00111111011011", -- t[4059] = 0
      "0000" when "00111111011100", -- t[4060] = 0
      "0000" when "00111111011101", -- t[4061] = 0
      "0000" when "00111111011110", -- t[4062] = 0
      "0000" when "00111111011111", -- t[4063] = 0
      "0000" when "00111111100000", -- t[4064] = 0
      "0000" when "00111111100001", -- t[4065] = 0
      "0000" when "00111111100010", -- t[4066] = 0
      "0000" when "00111111100011", -- t[4067] = 0
      "0000" when "00111111100100", -- t[4068] = 0
      "0000" when "00111111100101", -- t[4069] = 0
      "0000" when "00111111100110", -- t[4070] = 0
      "0000" when "00111111100111", -- t[4071] = 0
      "0000" when "00111111101000", -- t[4072] = 0
      "0000" when "00111111101001", -- t[4073] = 0
      "0000" when "00111111101010", -- t[4074] = 0
      "0000" when "00111111101011", -- t[4075] = 0
      "0000" when "00111111101100", -- t[4076] = 0
      "0000" when "00111111101101", -- t[4077] = 0
      "0000" when "00111111101110", -- t[4078] = 0
      "0000" when "00111111101111", -- t[4079] = 0
      "0000" when "00111111110000", -- t[4080] = 0
      "0000" when "00111111110001", -- t[4081] = 0
      "0000" when "00111111110010", -- t[4082] = 0
      "0000" when "00111111110011", -- t[4083] = 0
      "0000" when "00111111110100", -- t[4084] = 0
      "0000" when "00111111110101", -- t[4085] = 0
      "0000" when "00111111110110", -- t[4086] = 0
      "0000" when "00111111110111", -- t[4087] = 0
      "0000" when "00111111111000", -- t[4088] = 0
      "0000" when "00111111111001", -- t[4089] = 0
      "0000" when "00111111111010", -- t[4090] = 0
      "0000" when "00111111111011", -- t[4091] = 0
      "0000" when "00111111111100", -- t[4092] = 0
      "0000" when "00111111111101", -- t[4093] = 0
      "0000" when "00111111111110", -- t[4094] = 0
      "0000" when "00111111111111", -- t[4095] = 0
      "0000" when "01000000000000", -- t[4096] = 0
      "0000" when "01000000000001", -- t[4097] = 0
      "0000" when "01000000000010", -- t[4098] = 0
      "0000" when "01000000000011", -- t[4099] = 0
      "0000" when "01000000000100", -- t[4100] = 0
      "0000" when "01000000000101", -- t[4101] = 0
      "0000" when "01000000000110", -- t[4102] = 0
      "0000" when "01000000000111", -- t[4103] = 0
      "0000" when "01000000001000", -- t[4104] = 0
      "0000" when "01000000001001", -- t[4105] = 0
      "0000" when "01000000001010", -- t[4106] = 0
      "0000" when "01000000001011", -- t[4107] = 0
      "0000" when "01000000001100", -- t[4108] = 0
      "0000" when "01000000001101", -- t[4109] = 0
      "0000" when "01000000001110", -- t[4110] = 0
      "0000" when "01000000001111", -- t[4111] = 0
      "0000" when "01000000010000", -- t[4112] = 0
      "0000" when "01000000010001", -- t[4113] = 0
      "0000" when "01000000010010", -- t[4114] = 0
      "0000" when "01000000010011", -- t[4115] = 0
      "0000" when "01000000010100", -- t[4116] = 0
      "0000" when "01000000010101", -- t[4117] = 0
      "0000" when "01000000010110", -- t[4118] = 0
      "0000" when "01000000010111", -- t[4119] = 0
      "0000" when "01000000011000", -- t[4120] = 0
      "0000" when "01000000011001", -- t[4121] = 0
      "0000" when "01000000011010", -- t[4122] = 0
      "0000" when "01000000011011", -- t[4123] = 0
      "0000" when "01000000011100", -- t[4124] = 0
      "0000" when "01000000011101", -- t[4125] = 0
      "0000" when "01000000011110", -- t[4126] = 0
      "0000" when "01000000011111", -- t[4127] = 0
      "0000" when "01000000100000", -- t[4128] = 0
      "0000" when "01000000100001", -- t[4129] = 0
      "0000" when "01000000100010", -- t[4130] = 0
      "0000" when "01000000100011", -- t[4131] = 0
      "0000" when "01000000100100", -- t[4132] = 0
      "0000" when "01000000100101", -- t[4133] = 0
      "0000" when "01000000100110", -- t[4134] = 0
      "0000" when "01000000100111", -- t[4135] = 0
      "0000" when "01000000101000", -- t[4136] = 0
      "0000" when "01000000101001", -- t[4137] = 0
      "0000" when "01000000101010", -- t[4138] = 0
      "0000" when "01000000101011", -- t[4139] = 0
      "0000" when "01000000101100", -- t[4140] = 0
      "0000" when "01000000101101", -- t[4141] = 0
      "0000" when "01000000101110", -- t[4142] = 0
      "0000" when "01000000101111", -- t[4143] = 0
      "0000" when "01000000110000", -- t[4144] = 0
      "0000" when "01000000110001", -- t[4145] = 0
      "0000" when "01000000110010", -- t[4146] = 0
      "0000" when "01000000110011", -- t[4147] = 0
      "0000" when "01000000110100", -- t[4148] = 0
      "0000" when "01000000110101", -- t[4149] = 0
      "0000" when "01000000110110", -- t[4150] = 0
      "0000" when "01000000110111", -- t[4151] = 0
      "0000" when "01000000111000", -- t[4152] = 0
      "0000" when "01000000111001", -- t[4153] = 0
      "0000" when "01000000111010", -- t[4154] = 0
      "0000" when "01000000111011", -- t[4155] = 0
      "0000" when "01000000111100", -- t[4156] = 0
      "0000" when "01000000111101", -- t[4157] = 0
      "0000" when "01000000111110", -- t[4158] = 0
      "0000" when "01000000111111", -- t[4159] = 0
      "0000" when "01000001000000", -- t[4160] = 0
      "0000" when "01000001000001", -- t[4161] = 0
      "0000" when "01000001000010", -- t[4162] = 0
      "0000" when "01000001000011", -- t[4163] = 0
      "0000" when "01000001000100", -- t[4164] = 0
      "0000" when "01000001000101", -- t[4165] = 0
      "0000" when "01000001000110", -- t[4166] = 0
      "0000" when "01000001000111", -- t[4167] = 0
      "0000" when "01000001001000", -- t[4168] = 0
      "0000" when "01000001001001", -- t[4169] = 0
      "0000" when "01000001001010", -- t[4170] = 0
      "0000" when "01000001001011", -- t[4171] = 0
      "0000" when "01000001001100", -- t[4172] = 0
      "0000" when "01000001001101", -- t[4173] = 0
      "0000" when "01000001001110", -- t[4174] = 0
      "0000" when "01000001001111", -- t[4175] = 0
      "0000" when "01000001010000", -- t[4176] = 0
      "0000" when "01000001010001", -- t[4177] = 0
      "0000" when "01000001010010", -- t[4178] = 0
      "0000" when "01000001010011", -- t[4179] = 0
      "0000" when "01000001010100", -- t[4180] = 0
      "0000" when "01000001010101", -- t[4181] = 0
      "0000" when "01000001010110", -- t[4182] = 0
      "0000" when "01000001010111", -- t[4183] = 0
      "0000" when "01000001011000", -- t[4184] = 0
      "0000" when "01000001011001", -- t[4185] = 0
      "0000" when "01000001011010", -- t[4186] = 0
      "0000" when "01000001011011", -- t[4187] = 0
      "0000" when "01000001011100", -- t[4188] = 0
      "0000" when "01000001011101", -- t[4189] = 0
      "0000" when "01000001011110", -- t[4190] = 0
      "0000" when "01000001011111", -- t[4191] = 0
      "0000" when "01000001100000", -- t[4192] = 0
      "0000" when "01000001100001", -- t[4193] = 0
      "0000" when "01000001100010", -- t[4194] = 0
      "0000" when "01000001100011", -- t[4195] = 0
      "0000" when "01000001100100", -- t[4196] = 0
      "0000" when "01000001100101", -- t[4197] = 0
      "0000" when "01000001100110", -- t[4198] = 0
      "0000" when "01000001100111", -- t[4199] = 0
      "0000" when "01000001101000", -- t[4200] = 0
      "0000" when "01000001101001", -- t[4201] = 0
      "0000" when "01000001101010", -- t[4202] = 0
      "0000" when "01000001101011", -- t[4203] = 0
      "0000" when "01000001101100", -- t[4204] = 0
      "0000" when "01000001101101", -- t[4205] = 0
      "0000" when "01000001101110", -- t[4206] = 0
      "0000" when "01000001101111", -- t[4207] = 0
      "0000" when "01000001110000", -- t[4208] = 0
      "0000" when "01000001110001", -- t[4209] = 0
      "0000" when "01000001110010", -- t[4210] = 0
      "0000" when "01000001110011", -- t[4211] = 0
      "0000" when "01000001110100", -- t[4212] = 0
      "0000" when "01000001110101", -- t[4213] = 0
      "0000" when "01000001110110", -- t[4214] = 0
      "0000" when "01000001110111", -- t[4215] = 0
      "0000" when "01000001111000", -- t[4216] = 0
      "0000" when "01000001111001", -- t[4217] = 0
      "0000" when "01000001111010", -- t[4218] = 0
      "0000" when "01000001111011", -- t[4219] = 0
      "0000" when "01000001111100", -- t[4220] = 0
      "0000" when "01000001111101", -- t[4221] = 0
      "0000" when "01000001111110", -- t[4222] = 0
      "0000" when "01000001111111", -- t[4223] = 0
      "0000" when "01000010000000", -- t[4224] = 0
      "0000" when "01000010000001", -- t[4225] = 0
      "0000" when "01000010000010", -- t[4226] = 0
      "0000" when "01000010000011", -- t[4227] = 0
      "0000" when "01000010000100", -- t[4228] = 0
      "0000" when "01000010000101", -- t[4229] = 0
      "0000" when "01000010000110", -- t[4230] = 0
      "0000" when "01000010000111", -- t[4231] = 0
      "0000" when "01000010001000", -- t[4232] = 0
      "0000" when "01000010001001", -- t[4233] = 0
      "0000" when "01000010001010", -- t[4234] = 0
      "0000" when "01000010001011", -- t[4235] = 0
      "0000" when "01000010001100", -- t[4236] = 0
      "0000" when "01000010001101", -- t[4237] = 0
      "0000" when "01000010001110", -- t[4238] = 0
      "0000" when "01000010001111", -- t[4239] = 0
      "0000" when "01000010010000", -- t[4240] = 0
      "0000" when "01000010010001", -- t[4241] = 0
      "0000" when "01000010010010", -- t[4242] = 0
      "0000" when "01000010010011", -- t[4243] = 0
      "0000" when "01000010010100", -- t[4244] = 0
      "0000" when "01000010010101", -- t[4245] = 0
      "0000" when "01000010010110", -- t[4246] = 0
      "0000" when "01000010010111", -- t[4247] = 0
      "0000" when "01000010011000", -- t[4248] = 0
      "0000" when "01000010011001", -- t[4249] = 0
      "0000" when "01000010011010", -- t[4250] = 0
      "0000" when "01000010011011", -- t[4251] = 0
      "0000" when "01000010011100", -- t[4252] = 0
      "0000" when "01000010011101", -- t[4253] = 0
      "0000" when "01000010011110", -- t[4254] = 0
      "0000" when "01000010011111", -- t[4255] = 0
      "0000" when "01000010100000", -- t[4256] = 0
      "0000" when "01000010100001", -- t[4257] = 0
      "0000" when "01000010100010", -- t[4258] = 0
      "0000" when "01000010100011", -- t[4259] = 0
      "0000" when "01000010100100", -- t[4260] = 0
      "0000" when "01000010100101", -- t[4261] = 0
      "0000" when "01000010100110", -- t[4262] = 0
      "0000" when "01000010100111", -- t[4263] = 0
      "0000" when "01000010101000", -- t[4264] = 0
      "0000" when "01000010101001", -- t[4265] = 0
      "0000" when "01000010101010", -- t[4266] = 0
      "0000" when "01000010101011", -- t[4267] = 0
      "0000" when "01000010101100", -- t[4268] = 0
      "0000" when "01000010101101", -- t[4269] = 0
      "0000" when "01000010101110", -- t[4270] = 0
      "0000" when "01000010101111", -- t[4271] = 0
      "0000" when "01000010110000", -- t[4272] = 0
      "0000" when "01000010110001", -- t[4273] = 0
      "0000" when "01000010110010", -- t[4274] = 0
      "0000" when "01000010110011", -- t[4275] = 0
      "0000" when "01000010110100", -- t[4276] = 0
      "0000" when "01000010110101", -- t[4277] = 0
      "0000" when "01000010110110", -- t[4278] = 0
      "0000" when "01000010110111", -- t[4279] = 0
      "0000" when "01000010111000", -- t[4280] = 0
      "0000" when "01000010111001", -- t[4281] = 0
      "0000" when "01000010111010", -- t[4282] = 0
      "0000" when "01000010111011", -- t[4283] = 0
      "0000" when "01000010111100", -- t[4284] = 0
      "0000" when "01000010111101", -- t[4285] = 0
      "0000" when "01000010111110", -- t[4286] = 0
      "0000" when "01000010111111", -- t[4287] = 0
      "0000" when "01000011000000", -- t[4288] = 0
      "0000" when "01000011000001", -- t[4289] = 0
      "0000" when "01000011000010", -- t[4290] = 0
      "0000" when "01000011000011", -- t[4291] = 0
      "0000" when "01000011000100", -- t[4292] = 0
      "0000" when "01000011000101", -- t[4293] = 0
      "0000" when "01000011000110", -- t[4294] = 0
      "0000" when "01000011000111", -- t[4295] = 0
      "0000" when "01000011001000", -- t[4296] = 0
      "0000" when "01000011001001", -- t[4297] = 0
      "0000" when "01000011001010", -- t[4298] = 0
      "0000" when "01000011001011", -- t[4299] = 0
      "0000" when "01000011001100", -- t[4300] = 0
      "0000" when "01000011001101", -- t[4301] = 0
      "0000" when "01000011001110", -- t[4302] = 0
      "0000" when "01000011001111", -- t[4303] = 0
      "0000" when "01000011010000", -- t[4304] = 0
      "0000" when "01000011010001", -- t[4305] = 0
      "0000" when "01000011010010", -- t[4306] = 0
      "0000" when "01000011010011", -- t[4307] = 0
      "0000" when "01000011010100", -- t[4308] = 0
      "0000" when "01000011010101", -- t[4309] = 0
      "0000" when "01000011010110", -- t[4310] = 0
      "0000" when "01000011010111", -- t[4311] = 0
      "0000" when "01000011011000", -- t[4312] = 0
      "0000" when "01000011011001", -- t[4313] = 0
      "0000" when "01000011011010", -- t[4314] = 0
      "0000" when "01000011011011", -- t[4315] = 0
      "0000" when "01000011011100", -- t[4316] = 0
      "0000" when "01000011011101", -- t[4317] = 0
      "0000" when "01000011011110", -- t[4318] = 0
      "0000" when "01000011011111", -- t[4319] = 0
      "0000" when "01000011100000", -- t[4320] = 0
      "0000" when "01000011100001", -- t[4321] = 0
      "0000" when "01000011100010", -- t[4322] = 0
      "0000" when "01000011100011", -- t[4323] = 0
      "0000" when "01000011100100", -- t[4324] = 0
      "0000" when "01000011100101", -- t[4325] = 0
      "0000" when "01000011100110", -- t[4326] = 0
      "0000" when "01000011100111", -- t[4327] = 0
      "0000" when "01000011101000", -- t[4328] = 0
      "0000" when "01000011101001", -- t[4329] = 0
      "0000" when "01000011101010", -- t[4330] = 0
      "0000" when "01000011101011", -- t[4331] = 0
      "0000" when "01000011101100", -- t[4332] = 0
      "0000" when "01000011101101", -- t[4333] = 0
      "0000" when "01000011101110", -- t[4334] = 0
      "0000" when "01000011101111", -- t[4335] = 0
      "0000" when "01000011110000", -- t[4336] = 0
      "0000" when "01000011110001", -- t[4337] = 0
      "0000" when "01000011110010", -- t[4338] = 0
      "0000" when "01000011110011", -- t[4339] = 0
      "0000" when "01000011110100", -- t[4340] = 0
      "0000" when "01000011110101", -- t[4341] = 0
      "0000" when "01000011110110", -- t[4342] = 0
      "0000" when "01000011110111", -- t[4343] = 0
      "0000" when "01000011111000", -- t[4344] = 0
      "0000" when "01000011111001", -- t[4345] = 0
      "0000" when "01000011111010", -- t[4346] = 0
      "0000" when "01000011111011", -- t[4347] = 0
      "0000" when "01000011111100", -- t[4348] = 0
      "0000" when "01000011111101", -- t[4349] = 0
      "0000" when "01000011111110", -- t[4350] = 0
      "0000" when "01000011111111", -- t[4351] = 0
      "0000" when "01000100000000", -- t[4352] = 0
      "0000" when "01000100000001", -- t[4353] = 0
      "0000" when "01000100000010", -- t[4354] = 0
      "0000" when "01000100000011", -- t[4355] = 0
      "0000" when "01000100000100", -- t[4356] = 0
      "0000" when "01000100000101", -- t[4357] = 0
      "0000" when "01000100000110", -- t[4358] = 0
      "0000" when "01000100000111", -- t[4359] = 0
      "0000" when "01000100001000", -- t[4360] = 0
      "0000" when "01000100001001", -- t[4361] = 0
      "0000" when "01000100001010", -- t[4362] = 0
      "0000" when "01000100001011", -- t[4363] = 0
      "0000" when "01000100001100", -- t[4364] = 0
      "0000" when "01000100001101", -- t[4365] = 0
      "0000" when "01000100001110", -- t[4366] = 0
      "0000" when "01000100001111", -- t[4367] = 0
      "0000" when "01000100010000", -- t[4368] = 0
      "0000" when "01000100010001", -- t[4369] = 0
      "0000" when "01000100010010", -- t[4370] = 0
      "0000" when "01000100010011", -- t[4371] = 0
      "0000" when "01000100010100", -- t[4372] = 0
      "0000" when "01000100010101", -- t[4373] = 0
      "0000" when "01000100010110", -- t[4374] = 0
      "0000" when "01000100010111", -- t[4375] = 0
      "0000" when "01000100011000", -- t[4376] = 0
      "0000" when "01000100011001", -- t[4377] = 0
      "0000" when "01000100011010", -- t[4378] = 0
      "0000" when "01000100011011", -- t[4379] = 0
      "0000" when "01000100011100", -- t[4380] = 0
      "0000" when "01000100011101", -- t[4381] = 0
      "0000" when "01000100011110", -- t[4382] = 0
      "0000" when "01000100011111", -- t[4383] = 0
      "0000" when "01000100100000", -- t[4384] = 0
      "0000" when "01000100100001", -- t[4385] = 0
      "0000" when "01000100100010", -- t[4386] = 0
      "0000" when "01000100100011", -- t[4387] = 0
      "0000" when "01000100100100", -- t[4388] = 0
      "0000" when "01000100100101", -- t[4389] = 0
      "0000" when "01000100100110", -- t[4390] = 0
      "0000" when "01000100100111", -- t[4391] = 0
      "0000" when "01000100101000", -- t[4392] = 0
      "0000" when "01000100101001", -- t[4393] = 0
      "0000" when "01000100101010", -- t[4394] = 0
      "0000" when "01000100101011", -- t[4395] = 0
      "0000" when "01000100101100", -- t[4396] = 0
      "0000" when "01000100101101", -- t[4397] = 0
      "0000" when "01000100101110", -- t[4398] = 0
      "0000" when "01000100101111", -- t[4399] = 0
      "0000" when "01000100110000", -- t[4400] = 0
      "0000" when "01000100110001", -- t[4401] = 0
      "0000" when "01000100110010", -- t[4402] = 0
      "0000" when "01000100110011", -- t[4403] = 0
      "0000" when "01000100110100", -- t[4404] = 0
      "0000" when "01000100110101", -- t[4405] = 0
      "0000" when "01000100110110", -- t[4406] = 0
      "0000" when "01000100110111", -- t[4407] = 0
      "0000" when "01000100111000", -- t[4408] = 0
      "0000" when "01000100111001", -- t[4409] = 0
      "0000" when "01000100111010", -- t[4410] = 0
      "0000" when "01000100111011", -- t[4411] = 0
      "0000" when "01000100111100", -- t[4412] = 0
      "0000" when "01000100111101", -- t[4413] = 0
      "0000" when "01000100111110", -- t[4414] = 0
      "0000" when "01000100111111", -- t[4415] = 0
      "0000" when "01000101000000", -- t[4416] = 0
      "0000" when "01000101000001", -- t[4417] = 0
      "0000" when "01000101000010", -- t[4418] = 0
      "0000" when "01000101000011", -- t[4419] = 0
      "0000" when "01000101000100", -- t[4420] = 0
      "0000" when "01000101000101", -- t[4421] = 0
      "0000" when "01000101000110", -- t[4422] = 0
      "0000" when "01000101000111", -- t[4423] = 0
      "0000" when "01000101001000", -- t[4424] = 0
      "0000" when "01000101001001", -- t[4425] = 0
      "0000" when "01000101001010", -- t[4426] = 0
      "0000" when "01000101001011", -- t[4427] = 0
      "0000" when "01000101001100", -- t[4428] = 0
      "0000" when "01000101001101", -- t[4429] = 0
      "0000" when "01000101001110", -- t[4430] = 0
      "0000" when "01000101001111", -- t[4431] = 0
      "0000" when "01000101010000", -- t[4432] = 0
      "0000" when "01000101010001", -- t[4433] = 0
      "0000" when "01000101010010", -- t[4434] = 0
      "0000" when "01000101010011", -- t[4435] = 0
      "0000" when "01000101010100", -- t[4436] = 0
      "0000" when "01000101010101", -- t[4437] = 0
      "0000" when "01000101010110", -- t[4438] = 0
      "0000" when "01000101010111", -- t[4439] = 0
      "0000" when "01000101011000", -- t[4440] = 0
      "0000" when "01000101011001", -- t[4441] = 0
      "0000" when "01000101011010", -- t[4442] = 0
      "0000" when "01000101011011", -- t[4443] = 0
      "0000" when "01000101011100", -- t[4444] = 0
      "0000" when "01000101011101", -- t[4445] = 0
      "0000" when "01000101011110", -- t[4446] = 0
      "0000" when "01000101011111", -- t[4447] = 0
      "0000" when "01000101100000", -- t[4448] = 0
      "0000" when "01000101100001", -- t[4449] = 0
      "0000" when "01000101100010", -- t[4450] = 0
      "0000" when "01000101100011", -- t[4451] = 0
      "0000" when "01000101100100", -- t[4452] = 0
      "0000" when "01000101100101", -- t[4453] = 0
      "0000" when "01000101100110", -- t[4454] = 0
      "0000" when "01000101100111", -- t[4455] = 0
      "0000" when "01000101101000", -- t[4456] = 0
      "0000" when "01000101101001", -- t[4457] = 0
      "0000" when "01000101101010", -- t[4458] = 0
      "0000" when "01000101101011", -- t[4459] = 0
      "0000" when "01000101101100", -- t[4460] = 0
      "0000" when "01000101101101", -- t[4461] = 0
      "0000" when "01000101101110", -- t[4462] = 0
      "0000" when "01000101101111", -- t[4463] = 0
      "0000" when "01000101110000", -- t[4464] = 0
      "0000" when "01000101110001", -- t[4465] = 0
      "0000" when "01000101110010", -- t[4466] = 0
      "0000" when "01000101110011", -- t[4467] = 0
      "0000" when "01000101110100", -- t[4468] = 0
      "0000" when "01000101110101", -- t[4469] = 0
      "0000" when "01000101110110", -- t[4470] = 0
      "0000" when "01000101110111", -- t[4471] = 0
      "0000" when "01000101111000", -- t[4472] = 0
      "0000" when "01000101111001", -- t[4473] = 0
      "0000" when "01000101111010", -- t[4474] = 0
      "0000" when "01000101111011", -- t[4475] = 0
      "0000" when "01000101111100", -- t[4476] = 0
      "0000" when "01000101111101", -- t[4477] = 0
      "0000" when "01000101111110", -- t[4478] = 0
      "0000" when "01000101111111", -- t[4479] = 0
      "0000" when "01000110000000", -- t[4480] = 0
      "0000" when "01000110000001", -- t[4481] = 0
      "0000" when "01000110000010", -- t[4482] = 0
      "0000" when "01000110000011", -- t[4483] = 0
      "0000" when "01000110000100", -- t[4484] = 0
      "0000" when "01000110000101", -- t[4485] = 0
      "0000" when "01000110000110", -- t[4486] = 0
      "0000" when "01000110000111", -- t[4487] = 0
      "0000" when "01000110001000", -- t[4488] = 0
      "0000" when "01000110001001", -- t[4489] = 0
      "0000" when "01000110001010", -- t[4490] = 0
      "0000" when "01000110001011", -- t[4491] = 0
      "0000" when "01000110001100", -- t[4492] = 0
      "0000" when "01000110001101", -- t[4493] = 0
      "0000" when "01000110001110", -- t[4494] = 0
      "0000" when "01000110001111", -- t[4495] = 0
      "0000" when "01000110010000", -- t[4496] = 0
      "0000" when "01000110010001", -- t[4497] = 0
      "0000" when "01000110010010", -- t[4498] = 0
      "0000" when "01000110010011", -- t[4499] = 0
      "0000" when "01000110010100", -- t[4500] = 0
      "0000" when "01000110010101", -- t[4501] = 0
      "0000" when "01000110010110", -- t[4502] = 0
      "0000" when "01000110010111", -- t[4503] = 0
      "0000" when "01000110011000", -- t[4504] = 0
      "0000" when "01000110011001", -- t[4505] = 0
      "0000" when "01000110011010", -- t[4506] = 0
      "0000" when "01000110011011", -- t[4507] = 0
      "0000" when "01000110011100", -- t[4508] = 0
      "0000" when "01000110011101", -- t[4509] = 0
      "0000" when "01000110011110", -- t[4510] = 0
      "0000" when "01000110011111", -- t[4511] = 0
      "0000" when "01000110100000", -- t[4512] = 0
      "0000" when "01000110100001", -- t[4513] = 0
      "0000" when "01000110100010", -- t[4514] = 0
      "0000" when "01000110100011", -- t[4515] = 0
      "0000" when "01000110100100", -- t[4516] = 0
      "0000" when "01000110100101", -- t[4517] = 0
      "0000" when "01000110100110", -- t[4518] = 0
      "0000" when "01000110100111", -- t[4519] = 0
      "0000" when "01000110101000", -- t[4520] = 0
      "0000" when "01000110101001", -- t[4521] = 0
      "0000" when "01000110101010", -- t[4522] = 0
      "0000" when "01000110101011", -- t[4523] = 0
      "0000" when "01000110101100", -- t[4524] = 0
      "0000" when "01000110101101", -- t[4525] = 0
      "0000" when "01000110101110", -- t[4526] = 0
      "0000" when "01000110101111", -- t[4527] = 0
      "0000" when "01000110110000", -- t[4528] = 0
      "0000" when "01000110110001", -- t[4529] = 0
      "0000" when "01000110110010", -- t[4530] = 0
      "0000" when "01000110110011", -- t[4531] = 0
      "0000" when "01000110110100", -- t[4532] = 0
      "0000" when "01000110110101", -- t[4533] = 0
      "0000" when "01000110110110", -- t[4534] = 0
      "0000" when "01000110110111", -- t[4535] = 0
      "0000" when "01000110111000", -- t[4536] = 0
      "0000" when "01000110111001", -- t[4537] = 0
      "0000" when "01000110111010", -- t[4538] = 0
      "0000" when "01000110111011", -- t[4539] = 0
      "0000" when "01000110111100", -- t[4540] = 0
      "0000" when "01000110111101", -- t[4541] = 0
      "0000" when "01000110111110", -- t[4542] = 0
      "0000" when "01000110111111", -- t[4543] = 0
      "0000" when "01000111000000", -- t[4544] = 0
      "0000" when "01000111000001", -- t[4545] = 0
      "0000" when "01000111000010", -- t[4546] = 0
      "0000" when "01000111000011", -- t[4547] = 0
      "0000" when "01000111000100", -- t[4548] = 0
      "0000" when "01000111000101", -- t[4549] = 0
      "0000" when "01000111000110", -- t[4550] = 0
      "0000" when "01000111000111", -- t[4551] = 0
      "0000" when "01000111001000", -- t[4552] = 0
      "0000" when "01000111001001", -- t[4553] = 0
      "0000" when "01000111001010", -- t[4554] = 0
      "0000" when "01000111001011", -- t[4555] = 0
      "0000" when "01000111001100", -- t[4556] = 0
      "0000" when "01000111001101", -- t[4557] = 0
      "0000" when "01000111001110", -- t[4558] = 0
      "0000" when "01000111001111", -- t[4559] = 0
      "0000" when "01000111010000", -- t[4560] = 0
      "0000" when "01000111010001", -- t[4561] = 0
      "0000" when "01000111010010", -- t[4562] = 0
      "0000" when "01000111010011", -- t[4563] = 0
      "0000" when "01000111010100", -- t[4564] = 0
      "0000" when "01000111010101", -- t[4565] = 0
      "0000" when "01000111010110", -- t[4566] = 0
      "0000" when "01000111010111", -- t[4567] = 0
      "0000" when "01000111011000", -- t[4568] = 0
      "0000" when "01000111011001", -- t[4569] = 0
      "0000" when "01000111011010", -- t[4570] = 0
      "0000" when "01000111011011", -- t[4571] = 0
      "0000" when "01000111011100", -- t[4572] = 0
      "0000" when "01000111011101", -- t[4573] = 0
      "0000" when "01000111011110", -- t[4574] = 0
      "0000" when "01000111011111", -- t[4575] = 0
      "0000" when "01000111100000", -- t[4576] = 0
      "0000" when "01000111100001", -- t[4577] = 0
      "0000" when "01000111100010", -- t[4578] = 0
      "0001" when "01000111100011", -- t[4579] = 1
      "0001" when "01000111100100", -- t[4580] = 1
      "0001" when "01000111100101", -- t[4581] = 1
      "0001" when "01000111100110", -- t[4582] = 1
      "0001" when "01000111100111", -- t[4583] = 1
      "0001" when "01000111101000", -- t[4584] = 1
      "0001" when "01000111101001", -- t[4585] = 1
      "0001" when "01000111101010", -- t[4586] = 1
      "0001" when "01000111101011", -- t[4587] = 1
      "0001" when "01000111101100", -- t[4588] = 1
      "0001" when "01000111101101", -- t[4589] = 1
      "0001" when "01000111101110", -- t[4590] = 1
      "0001" when "01000111101111", -- t[4591] = 1
      "0001" when "01000111110000", -- t[4592] = 1
      "0001" when "01000111110001", -- t[4593] = 1
      "0001" when "01000111110010", -- t[4594] = 1
      "0001" when "01000111110011", -- t[4595] = 1
      "0001" when "01000111110100", -- t[4596] = 1
      "0001" when "01000111110101", -- t[4597] = 1
      "0001" when "01000111110110", -- t[4598] = 1
      "0001" when "01000111110111", -- t[4599] = 1
      "0001" when "01000111111000", -- t[4600] = 1
      "0001" when "01000111111001", -- t[4601] = 1
      "0001" when "01000111111010", -- t[4602] = 1
      "0001" when "01000111111011", -- t[4603] = 1
      "0001" when "01000111111100", -- t[4604] = 1
      "0001" when "01000111111101", -- t[4605] = 1
      "0001" when "01000111111110", -- t[4606] = 1
      "0001" when "01000111111111", -- t[4607] = 1
      "0001" when "01001000000000", -- t[4608] = 1
      "0001" when "01001000000001", -- t[4609] = 1
      "0001" when "01001000000010", -- t[4610] = 1
      "0001" when "01001000000011", -- t[4611] = 1
      "0001" when "01001000000100", -- t[4612] = 1
      "0001" when "01001000000101", -- t[4613] = 1
      "0001" when "01001000000110", -- t[4614] = 1
      "0001" when "01001000000111", -- t[4615] = 1
      "0001" when "01001000001000", -- t[4616] = 1
      "0001" when "01001000001001", -- t[4617] = 1
      "0001" when "01001000001010", -- t[4618] = 1
      "0001" when "01001000001011", -- t[4619] = 1
      "0001" when "01001000001100", -- t[4620] = 1
      "0001" when "01001000001101", -- t[4621] = 1
      "0001" when "01001000001110", -- t[4622] = 1
      "0001" when "01001000001111", -- t[4623] = 1
      "0001" when "01001000010000", -- t[4624] = 1
      "0001" when "01001000010001", -- t[4625] = 1
      "0001" when "01001000010010", -- t[4626] = 1
      "0001" when "01001000010011", -- t[4627] = 1
      "0001" when "01001000010100", -- t[4628] = 1
      "0001" when "01001000010101", -- t[4629] = 1
      "0001" when "01001000010110", -- t[4630] = 1
      "0001" when "01001000010111", -- t[4631] = 1
      "0001" when "01001000011000", -- t[4632] = 1
      "0001" when "01001000011001", -- t[4633] = 1
      "0001" when "01001000011010", -- t[4634] = 1
      "0001" when "01001000011011", -- t[4635] = 1
      "0001" when "01001000011100", -- t[4636] = 1
      "0001" when "01001000011101", -- t[4637] = 1
      "0001" when "01001000011110", -- t[4638] = 1
      "0001" when "01001000011111", -- t[4639] = 1
      "0001" when "01001000100000", -- t[4640] = 1
      "0001" when "01001000100001", -- t[4641] = 1
      "0001" when "01001000100010", -- t[4642] = 1
      "0001" when "01001000100011", -- t[4643] = 1
      "0001" when "01001000100100", -- t[4644] = 1
      "0001" when "01001000100101", -- t[4645] = 1
      "0001" when "01001000100110", -- t[4646] = 1
      "0001" when "01001000100111", -- t[4647] = 1
      "0001" when "01001000101000", -- t[4648] = 1
      "0001" when "01001000101001", -- t[4649] = 1
      "0001" when "01001000101010", -- t[4650] = 1
      "0001" when "01001000101011", -- t[4651] = 1
      "0001" when "01001000101100", -- t[4652] = 1
      "0001" when "01001000101101", -- t[4653] = 1
      "0001" when "01001000101110", -- t[4654] = 1
      "0001" when "01001000101111", -- t[4655] = 1
      "0001" when "01001000110000", -- t[4656] = 1
      "0001" when "01001000110001", -- t[4657] = 1
      "0001" when "01001000110010", -- t[4658] = 1
      "0001" when "01001000110011", -- t[4659] = 1
      "0001" when "01001000110100", -- t[4660] = 1
      "0001" when "01001000110101", -- t[4661] = 1
      "0001" when "01001000110110", -- t[4662] = 1
      "0001" when "01001000110111", -- t[4663] = 1
      "0001" when "01001000111000", -- t[4664] = 1
      "0001" when "01001000111001", -- t[4665] = 1
      "0001" when "01001000111010", -- t[4666] = 1
      "0001" when "01001000111011", -- t[4667] = 1
      "0001" when "01001000111100", -- t[4668] = 1
      "0001" when "01001000111101", -- t[4669] = 1
      "0001" when "01001000111110", -- t[4670] = 1
      "0001" when "01001000111111", -- t[4671] = 1
      "0001" when "01001001000000", -- t[4672] = 1
      "0001" when "01001001000001", -- t[4673] = 1
      "0001" when "01001001000010", -- t[4674] = 1
      "0001" when "01001001000011", -- t[4675] = 1
      "0001" when "01001001000100", -- t[4676] = 1
      "0001" when "01001001000101", -- t[4677] = 1
      "0001" when "01001001000110", -- t[4678] = 1
      "0001" when "01001001000111", -- t[4679] = 1
      "0001" when "01001001001000", -- t[4680] = 1
      "0001" when "01001001001001", -- t[4681] = 1
      "0001" when "01001001001010", -- t[4682] = 1
      "0001" when "01001001001011", -- t[4683] = 1
      "0001" when "01001001001100", -- t[4684] = 1
      "0001" when "01001001001101", -- t[4685] = 1
      "0001" when "01001001001110", -- t[4686] = 1
      "0001" when "01001001001111", -- t[4687] = 1
      "0001" when "01001001010000", -- t[4688] = 1
      "0001" when "01001001010001", -- t[4689] = 1
      "0001" when "01001001010010", -- t[4690] = 1
      "0001" when "01001001010011", -- t[4691] = 1
      "0001" when "01001001010100", -- t[4692] = 1
      "0001" when "01001001010101", -- t[4693] = 1
      "0001" when "01001001010110", -- t[4694] = 1
      "0001" when "01001001010111", -- t[4695] = 1
      "0001" when "01001001011000", -- t[4696] = 1
      "0001" when "01001001011001", -- t[4697] = 1
      "0001" when "01001001011010", -- t[4698] = 1
      "0001" when "01001001011011", -- t[4699] = 1
      "0001" when "01001001011100", -- t[4700] = 1
      "0001" when "01001001011101", -- t[4701] = 1
      "0001" when "01001001011110", -- t[4702] = 1
      "0001" when "01001001011111", -- t[4703] = 1
      "0001" when "01001001100000", -- t[4704] = 1
      "0001" when "01001001100001", -- t[4705] = 1
      "0001" when "01001001100010", -- t[4706] = 1
      "0001" when "01001001100011", -- t[4707] = 1
      "0001" when "01001001100100", -- t[4708] = 1
      "0001" when "01001001100101", -- t[4709] = 1
      "0001" when "01001001100110", -- t[4710] = 1
      "0001" when "01001001100111", -- t[4711] = 1
      "0001" when "01001001101000", -- t[4712] = 1
      "0001" when "01001001101001", -- t[4713] = 1
      "0001" when "01001001101010", -- t[4714] = 1
      "0001" when "01001001101011", -- t[4715] = 1
      "0001" when "01001001101100", -- t[4716] = 1
      "0001" when "01001001101101", -- t[4717] = 1
      "0001" when "01001001101110", -- t[4718] = 1
      "0001" when "01001001101111", -- t[4719] = 1
      "0001" when "01001001110000", -- t[4720] = 1
      "0001" when "01001001110001", -- t[4721] = 1
      "0001" when "01001001110010", -- t[4722] = 1
      "0001" when "01001001110011", -- t[4723] = 1
      "0001" when "01001001110100", -- t[4724] = 1
      "0001" when "01001001110101", -- t[4725] = 1
      "0001" when "01001001110110", -- t[4726] = 1
      "0001" when "01001001110111", -- t[4727] = 1
      "0001" when "01001001111000", -- t[4728] = 1
      "0001" when "01001001111001", -- t[4729] = 1
      "0001" when "01001001111010", -- t[4730] = 1
      "0001" when "01001001111011", -- t[4731] = 1
      "0001" when "01001001111100", -- t[4732] = 1
      "0001" when "01001001111101", -- t[4733] = 1
      "0001" when "01001001111110", -- t[4734] = 1
      "0001" when "01001001111111", -- t[4735] = 1
      "0001" when "01001010000000", -- t[4736] = 1
      "0001" when "01001010000001", -- t[4737] = 1
      "0001" when "01001010000010", -- t[4738] = 1
      "0001" when "01001010000011", -- t[4739] = 1
      "0001" when "01001010000100", -- t[4740] = 1
      "0001" when "01001010000101", -- t[4741] = 1
      "0001" when "01001010000110", -- t[4742] = 1
      "0001" when "01001010000111", -- t[4743] = 1
      "0001" when "01001010001000", -- t[4744] = 1
      "0001" when "01001010001001", -- t[4745] = 1
      "0001" when "01001010001010", -- t[4746] = 1
      "0001" when "01001010001011", -- t[4747] = 1
      "0001" when "01001010001100", -- t[4748] = 1
      "0001" when "01001010001101", -- t[4749] = 1
      "0001" when "01001010001110", -- t[4750] = 1
      "0001" when "01001010001111", -- t[4751] = 1
      "0001" when "01001010010000", -- t[4752] = 1
      "0001" when "01001010010001", -- t[4753] = 1
      "0001" when "01001010010010", -- t[4754] = 1
      "0001" when "01001010010011", -- t[4755] = 1
      "0001" when "01001010010100", -- t[4756] = 1
      "0001" when "01001010010101", -- t[4757] = 1
      "0001" when "01001010010110", -- t[4758] = 1
      "0001" when "01001010010111", -- t[4759] = 1
      "0001" when "01001010011000", -- t[4760] = 1
      "0001" when "01001010011001", -- t[4761] = 1
      "0001" when "01001010011010", -- t[4762] = 1
      "0001" when "01001010011011", -- t[4763] = 1
      "0001" when "01001010011100", -- t[4764] = 1
      "0001" when "01001010011101", -- t[4765] = 1
      "0001" when "01001010011110", -- t[4766] = 1
      "0001" when "01001010011111", -- t[4767] = 1
      "0001" when "01001010100000", -- t[4768] = 1
      "0001" when "01001010100001", -- t[4769] = 1
      "0001" when "01001010100010", -- t[4770] = 1
      "0001" when "01001010100011", -- t[4771] = 1
      "0001" when "01001010100100", -- t[4772] = 1
      "0001" when "01001010100101", -- t[4773] = 1
      "0001" when "01001010100110", -- t[4774] = 1
      "0001" when "01001010100111", -- t[4775] = 1
      "0001" when "01001010101000", -- t[4776] = 1
      "0001" when "01001010101001", -- t[4777] = 1
      "0001" when "01001010101010", -- t[4778] = 1
      "0001" when "01001010101011", -- t[4779] = 1
      "0001" when "01001010101100", -- t[4780] = 1
      "0001" when "01001010101101", -- t[4781] = 1
      "0001" when "01001010101110", -- t[4782] = 1
      "0001" when "01001010101111", -- t[4783] = 1
      "0001" when "01001010110000", -- t[4784] = 1
      "0001" when "01001010110001", -- t[4785] = 1
      "0001" when "01001010110010", -- t[4786] = 1
      "0001" when "01001010110011", -- t[4787] = 1
      "0001" when "01001010110100", -- t[4788] = 1
      "0001" when "01001010110101", -- t[4789] = 1
      "0001" when "01001010110110", -- t[4790] = 1
      "0001" when "01001010110111", -- t[4791] = 1
      "0001" when "01001010111000", -- t[4792] = 1
      "0001" when "01001010111001", -- t[4793] = 1
      "0001" when "01001010111010", -- t[4794] = 1
      "0001" when "01001010111011", -- t[4795] = 1
      "0001" when "01001010111100", -- t[4796] = 1
      "0001" when "01001010111101", -- t[4797] = 1
      "0001" when "01001010111110", -- t[4798] = 1
      "0001" when "01001010111111", -- t[4799] = 1
      "0001" when "01001011000000", -- t[4800] = 1
      "0001" when "01001011000001", -- t[4801] = 1
      "0001" when "01001011000010", -- t[4802] = 1
      "0001" when "01001011000011", -- t[4803] = 1
      "0001" when "01001011000100", -- t[4804] = 1
      "0001" when "01001011000101", -- t[4805] = 1
      "0001" when "01001011000110", -- t[4806] = 1
      "0001" when "01001011000111", -- t[4807] = 1
      "0001" when "01001011001000", -- t[4808] = 1
      "0001" when "01001011001001", -- t[4809] = 1
      "0001" when "01001011001010", -- t[4810] = 1
      "0001" when "01001011001011", -- t[4811] = 1
      "0001" when "01001011001100", -- t[4812] = 1
      "0001" when "01001011001101", -- t[4813] = 1
      "0001" when "01001011001110", -- t[4814] = 1
      "0001" when "01001011001111", -- t[4815] = 1
      "0001" when "01001011010000", -- t[4816] = 1
      "0001" when "01001011010001", -- t[4817] = 1
      "0001" when "01001011010010", -- t[4818] = 1
      "0001" when "01001011010011", -- t[4819] = 1
      "0001" when "01001011010100", -- t[4820] = 1
      "0001" when "01001011010101", -- t[4821] = 1
      "0001" when "01001011010110", -- t[4822] = 1
      "0001" when "01001011010111", -- t[4823] = 1
      "0001" when "01001011011000", -- t[4824] = 1
      "0001" when "01001011011001", -- t[4825] = 1
      "0001" when "01001011011010", -- t[4826] = 1
      "0001" when "01001011011011", -- t[4827] = 1
      "0001" when "01001011011100", -- t[4828] = 1
      "0001" when "01001011011101", -- t[4829] = 1
      "0001" when "01001011011110", -- t[4830] = 1
      "0001" when "01001011011111", -- t[4831] = 1
      "0001" when "01001011100000", -- t[4832] = 1
      "0001" when "01001011100001", -- t[4833] = 1
      "0001" when "01001011100010", -- t[4834] = 1
      "0001" when "01001011100011", -- t[4835] = 1
      "0001" when "01001011100100", -- t[4836] = 1
      "0001" when "01001011100101", -- t[4837] = 1
      "0001" when "01001011100110", -- t[4838] = 1
      "0001" when "01001011100111", -- t[4839] = 1
      "0001" when "01001011101000", -- t[4840] = 1
      "0001" when "01001011101001", -- t[4841] = 1
      "0001" when "01001011101010", -- t[4842] = 1
      "0001" when "01001011101011", -- t[4843] = 1
      "0001" when "01001011101100", -- t[4844] = 1
      "0001" when "01001011101101", -- t[4845] = 1
      "0001" when "01001011101110", -- t[4846] = 1
      "0001" when "01001011101111", -- t[4847] = 1
      "0001" when "01001011110000", -- t[4848] = 1
      "0001" when "01001011110001", -- t[4849] = 1
      "0001" when "01001011110010", -- t[4850] = 1
      "0001" when "01001011110011", -- t[4851] = 1
      "0001" when "01001011110100", -- t[4852] = 1
      "0001" when "01001011110101", -- t[4853] = 1
      "0001" when "01001011110110", -- t[4854] = 1
      "0001" when "01001011110111", -- t[4855] = 1
      "0001" when "01001011111000", -- t[4856] = 1
      "0001" when "01001011111001", -- t[4857] = 1
      "0001" when "01001011111010", -- t[4858] = 1
      "0001" when "01001011111011", -- t[4859] = 1
      "0001" when "01001011111100", -- t[4860] = 1
      "0001" when "01001011111101", -- t[4861] = 1
      "0001" when "01001011111110", -- t[4862] = 1
      "0001" when "01001011111111", -- t[4863] = 1
      "0001" when "01001100000000", -- t[4864] = 1
      "0001" when "01001100000001", -- t[4865] = 1
      "0001" when "01001100000010", -- t[4866] = 1
      "0001" when "01001100000011", -- t[4867] = 1
      "0001" when "01001100000100", -- t[4868] = 1
      "0001" when "01001100000101", -- t[4869] = 1
      "0001" when "01001100000110", -- t[4870] = 1
      "0001" when "01001100000111", -- t[4871] = 1
      "0001" when "01001100001000", -- t[4872] = 1
      "0001" when "01001100001001", -- t[4873] = 1
      "0001" when "01001100001010", -- t[4874] = 1
      "0001" when "01001100001011", -- t[4875] = 1
      "0001" when "01001100001100", -- t[4876] = 1
      "0001" when "01001100001101", -- t[4877] = 1
      "0001" when "01001100001110", -- t[4878] = 1
      "0001" when "01001100001111", -- t[4879] = 1
      "0001" when "01001100010000", -- t[4880] = 1
      "0001" when "01001100010001", -- t[4881] = 1
      "0001" when "01001100010010", -- t[4882] = 1
      "0001" when "01001100010011", -- t[4883] = 1
      "0001" when "01001100010100", -- t[4884] = 1
      "0001" when "01001100010101", -- t[4885] = 1
      "0001" when "01001100010110", -- t[4886] = 1
      "0001" when "01001100010111", -- t[4887] = 1
      "0001" when "01001100011000", -- t[4888] = 1
      "0001" when "01001100011001", -- t[4889] = 1
      "0001" when "01001100011010", -- t[4890] = 1
      "0001" when "01001100011011", -- t[4891] = 1
      "0001" when "01001100011100", -- t[4892] = 1
      "0001" when "01001100011101", -- t[4893] = 1
      "0001" when "01001100011110", -- t[4894] = 1
      "0001" when "01001100011111", -- t[4895] = 1
      "0001" when "01001100100000", -- t[4896] = 1
      "0001" when "01001100100001", -- t[4897] = 1
      "0001" when "01001100100010", -- t[4898] = 1
      "0001" when "01001100100011", -- t[4899] = 1
      "0001" when "01001100100100", -- t[4900] = 1
      "0001" when "01001100100101", -- t[4901] = 1
      "0001" when "01001100100110", -- t[4902] = 1
      "0001" when "01001100100111", -- t[4903] = 1
      "0001" when "01001100101000", -- t[4904] = 1
      "0001" when "01001100101001", -- t[4905] = 1
      "0001" when "01001100101010", -- t[4906] = 1
      "0001" when "01001100101011", -- t[4907] = 1
      "0001" when "01001100101100", -- t[4908] = 1
      "0001" when "01001100101101", -- t[4909] = 1
      "0001" when "01001100101110", -- t[4910] = 1
      "0001" when "01001100101111", -- t[4911] = 1
      "0001" when "01001100110000", -- t[4912] = 1
      "0001" when "01001100110001", -- t[4913] = 1
      "0001" when "01001100110010", -- t[4914] = 1
      "0001" when "01001100110011", -- t[4915] = 1
      "0001" when "01001100110100", -- t[4916] = 1
      "0001" when "01001100110101", -- t[4917] = 1
      "0001" when "01001100110110", -- t[4918] = 1
      "0001" when "01001100110111", -- t[4919] = 1
      "0001" when "01001100111000", -- t[4920] = 1
      "0001" when "01001100111001", -- t[4921] = 1
      "0001" when "01001100111010", -- t[4922] = 1
      "0001" when "01001100111011", -- t[4923] = 1
      "0001" when "01001100111100", -- t[4924] = 1
      "0001" when "01001100111101", -- t[4925] = 1
      "0001" when "01001100111110", -- t[4926] = 1
      "0001" when "01001100111111", -- t[4927] = 1
      "0001" when "01001101000000", -- t[4928] = 1
      "0001" when "01001101000001", -- t[4929] = 1
      "0001" when "01001101000010", -- t[4930] = 1
      "0001" when "01001101000011", -- t[4931] = 1
      "0001" when "01001101000100", -- t[4932] = 1
      "0001" when "01001101000101", -- t[4933] = 1
      "0001" when "01001101000110", -- t[4934] = 1
      "0001" when "01001101000111", -- t[4935] = 1
      "0001" when "01001101001000", -- t[4936] = 1
      "0001" when "01001101001001", -- t[4937] = 1
      "0001" when "01001101001010", -- t[4938] = 1
      "0001" when "01001101001011", -- t[4939] = 1
      "0001" when "01001101001100", -- t[4940] = 1
      "0001" when "01001101001101", -- t[4941] = 1
      "0001" when "01001101001110", -- t[4942] = 1
      "0001" when "01001101001111", -- t[4943] = 1
      "0001" when "01001101010000", -- t[4944] = 1
      "0001" when "01001101010001", -- t[4945] = 1
      "0001" when "01001101010010", -- t[4946] = 1
      "0001" when "01001101010011", -- t[4947] = 1
      "0001" when "01001101010100", -- t[4948] = 1
      "0001" when "01001101010101", -- t[4949] = 1
      "0001" when "01001101010110", -- t[4950] = 1
      "0001" when "01001101010111", -- t[4951] = 1
      "0001" when "01001101011000", -- t[4952] = 1
      "0001" when "01001101011001", -- t[4953] = 1
      "0001" when "01001101011010", -- t[4954] = 1
      "0001" when "01001101011011", -- t[4955] = 1
      "0001" when "01001101011100", -- t[4956] = 1
      "0001" when "01001101011101", -- t[4957] = 1
      "0001" when "01001101011110", -- t[4958] = 1
      "0001" when "01001101011111", -- t[4959] = 1
      "0001" when "01001101100000", -- t[4960] = 1
      "0001" when "01001101100001", -- t[4961] = 1
      "0001" when "01001101100010", -- t[4962] = 1
      "0001" when "01001101100011", -- t[4963] = 1
      "0001" when "01001101100100", -- t[4964] = 1
      "0001" when "01001101100101", -- t[4965] = 1
      "0001" when "01001101100110", -- t[4966] = 1
      "0001" when "01001101100111", -- t[4967] = 1
      "0001" when "01001101101000", -- t[4968] = 1
      "0001" when "01001101101001", -- t[4969] = 1
      "0001" when "01001101101010", -- t[4970] = 1
      "0001" when "01001101101011", -- t[4971] = 1
      "0001" when "01001101101100", -- t[4972] = 1
      "0001" when "01001101101101", -- t[4973] = 1
      "0001" when "01001101101110", -- t[4974] = 1
      "0001" when "01001101101111", -- t[4975] = 1
      "0001" when "01001101110000", -- t[4976] = 1
      "0001" when "01001101110001", -- t[4977] = 1
      "0001" when "01001101110010", -- t[4978] = 1
      "0001" when "01001101110011", -- t[4979] = 1
      "0001" when "01001101110100", -- t[4980] = 1
      "0001" when "01001101110101", -- t[4981] = 1
      "0001" when "01001101110110", -- t[4982] = 1
      "0001" when "01001101110111", -- t[4983] = 1
      "0001" when "01001101111000", -- t[4984] = 1
      "0001" when "01001101111001", -- t[4985] = 1
      "0001" when "01001101111010", -- t[4986] = 1
      "0001" when "01001101111011", -- t[4987] = 1
      "0001" when "01001101111100", -- t[4988] = 1
      "0001" when "01001101111101", -- t[4989] = 1
      "0001" when "01001101111110", -- t[4990] = 1
      "0001" when "01001101111111", -- t[4991] = 1
      "0001" when "01001110000000", -- t[4992] = 1
      "0001" when "01001110000001", -- t[4993] = 1
      "0001" when "01001110000010", -- t[4994] = 1
      "0001" when "01001110000011", -- t[4995] = 1
      "0001" when "01001110000100", -- t[4996] = 1
      "0001" when "01001110000101", -- t[4997] = 1
      "0001" when "01001110000110", -- t[4998] = 1
      "0001" when "01001110000111", -- t[4999] = 1
      "0001" when "01001110001000", -- t[5000] = 1
      "0001" when "01001110001001", -- t[5001] = 1
      "0001" when "01001110001010", -- t[5002] = 1
      "0001" when "01001110001011", -- t[5003] = 1
      "0001" when "01001110001100", -- t[5004] = 1
      "0001" when "01001110001101", -- t[5005] = 1
      "0001" when "01001110001110", -- t[5006] = 1
      "0001" when "01001110001111", -- t[5007] = 1
      "0001" when "01001110010000", -- t[5008] = 1
      "0001" when "01001110010001", -- t[5009] = 1
      "0001" when "01001110010010", -- t[5010] = 1
      "0001" when "01001110010011", -- t[5011] = 1
      "0001" when "01001110010100", -- t[5012] = 1
      "0001" when "01001110010101", -- t[5013] = 1
      "0001" when "01001110010110", -- t[5014] = 1
      "0001" when "01001110010111", -- t[5015] = 1
      "0001" when "01001110011000", -- t[5016] = 1
      "0001" when "01001110011001", -- t[5017] = 1
      "0001" when "01001110011010", -- t[5018] = 1
      "0001" when "01001110011011", -- t[5019] = 1
      "0001" when "01001110011100", -- t[5020] = 1
      "0001" when "01001110011101", -- t[5021] = 1
      "0001" when "01001110011110", -- t[5022] = 1
      "0001" when "01001110011111", -- t[5023] = 1
      "0001" when "01001110100000", -- t[5024] = 1
      "0001" when "01001110100001", -- t[5025] = 1
      "0001" when "01001110100010", -- t[5026] = 1
      "0001" when "01001110100011", -- t[5027] = 1
      "0001" when "01001110100100", -- t[5028] = 1
      "0001" when "01001110100101", -- t[5029] = 1
      "0001" when "01001110100110", -- t[5030] = 1
      "0001" when "01001110100111", -- t[5031] = 1
      "0001" when "01001110101000", -- t[5032] = 1
      "0001" when "01001110101001", -- t[5033] = 1
      "0001" when "01001110101010", -- t[5034] = 1
      "0001" when "01001110101011", -- t[5035] = 1
      "0001" when "01001110101100", -- t[5036] = 1
      "0001" when "01001110101101", -- t[5037] = 1
      "0001" when "01001110101110", -- t[5038] = 1
      "0001" when "01001110101111", -- t[5039] = 1
      "0001" when "01001110110000", -- t[5040] = 1
      "0001" when "01001110110001", -- t[5041] = 1
      "0001" when "01001110110010", -- t[5042] = 1
      "0001" when "01001110110011", -- t[5043] = 1
      "0001" when "01001110110100", -- t[5044] = 1
      "0001" when "01001110110101", -- t[5045] = 1
      "0001" when "01001110110110", -- t[5046] = 1
      "0001" when "01001110110111", -- t[5047] = 1
      "0001" when "01001110111000", -- t[5048] = 1
      "0001" when "01001110111001", -- t[5049] = 1
      "0001" when "01001110111010", -- t[5050] = 1
      "0001" when "01001110111011", -- t[5051] = 1
      "0001" when "01001110111100", -- t[5052] = 1
      "0001" when "01001110111101", -- t[5053] = 1
      "0001" when "01001110111110", -- t[5054] = 1
      "0001" when "01001110111111", -- t[5055] = 1
      "0001" when "01001111000000", -- t[5056] = 1
      "0001" when "01001111000001", -- t[5057] = 1
      "0001" when "01001111000010", -- t[5058] = 1
      "0001" when "01001111000011", -- t[5059] = 1
      "0001" when "01001111000100", -- t[5060] = 1
      "0001" when "01001111000101", -- t[5061] = 1
      "0001" when "01001111000110", -- t[5062] = 1
      "0001" when "01001111000111", -- t[5063] = 1
      "0001" when "01001111001000", -- t[5064] = 1
      "0001" when "01001111001001", -- t[5065] = 1
      "0001" when "01001111001010", -- t[5066] = 1
      "0001" when "01001111001011", -- t[5067] = 1
      "0001" when "01001111001100", -- t[5068] = 1
      "0001" when "01001111001101", -- t[5069] = 1
      "0001" when "01001111001110", -- t[5070] = 1
      "0001" when "01001111001111", -- t[5071] = 1
      "0001" when "01001111010000", -- t[5072] = 1
      "0001" when "01001111010001", -- t[5073] = 1
      "0001" when "01001111010010", -- t[5074] = 1
      "0001" when "01001111010011", -- t[5075] = 1
      "0001" when "01001111010100", -- t[5076] = 1
      "0001" when "01001111010101", -- t[5077] = 1
      "0001" when "01001111010110", -- t[5078] = 1
      "0001" when "01001111010111", -- t[5079] = 1
      "0001" when "01001111011000", -- t[5080] = 1
      "0001" when "01001111011001", -- t[5081] = 1
      "0001" when "01001111011010", -- t[5082] = 1
      "0001" when "01001111011011", -- t[5083] = 1
      "0001" when "01001111011100", -- t[5084] = 1
      "0001" when "01001111011101", -- t[5085] = 1
      "0001" when "01001111011110", -- t[5086] = 1
      "0001" when "01001111011111", -- t[5087] = 1
      "0001" when "01001111100000", -- t[5088] = 1
      "0001" when "01001111100001", -- t[5089] = 1
      "0001" when "01001111100010", -- t[5090] = 1
      "0001" when "01001111100011", -- t[5091] = 1
      "0001" when "01001111100100", -- t[5092] = 1
      "0001" when "01001111100101", -- t[5093] = 1
      "0001" when "01001111100110", -- t[5094] = 1
      "0001" when "01001111100111", -- t[5095] = 1
      "0001" when "01001111101000", -- t[5096] = 1
      "0001" when "01001111101001", -- t[5097] = 1
      "0001" when "01001111101010", -- t[5098] = 1
      "0001" when "01001111101011", -- t[5099] = 1
      "0001" when "01001111101100", -- t[5100] = 1
      "0001" when "01001111101101", -- t[5101] = 1
      "0001" when "01001111101110", -- t[5102] = 1
      "0001" when "01001111101111", -- t[5103] = 1
      "0001" when "01001111110000", -- t[5104] = 1
      "0001" when "01001111110001", -- t[5105] = 1
      "0001" when "01001111110010", -- t[5106] = 1
      "0001" when "01001111110011", -- t[5107] = 1
      "0001" when "01001111110100", -- t[5108] = 1
      "0001" when "01001111110101", -- t[5109] = 1
      "0001" when "01001111110110", -- t[5110] = 1
      "0001" when "01001111110111", -- t[5111] = 1
      "0001" when "01001111111000", -- t[5112] = 1
      "0001" when "01001111111001", -- t[5113] = 1
      "0001" when "01001111111010", -- t[5114] = 1
      "0001" when "01001111111011", -- t[5115] = 1
      "0001" when "01001111111100", -- t[5116] = 1
      "0001" when "01001111111101", -- t[5117] = 1
      "0001" when "01001111111110", -- t[5118] = 1
      "0001" when "01001111111111", -- t[5119] = 1
      "0001" when "01010000000000", -- t[5120] = 1
      "0001" when "01010000000001", -- t[5121] = 1
      "0001" when "01010000000010", -- t[5122] = 1
      "0001" when "01010000000011", -- t[5123] = 1
      "0001" when "01010000000100", -- t[5124] = 1
      "0001" when "01010000000101", -- t[5125] = 1
      "0001" when "01010000000110", -- t[5126] = 1
      "0001" when "01010000000111", -- t[5127] = 1
      "0001" when "01010000001000", -- t[5128] = 1
      "0001" when "01010000001001", -- t[5129] = 1
      "0001" when "01010000001010", -- t[5130] = 1
      "0001" when "01010000001011", -- t[5131] = 1
      "0001" when "01010000001100", -- t[5132] = 1
      "0001" when "01010000001101", -- t[5133] = 1
      "0001" when "01010000001110", -- t[5134] = 1
      "0001" when "01010000001111", -- t[5135] = 1
      "0001" when "01010000010000", -- t[5136] = 1
      "0001" when "01010000010001", -- t[5137] = 1
      "0001" when "01010000010010", -- t[5138] = 1
      "0001" when "01010000010011", -- t[5139] = 1
      "0001" when "01010000010100", -- t[5140] = 1
      "0001" when "01010000010101", -- t[5141] = 1
      "0001" when "01010000010110", -- t[5142] = 1
      "0001" when "01010000010111", -- t[5143] = 1
      "0001" when "01010000011000", -- t[5144] = 1
      "0001" when "01010000011001", -- t[5145] = 1
      "0001" when "01010000011010", -- t[5146] = 1
      "0001" when "01010000011011", -- t[5147] = 1
      "0001" when "01010000011100", -- t[5148] = 1
      "0001" when "01010000011101", -- t[5149] = 1
      "0001" when "01010000011110", -- t[5150] = 1
      "0001" when "01010000011111", -- t[5151] = 1
      "0001" when "01010000100000", -- t[5152] = 1
      "0001" when "01010000100001", -- t[5153] = 1
      "0001" when "01010000100010", -- t[5154] = 1
      "0001" when "01010000100011", -- t[5155] = 1
      "0001" when "01010000100100", -- t[5156] = 1
      "0001" when "01010000100101", -- t[5157] = 1
      "0001" when "01010000100110", -- t[5158] = 1
      "0001" when "01010000100111", -- t[5159] = 1
      "0001" when "01010000101000", -- t[5160] = 1
      "0001" when "01010000101001", -- t[5161] = 1
      "0001" when "01010000101010", -- t[5162] = 1
      "0001" when "01010000101011", -- t[5163] = 1
      "0001" when "01010000101100", -- t[5164] = 1
      "0001" when "01010000101101", -- t[5165] = 1
      "0001" when "01010000101110", -- t[5166] = 1
      "0001" when "01010000101111", -- t[5167] = 1
      "0001" when "01010000110000", -- t[5168] = 1
      "0001" when "01010000110001", -- t[5169] = 1
      "0001" when "01010000110010", -- t[5170] = 1
      "0001" when "01010000110011", -- t[5171] = 1
      "0001" when "01010000110100", -- t[5172] = 1
      "0001" when "01010000110101", -- t[5173] = 1
      "0001" when "01010000110110", -- t[5174] = 1
      "0001" when "01010000110111", -- t[5175] = 1
      "0001" when "01010000111000", -- t[5176] = 1
      "0001" when "01010000111001", -- t[5177] = 1
      "0001" when "01010000111010", -- t[5178] = 1
      "0001" when "01010000111011", -- t[5179] = 1
      "0001" when "01010000111100", -- t[5180] = 1
      "0001" when "01010000111101", -- t[5181] = 1
      "0001" when "01010000111110", -- t[5182] = 1
      "0001" when "01010000111111", -- t[5183] = 1
      "0001" when "01010001000000", -- t[5184] = 1
      "0001" when "01010001000001", -- t[5185] = 1
      "0001" when "01010001000010", -- t[5186] = 1
      "0001" when "01010001000011", -- t[5187] = 1
      "0001" when "01010001000100", -- t[5188] = 1
      "0001" when "01010001000101", -- t[5189] = 1
      "0001" when "01010001000110", -- t[5190] = 1
      "0001" when "01010001000111", -- t[5191] = 1
      "0001" when "01010001001000", -- t[5192] = 1
      "0001" when "01010001001001", -- t[5193] = 1
      "0001" when "01010001001010", -- t[5194] = 1
      "0001" when "01010001001011", -- t[5195] = 1
      "0001" when "01010001001100", -- t[5196] = 1
      "0001" when "01010001001101", -- t[5197] = 1
      "0001" when "01010001001110", -- t[5198] = 1
      "0001" when "01010001001111", -- t[5199] = 1
      "0001" when "01010001010000", -- t[5200] = 1
      "0001" when "01010001010001", -- t[5201] = 1
      "0001" when "01010001010010", -- t[5202] = 1
      "0001" when "01010001010011", -- t[5203] = 1
      "0001" when "01010001010100", -- t[5204] = 1
      "0001" when "01010001010101", -- t[5205] = 1
      "0001" when "01010001010110", -- t[5206] = 1
      "0001" when "01010001010111", -- t[5207] = 1
      "0001" when "01010001011000", -- t[5208] = 1
      "0001" when "01010001011001", -- t[5209] = 1
      "0001" when "01010001011010", -- t[5210] = 1
      "0001" when "01010001011011", -- t[5211] = 1
      "0001" when "01010001011100", -- t[5212] = 1
      "0001" when "01010001011101", -- t[5213] = 1
      "0001" when "01010001011110", -- t[5214] = 1
      "0001" when "01010001011111", -- t[5215] = 1
      "0001" when "01010001100000", -- t[5216] = 1
      "0001" when "01010001100001", -- t[5217] = 1
      "0001" when "01010001100010", -- t[5218] = 1
      "0001" when "01010001100011", -- t[5219] = 1
      "0001" when "01010001100100", -- t[5220] = 1
      "0001" when "01010001100101", -- t[5221] = 1
      "0001" when "01010001100110", -- t[5222] = 1
      "0001" when "01010001100111", -- t[5223] = 1
      "0001" when "01010001101000", -- t[5224] = 1
      "0001" when "01010001101001", -- t[5225] = 1
      "0001" when "01010001101010", -- t[5226] = 1
      "0001" when "01010001101011", -- t[5227] = 1
      "0001" when "01010001101100", -- t[5228] = 1
      "0001" when "01010001101101", -- t[5229] = 1
      "0001" when "01010001101110", -- t[5230] = 1
      "0001" when "01010001101111", -- t[5231] = 1
      "0001" when "01010001110000", -- t[5232] = 1
      "0001" when "01010001110001", -- t[5233] = 1
      "0001" when "01010001110010", -- t[5234] = 1
      "0001" when "01010001110011", -- t[5235] = 1
      "0001" when "01010001110100", -- t[5236] = 1
      "0001" when "01010001110101", -- t[5237] = 1
      "0001" when "01010001110110", -- t[5238] = 1
      "0001" when "01010001110111", -- t[5239] = 1
      "0001" when "01010001111000", -- t[5240] = 1
      "0001" when "01010001111001", -- t[5241] = 1
      "0001" when "01010001111010", -- t[5242] = 1
      "0001" when "01010001111011", -- t[5243] = 1
      "0001" when "01010001111100", -- t[5244] = 1
      "0001" when "01010001111101", -- t[5245] = 1
      "0001" when "01010001111110", -- t[5246] = 1
      "0001" when "01010001111111", -- t[5247] = 1
      "0001" when "01010010000000", -- t[5248] = 1
      "0001" when "01010010000001", -- t[5249] = 1
      "0001" when "01010010000010", -- t[5250] = 1
      "0001" when "01010010000011", -- t[5251] = 1
      "0001" when "01010010000100", -- t[5252] = 1
      "0001" when "01010010000101", -- t[5253] = 1
      "0001" when "01010010000110", -- t[5254] = 1
      "0001" when "01010010000111", -- t[5255] = 1
      "0001" when "01010010001000", -- t[5256] = 1
      "0001" when "01010010001001", -- t[5257] = 1
      "0001" when "01010010001010", -- t[5258] = 1
      "0001" when "01010010001011", -- t[5259] = 1
      "0001" when "01010010001100", -- t[5260] = 1
      "0001" when "01010010001101", -- t[5261] = 1
      "0001" when "01010010001110", -- t[5262] = 1
      "0001" when "01010010001111", -- t[5263] = 1
      "0001" when "01010010010000", -- t[5264] = 1
      "0001" when "01010010010001", -- t[5265] = 1
      "0001" when "01010010010010", -- t[5266] = 1
      "0001" when "01010010010011", -- t[5267] = 1
      "0001" when "01010010010100", -- t[5268] = 1
      "0001" when "01010010010101", -- t[5269] = 1
      "0001" when "01010010010110", -- t[5270] = 1
      "0001" when "01010010010111", -- t[5271] = 1
      "0001" when "01010010011000", -- t[5272] = 1
      "0001" when "01010010011001", -- t[5273] = 1
      "0001" when "01010010011010", -- t[5274] = 1
      "0001" when "01010010011011", -- t[5275] = 1
      "0001" when "01010010011100", -- t[5276] = 1
      "0001" when "01010010011101", -- t[5277] = 1
      "0001" when "01010010011110", -- t[5278] = 1
      "0001" when "01010010011111", -- t[5279] = 1
      "0001" when "01010010100000", -- t[5280] = 1
      "0001" when "01010010100001", -- t[5281] = 1
      "0001" when "01010010100010", -- t[5282] = 1
      "0001" when "01010010100011", -- t[5283] = 1
      "0001" when "01010010100100", -- t[5284] = 1
      "0001" when "01010010100101", -- t[5285] = 1
      "0001" when "01010010100110", -- t[5286] = 1
      "0001" when "01010010100111", -- t[5287] = 1
      "0001" when "01010010101000", -- t[5288] = 1
      "0001" when "01010010101001", -- t[5289] = 1
      "0001" when "01010010101010", -- t[5290] = 1
      "0001" when "01010010101011", -- t[5291] = 1
      "0001" when "01010010101100", -- t[5292] = 1
      "0001" when "01010010101101", -- t[5293] = 1
      "0001" when "01010010101110", -- t[5294] = 1
      "0001" when "01010010101111", -- t[5295] = 1
      "0001" when "01010010110000", -- t[5296] = 1
      "0001" when "01010010110001", -- t[5297] = 1
      "0001" when "01010010110010", -- t[5298] = 1
      "0001" when "01010010110011", -- t[5299] = 1
      "0001" when "01010010110100", -- t[5300] = 1
      "0001" when "01010010110101", -- t[5301] = 1
      "0001" when "01010010110110", -- t[5302] = 1
      "0001" when "01010010110111", -- t[5303] = 1
      "0001" when "01010010111000", -- t[5304] = 1
      "0001" when "01010010111001", -- t[5305] = 1
      "0001" when "01010010111010", -- t[5306] = 1
      "0001" when "01010010111011", -- t[5307] = 1
      "0001" when "01010010111100", -- t[5308] = 1
      "0001" when "01010010111101", -- t[5309] = 1
      "0001" when "01010010111110", -- t[5310] = 1
      "0001" when "01010010111111", -- t[5311] = 1
      "0001" when "01010011000000", -- t[5312] = 1
      "0001" when "01010011000001", -- t[5313] = 1
      "0001" when "01010011000010", -- t[5314] = 1
      "0001" when "01010011000011", -- t[5315] = 1
      "0001" when "01010011000100", -- t[5316] = 1
      "0001" when "01010011000101", -- t[5317] = 1
      "0001" when "01010011000110", -- t[5318] = 1
      "0001" when "01010011000111", -- t[5319] = 1
      "0001" when "01010011001000", -- t[5320] = 1
      "0001" when "01010011001001", -- t[5321] = 1
      "0001" when "01010011001010", -- t[5322] = 1
      "0001" when "01010011001011", -- t[5323] = 1
      "0001" when "01010011001100", -- t[5324] = 1
      "0001" when "01010011001101", -- t[5325] = 1
      "0001" when "01010011001110", -- t[5326] = 1
      "0001" when "01010011001111", -- t[5327] = 1
      "0001" when "01010011010000", -- t[5328] = 1
      "0001" when "01010011010001", -- t[5329] = 1
      "0001" when "01010011010010", -- t[5330] = 1
      "0001" when "01010011010011", -- t[5331] = 1
      "0001" when "01010011010100", -- t[5332] = 1
      "0001" when "01010011010101", -- t[5333] = 1
      "0001" when "01010011010110", -- t[5334] = 1
      "0001" when "01010011010111", -- t[5335] = 1
      "0001" when "01010011011000", -- t[5336] = 1
      "0001" when "01010011011001", -- t[5337] = 1
      "0001" when "01010011011010", -- t[5338] = 1
      "0001" when "01010011011011", -- t[5339] = 1
      "0001" when "01010011011100", -- t[5340] = 1
      "0001" when "01010011011101", -- t[5341] = 1
      "0001" when "01010011011110", -- t[5342] = 1
      "0001" when "01010011011111", -- t[5343] = 1
      "0001" when "01010011100000", -- t[5344] = 1
      "0001" when "01010011100001", -- t[5345] = 1
      "0001" when "01010011100010", -- t[5346] = 1
      "0001" when "01010011100011", -- t[5347] = 1
      "0001" when "01010011100100", -- t[5348] = 1
      "0001" when "01010011100101", -- t[5349] = 1
      "0001" when "01010011100110", -- t[5350] = 1
      "0001" when "01010011100111", -- t[5351] = 1
      "0001" when "01010011101000", -- t[5352] = 1
      "0001" when "01010011101001", -- t[5353] = 1
      "0001" when "01010011101010", -- t[5354] = 1
      "0001" when "01010011101011", -- t[5355] = 1
      "0001" when "01010011101100", -- t[5356] = 1
      "0001" when "01010011101101", -- t[5357] = 1
      "0001" when "01010011101110", -- t[5358] = 1
      "0001" when "01010011101111", -- t[5359] = 1
      "0001" when "01010011110000", -- t[5360] = 1
      "0001" when "01010011110001", -- t[5361] = 1
      "0001" when "01010011110010", -- t[5362] = 1
      "0001" when "01010011110011", -- t[5363] = 1
      "0001" when "01010011110100", -- t[5364] = 1
      "0001" when "01010011110101", -- t[5365] = 1
      "0001" when "01010011110110", -- t[5366] = 1
      "0001" when "01010011110111", -- t[5367] = 1
      "0001" when "01010011111000", -- t[5368] = 1
      "0001" when "01010011111001", -- t[5369] = 1
      "0001" when "01010011111010", -- t[5370] = 1
      "0001" when "01010011111011", -- t[5371] = 1
      "0001" when "01010011111100", -- t[5372] = 1
      "0001" when "01010011111101", -- t[5373] = 1
      "0001" when "01010011111110", -- t[5374] = 1
      "0001" when "01010011111111", -- t[5375] = 1
      "0001" when "01010100000000", -- t[5376] = 1
      "0001" when "01010100000001", -- t[5377] = 1
      "0001" when "01010100000010", -- t[5378] = 1
      "0001" when "01010100000011", -- t[5379] = 1
      "0001" when "01010100000100", -- t[5380] = 1
      "0001" when "01010100000101", -- t[5381] = 1
      "0001" when "01010100000110", -- t[5382] = 1
      "0001" when "01010100000111", -- t[5383] = 1
      "0001" when "01010100001000", -- t[5384] = 1
      "0001" when "01010100001001", -- t[5385] = 1
      "0001" when "01010100001010", -- t[5386] = 1
      "0001" when "01010100001011", -- t[5387] = 1
      "0001" when "01010100001100", -- t[5388] = 1
      "0001" when "01010100001101", -- t[5389] = 1
      "0001" when "01010100001110", -- t[5390] = 1
      "0001" when "01010100001111", -- t[5391] = 1
      "0001" when "01010100010000", -- t[5392] = 1
      "0001" when "01010100010001", -- t[5393] = 1
      "0001" when "01010100010010", -- t[5394] = 1
      "0001" when "01010100010011", -- t[5395] = 1
      "0001" when "01010100010100", -- t[5396] = 1
      "0001" when "01010100010101", -- t[5397] = 1
      "0001" when "01010100010110", -- t[5398] = 1
      "0001" when "01010100010111", -- t[5399] = 1
      "0001" when "01010100011000", -- t[5400] = 1
      "0001" when "01010100011001", -- t[5401] = 1
      "0001" when "01010100011010", -- t[5402] = 1
      "0001" when "01010100011011", -- t[5403] = 1
      "0001" when "01010100011100", -- t[5404] = 1
      "0001" when "01010100011101", -- t[5405] = 1
      "0001" when "01010100011110", -- t[5406] = 1
      "0001" when "01010100011111", -- t[5407] = 1
      "0001" when "01010100100000", -- t[5408] = 1
      "0001" when "01010100100001", -- t[5409] = 1
      "0001" when "01010100100010", -- t[5410] = 1
      "0001" when "01010100100011", -- t[5411] = 1
      "0001" when "01010100100100", -- t[5412] = 1
      "0001" when "01010100100101", -- t[5413] = 1
      "0001" when "01010100100110", -- t[5414] = 1
      "0001" when "01010100100111", -- t[5415] = 1
      "0001" when "01010100101000", -- t[5416] = 1
      "0001" when "01010100101001", -- t[5417] = 1
      "0001" when "01010100101010", -- t[5418] = 1
      "0001" when "01010100101011", -- t[5419] = 1
      "0001" when "01010100101100", -- t[5420] = 1
      "0001" when "01010100101101", -- t[5421] = 1
      "0001" when "01010100101110", -- t[5422] = 1
      "0001" when "01010100101111", -- t[5423] = 1
      "0001" when "01010100110000", -- t[5424] = 1
      "0001" when "01010100110001", -- t[5425] = 1
      "0001" when "01010100110010", -- t[5426] = 1
      "0001" when "01010100110011", -- t[5427] = 1
      "0001" when "01010100110100", -- t[5428] = 1
      "0001" when "01010100110101", -- t[5429] = 1
      "0001" when "01010100110110", -- t[5430] = 1
      "0001" when "01010100110111", -- t[5431] = 1
      "0001" when "01010100111000", -- t[5432] = 1
      "0001" when "01010100111001", -- t[5433] = 1
      "0001" when "01010100111010", -- t[5434] = 1
      "0001" when "01010100111011", -- t[5435] = 1
      "0001" when "01010100111100", -- t[5436] = 1
      "0001" when "01010100111101", -- t[5437] = 1
      "0001" when "01010100111110", -- t[5438] = 1
      "0001" when "01010100111111", -- t[5439] = 1
      "0001" when "01010101000000", -- t[5440] = 1
      "0001" when "01010101000001", -- t[5441] = 1
      "0001" when "01010101000010", -- t[5442] = 1
      "0001" when "01010101000011", -- t[5443] = 1
      "0001" when "01010101000100", -- t[5444] = 1
      "0001" when "01010101000101", -- t[5445] = 1
      "0001" when "01010101000110", -- t[5446] = 1
      "0001" when "01010101000111", -- t[5447] = 1
      "0001" when "01010101001000", -- t[5448] = 1
      "0001" when "01010101001001", -- t[5449] = 1
      "0001" when "01010101001010", -- t[5450] = 1
      "0001" when "01010101001011", -- t[5451] = 1
      "0001" when "01010101001100", -- t[5452] = 1
      "0001" when "01010101001101", -- t[5453] = 1
      "0001" when "01010101001110", -- t[5454] = 1
      "0001" when "01010101001111", -- t[5455] = 1
      "0001" when "01010101010000", -- t[5456] = 1
      "0001" when "01010101010001", -- t[5457] = 1
      "0001" when "01010101010010", -- t[5458] = 1
      "0001" when "01010101010011", -- t[5459] = 1
      "0001" when "01010101010100", -- t[5460] = 1
      "0001" when "01010101010101", -- t[5461] = 1
      "0001" when "01010101010110", -- t[5462] = 1
      "0001" when "01010101010111", -- t[5463] = 1
      "0001" when "01010101011000", -- t[5464] = 1
      "0001" when "01010101011001", -- t[5465] = 1
      "0001" when "01010101011010", -- t[5466] = 1
      "0001" when "01010101011011", -- t[5467] = 1
      "0001" when "01010101011100", -- t[5468] = 1
      "0001" when "01010101011101", -- t[5469] = 1
      "0001" when "01010101011110", -- t[5470] = 1
      "0001" when "01010101011111", -- t[5471] = 1
      "0001" when "01010101100000", -- t[5472] = 1
      "0001" when "01010101100001", -- t[5473] = 1
      "0001" when "01010101100010", -- t[5474] = 1
      "0001" when "01010101100011", -- t[5475] = 1
      "0001" when "01010101100100", -- t[5476] = 1
      "0001" when "01010101100101", -- t[5477] = 1
      "0001" when "01010101100110", -- t[5478] = 1
      "0001" when "01010101100111", -- t[5479] = 1
      "0001" when "01010101101000", -- t[5480] = 1
      "0001" when "01010101101001", -- t[5481] = 1
      "0001" when "01010101101010", -- t[5482] = 1
      "0001" when "01010101101011", -- t[5483] = 1
      "0001" when "01010101101100", -- t[5484] = 1
      "0001" when "01010101101101", -- t[5485] = 1
      "0001" when "01010101101110", -- t[5486] = 1
      "0001" when "01010101101111", -- t[5487] = 1
      "0001" when "01010101110000", -- t[5488] = 1
      "0001" when "01010101110001", -- t[5489] = 1
      "0001" when "01010101110010", -- t[5490] = 1
      "0001" when "01010101110011", -- t[5491] = 1
      "0001" when "01010101110100", -- t[5492] = 1
      "0001" when "01010101110101", -- t[5493] = 1
      "0001" when "01010101110110", -- t[5494] = 1
      "0001" when "01010101110111", -- t[5495] = 1
      "0001" when "01010101111000", -- t[5496] = 1
      "0001" when "01010101111001", -- t[5497] = 1
      "0001" when "01010101111010", -- t[5498] = 1
      "0001" when "01010101111011", -- t[5499] = 1
      "0001" when "01010101111100", -- t[5500] = 1
      "0001" when "01010101111101", -- t[5501] = 1
      "0001" when "01010101111110", -- t[5502] = 1
      "0001" when "01010101111111", -- t[5503] = 1
      "0001" when "01010110000000", -- t[5504] = 1
      "0001" when "01010110000001", -- t[5505] = 1
      "0001" when "01010110000010", -- t[5506] = 1
      "0001" when "01010110000011", -- t[5507] = 1
      "0001" when "01010110000100", -- t[5508] = 1
      "0001" when "01010110000101", -- t[5509] = 1
      "0001" when "01010110000110", -- t[5510] = 1
      "0001" when "01010110000111", -- t[5511] = 1
      "0001" when "01010110001000", -- t[5512] = 1
      "0001" when "01010110001001", -- t[5513] = 1
      "0001" when "01010110001010", -- t[5514] = 1
      "0001" when "01010110001011", -- t[5515] = 1
      "0001" when "01010110001100", -- t[5516] = 1
      "0001" when "01010110001101", -- t[5517] = 1
      "0001" when "01010110001110", -- t[5518] = 1
      "0001" when "01010110001111", -- t[5519] = 1
      "0001" when "01010110010000", -- t[5520] = 1
      "0001" when "01010110010001", -- t[5521] = 1
      "0001" when "01010110010010", -- t[5522] = 1
      "0001" when "01010110010011", -- t[5523] = 1
      "0001" when "01010110010100", -- t[5524] = 1
      "0001" when "01010110010101", -- t[5525] = 1
      "0001" when "01010110010110", -- t[5526] = 1
      "0001" when "01010110010111", -- t[5527] = 1
      "0001" when "01010110011000", -- t[5528] = 1
      "0001" when "01010110011001", -- t[5529] = 1
      "0001" when "01010110011010", -- t[5530] = 1
      "0001" when "01010110011011", -- t[5531] = 1
      "0001" when "01010110011100", -- t[5532] = 1
      "0001" when "01010110011101", -- t[5533] = 1
      "0001" when "01010110011110", -- t[5534] = 1
      "0001" when "01010110011111", -- t[5535] = 1
      "0001" when "01010110100000", -- t[5536] = 1
      "0001" when "01010110100001", -- t[5537] = 1
      "0001" when "01010110100010", -- t[5538] = 1
      "0001" when "01010110100011", -- t[5539] = 1
      "0001" when "01010110100100", -- t[5540] = 1
      "0001" when "01010110100101", -- t[5541] = 1
      "0001" when "01010110100110", -- t[5542] = 1
      "0001" when "01010110100111", -- t[5543] = 1
      "0001" when "01010110101000", -- t[5544] = 1
      "0001" when "01010110101001", -- t[5545] = 1
      "0001" when "01010110101010", -- t[5546] = 1
      "0001" when "01010110101011", -- t[5547] = 1
      "0001" when "01010110101100", -- t[5548] = 1
      "0001" when "01010110101101", -- t[5549] = 1
      "0001" when "01010110101110", -- t[5550] = 1
      "0001" when "01010110101111", -- t[5551] = 1
      "0001" when "01010110110000", -- t[5552] = 1
      "0001" when "01010110110001", -- t[5553] = 1
      "0001" when "01010110110010", -- t[5554] = 1
      "0001" when "01010110110011", -- t[5555] = 1
      "0001" when "01010110110100", -- t[5556] = 1
      "0001" when "01010110110101", -- t[5557] = 1
      "0001" when "01010110110110", -- t[5558] = 1
      "0001" when "01010110110111", -- t[5559] = 1
      "0001" when "01010110111000", -- t[5560] = 1
      "0001" when "01010110111001", -- t[5561] = 1
      "0001" when "01010110111010", -- t[5562] = 1
      "0001" when "01010110111011", -- t[5563] = 1
      "0001" when "01010110111100", -- t[5564] = 1
      "0001" when "01010110111101", -- t[5565] = 1
      "0001" when "01010110111110", -- t[5566] = 1
      "0001" when "01010110111111", -- t[5567] = 1
      "0001" when "01010111000000", -- t[5568] = 1
      "0001" when "01010111000001", -- t[5569] = 1
      "0001" when "01010111000010", -- t[5570] = 1
      "0001" when "01010111000011", -- t[5571] = 1
      "0001" when "01010111000100", -- t[5572] = 1
      "0001" when "01010111000101", -- t[5573] = 1
      "0001" when "01010111000110", -- t[5574] = 1
      "0001" when "01010111000111", -- t[5575] = 1
      "0001" when "01010111001000", -- t[5576] = 1
      "0001" when "01010111001001", -- t[5577] = 1
      "0001" when "01010111001010", -- t[5578] = 1
      "0001" when "01010111001011", -- t[5579] = 1
      "0001" when "01010111001100", -- t[5580] = 1
      "0001" when "01010111001101", -- t[5581] = 1
      "0001" when "01010111001110", -- t[5582] = 1
      "0001" when "01010111001111", -- t[5583] = 1
      "0001" when "01010111010000", -- t[5584] = 1
      "0001" when "01010111010001", -- t[5585] = 1
      "0001" when "01010111010010", -- t[5586] = 1
      "0001" when "01010111010011", -- t[5587] = 1
      "0001" when "01010111010100", -- t[5588] = 1
      "0001" when "01010111010101", -- t[5589] = 1
      "0001" when "01010111010110", -- t[5590] = 1
      "0001" when "01010111010111", -- t[5591] = 1
      "0001" when "01010111011000", -- t[5592] = 1
      "0001" when "01010111011001", -- t[5593] = 1
      "0001" when "01010111011010", -- t[5594] = 1
      "0001" when "01010111011011", -- t[5595] = 1
      "0001" when "01010111011100", -- t[5596] = 1
      "0001" when "01010111011101", -- t[5597] = 1
      "0001" when "01010111011110", -- t[5598] = 1
      "0001" when "01010111011111", -- t[5599] = 1
      "0001" when "01010111100000", -- t[5600] = 1
      "0001" when "01010111100001", -- t[5601] = 1
      "0001" when "01010111100010", -- t[5602] = 1
      "0001" when "01010111100011", -- t[5603] = 1
      "0001" when "01010111100100", -- t[5604] = 1
      "0001" when "01010111100101", -- t[5605] = 1
      "0001" when "01010111100110", -- t[5606] = 1
      "0001" when "01010111100111", -- t[5607] = 1
      "0001" when "01010111101000", -- t[5608] = 1
      "0001" when "01010111101001", -- t[5609] = 1
      "0001" when "01010111101010", -- t[5610] = 1
      "0001" when "01010111101011", -- t[5611] = 1
      "0001" when "01010111101100", -- t[5612] = 1
      "0001" when "01010111101101", -- t[5613] = 1
      "0001" when "01010111101110", -- t[5614] = 1
      "0001" when "01010111101111", -- t[5615] = 1
      "0001" when "01010111110000", -- t[5616] = 1
      "0001" when "01010111110001", -- t[5617] = 1
      "0001" when "01010111110010", -- t[5618] = 1
      "0001" when "01010111110011", -- t[5619] = 1
      "0001" when "01010111110100", -- t[5620] = 1
      "0001" when "01010111110101", -- t[5621] = 1
      "0001" when "01010111110110", -- t[5622] = 1
      "0001" when "01010111110111", -- t[5623] = 1
      "0001" when "01010111111000", -- t[5624] = 1
      "0001" when "01010111111001", -- t[5625] = 1
      "0001" when "01010111111010", -- t[5626] = 1
      "0001" when "01010111111011", -- t[5627] = 1
      "0001" when "01010111111100", -- t[5628] = 1
      "0001" when "01010111111101", -- t[5629] = 1
      "0001" when "01010111111110", -- t[5630] = 1
      "0001" when "01010111111111", -- t[5631] = 1
      "0001" when "01011000000000", -- t[5632] = 1
      "0001" when "01011000000001", -- t[5633] = 1
      "0001" when "01011000000010", -- t[5634] = 1
      "0001" when "01011000000011", -- t[5635] = 1
      "0001" when "01011000000100", -- t[5636] = 1
      "0001" when "01011000000101", -- t[5637] = 1
      "0001" when "01011000000110", -- t[5638] = 1
      "0001" when "01011000000111", -- t[5639] = 1
      "0001" when "01011000001000", -- t[5640] = 1
      "0001" when "01011000001001", -- t[5641] = 1
      "0001" when "01011000001010", -- t[5642] = 1
      "0001" when "01011000001011", -- t[5643] = 1
      "0001" when "01011000001100", -- t[5644] = 1
      "0001" when "01011000001101", -- t[5645] = 1
      "0001" when "01011000001110", -- t[5646] = 1
      "0001" when "01011000001111", -- t[5647] = 1
      "0001" when "01011000010000", -- t[5648] = 1
      "0001" when "01011000010001", -- t[5649] = 1
      "0001" when "01011000010010", -- t[5650] = 1
      "0001" when "01011000010011", -- t[5651] = 1
      "0001" when "01011000010100", -- t[5652] = 1
      "0001" when "01011000010101", -- t[5653] = 1
      "0001" when "01011000010110", -- t[5654] = 1
      "0001" when "01011000010111", -- t[5655] = 1
      "0001" when "01011000011000", -- t[5656] = 1
      "0001" when "01011000011001", -- t[5657] = 1
      "0001" when "01011000011010", -- t[5658] = 1
      "0001" when "01011000011011", -- t[5659] = 1
      "0001" when "01011000011100", -- t[5660] = 1
      "0001" when "01011000011101", -- t[5661] = 1
      "0001" when "01011000011110", -- t[5662] = 1
      "0001" when "01011000011111", -- t[5663] = 1
      "0001" when "01011000100000", -- t[5664] = 1
      "0001" when "01011000100001", -- t[5665] = 1
      "0001" when "01011000100010", -- t[5666] = 1
      "0001" when "01011000100011", -- t[5667] = 1
      "0001" when "01011000100100", -- t[5668] = 1
      "0001" when "01011000100101", -- t[5669] = 1
      "0001" when "01011000100110", -- t[5670] = 1
      "0001" when "01011000100111", -- t[5671] = 1
      "0001" when "01011000101000", -- t[5672] = 1
      "0001" when "01011000101001", -- t[5673] = 1
      "0001" when "01011000101010", -- t[5674] = 1
      "0001" when "01011000101011", -- t[5675] = 1
      "0001" when "01011000101100", -- t[5676] = 1
      "0001" when "01011000101101", -- t[5677] = 1
      "0001" when "01011000101110", -- t[5678] = 1
      "0001" when "01011000101111", -- t[5679] = 1
      "0001" when "01011000110000", -- t[5680] = 1
      "0001" when "01011000110001", -- t[5681] = 1
      "0001" when "01011000110010", -- t[5682] = 1
      "0001" when "01011000110011", -- t[5683] = 1
      "0001" when "01011000110100", -- t[5684] = 1
      "0001" when "01011000110101", -- t[5685] = 1
      "0001" when "01011000110110", -- t[5686] = 1
      "0001" when "01011000110111", -- t[5687] = 1
      "0001" when "01011000111000", -- t[5688] = 1
      "0001" when "01011000111001", -- t[5689] = 1
      "0001" when "01011000111010", -- t[5690] = 1
      "0001" when "01011000111011", -- t[5691] = 1
      "0001" when "01011000111100", -- t[5692] = 1
      "0001" when "01011000111101", -- t[5693] = 1
      "0001" when "01011000111110", -- t[5694] = 1
      "0001" when "01011000111111", -- t[5695] = 1
      "0001" when "01011001000000", -- t[5696] = 1
      "0001" when "01011001000001", -- t[5697] = 1
      "0001" when "01011001000010", -- t[5698] = 1
      "0001" when "01011001000011", -- t[5699] = 1
      "0001" when "01011001000100", -- t[5700] = 1
      "0001" when "01011001000101", -- t[5701] = 1
      "0001" when "01011001000110", -- t[5702] = 1
      "0001" when "01011001000111", -- t[5703] = 1
      "0001" when "01011001001000", -- t[5704] = 1
      "0001" when "01011001001001", -- t[5705] = 1
      "0001" when "01011001001010", -- t[5706] = 1
      "0001" when "01011001001011", -- t[5707] = 1
      "0001" when "01011001001100", -- t[5708] = 1
      "0001" when "01011001001101", -- t[5709] = 1
      "0001" when "01011001001110", -- t[5710] = 1
      "0001" when "01011001001111", -- t[5711] = 1
      "0001" when "01011001010000", -- t[5712] = 1
      "0001" when "01011001010001", -- t[5713] = 1
      "0001" when "01011001010010", -- t[5714] = 1
      "0001" when "01011001010011", -- t[5715] = 1
      "0001" when "01011001010100", -- t[5716] = 1
      "0001" when "01011001010101", -- t[5717] = 1
      "0001" when "01011001010110", -- t[5718] = 1
      "0001" when "01011001010111", -- t[5719] = 1
      "0001" when "01011001011000", -- t[5720] = 1
      "0001" when "01011001011001", -- t[5721] = 1
      "0001" when "01011001011010", -- t[5722] = 1
      "0001" when "01011001011011", -- t[5723] = 1
      "0001" when "01011001011100", -- t[5724] = 1
      "0001" when "01011001011101", -- t[5725] = 1
      "0001" when "01011001011110", -- t[5726] = 1
      "0001" when "01011001011111", -- t[5727] = 1
      "0001" when "01011001100000", -- t[5728] = 1
      "0001" when "01011001100001", -- t[5729] = 1
      "0001" when "01011001100010", -- t[5730] = 1
      "0001" when "01011001100011", -- t[5731] = 1
      "0001" when "01011001100100", -- t[5732] = 1
      "0001" when "01011001100101", -- t[5733] = 1
      "0001" when "01011001100110", -- t[5734] = 1
      "0001" when "01011001100111", -- t[5735] = 1
      "0001" when "01011001101000", -- t[5736] = 1
      "0001" when "01011001101001", -- t[5737] = 1
      "0001" when "01011001101010", -- t[5738] = 1
      "0001" when "01011001101011", -- t[5739] = 1
      "0001" when "01011001101100", -- t[5740] = 1
      "0001" when "01011001101101", -- t[5741] = 1
      "0001" when "01011001101110", -- t[5742] = 1
      "0001" when "01011001101111", -- t[5743] = 1
      "0001" when "01011001110000", -- t[5744] = 1
      "0001" when "01011001110001", -- t[5745] = 1
      "0001" when "01011001110010", -- t[5746] = 1
      "0001" when "01011001110011", -- t[5747] = 1
      "0001" when "01011001110100", -- t[5748] = 1
      "0001" when "01011001110101", -- t[5749] = 1
      "0001" when "01011001110110", -- t[5750] = 1
      "0001" when "01011001110111", -- t[5751] = 1
      "0001" when "01011001111000", -- t[5752] = 1
      "0001" when "01011001111001", -- t[5753] = 1
      "0001" when "01011001111010", -- t[5754] = 1
      "0001" when "01011001111011", -- t[5755] = 1
      "0001" when "01011001111100", -- t[5756] = 1
      "0001" when "01011001111101", -- t[5757] = 1
      "0001" when "01011001111110", -- t[5758] = 1
      "0001" when "01011001111111", -- t[5759] = 1
      "0001" when "01011010000000", -- t[5760] = 1
      "0001" when "01011010000001", -- t[5761] = 1
      "0001" when "01011010000010", -- t[5762] = 1
      "0001" when "01011010000011", -- t[5763] = 1
      "0001" when "01011010000100", -- t[5764] = 1
      "0001" when "01011010000101", -- t[5765] = 1
      "0001" when "01011010000110", -- t[5766] = 1
      "0001" when "01011010000111", -- t[5767] = 1
      "0001" when "01011010001000", -- t[5768] = 1
      "0001" when "01011010001001", -- t[5769] = 1
      "0001" when "01011010001010", -- t[5770] = 1
      "0001" when "01011010001011", -- t[5771] = 1
      "0001" when "01011010001100", -- t[5772] = 1
      "0001" when "01011010001101", -- t[5773] = 1
      "0001" when "01011010001110", -- t[5774] = 1
      "0001" when "01011010001111", -- t[5775] = 1
      "0001" when "01011010010000", -- t[5776] = 1
      "0001" when "01011010010001", -- t[5777] = 1
      "0001" when "01011010010010", -- t[5778] = 1
      "0001" when "01011010010011", -- t[5779] = 1
      "0001" when "01011010010100", -- t[5780] = 1
      "0001" when "01011010010101", -- t[5781] = 1
      "0001" when "01011010010110", -- t[5782] = 1
      "0001" when "01011010010111", -- t[5783] = 1
      "0001" when "01011010011000", -- t[5784] = 1
      "0001" when "01011010011001", -- t[5785] = 1
      "0001" when "01011010011010", -- t[5786] = 1
      "0001" when "01011010011011", -- t[5787] = 1
      "0001" when "01011010011100", -- t[5788] = 1
      "0001" when "01011010011101", -- t[5789] = 1
      "0001" when "01011010011110", -- t[5790] = 1
      "0001" when "01011010011111", -- t[5791] = 1
      "0001" when "01011010100000", -- t[5792] = 1
      "0001" when "01011010100001", -- t[5793] = 1
      "0001" when "01011010100010", -- t[5794] = 1
      "0001" when "01011010100011", -- t[5795] = 1
      "0001" when "01011010100100", -- t[5796] = 1
      "0001" when "01011010100101", -- t[5797] = 1
      "0001" when "01011010100110", -- t[5798] = 1
      "0001" when "01011010100111", -- t[5799] = 1
      "0001" when "01011010101000", -- t[5800] = 1
      "0001" when "01011010101001", -- t[5801] = 1
      "0001" when "01011010101010", -- t[5802] = 1
      "0001" when "01011010101011", -- t[5803] = 1
      "0001" when "01011010101100", -- t[5804] = 1
      "0001" when "01011010101101", -- t[5805] = 1
      "0001" when "01011010101110", -- t[5806] = 1
      "0001" when "01011010101111", -- t[5807] = 1
      "0001" when "01011010110000", -- t[5808] = 1
      "0001" when "01011010110001", -- t[5809] = 1
      "0001" when "01011010110010", -- t[5810] = 1
      "0001" when "01011010110011", -- t[5811] = 1
      "0001" when "01011010110100", -- t[5812] = 1
      "0001" when "01011010110101", -- t[5813] = 1
      "0001" when "01011010110110", -- t[5814] = 1
      "0001" when "01011010110111", -- t[5815] = 1
      "0001" when "01011010111000", -- t[5816] = 1
      "0001" when "01011010111001", -- t[5817] = 1
      "0001" when "01011010111010", -- t[5818] = 1
      "0001" when "01011010111011", -- t[5819] = 1
      "0001" when "01011010111100", -- t[5820] = 1
      "0001" when "01011010111101", -- t[5821] = 1
      "0001" when "01011010111110", -- t[5822] = 1
      "0001" when "01011010111111", -- t[5823] = 1
      "0001" when "01011011000000", -- t[5824] = 1
      "0001" when "01011011000001", -- t[5825] = 1
      "0001" when "01011011000010", -- t[5826] = 1
      "0001" when "01011011000011", -- t[5827] = 1
      "0001" when "01011011000100", -- t[5828] = 1
      "0001" when "01011011000101", -- t[5829] = 1
      "0001" when "01011011000110", -- t[5830] = 1
      "0001" when "01011011000111", -- t[5831] = 1
      "0001" when "01011011001000", -- t[5832] = 1
      "0001" when "01011011001001", -- t[5833] = 1
      "0001" when "01011011001010", -- t[5834] = 1
      "0001" when "01011011001011", -- t[5835] = 1
      "0001" when "01011011001100", -- t[5836] = 1
      "0001" when "01011011001101", -- t[5837] = 1
      "0001" when "01011011001110", -- t[5838] = 1
      "0001" when "01011011001111", -- t[5839] = 1
      "0001" when "01011011010000", -- t[5840] = 1
      "0001" when "01011011010001", -- t[5841] = 1
      "0001" when "01011011010010", -- t[5842] = 1
      "0001" when "01011011010011", -- t[5843] = 1
      "0001" when "01011011010100", -- t[5844] = 1
      "0001" when "01011011010101", -- t[5845] = 1
      "0001" when "01011011010110", -- t[5846] = 1
      "0001" when "01011011010111", -- t[5847] = 1
      "0001" when "01011011011000", -- t[5848] = 1
      "0001" when "01011011011001", -- t[5849] = 1
      "0001" when "01011011011010", -- t[5850] = 1
      "0001" when "01011011011011", -- t[5851] = 1
      "0001" when "01011011011100", -- t[5852] = 1
      "0001" when "01011011011101", -- t[5853] = 1
      "0001" when "01011011011110", -- t[5854] = 1
      "0001" when "01011011011111", -- t[5855] = 1
      "0001" when "01011011100000", -- t[5856] = 1
      "0001" when "01011011100001", -- t[5857] = 1
      "0001" when "01011011100010", -- t[5858] = 1
      "0001" when "01011011100011", -- t[5859] = 1
      "0001" when "01011011100100", -- t[5860] = 1
      "0001" when "01011011100101", -- t[5861] = 1
      "0001" when "01011011100110", -- t[5862] = 1
      "0001" when "01011011100111", -- t[5863] = 1
      "0001" when "01011011101000", -- t[5864] = 1
      "0001" when "01011011101001", -- t[5865] = 1
      "0001" when "01011011101010", -- t[5866] = 1
      "0001" when "01011011101011", -- t[5867] = 1
      "0001" when "01011011101100", -- t[5868] = 1
      "0001" when "01011011101101", -- t[5869] = 1
      "0001" when "01011011101110", -- t[5870] = 1
      "0001" when "01011011101111", -- t[5871] = 1
      "0001" when "01011011110000", -- t[5872] = 1
      "0001" when "01011011110001", -- t[5873] = 1
      "0001" when "01011011110010", -- t[5874] = 1
      "0001" when "01011011110011", -- t[5875] = 1
      "0001" when "01011011110100", -- t[5876] = 1
      "0001" when "01011011110101", -- t[5877] = 1
      "0001" when "01011011110110", -- t[5878] = 1
      "0001" when "01011011110111", -- t[5879] = 1
      "0001" when "01011011111000", -- t[5880] = 1
      "0001" when "01011011111001", -- t[5881] = 1
      "0001" when "01011011111010", -- t[5882] = 1
      "0001" when "01011011111011", -- t[5883] = 1
      "0001" when "01011011111100", -- t[5884] = 1
      "0001" when "01011011111101", -- t[5885] = 1
      "0001" when "01011011111110", -- t[5886] = 1
      "0001" when "01011011111111", -- t[5887] = 1
      "0001" when "01011100000000", -- t[5888] = 1
      "0001" when "01011100000001", -- t[5889] = 1
      "0001" when "01011100000010", -- t[5890] = 1
      "0001" when "01011100000011", -- t[5891] = 1
      "0001" when "01011100000100", -- t[5892] = 1
      "0001" when "01011100000101", -- t[5893] = 1
      "0001" when "01011100000110", -- t[5894] = 1
      "0001" when "01011100000111", -- t[5895] = 1
      "0001" when "01011100001000", -- t[5896] = 1
      "0001" when "01011100001001", -- t[5897] = 1
      "0001" when "01011100001010", -- t[5898] = 1
      "0001" when "01011100001011", -- t[5899] = 1
      "0001" when "01011100001100", -- t[5900] = 1
      "0001" when "01011100001101", -- t[5901] = 1
      "0001" when "01011100001110", -- t[5902] = 1
      "0001" when "01011100001111", -- t[5903] = 1
      "0001" when "01011100010000", -- t[5904] = 1
      "0001" when "01011100010001", -- t[5905] = 1
      "0001" when "01011100010010", -- t[5906] = 1
      "0001" when "01011100010011", -- t[5907] = 1
      "0001" when "01011100010100", -- t[5908] = 1
      "0001" when "01011100010101", -- t[5909] = 1
      "0001" when "01011100010110", -- t[5910] = 1
      "0001" when "01011100010111", -- t[5911] = 1
      "0001" when "01011100011000", -- t[5912] = 1
      "0001" when "01011100011001", -- t[5913] = 1
      "0001" when "01011100011010", -- t[5914] = 1
      "0001" when "01011100011011", -- t[5915] = 1
      "0001" when "01011100011100", -- t[5916] = 1
      "0001" when "01011100011101", -- t[5917] = 1
      "0001" when "01011100011110", -- t[5918] = 1
      "0001" when "01011100011111", -- t[5919] = 1
      "0001" when "01011100100000", -- t[5920] = 1
      "0001" when "01011100100001", -- t[5921] = 1
      "0001" when "01011100100010", -- t[5922] = 1
      "0001" when "01011100100011", -- t[5923] = 1
      "0001" when "01011100100100", -- t[5924] = 1
      "0001" when "01011100100101", -- t[5925] = 1
      "0001" when "01011100100110", -- t[5926] = 1
      "0001" when "01011100100111", -- t[5927] = 1
      "0001" when "01011100101000", -- t[5928] = 1
      "0001" when "01011100101001", -- t[5929] = 1
      "0001" when "01011100101010", -- t[5930] = 1
      "0001" when "01011100101011", -- t[5931] = 1
      "0001" when "01011100101100", -- t[5932] = 1
      "0001" when "01011100101101", -- t[5933] = 1
      "0001" when "01011100101110", -- t[5934] = 1
      "0001" when "01011100101111", -- t[5935] = 1
      "0001" when "01011100110000", -- t[5936] = 1
      "0001" when "01011100110001", -- t[5937] = 1
      "0001" when "01011100110010", -- t[5938] = 1
      "0001" when "01011100110011", -- t[5939] = 1
      "0001" when "01011100110100", -- t[5940] = 1
      "0001" when "01011100110101", -- t[5941] = 1
      "0001" when "01011100110110", -- t[5942] = 1
      "0001" when "01011100110111", -- t[5943] = 1
      "0001" when "01011100111000", -- t[5944] = 1
      "0001" when "01011100111001", -- t[5945] = 1
      "0001" when "01011100111010", -- t[5946] = 1
      "0001" when "01011100111011", -- t[5947] = 1
      "0001" when "01011100111100", -- t[5948] = 1
      "0001" when "01011100111101", -- t[5949] = 1
      "0001" when "01011100111110", -- t[5950] = 1
      "0001" when "01011100111111", -- t[5951] = 1
      "0001" when "01011101000000", -- t[5952] = 1
      "0001" when "01011101000001", -- t[5953] = 1
      "0001" when "01011101000010", -- t[5954] = 1
      "0001" when "01011101000011", -- t[5955] = 1
      "0001" when "01011101000100", -- t[5956] = 1
      "0001" when "01011101000101", -- t[5957] = 1
      "0001" when "01011101000110", -- t[5958] = 1
      "0001" when "01011101000111", -- t[5959] = 1
      "0001" when "01011101001000", -- t[5960] = 1
      "0001" when "01011101001001", -- t[5961] = 1
      "0001" when "01011101001010", -- t[5962] = 1
      "0001" when "01011101001011", -- t[5963] = 1
      "0001" when "01011101001100", -- t[5964] = 1
      "0001" when "01011101001101", -- t[5965] = 1
      "0001" when "01011101001110", -- t[5966] = 1
      "0001" when "01011101001111", -- t[5967] = 1
      "0001" when "01011101010000", -- t[5968] = 1
      "0001" when "01011101010001", -- t[5969] = 1
      "0001" when "01011101010010", -- t[5970] = 1
      "0001" when "01011101010011", -- t[5971] = 1
      "0001" when "01011101010100", -- t[5972] = 1
      "0001" when "01011101010101", -- t[5973] = 1
      "0001" when "01011101010110", -- t[5974] = 1
      "0001" when "01011101010111", -- t[5975] = 1
      "0001" when "01011101011000", -- t[5976] = 1
      "0001" when "01011101011001", -- t[5977] = 1
      "0001" when "01011101011010", -- t[5978] = 1
      "0001" when "01011101011011", -- t[5979] = 1
      "0001" when "01011101011100", -- t[5980] = 1
      "0001" when "01011101011101", -- t[5981] = 1
      "0001" when "01011101011110", -- t[5982] = 1
      "0001" when "01011101011111", -- t[5983] = 1
      "0001" when "01011101100000", -- t[5984] = 1
      "0001" when "01011101100001", -- t[5985] = 1
      "0001" when "01011101100010", -- t[5986] = 1
      "0001" when "01011101100011", -- t[5987] = 1
      "0001" when "01011101100100", -- t[5988] = 1
      "0001" when "01011101100101", -- t[5989] = 1
      "0001" when "01011101100110", -- t[5990] = 1
      "0001" when "01011101100111", -- t[5991] = 1
      "0001" when "01011101101000", -- t[5992] = 1
      "0001" when "01011101101001", -- t[5993] = 1
      "0001" when "01011101101010", -- t[5994] = 1
      "0001" when "01011101101011", -- t[5995] = 1
      "0001" when "01011101101100", -- t[5996] = 1
      "0001" when "01011101101101", -- t[5997] = 1
      "0001" when "01011101101110", -- t[5998] = 1
      "0001" when "01011101101111", -- t[5999] = 1
      "0001" when "01011101110000", -- t[6000] = 1
      "0001" when "01011101110001", -- t[6001] = 1
      "0001" when "01011101110010", -- t[6002] = 1
      "0001" when "01011101110011", -- t[6003] = 1
      "0001" when "01011101110100", -- t[6004] = 1
      "0001" when "01011101110101", -- t[6005] = 1
      "0001" when "01011101110110", -- t[6006] = 1
      "0001" when "01011101110111", -- t[6007] = 1
      "0001" when "01011101111000", -- t[6008] = 1
      "0001" when "01011101111001", -- t[6009] = 1
      "0001" when "01011101111010", -- t[6010] = 1
      "0001" when "01011101111011", -- t[6011] = 1
      "0001" when "01011101111100", -- t[6012] = 1
      "0001" when "01011101111101", -- t[6013] = 1
      "0001" when "01011101111110", -- t[6014] = 1
      "0001" when "01011101111111", -- t[6015] = 1
      "0001" when "01011110000000", -- t[6016] = 1
      "0001" when "01011110000001", -- t[6017] = 1
      "0001" when "01011110000010", -- t[6018] = 1
      "0001" when "01011110000011", -- t[6019] = 1
      "0001" when "01011110000100", -- t[6020] = 1
      "0001" when "01011110000101", -- t[6021] = 1
      "0001" when "01011110000110", -- t[6022] = 1
      "0001" when "01011110000111", -- t[6023] = 1
      "0001" when "01011110001000", -- t[6024] = 1
      "0001" when "01011110001001", -- t[6025] = 1
      "0001" when "01011110001010", -- t[6026] = 1
      "0001" when "01011110001011", -- t[6027] = 1
      "0001" when "01011110001100", -- t[6028] = 1
      "0001" when "01011110001101", -- t[6029] = 1
      "0001" when "01011110001110", -- t[6030] = 1
      "0001" when "01011110001111", -- t[6031] = 1
      "0001" when "01011110010000", -- t[6032] = 1
      "0001" when "01011110010001", -- t[6033] = 1
      "0001" when "01011110010010", -- t[6034] = 1
      "0001" when "01011110010011", -- t[6035] = 1
      "0001" when "01011110010100", -- t[6036] = 1
      "0001" when "01011110010101", -- t[6037] = 1
      "0001" when "01011110010110", -- t[6038] = 1
      "0001" when "01011110010111", -- t[6039] = 1
      "0001" when "01011110011000", -- t[6040] = 1
      "0001" when "01011110011001", -- t[6041] = 1
      "0001" when "01011110011010", -- t[6042] = 1
      "0001" when "01011110011011", -- t[6043] = 1
      "0001" when "01011110011100", -- t[6044] = 1
      "0001" when "01011110011101", -- t[6045] = 1
      "0001" when "01011110011110", -- t[6046] = 1
      "0001" when "01011110011111", -- t[6047] = 1
      "0001" when "01011110100000", -- t[6048] = 1
      "0001" when "01011110100001", -- t[6049] = 1
      "0001" when "01011110100010", -- t[6050] = 1
      "0001" when "01011110100011", -- t[6051] = 1
      "0001" when "01011110100100", -- t[6052] = 1
      "0001" when "01011110100101", -- t[6053] = 1
      "0001" when "01011110100110", -- t[6054] = 1
      "0001" when "01011110100111", -- t[6055] = 1
      "0001" when "01011110101000", -- t[6056] = 1
      "0001" when "01011110101001", -- t[6057] = 1
      "0001" when "01011110101010", -- t[6058] = 1
      "0001" when "01011110101011", -- t[6059] = 1
      "0001" when "01011110101100", -- t[6060] = 1
      "0001" when "01011110101101", -- t[6061] = 1
      "0001" when "01011110101110", -- t[6062] = 1
      "0001" when "01011110101111", -- t[6063] = 1
      "0001" when "01011110110000", -- t[6064] = 1
      "0001" when "01011110110001", -- t[6065] = 1
      "0001" when "01011110110010", -- t[6066] = 1
      "0001" when "01011110110011", -- t[6067] = 1
      "0001" when "01011110110100", -- t[6068] = 1
      "0001" when "01011110110101", -- t[6069] = 1
      "0001" when "01011110110110", -- t[6070] = 1
      "0001" when "01011110110111", -- t[6071] = 1
      "0001" when "01011110111000", -- t[6072] = 1
      "0001" when "01011110111001", -- t[6073] = 1
      "0001" when "01011110111010", -- t[6074] = 1
      "0001" when "01011110111011", -- t[6075] = 1
      "0001" when "01011110111100", -- t[6076] = 1
      "0001" when "01011110111101", -- t[6077] = 1
      "0001" when "01011110111110", -- t[6078] = 1
      "0001" when "01011110111111", -- t[6079] = 1
      "0001" when "01011111000000", -- t[6080] = 1
      "0001" when "01011111000001", -- t[6081] = 1
      "0001" when "01011111000010", -- t[6082] = 1
      "0001" when "01011111000011", -- t[6083] = 1
      "0001" when "01011111000100", -- t[6084] = 1
      "0001" when "01011111000101", -- t[6085] = 1
      "0001" when "01011111000110", -- t[6086] = 1
      "0001" when "01011111000111", -- t[6087] = 1
      "0001" when "01011111001000", -- t[6088] = 1
      "0001" when "01011111001001", -- t[6089] = 1
      "0001" when "01011111001010", -- t[6090] = 1
      "0001" when "01011111001011", -- t[6091] = 1
      "0001" when "01011111001100", -- t[6092] = 1
      "0001" when "01011111001101", -- t[6093] = 1
      "0001" when "01011111001110", -- t[6094] = 1
      "0001" when "01011111001111", -- t[6095] = 1
      "0001" when "01011111010000", -- t[6096] = 1
      "0001" when "01011111010001", -- t[6097] = 1
      "0001" when "01011111010010", -- t[6098] = 1
      "0001" when "01011111010011", -- t[6099] = 1
      "0001" when "01011111010100", -- t[6100] = 1
      "0001" when "01011111010101", -- t[6101] = 1
      "0001" when "01011111010110", -- t[6102] = 1
      "0001" when "01011111010111", -- t[6103] = 1
      "0001" when "01011111011000", -- t[6104] = 1
      "0001" when "01011111011001", -- t[6105] = 1
      "0001" when "01011111011010", -- t[6106] = 1
      "0001" when "01011111011011", -- t[6107] = 1
      "0001" when "01011111011100", -- t[6108] = 1
      "0001" when "01011111011101", -- t[6109] = 1
      "0001" when "01011111011110", -- t[6110] = 1
      "0001" when "01011111011111", -- t[6111] = 1
      "0001" when "01011111100000", -- t[6112] = 1
      "0001" when "01011111100001", -- t[6113] = 1
      "0001" when "01011111100010", -- t[6114] = 1
      "0001" when "01011111100011", -- t[6115] = 1
      "0001" when "01011111100100", -- t[6116] = 1
      "0001" when "01011111100101", -- t[6117] = 1
      "0001" when "01011111100110", -- t[6118] = 1
      "0001" when "01011111100111", -- t[6119] = 1
      "0001" when "01011111101000", -- t[6120] = 1
      "0001" when "01011111101001", -- t[6121] = 1
      "0001" when "01011111101010", -- t[6122] = 1
      "0001" when "01011111101011", -- t[6123] = 1
      "0001" when "01011111101100", -- t[6124] = 1
      "0001" when "01011111101101", -- t[6125] = 1
      "0001" when "01011111101110", -- t[6126] = 1
      "0001" when "01011111101111", -- t[6127] = 1
      "0001" when "01011111110000", -- t[6128] = 1
      "0001" when "01011111110001", -- t[6129] = 1
      "0001" when "01011111110010", -- t[6130] = 1
      "0001" when "01011111110011", -- t[6131] = 1
      "0001" when "01011111110100", -- t[6132] = 1
      "0001" when "01011111110101", -- t[6133] = 1
      "0001" when "01011111110110", -- t[6134] = 1
      "0001" when "01011111110111", -- t[6135] = 1
      "0001" when "01011111111000", -- t[6136] = 1
      "0001" when "01011111111001", -- t[6137] = 1
      "0001" when "01011111111010", -- t[6138] = 1
      "0001" when "01011111111011", -- t[6139] = 1
      "0001" when "01011111111100", -- t[6140] = 1
      "0001" when "01011111111101", -- t[6141] = 1
      "0001" when "01011111111110", -- t[6142] = 1
      "0001" when "01011111111111", -- t[6143] = 1
      "0001" when "01100000000000", -- t[6144] = 1
      "0001" when "01100000000001", -- t[6145] = 1
      "0001" when "01100000000010", -- t[6146] = 1
      "0001" when "01100000000011", -- t[6147] = 1
      "0001" when "01100000000100", -- t[6148] = 1
      "0001" when "01100000000101", -- t[6149] = 1
      "0001" when "01100000000110", -- t[6150] = 1
      "0001" when "01100000000111", -- t[6151] = 1
      "0001" when "01100000001000", -- t[6152] = 1
      "0001" when "01100000001001", -- t[6153] = 1
      "0001" when "01100000001010", -- t[6154] = 1
      "0001" when "01100000001011", -- t[6155] = 1
      "0001" when "01100000001100", -- t[6156] = 1
      "0001" when "01100000001101", -- t[6157] = 1
      "0001" when "01100000001110", -- t[6158] = 1
      "0001" when "01100000001111", -- t[6159] = 1
      "0001" when "01100000010000", -- t[6160] = 1
      "0001" when "01100000010001", -- t[6161] = 1
      "0001" when "01100000010010", -- t[6162] = 1
      "0001" when "01100000010011", -- t[6163] = 1
      "0001" when "01100000010100", -- t[6164] = 1
      "0001" when "01100000010101", -- t[6165] = 1
      "0001" when "01100000010110", -- t[6166] = 1
      "0001" when "01100000010111", -- t[6167] = 1
      "0001" when "01100000011000", -- t[6168] = 1
      "0001" when "01100000011001", -- t[6169] = 1
      "0001" when "01100000011010", -- t[6170] = 1
      "0001" when "01100000011011", -- t[6171] = 1
      "0001" when "01100000011100", -- t[6172] = 1
      "0001" when "01100000011101", -- t[6173] = 1
      "0001" when "01100000011110", -- t[6174] = 1
      "0001" when "01100000011111", -- t[6175] = 1
      "0001" when "01100000100000", -- t[6176] = 1
      "0001" when "01100000100001", -- t[6177] = 1
      "0001" when "01100000100010", -- t[6178] = 1
      "0001" when "01100000100011", -- t[6179] = 1
      "0001" when "01100000100100", -- t[6180] = 1
      "0001" when "01100000100101", -- t[6181] = 1
      "0001" when "01100000100110", -- t[6182] = 1
      "0001" when "01100000100111", -- t[6183] = 1
      "0001" when "01100000101000", -- t[6184] = 1
      "0001" when "01100000101001", -- t[6185] = 1
      "0001" when "01100000101010", -- t[6186] = 1
      "0001" when "01100000101011", -- t[6187] = 1
      "0001" when "01100000101100", -- t[6188] = 1
      "0001" when "01100000101101", -- t[6189] = 1
      "0001" when "01100000101110", -- t[6190] = 1
      "0001" when "01100000101111", -- t[6191] = 1
      "0001" when "01100000110000", -- t[6192] = 1
      "0001" when "01100000110001", -- t[6193] = 1
      "0001" when "01100000110010", -- t[6194] = 1
      "0001" when "01100000110011", -- t[6195] = 1
      "0001" when "01100000110100", -- t[6196] = 1
      "0001" when "01100000110101", -- t[6197] = 1
      "0001" when "01100000110110", -- t[6198] = 1
      "0001" when "01100000110111", -- t[6199] = 1
      "0001" when "01100000111000", -- t[6200] = 1
      "0010" when "01100000111001", -- t[6201] = 2
      "0010" when "01100000111010", -- t[6202] = 2
      "0010" when "01100000111011", -- t[6203] = 2
      "0010" when "01100000111100", -- t[6204] = 2
      "0010" when "01100000111101", -- t[6205] = 2
      "0010" when "01100000111110", -- t[6206] = 2
      "0010" when "01100000111111", -- t[6207] = 2
      "0010" when "01100001000000", -- t[6208] = 2
      "0010" when "01100001000001", -- t[6209] = 2
      "0010" when "01100001000010", -- t[6210] = 2
      "0010" when "01100001000011", -- t[6211] = 2
      "0010" when "01100001000100", -- t[6212] = 2
      "0010" when "01100001000101", -- t[6213] = 2
      "0010" when "01100001000110", -- t[6214] = 2
      "0010" when "01100001000111", -- t[6215] = 2
      "0010" when "01100001001000", -- t[6216] = 2
      "0010" when "01100001001001", -- t[6217] = 2
      "0010" when "01100001001010", -- t[6218] = 2
      "0010" when "01100001001011", -- t[6219] = 2
      "0010" when "01100001001100", -- t[6220] = 2
      "0010" when "01100001001101", -- t[6221] = 2
      "0010" when "01100001001110", -- t[6222] = 2
      "0010" when "01100001001111", -- t[6223] = 2
      "0010" when "01100001010000", -- t[6224] = 2
      "0010" when "01100001010001", -- t[6225] = 2
      "0010" when "01100001010010", -- t[6226] = 2
      "0010" when "01100001010011", -- t[6227] = 2
      "0010" when "01100001010100", -- t[6228] = 2
      "0010" when "01100001010101", -- t[6229] = 2
      "0010" when "01100001010110", -- t[6230] = 2
      "0010" when "01100001010111", -- t[6231] = 2
      "0010" when "01100001011000", -- t[6232] = 2
      "0010" when "01100001011001", -- t[6233] = 2
      "0010" when "01100001011010", -- t[6234] = 2
      "0010" when "01100001011011", -- t[6235] = 2
      "0010" when "01100001011100", -- t[6236] = 2
      "0010" when "01100001011101", -- t[6237] = 2
      "0010" when "01100001011110", -- t[6238] = 2
      "0010" when "01100001011111", -- t[6239] = 2
      "0010" when "01100001100000", -- t[6240] = 2
      "0010" when "01100001100001", -- t[6241] = 2
      "0010" when "01100001100010", -- t[6242] = 2
      "0010" when "01100001100011", -- t[6243] = 2
      "0010" when "01100001100100", -- t[6244] = 2
      "0010" when "01100001100101", -- t[6245] = 2
      "0010" when "01100001100110", -- t[6246] = 2
      "0010" when "01100001100111", -- t[6247] = 2
      "0010" when "01100001101000", -- t[6248] = 2
      "0010" when "01100001101001", -- t[6249] = 2
      "0010" when "01100001101010", -- t[6250] = 2
      "0010" when "01100001101011", -- t[6251] = 2
      "0010" when "01100001101100", -- t[6252] = 2
      "0010" when "01100001101101", -- t[6253] = 2
      "0010" when "01100001101110", -- t[6254] = 2
      "0010" when "01100001101111", -- t[6255] = 2
      "0010" when "01100001110000", -- t[6256] = 2
      "0010" when "01100001110001", -- t[6257] = 2
      "0010" when "01100001110010", -- t[6258] = 2
      "0010" when "01100001110011", -- t[6259] = 2
      "0010" when "01100001110100", -- t[6260] = 2
      "0010" when "01100001110101", -- t[6261] = 2
      "0010" when "01100001110110", -- t[6262] = 2
      "0010" when "01100001110111", -- t[6263] = 2
      "0010" when "01100001111000", -- t[6264] = 2
      "0010" when "01100001111001", -- t[6265] = 2
      "0010" when "01100001111010", -- t[6266] = 2
      "0010" when "01100001111011", -- t[6267] = 2
      "0010" when "01100001111100", -- t[6268] = 2
      "0010" when "01100001111101", -- t[6269] = 2
      "0010" when "01100001111110", -- t[6270] = 2
      "0010" when "01100001111111", -- t[6271] = 2
      "0010" when "01100010000000", -- t[6272] = 2
      "0010" when "01100010000001", -- t[6273] = 2
      "0010" when "01100010000010", -- t[6274] = 2
      "0010" when "01100010000011", -- t[6275] = 2
      "0010" when "01100010000100", -- t[6276] = 2
      "0010" when "01100010000101", -- t[6277] = 2
      "0010" when "01100010000110", -- t[6278] = 2
      "0010" when "01100010000111", -- t[6279] = 2
      "0010" when "01100010001000", -- t[6280] = 2
      "0010" when "01100010001001", -- t[6281] = 2
      "0010" when "01100010001010", -- t[6282] = 2
      "0010" when "01100010001011", -- t[6283] = 2
      "0010" when "01100010001100", -- t[6284] = 2
      "0010" when "01100010001101", -- t[6285] = 2
      "0010" when "01100010001110", -- t[6286] = 2
      "0010" when "01100010001111", -- t[6287] = 2
      "0010" when "01100010010000", -- t[6288] = 2
      "0010" when "01100010010001", -- t[6289] = 2
      "0010" when "01100010010010", -- t[6290] = 2
      "0010" when "01100010010011", -- t[6291] = 2
      "0010" when "01100010010100", -- t[6292] = 2
      "0010" when "01100010010101", -- t[6293] = 2
      "0010" when "01100010010110", -- t[6294] = 2
      "0010" when "01100010010111", -- t[6295] = 2
      "0010" when "01100010011000", -- t[6296] = 2
      "0010" when "01100010011001", -- t[6297] = 2
      "0010" when "01100010011010", -- t[6298] = 2
      "0010" when "01100010011011", -- t[6299] = 2
      "0010" when "01100010011100", -- t[6300] = 2
      "0010" when "01100010011101", -- t[6301] = 2
      "0010" when "01100010011110", -- t[6302] = 2
      "0010" when "01100010011111", -- t[6303] = 2
      "0010" when "01100010100000", -- t[6304] = 2
      "0010" when "01100010100001", -- t[6305] = 2
      "0010" when "01100010100010", -- t[6306] = 2
      "0010" when "01100010100011", -- t[6307] = 2
      "0010" when "01100010100100", -- t[6308] = 2
      "0010" when "01100010100101", -- t[6309] = 2
      "0010" when "01100010100110", -- t[6310] = 2
      "0010" when "01100010100111", -- t[6311] = 2
      "0010" when "01100010101000", -- t[6312] = 2
      "0010" when "01100010101001", -- t[6313] = 2
      "0010" when "01100010101010", -- t[6314] = 2
      "0010" when "01100010101011", -- t[6315] = 2
      "0010" when "01100010101100", -- t[6316] = 2
      "0010" when "01100010101101", -- t[6317] = 2
      "0010" when "01100010101110", -- t[6318] = 2
      "0010" when "01100010101111", -- t[6319] = 2
      "0010" when "01100010110000", -- t[6320] = 2
      "0010" when "01100010110001", -- t[6321] = 2
      "0010" when "01100010110010", -- t[6322] = 2
      "0010" when "01100010110011", -- t[6323] = 2
      "0010" when "01100010110100", -- t[6324] = 2
      "0010" when "01100010110101", -- t[6325] = 2
      "0010" when "01100010110110", -- t[6326] = 2
      "0010" when "01100010110111", -- t[6327] = 2
      "0010" when "01100010111000", -- t[6328] = 2
      "0010" when "01100010111001", -- t[6329] = 2
      "0010" when "01100010111010", -- t[6330] = 2
      "0010" when "01100010111011", -- t[6331] = 2
      "0010" when "01100010111100", -- t[6332] = 2
      "0010" when "01100010111101", -- t[6333] = 2
      "0010" when "01100010111110", -- t[6334] = 2
      "0010" when "01100010111111", -- t[6335] = 2
      "0010" when "01100011000000", -- t[6336] = 2
      "0010" when "01100011000001", -- t[6337] = 2
      "0010" when "01100011000010", -- t[6338] = 2
      "0010" when "01100011000011", -- t[6339] = 2
      "0010" when "01100011000100", -- t[6340] = 2
      "0010" when "01100011000101", -- t[6341] = 2
      "0010" when "01100011000110", -- t[6342] = 2
      "0010" when "01100011000111", -- t[6343] = 2
      "0010" when "01100011001000", -- t[6344] = 2
      "0010" when "01100011001001", -- t[6345] = 2
      "0010" when "01100011001010", -- t[6346] = 2
      "0010" when "01100011001011", -- t[6347] = 2
      "0010" when "01100011001100", -- t[6348] = 2
      "0010" when "01100011001101", -- t[6349] = 2
      "0010" when "01100011001110", -- t[6350] = 2
      "0010" when "01100011001111", -- t[6351] = 2
      "0010" when "01100011010000", -- t[6352] = 2
      "0010" when "01100011010001", -- t[6353] = 2
      "0010" when "01100011010010", -- t[6354] = 2
      "0010" when "01100011010011", -- t[6355] = 2
      "0010" when "01100011010100", -- t[6356] = 2
      "0010" when "01100011010101", -- t[6357] = 2
      "0010" when "01100011010110", -- t[6358] = 2
      "0010" when "01100011010111", -- t[6359] = 2
      "0010" when "01100011011000", -- t[6360] = 2
      "0010" when "01100011011001", -- t[6361] = 2
      "0010" when "01100011011010", -- t[6362] = 2
      "0010" when "01100011011011", -- t[6363] = 2
      "0010" when "01100011011100", -- t[6364] = 2
      "0010" when "01100011011101", -- t[6365] = 2
      "0010" when "01100011011110", -- t[6366] = 2
      "0010" when "01100011011111", -- t[6367] = 2
      "0010" when "01100011100000", -- t[6368] = 2
      "0010" when "01100011100001", -- t[6369] = 2
      "0010" when "01100011100010", -- t[6370] = 2
      "0010" when "01100011100011", -- t[6371] = 2
      "0010" when "01100011100100", -- t[6372] = 2
      "0010" when "01100011100101", -- t[6373] = 2
      "0010" when "01100011100110", -- t[6374] = 2
      "0010" when "01100011100111", -- t[6375] = 2
      "0010" when "01100011101000", -- t[6376] = 2
      "0010" when "01100011101001", -- t[6377] = 2
      "0010" when "01100011101010", -- t[6378] = 2
      "0010" when "01100011101011", -- t[6379] = 2
      "0010" when "01100011101100", -- t[6380] = 2
      "0010" when "01100011101101", -- t[6381] = 2
      "0010" when "01100011101110", -- t[6382] = 2
      "0010" when "01100011101111", -- t[6383] = 2
      "0010" when "01100011110000", -- t[6384] = 2
      "0010" when "01100011110001", -- t[6385] = 2
      "0010" when "01100011110010", -- t[6386] = 2
      "0010" when "01100011110011", -- t[6387] = 2
      "0010" when "01100011110100", -- t[6388] = 2
      "0010" when "01100011110101", -- t[6389] = 2
      "0010" when "01100011110110", -- t[6390] = 2
      "0010" when "01100011110111", -- t[6391] = 2
      "0010" when "01100011111000", -- t[6392] = 2
      "0010" when "01100011111001", -- t[6393] = 2
      "0010" when "01100011111010", -- t[6394] = 2
      "0010" when "01100011111011", -- t[6395] = 2
      "0010" when "01100011111100", -- t[6396] = 2
      "0010" when "01100011111101", -- t[6397] = 2
      "0010" when "01100011111110", -- t[6398] = 2
      "0010" when "01100011111111", -- t[6399] = 2
      "0010" when "01100100000000", -- t[6400] = 2
      "0010" when "01100100000001", -- t[6401] = 2
      "0010" when "01100100000010", -- t[6402] = 2
      "0010" when "01100100000011", -- t[6403] = 2
      "0010" when "01100100000100", -- t[6404] = 2
      "0010" when "01100100000101", -- t[6405] = 2
      "0010" when "01100100000110", -- t[6406] = 2
      "0010" when "01100100000111", -- t[6407] = 2
      "0010" when "01100100001000", -- t[6408] = 2
      "0010" when "01100100001001", -- t[6409] = 2
      "0010" when "01100100001010", -- t[6410] = 2
      "0010" when "01100100001011", -- t[6411] = 2
      "0010" when "01100100001100", -- t[6412] = 2
      "0010" when "01100100001101", -- t[6413] = 2
      "0010" when "01100100001110", -- t[6414] = 2
      "0010" when "01100100001111", -- t[6415] = 2
      "0010" when "01100100010000", -- t[6416] = 2
      "0010" when "01100100010001", -- t[6417] = 2
      "0010" when "01100100010010", -- t[6418] = 2
      "0010" when "01100100010011", -- t[6419] = 2
      "0010" when "01100100010100", -- t[6420] = 2
      "0010" when "01100100010101", -- t[6421] = 2
      "0010" when "01100100010110", -- t[6422] = 2
      "0010" when "01100100010111", -- t[6423] = 2
      "0010" when "01100100011000", -- t[6424] = 2
      "0010" when "01100100011001", -- t[6425] = 2
      "0010" when "01100100011010", -- t[6426] = 2
      "0010" when "01100100011011", -- t[6427] = 2
      "0010" when "01100100011100", -- t[6428] = 2
      "0010" when "01100100011101", -- t[6429] = 2
      "0010" when "01100100011110", -- t[6430] = 2
      "0010" when "01100100011111", -- t[6431] = 2
      "0010" when "01100100100000", -- t[6432] = 2
      "0010" when "01100100100001", -- t[6433] = 2
      "0010" when "01100100100010", -- t[6434] = 2
      "0010" when "01100100100011", -- t[6435] = 2
      "0010" when "01100100100100", -- t[6436] = 2
      "0010" when "01100100100101", -- t[6437] = 2
      "0010" when "01100100100110", -- t[6438] = 2
      "0010" when "01100100100111", -- t[6439] = 2
      "0010" when "01100100101000", -- t[6440] = 2
      "0010" when "01100100101001", -- t[6441] = 2
      "0010" when "01100100101010", -- t[6442] = 2
      "0010" when "01100100101011", -- t[6443] = 2
      "0010" when "01100100101100", -- t[6444] = 2
      "0010" when "01100100101101", -- t[6445] = 2
      "0010" when "01100100101110", -- t[6446] = 2
      "0010" when "01100100101111", -- t[6447] = 2
      "0010" when "01100100110000", -- t[6448] = 2
      "0010" when "01100100110001", -- t[6449] = 2
      "0010" when "01100100110010", -- t[6450] = 2
      "0010" when "01100100110011", -- t[6451] = 2
      "0010" when "01100100110100", -- t[6452] = 2
      "0010" when "01100100110101", -- t[6453] = 2
      "0010" when "01100100110110", -- t[6454] = 2
      "0010" when "01100100110111", -- t[6455] = 2
      "0010" when "01100100111000", -- t[6456] = 2
      "0010" when "01100100111001", -- t[6457] = 2
      "0010" when "01100100111010", -- t[6458] = 2
      "0010" when "01100100111011", -- t[6459] = 2
      "0010" when "01100100111100", -- t[6460] = 2
      "0010" when "01100100111101", -- t[6461] = 2
      "0010" when "01100100111110", -- t[6462] = 2
      "0010" when "01100100111111", -- t[6463] = 2
      "0010" when "01100101000000", -- t[6464] = 2
      "0010" when "01100101000001", -- t[6465] = 2
      "0010" when "01100101000010", -- t[6466] = 2
      "0010" when "01100101000011", -- t[6467] = 2
      "0010" when "01100101000100", -- t[6468] = 2
      "0010" when "01100101000101", -- t[6469] = 2
      "0010" when "01100101000110", -- t[6470] = 2
      "0010" when "01100101000111", -- t[6471] = 2
      "0010" when "01100101001000", -- t[6472] = 2
      "0010" when "01100101001001", -- t[6473] = 2
      "0010" when "01100101001010", -- t[6474] = 2
      "0010" when "01100101001011", -- t[6475] = 2
      "0010" when "01100101001100", -- t[6476] = 2
      "0010" when "01100101001101", -- t[6477] = 2
      "0010" when "01100101001110", -- t[6478] = 2
      "0010" when "01100101001111", -- t[6479] = 2
      "0010" when "01100101010000", -- t[6480] = 2
      "0010" when "01100101010001", -- t[6481] = 2
      "0010" when "01100101010010", -- t[6482] = 2
      "0010" when "01100101010011", -- t[6483] = 2
      "0010" when "01100101010100", -- t[6484] = 2
      "0010" when "01100101010101", -- t[6485] = 2
      "0010" when "01100101010110", -- t[6486] = 2
      "0010" when "01100101010111", -- t[6487] = 2
      "0010" when "01100101011000", -- t[6488] = 2
      "0010" when "01100101011001", -- t[6489] = 2
      "0010" when "01100101011010", -- t[6490] = 2
      "0010" when "01100101011011", -- t[6491] = 2
      "0010" when "01100101011100", -- t[6492] = 2
      "0010" when "01100101011101", -- t[6493] = 2
      "0010" when "01100101011110", -- t[6494] = 2
      "0010" when "01100101011111", -- t[6495] = 2
      "0010" when "01100101100000", -- t[6496] = 2
      "0010" when "01100101100001", -- t[6497] = 2
      "0010" when "01100101100010", -- t[6498] = 2
      "0010" when "01100101100011", -- t[6499] = 2
      "0010" when "01100101100100", -- t[6500] = 2
      "0010" when "01100101100101", -- t[6501] = 2
      "0010" when "01100101100110", -- t[6502] = 2
      "0010" when "01100101100111", -- t[6503] = 2
      "0010" when "01100101101000", -- t[6504] = 2
      "0010" when "01100101101001", -- t[6505] = 2
      "0010" when "01100101101010", -- t[6506] = 2
      "0010" when "01100101101011", -- t[6507] = 2
      "0010" when "01100101101100", -- t[6508] = 2
      "0010" when "01100101101101", -- t[6509] = 2
      "0010" when "01100101101110", -- t[6510] = 2
      "0010" when "01100101101111", -- t[6511] = 2
      "0010" when "01100101110000", -- t[6512] = 2
      "0010" when "01100101110001", -- t[6513] = 2
      "0010" when "01100101110010", -- t[6514] = 2
      "0010" when "01100101110011", -- t[6515] = 2
      "0010" when "01100101110100", -- t[6516] = 2
      "0010" when "01100101110101", -- t[6517] = 2
      "0010" when "01100101110110", -- t[6518] = 2
      "0010" when "01100101110111", -- t[6519] = 2
      "0010" when "01100101111000", -- t[6520] = 2
      "0010" when "01100101111001", -- t[6521] = 2
      "0010" when "01100101111010", -- t[6522] = 2
      "0010" when "01100101111011", -- t[6523] = 2
      "0010" when "01100101111100", -- t[6524] = 2
      "0010" when "01100101111101", -- t[6525] = 2
      "0010" when "01100101111110", -- t[6526] = 2
      "0010" when "01100101111111", -- t[6527] = 2
      "0010" when "01100110000000", -- t[6528] = 2
      "0010" when "01100110000001", -- t[6529] = 2
      "0010" when "01100110000010", -- t[6530] = 2
      "0010" when "01100110000011", -- t[6531] = 2
      "0010" when "01100110000100", -- t[6532] = 2
      "0010" when "01100110000101", -- t[6533] = 2
      "0010" when "01100110000110", -- t[6534] = 2
      "0010" when "01100110000111", -- t[6535] = 2
      "0010" when "01100110001000", -- t[6536] = 2
      "0010" when "01100110001001", -- t[6537] = 2
      "0010" when "01100110001010", -- t[6538] = 2
      "0010" when "01100110001011", -- t[6539] = 2
      "0010" when "01100110001100", -- t[6540] = 2
      "0010" when "01100110001101", -- t[6541] = 2
      "0010" when "01100110001110", -- t[6542] = 2
      "0010" when "01100110001111", -- t[6543] = 2
      "0010" when "01100110010000", -- t[6544] = 2
      "0010" when "01100110010001", -- t[6545] = 2
      "0010" when "01100110010010", -- t[6546] = 2
      "0010" when "01100110010011", -- t[6547] = 2
      "0010" when "01100110010100", -- t[6548] = 2
      "0010" when "01100110010101", -- t[6549] = 2
      "0010" when "01100110010110", -- t[6550] = 2
      "0010" when "01100110010111", -- t[6551] = 2
      "0010" when "01100110011000", -- t[6552] = 2
      "0010" when "01100110011001", -- t[6553] = 2
      "0010" when "01100110011010", -- t[6554] = 2
      "0010" when "01100110011011", -- t[6555] = 2
      "0010" when "01100110011100", -- t[6556] = 2
      "0010" when "01100110011101", -- t[6557] = 2
      "0010" when "01100110011110", -- t[6558] = 2
      "0010" when "01100110011111", -- t[6559] = 2
      "0010" when "01100110100000", -- t[6560] = 2
      "0010" when "01100110100001", -- t[6561] = 2
      "0010" when "01100110100010", -- t[6562] = 2
      "0010" when "01100110100011", -- t[6563] = 2
      "0010" when "01100110100100", -- t[6564] = 2
      "0010" when "01100110100101", -- t[6565] = 2
      "0010" when "01100110100110", -- t[6566] = 2
      "0010" when "01100110100111", -- t[6567] = 2
      "0010" when "01100110101000", -- t[6568] = 2
      "0010" when "01100110101001", -- t[6569] = 2
      "0010" when "01100110101010", -- t[6570] = 2
      "0010" when "01100110101011", -- t[6571] = 2
      "0010" when "01100110101100", -- t[6572] = 2
      "0010" when "01100110101101", -- t[6573] = 2
      "0010" when "01100110101110", -- t[6574] = 2
      "0010" when "01100110101111", -- t[6575] = 2
      "0010" when "01100110110000", -- t[6576] = 2
      "0010" when "01100110110001", -- t[6577] = 2
      "0010" when "01100110110010", -- t[6578] = 2
      "0010" when "01100110110011", -- t[6579] = 2
      "0010" when "01100110110100", -- t[6580] = 2
      "0010" when "01100110110101", -- t[6581] = 2
      "0010" when "01100110110110", -- t[6582] = 2
      "0010" when "01100110110111", -- t[6583] = 2
      "0010" when "01100110111000", -- t[6584] = 2
      "0010" when "01100110111001", -- t[6585] = 2
      "0010" when "01100110111010", -- t[6586] = 2
      "0010" when "01100110111011", -- t[6587] = 2
      "0010" when "01100110111100", -- t[6588] = 2
      "0010" when "01100110111101", -- t[6589] = 2
      "0010" when "01100110111110", -- t[6590] = 2
      "0010" when "01100110111111", -- t[6591] = 2
      "0010" when "01100111000000", -- t[6592] = 2
      "0010" when "01100111000001", -- t[6593] = 2
      "0010" when "01100111000010", -- t[6594] = 2
      "0010" when "01100111000011", -- t[6595] = 2
      "0010" when "01100111000100", -- t[6596] = 2
      "0010" when "01100111000101", -- t[6597] = 2
      "0010" when "01100111000110", -- t[6598] = 2
      "0010" when "01100111000111", -- t[6599] = 2
      "0010" when "01100111001000", -- t[6600] = 2
      "0010" when "01100111001001", -- t[6601] = 2
      "0010" when "01100111001010", -- t[6602] = 2
      "0010" when "01100111001011", -- t[6603] = 2
      "0010" when "01100111001100", -- t[6604] = 2
      "0010" when "01100111001101", -- t[6605] = 2
      "0010" when "01100111001110", -- t[6606] = 2
      "0010" when "01100111001111", -- t[6607] = 2
      "0010" when "01100111010000", -- t[6608] = 2
      "0010" when "01100111010001", -- t[6609] = 2
      "0010" when "01100111010010", -- t[6610] = 2
      "0010" when "01100111010011", -- t[6611] = 2
      "0010" when "01100111010100", -- t[6612] = 2
      "0010" when "01100111010101", -- t[6613] = 2
      "0010" when "01100111010110", -- t[6614] = 2
      "0010" when "01100111010111", -- t[6615] = 2
      "0010" when "01100111011000", -- t[6616] = 2
      "0010" when "01100111011001", -- t[6617] = 2
      "0010" when "01100111011010", -- t[6618] = 2
      "0010" when "01100111011011", -- t[6619] = 2
      "0010" when "01100111011100", -- t[6620] = 2
      "0010" when "01100111011101", -- t[6621] = 2
      "0010" when "01100111011110", -- t[6622] = 2
      "0010" when "01100111011111", -- t[6623] = 2
      "0010" when "01100111100000", -- t[6624] = 2
      "0010" when "01100111100001", -- t[6625] = 2
      "0010" when "01100111100010", -- t[6626] = 2
      "0010" when "01100111100011", -- t[6627] = 2
      "0010" when "01100111100100", -- t[6628] = 2
      "0010" when "01100111100101", -- t[6629] = 2
      "0010" when "01100111100110", -- t[6630] = 2
      "0010" when "01100111100111", -- t[6631] = 2
      "0010" when "01100111101000", -- t[6632] = 2
      "0010" when "01100111101001", -- t[6633] = 2
      "0010" when "01100111101010", -- t[6634] = 2
      "0010" when "01100111101011", -- t[6635] = 2
      "0010" when "01100111101100", -- t[6636] = 2
      "0010" when "01100111101101", -- t[6637] = 2
      "0010" when "01100111101110", -- t[6638] = 2
      "0010" when "01100111101111", -- t[6639] = 2
      "0010" when "01100111110000", -- t[6640] = 2
      "0010" when "01100111110001", -- t[6641] = 2
      "0010" when "01100111110010", -- t[6642] = 2
      "0010" when "01100111110011", -- t[6643] = 2
      "0010" when "01100111110100", -- t[6644] = 2
      "0010" when "01100111110101", -- t[6645] = 2
      "0010" when "01100111110110", -- t[6646] = 2
      "0010" when "01100111110111", -- t[6647] = 2
      "0010" when "01100111111000", -- t[6648] = 2
      "0010" when "01100111111001", -- t[6649] = 2
      "0010" when "01100111111010", -- t[6650] = 2
      "0010" when "01100111111011", -- t[6651] = 2
      "0010" when "01100111111100", -- t[6652] = 2
      "0010" when "01100111111101", -- t[6653] = 2
      "0010" when "01100111111110", -- t[6654] = 2
      "0010" when "01100111111111", -- t[6655] = 2
      "0010" when "01101000000000", -- t[6656] = 2
      "0010" when "01101000000001", -- t[6657] = 2
      "0010" when "01101000000010", -- t[6658] = 2
      "0010" when "01101000000011", -- t[6659] = 2
      "0010" when "01101000000100", -- t[6660] = 2
      "0010" when "01101000000101", -- t[6661] = 2
      "0010" when "01101000000110", -- t[6662] = 2
      "0010" when "01101000000111", -- t[6663] = 2
      "0010" when "01101000001000", -- t[6664] = 2
      "0010" when "01101000001001", -- t[6665] = 2
      "0010" when "01101000001010", -- t[6666] = 2
      "0010" when "01101000001011", -- t[6667] = 2
      "0010" when "01101000001100", -- t[6668] = 2
      "0010" when "01101000001101", -- t[6669] = 2
      "0010" when "01101000001110", -- t[6670] = 2
      "0010" when "01101000001111", -- t[6671] = 2
      "0010" when "01101000010000", -- t[6672] = 2
      "0010" when "01101000010001", -- t[6673] = 2
      "0010" when "01101000010010", -- t[6674] = 2
      "0010" when "01101000010011", -- t[6675] = 2
      "0010" when "01101000010100", -- t[6676] = 2
      "0010" when "01101000010101", -- t[6677] = 2
      "0010" when "01101000010110", -- t[6678] = 2
      "0010" when "01101000010111", -- t[6679] = 2
      "0010" when "01101000011000", -- t[6680] = 2
      "0010" when "01101000011001", -- t[6681] = 2
      "0010" when "01101000011010", -- t[6682] = 2
      "0010" when "01101000011011", -- t[6683] = 2
      "0010" when "01101000011100", -- t[6684] = 2
      "0010" when "01101000011101", -- t[6685] = 2
      "0010" when "01101000011110", -- t[6686] = 2
      "0010" when "01101000011111", -- t[6687] = 2
      "0010" when "01101000100000", -- t[6688] = 2
      "0010" when "01101000100001", -- t[6689] = 2
      "0010" when "01101000100010", -- t[6690] = 2
      "0010" when "01101000100011", -- t[6691] = 2
      "0010" when "01101000100100", -- t[6692] = 2
      "0010" when "01101000100101", -- t[6693] = 2
      "0010" when "01101000100110", -- t[6694] = 2
      "0010" when "01101000100111", -- t[6695] = 2
      "0010" when "01101000101000", -- t[6696] = 2
      "0010" when "01101000101001", -- t[6697] = 2
      "0010" when "01101000101010", -- t[6698] = 2
      "0010" when "01101000101011", -- t[6699] = 2
      "0010" when "01101000101100", -- t[6700] = 2
      "0010" when "01101000101101", -- t[6701] = 2
      "0010" when "01101000101110", -- t[6702] = 2
      "0010" when "01101000101111", -- t[6703] = 2
      "0010" when "01101000110000", -- t[6704] = 2
      "0010" when "01101000110001", -- t[6705] = 2
      "0010" when "01101000110010", -- t[6706] = 2
      "0010" when "01101000110011", -- t[6707] = 2
      "0010" when "01101000110100", -- t[6708] = 2
      "0010" when "01101000110101", -- t[6709] = 2
      "0010" when "01101000110110", -- t[6710] = 2
      "0010" when "01101000110111", -- t[6711] = 2
      "0010" when "01101000111000", -- t[6712] = 2
      "0010" when "01101000111001", -- t[6713] = 2
      "0010" when "01101000111010", -- t[6714] = 2
      "0010" when "01101000111011", -- t[6715] = 2
      "0010" when "01101000111100", -- t[6716] = 2
      "0010" when "01101000111101", -- t[6717] = 2
      "0010" when "01101000111110", -- t[6718] = 2
      "0010" when "01101000111111", -- t[6719] = 2
      "0010" when "01101001000000", -- t[6720] = 2
      "0010" when "01101001000001", -- t[6721] = 2
      "0010" when "01101001000010", -- t[6722] = 2
      "0010" when "01101001000011", -- t[6723] = 2
      "0010" when "01101001000100", -- t[6724] = 2
      "0010" when "01101001000101", -- t[6725] = 2
      "0010" when "01101001000110", -- t[6726] = 2
      "0010" when "01101001000111", -- t[6727] = 2
      "0010" when "01101001001000", -- t[6728] = 2
      "0010" when "01101001001001", -- t[6729] = 2
      "0010" when "01101001001010", -- t[6730] = 2
      "0010" when "01101001001011", -- t[6731] = 2
      "0010" when "01101001001100", -- t[6732] = 2
      "0010" when "01101001001101", -- t[6733] = 2
      "0010" when "01101001001110", -- t[6734] = 2
      "0010" when "01101001001111", -- t[6735] = 2
      "0010" when "01101001010000", -- t[6736] = 2
      "0010" when "01101001010001", -- t[6737] = 2
      "0010" when "01101001010010", -- t[6738] = 2
      "0010" when "01101001010011", -- t[6739] = 2
      "0010" when "01101001010100", -- t[6740] = 2
      "0010" when "01101001010101", -- t[6741] = 2
      "0010" when "01101001010110", -- t[6742] = 2
      "0010" when "01101001010111", -- t[6743] = 2
      "0010" when "01101001011000", -- t[6744] = 2
      "0010" when "01101001011001", -- t[6745] = 2
      "0010" when "01101001011010", -- t[6746] = 2
      "0010" when "01101001011011", -- t[6747] = 2
      "0010" when "01101001011100", -- t[6748] = 2
      "0010" when "01101001011101", -- t[6749] = 2
      "0010" when "01101001011110", -- t[6750] = 2
      "0010" when "01101001011111", -- t[6751] = 2
      "0010" when "01101001100000", -- t[6752] = 2
      "0010" when "01101001100001", -- t[6753] = 2
      "0010" when "01101001100010", -- t[6754] = 2
      "0010" when "01101001100011", -- t[6755] = 2
      "0010" when "01101001100100", -- t[6756] = 2
      "0010" when "01101001100101", -- t[6757] = 2
      "0010" when "01101001100110", -- t[6758] = 2
      "0010" when "01101001100111", -- t[6759] = 2
      "0010" when "01101001101000", -- t[6760] = 2
      "0010" when "01101001101001", -- t[6761] = 2
      "0010" when "01101001101010", -- t[6762] = 2
      "0010" when "01101001101011", -- t[6763] = 2
      "0010" when "01101001101100", -- t[6764] = 2
      "0010" when "01101001101101", -- t[6765] = 2
      "0010" when "01101001101110", -- t[6766] = 2
      "0010" when "01101001101111", -- t[6767] = 2
      "0010" when "01101001110000", -- t[6768] = 2
      "0010" when "01101001110001", -- t[6769] = 2
      "0010" when "01101001110010", -- t[6770] = 2
      "0010" when "01101001110011", -- t[6771] = 2
      "0010" when "01101001110100", -- t[6772] = 2
      "0010" when "01101001110101", -- t[6773] = 2
      "0010" when "01101001110110", -- t[6774] = 2
      "0010" when "01101001110111", -- t[6775] = 2
      "0010" when "01101001111000", -- t[6776] = 2
      "0010" when "01101001111001", -- t[6777] = 2
      "0010" when "01101001111010", -- t[6778] = 2
      "0010" when "01101001111011", -- t[6779] = 2
      "0010" when "01101001111100", -- t[6780] = 2
      "0010" when "01101001111101", -- t[6781] = 2
      "0010" when "01101001111110", -- t[6782] = 2
      "0010" when "01101001111111", -- t[6783] = 2
      "0010" when "01101010000000", -- t[6784] = 2
      "0010" when "01101010000001", -- t[6785] = 2
      "0010" when "01101010000010", -- t[6786] = 2
      "0010" when "01101010000011", -- t[6787] = 2
      "0010" when "01101010000100", -- t[6788] = 2
      "0010" when "01101010000101", -- t[6789] = 2
      "0010" when "01101010000110", -- t[6790] = 2
      "0010" when "01101010000111", -- t[6791] = 2
      "0010" when "01101010001000", -- t[6792] = 2
      "0010" when "01101010001001", -- t[6793] = 2
      "0010" when "01101010001010", -- t[6794] = 2
      "0010" when "01101010001011", -- t[6795] = 2
      "0010" when "01101010001100", -- t[6796] = 2
      "0010" when "01101010001101", -- t[6797] = 2
      "0010" when "01101010001110", -- t[6798] = 2
      "0010" when "01101010001111", -- t[6799] = 2
      "0010" when "01101010010000", -- t[6800] = 2
      "0010" when "01101010010001", -- t[6801] = 2
      "0010" when "01101010010010", -- t[6802] = 2
      "0010" when "01101010010011", -- t[6803] = 2
      "0010" when "01101010010100", -- t[6804] = 2
      "0010" when "01101010010101", -- t[6805] = 2
      "0010" when "01101010010110", -- t[6806] = 2
      "0010" when "01101010010111", -- t[6807] = 2
      "0010" when "01101010011000", -- t[6808] = 2
      "0010" when "01101010011001", -- t[6809] = 2
      "0010" when "01101010011010", -- t[6810] = 2
      "0010" when "01101010011011", -- t[6811] = 2
      "0010" when "01101010011100", -- t[6812] = 2
      "0010" when "01101010011101", -- t[6813] = 2
      "0010" when "01101010011110", -- t[6814] = 2
      "0010" when "01101010011111", -- t[6815] = 2
      "0010" when "01101010100000", -- t[6816] = 2
      "0010" when "01101010100001", -- t[6817] = 2
      "0010" when "01101010100010", -- t[6818] = 2
      "0010" when "01101010100011", -- t[6819] = 2
      "0010" when "01101010100100", -- t[6820] = 2
      "0010" when "01101010100101", -- t[6821] = 2
      "0010" when "01101010100110", -- t[6822] = 2
      "0010" when "01101010100111", -- t[6823] = 2
      "0010" when "01101010101000", -- t[6824] = 2
      "0010" when "01101010101001", -- t[6825] = 2
      "0010" when "01101010101010", -- t[6826] = 2
      "0010" when "01101010101011", -- t[6827] = 2
      "0010" when "01101010101100", -- t[6828] = 2
      "0010" when "01101010101101", -- t[6829] = 2
      "0010" when "01101010101110", -- t[6830] = 2
      "0010" when "01101010101111", -- t[6831] = 2
      "0010" when "01101010110000", -- t[6832] = 2
      "0010" when "01101010110001", -- t[6833] = 2
      "0010" when "01101010110010", -- t[6834] = 2
      "0010" when "01101010110011", -- t[6835] = 2
      "0010" when "01101010110100", -- t[6836] = 2
      "0010" when "01101010110101", -- t[6837] = 2
      "0010" when "01101010110110", -- t[6838] = 2
      "0010" when "01101010110111", -- t[6839] = 2
      "0010" when "01101010111000", -- t[6840] = 2
      "0010" when "01101010111001", -- t[6841] = 2
      "0010" when "01101010111010", -- t[6842] = 2
      "0010" when "01101010111011", -- t[6843] = 2
      "0010" when "01101010111100", -- t[6844] = 2
      "0010" when "01101010111101", -- t[6845] = 2
      "0010" when "01101010111110", -- t[6846] = 2
      "0010" when "01101010111111", -- t[6847] = 2
      "0010" when "01101011000000", -- t[6848] = 2
      "0010" when "01101011000001", -- t[6849] = 2
      "0010" when "01101011000010", -- t[6850] = 2
      "0010" when "01101011000011", -- t[6851] = 2
      "0010" when "01101011000100", -- t[6852] = 2
      "0010" when "01101011000101", -- t[6853] = 2
      "0010" when "01101011000110", -- t[6854] = 2
      "0010" when "01101011000111", -- t[6855] = 2
      "0010" when "01101011001000", -- t[6856] = 2
      "0010" when "01101011001001", -- t[6857] = 2
      "0010" when "01101011001010", -- t[6858] = 2
      "0010" when "01101011001011", -- t[6859] = 2
      "0010" when "01101011001100", -- t[6860] = 2
      "0010" when "01101011001101", -- t[6861] = 2
      "0010" when "01101011001110", -- t[6862] = 2
      "0010" when "01101011001111", -- t[6863] = 2
      "0010" when "01101011010000", -- t[6864] = 2
      "0010" when "01101011010001", -- t[6865] = 2
      "0010" when "01101011010010", -- t[6866] = 2
      "0010" when "01101011010011", -- t[6867] = 2
      "0010" when "01101011010100", -- t[6868] = 2
      "0010" when "01101011010101", -- t[6869] = 2
      "0010" when "01101011010110", -- t[6870] = 2
      "0010" when "01101011010111", -- t[6871] = 2
      "0010" when "01101011011000", -- t[6872] = 2
      "0010" when "01101011011001", -- t[6873] = 2
      "0010" when "01101011011010", -- t[6874] = 2
      "0010" when "01101011011011", -- t[6875] = 2
      "0010" when "01101011011100", -- t[6876] = 2
      "0010" when "01101011011101", -- t[6877] = 2
      "0010" when "01101011011110", -- t[6878] = 2
      "0010" when "01101011011111", -- t[6879] = 2
      "0010" when "01101011100000", -- t[6880] = 2
      "0010" when "01101011100001", -- t[6881] = 2
      "0010" when "01101011100010", -- t[6882] = 2
      "0010" when "01101011100011", -- t[6883] = 2
      "0010" when "01101011100100", -- t[6884] = 2
      "0010" when "01101011100101", -- t[6885] = 2
      "0010" when "01101011100110", -- t[6886] = 2
      "0010" when "01101011100111", -- t[6887] = 2
      "0010" when "01101011101000", -- t[6888] = 2
      "0010" when "01101011101001", -- t[6889] = 2
      "0010" when "01101011101010", -- t[6890] = 2
      "0010" when "01101011101011", -- t[6891] = 2
      "0010" when "01101011101100", -- t[6892] = 2
      "0010" when "01101011101101", -- t[6893] = 2
      "0010" when "01101011101110", -- t[6894] = 2
      "0010" when "01101011101111", -- t[6895] = 2
      "0010" when "01101011110000", -- t[6896] = 2
      "0010" when "01101011110001", -- t[6897] = 2
      "0010" when "01101011110010", -- t[6898] = 2
      "0010" when "01101011110011", -- t[6899] = 2
      "0010" when "01101011110100", -- t[6900] = 2
      "0010" when "01101011110101", -- t[6901] = 2
      "0010" when "01101011110110", -- t[6902] = 2
      "0010" when "01101011110111", -- t[6903] = 2
      "0010" when "01101011111000", -- t[6904] = 2
      "0010" when "01101011111001", -- t[6905] = 2
      "0010" when "01101011111010", -- t[6906] = 2
      "0010" when "01101011111011", -- t[6907] = 2
      "0010" when "01101011111100", -- t[6908] = 2
      "0010" when "01101011111101", -- t[6909] = 2
      "0010" when "01101011111110", -- t[6910] = 2
      "0010" when "01101011111111", -- t[6911] = 2
      "0010" when "01101100000000", -- t[6912] = 2
      "0010" when "01101100000001", -- t[6913] = 2
      "0010" when "01101100000010", -- t[6914] = 2
      "0010" when "01101100000011", -- t[6915] = 2
      "0010" when "01101100000100", -- t[6916] = 2
      "0010" when "01101100000101", -- t[6917] = 2
      "0010" when "01101100000110", -- t[6918] = 2
      "0010" when "01101100000111", -- t[6919] = 2
      "0010" when "01101100001000", -- t[6920] = 2
      "0010" when "01101100001001", -- t[6921] = 2
      "0010" when "01101100001010", -- t[6922] = 2
      "0010" when "01101100001011", -- t[6923] = 2
      "0010" when "01101100001100", -- t[6924] = 2
      "0010" when "01101100001101", -- t[6925] = 2
      "0010" when "01101100001110", -- t[6926] = 2
      "0010" when "01101100001111", -- t[6927] = 2
      "0010" when "01101100010000", -- t[6928] = 2
      "0010" when "01101100010001", -- t[6929] = 2
      "0010" when "01101100010010", -- t[6930] = 2
      "0010" when "01101100010011", -- t[6931] = 2
      "0010" when "01101100010100", -- t[6932] = 2
      "0010" when "01101100010101", -- t[6933] = 2
      "0010" when "01101100010110", -- t[6934] = 2
      "0010" when "01101100010111", -- t[6935] = 2
      "0010" when "01101100011000", -- t[6936] = 2
      "0010" when "01101100011001", -- t[6937] = 2
      "0010" when "01101100011010", -- t[6938] = 2
      "0010" when "01101100011011", -- t[6939] = 2
      "0010" when "01101100011100", -- t[6940] = 2
      "0010" when "01101100011101", -- t[6941] = 2
      "0010" when "01101100011110", -- t[6942] = 2
      "0010" when "01101100011111", -- t[6943] = 2
      "0010" when "01101100100000", -- t[6944] = 2
      "0010" when "01101100100001", -- t[6945] = 2
      "0010" when "01101100100010", -- t[6946] = 2
      "0010" when "01101100100011", -- t[6947] = 2
      "0010" when "01101100100100", -- t[6948] = 2
      "0010" when "01101100100101", -- t[6949] = 2
      "0010" when "01101100100110", -- t[6950] = 2
      "0010" when "01101100100111", -- t[6951] = 2
      "0010" when "01101100101000", -- t[6952] = 2
      "0010" when "01101100101001", -- t[6953] = 2
      "0010" when "01101100101010", -- t[6954] = 2
      "0011" when "01101100101011", -- t[6955] = 3
      "0011" when "01101100101100", -- t[6956] = 3
      "0011" when "01101100101101", -- t[6957] = 3
      "0011" when "01101100101110", -- t[6958] = 3
      "0011" when "01101100101111", -- t[6959] = 3
      "0011" when "01101100110000", -- t[6960] = 3
      "0011" when "01101100110001", -- t[6961] = 3
      "0011" when "01101100110010", -- t[6962] = 3
      "0011" when "01101100110011", -- t[6963] = 3
      "0011" when "01101100110100", -- t[6964] = 3
      "0011" when "01101100110101", -- t[6965] = 3
      "0011" when "01101100110110", -- t[6966] = 3
      "0011" when "01101100110111", -- t[6967] = 3
      "0011" when "01101100111000", -- t[6968] = 3
      "0011" when "01101100111001", -- t[6969] = 3
      "0011" when "01101100111010", -- t[6970] = 3
      "0011" when "01101100111011", -- t[6971] = 3
      "0011" when "01101100111100", -- t[6972] = 3
      "0011" when "01101100111101", -- t[6973] = 3
      "0011" when "01101100111110", -- t[6974] = 3
      "0011" when "01101100111111", -- t[6975] = 3
      "0011" when "01101101000000", -- t[6976] = 3
      "0011" when "01101101000001", -- t[6977] = 3
      "0011" when "01101101000010", -- t[6978] = 3
      "0011" when "01101101000011", -- t[6979] = 3
      "0011" when "01101101000100", -- t[6980] = 3
      "0011" when "01101101000101", -- t[6981] = 3
      "0011" when "01101101000110", -- t[6982] = 3
      "0011" when "01101101000111", -- t[6983] = 3
      "0011" when "01101101001000", -- t[6984] = 3
      "0011" when "01101101001001", -- t[6985] = 3
      "0011" when "01101101001010", -- t[6986] = 3
      "0011" when "01101101001011", -- t[6987] = 3
      "0011" when "01101101001100", -- t[6988] = 3
      "0011" when "01101101001101", -- t[6989] = 3
      "0011" when "01101101001110", -- t[6990] = 3
      "0011" when "01101101001111", -- t[6991] = 3
      "0011" when "01101101010000", -- t[6992] = 3
      "0011" when "01101101010001", -- t[6993] = 3
      "0011" when "01101101010010", -- t[6994] = 3
      "0011" when "01101101010011", -- t[6995] = 3
      "0011" when "01101101010100", -- t[6996] = 3
      "0011" when "01101101010101", -- t[6997] = 3
      "0011" when "01101101010110", -- t[6998] = 3
      "0011" when "01101101010111", -- t[6999] = 3
      "0011" when "01101101011000", -- t[7000] = 3
      "0011" when "01101101011001", -- t[7001] = 3
      "0011" when "01101101011010", -- t[7002] = 3
      "0011" when "01101101011011", -- t[7003] = 3
      "0011" when "01101101011100", -- t[7004] = 3
      "0011" when "01101101011101", -- t[7005] = 3
      "0011" when "01101101011110", -- t[7006] = 3
      "0011" when "01101101011111", -- t[7007] = 3
      "0011" when "01101101100000", -- t[7008] = 3
      "0011" when "01101101100001", -- t[7009] = 3
      "0011" when "01101101100010", -- t[7010] = 3
      "0011" when "01101101100011", -- t[7011] = 3
      "0011" when "01101101100100", -- t[7012] = 3
      "0011" when "01101101100101", -- t[7013] = 3
      "0011" when "01101101100110", -- t[7014] = 3
      "0011" when "01101101100111", -- t[7015] = 3
      "0011" when "01101101101000", -- t[7016] = 3
      "0011" when "01101101101001", -- t[7017] = 3
      "0011" when "01101101101010", -- t[7018] = 3
      "0011" when "01101101101011", -- t[7019] = 3
      "0011" when "01101101101100", -- t[7020] = 3
      "0011" when "01101101101101", -- t[7021] = 3
      "0011" when "01101101101110", -- t[7022] = 3
      "0011" when "01101101101111", -- t[7023] = 3
      "0011" when "01101101110000", -- t[7024] = 3
      "0011" when "01101101110001", -- t[7025] = 3
      "0011" when "01101101110010", -- t[7026] = 3
      "0011" when "01101101110011", -- t[7027] = 3
      "0011" when "01101101110100", -- t[7028] = 3
      "0011" when "01101101110101", -- t[7029] = 3
      "0011" when "01101101110110", -- t[7030] = 3
      "0011" when "01101101110111", -- t[7031] = 3
      "0011" when "01101101111000", -- t[7032] = 3
      "0011" when "01101101111001", -- t[7033] = 3
      "0011" when "01101101111010", -- t[7034] = 3
      "0011" when "01101101111011", -- t[7035] = 3
      "0011" when "01101101111100", -- t[7036] = 3
      "0011" when "01101101111101", -- t[7037] = 3
      "0011" when "01101101111110", -- t[7038] = 3
      "0011" when "01101101111111", -- t[7039] = 3
      "0011" when "01101110000000", -- t[7040] = 3
      "0011" when "01101110000001", -- t[7041] = 3
      "0011" when "01101110000010", -- t[7042] = 3
      "0011" when "01101110000011", -- t[7043] = 3
      "0011" when "01101110000100", -- t[7044] = 3
      "0011" when "01101110000101", -- t[7045] = 3
      "0011" when "01101110000110", -- t[7046] = 3
      "0011" when "01101110000111", -- t[7047] = 3
      "0011" when "01101110001000", -- t[7048] = 3
      "0011" when "01101110001001", -- t[7049] = 3
      "0011" when "01101110001010", -- t[7050] = 3
      "0011" when "01101110001011", -- t[7051] = 3
      "0011" when "01101110001100", -- t[7052] = 3
      "0011" when "01101110001101", -- t[7053] = 3
      "0011" when "01101110001110", -- t[7054] = 3
      "0011" when "01101110001111", -- t[7055] = 3
      "0011" when "01101110010000", -- t[7056] = 3
      "0011" when "01101110010001", -- t[7057] = 3
      "0011" when "01101110010010", -- t[7058] = 3
      "0011" when "01101110010011", -- t[7059] = 3
      "0011" when "01101110010100", -- t[7060] = 3
      "0011" when "01101110010101", -- t[7061] = 3
      "0011" when "01101110010110", -- t[7062] = 3
      "0011" when "01101110010111", -- t[7063] = 3
      "0011" when "01101110011000", -- t[7064] = 3
      "0011" when "01101110011001", -- t[7065] = 3
      "0011" when "01101110011010", -- t[7066] = 3
      "0011" when "01101110011011", -- t[7067] = 3
      "0011" when "01101110011100", -- t[7068] = 3
      "0011" when "01101110011101", -- t[7069] = 3
      "0011" when "01101110011110", -- t[7070] = 3
      "0011" when "01101110011111", -- t[7071] = 3
      "0011" when "01101110100000", -- t[7072] = 3
      "0011" when "01101110100001", -- t[7073] = 3
      "0011" when "01101110100010", -- t[7074] = 3
      "0011" when "01101110100011", -- t[7075] = 3
      "0011" when "01101110100100", -- t[7076] = 3
      "0011" when "01101110100101", -- t[7077] = 3
      "0011" when "01101110100110", -- t[7078] = 3
      "0011" when "01101110100111", -- t[7079] = 3
      "0011" when "01101110101000", -- t[7080] = 3
      "0011" when "01101110101001", -- t[7081] = 3
      "0011" when "01101110101010", -- t[7082] = 3
      "0011" when "01101110101011", -- t[7083] = 3
      "0011" when "01101110101100", -- t[7084] = 3
      "0011" when "01101110101101", -- t[7085] = 3
      "0011" when "01101110101110", -- t[7086] = 3
      "0011" when "01101110101111", -- t[7087] = 3
      "0011" when "01101110110000", -- t[7088] = 3
      "0011" when "01101110110001", -- t[7089] = 3
      "0011" when "01101110110010", -- t[7090] = 3
      "0011" when "01101110110011", -- t[7091] = 3
      "0011" when "01101110110100", -- t[7092] = 3
      "0011" when "01101110110101", -- t[7093] = 3
      "0011" when "01101110110110", -- t[7094] = 3
      "0011" when "01101110110111", -- t[7095] = 3
      "0011" when "01101110111000", -- t[7096] = 3
      "0011" when "01101110111001", -- t[7097] = 3
      "0011" when "01101110111010", -- t[7098] = 3
      "0011" when "01101110111011", -- t[7099] = 3
      "0011" when "01101110111100", -- t[7100] = 3
      "0011" when "01101110111101", -- t[7101] = 3
      "0011" when "01101110111110", -- t[7102] = 3
      "0011" when "01101110111111", -- t[7103] = 3
      "0011" when "01101111000000", -- t[7104] = 3
      "0011" when "01101111000001", -- t[7105] = 3
      "0011" when "01101111000010", -- t[7106] = 3
      "0011" when "01101111000011", -- t[7107] = 3
      "0011" when "01101111000100", -- t[7108] = 3
      "0011" when "01101111000101", -- t[7109] = 3
      "0011" when "01101111000110", -- t[7110] = 3
      "0011" when "01101111000111", -- t[7111] = 3
      "0011" when "01101111001000", -- t[7112] = 3
      "0011" when "01101111001001", -- t[7113] = 3
      "0011" when "01101111001010", -- t[7114] = 3
      "0011" when "01101111001011", -- t[7115] = 3
      "0011" when "01101111001100", -- t[7116] = 3
      "0011" when "01101111001101", -- t[7117] = 3
      "0011" when "01101111001110", -- t[7118] = 3
      "0011" when "01101111001111", -- t[7119] = 3
      "0011" when "01101111010000", -- t[7120] = 3
      "0011" when "01101111010001", -- t[7121] = 3
      "0011" when "01101111010010", -- t[7122] = 3
      "0011" when "01101111010011", -- t[7123] = 3
      "0011" when "01101111010100", -- t[7124] = 3
      "0011" when "01101111010101", -- t[7125] = 3
      "0011" when "01101111010110", -- t[7126] = 3
      "0011" when "01101111010111", -- t[7127] = 3
      "0011" when "01101111011000", -- t[7128] = 3
      "0011" when "01101111011001", -- t[7129] = 3
      "0011" when "01101111011010", -- t[7130] = 3
      "0011" when "01101111011011", -- t[7131] = 3
      "0011" when "01101111011100", -- t[7132] = 3
      "0011" when "01101111011101", -- t[7133] = 3
      "0011" when "01101111011110", -- t[7134] = 3
      "0011" when "01101111011111", -- t[7135] = 3
      "0011" when "01101111100000", -- t[7136] = 3
      "0011" when "01101111100001", -- t[7137] = 3
      "0011" when "01101111100010", -- t[7138] = 3
      "0011" when "01101111100011", -- t[7139] = 3
      "0011" when "01101111100100", -- t[7140] = 3
      "0011" when "01101111100101", -- t[7141] = 3
      "0011" when "01101111100110", -- t[7142] = 3
      "0011" when "01101111100111", -- t[7143] = 3
      "0011" when "01101111101000", -- t[7144] = 3
      "0011" when "01101111101001", -- t[7145] = 3
      "0011" when "01101111101010", -- t[7146] = 3
      "0011" when "01101111101011", -- t[7147] = 3
      "0011" when "01101111101100", -- t[7148] = 3
      "0011" when "01101111101101", -- t[7149] = 3
      "0011" when "01101111101110", -- t[7150] = 3
      "0011" when "01101111101111", -- t[7151] = 3
      "0011" when "01101111110000", -- t[7152] = 3
      "0011" when "01101111110001", -- t[7153] = 3
      "0011" when "01101111110010", -- t[7154] = 3
      "0011" when "01101111110011", -- t[7155] = 3
      "0011" when "01101111110100", -- t[7156] = 3
      "0011" when "01101111110101", -- t[7157] = 3
      "0011" when "01101111110110", -- t[7158] = 3
      "0011" when "01101111110111", -- t[7159] = 3
      "0011" when "01101111111000", -- t[7160] = 3
      "0011" when "01101111111001", -- t[7161] = 3
      "0011" when "01101111111010", -- t[7162] = 3
      "0011" when "01101111111011", -- t[7163] = 3
      "0011" when "01101111111100", -- t[7164] = 3
      "0011" when "01101111111101", -- t[7165] = 3
      "0011" when "01101111111110", -- t[7166] = 3
      "0011" when "01101111111111", -- t[7167] = 3
      "0011" when "01110000000000", -- t[7168] = 3
      "0011" when "01110000000001", -- t[7169] = 3
      "0011" when "01110000000010", -- t[7170] = 3
      "0011" when "01110000000011", -- t[7171] = 3
      "0011" when "01110000000100", -- t[7172] = 3
      "0011" when "01110000000101", -- t[7173] = 3
      "0011" when "01110000000110", -- t[7174] = 3
      "0011" when "01110000000111", -- t[7175] = 3
      "0011" when "01110000001000", -- t[7176] = 3
      "0011" when "01110000001001", -- t[7177] = 3
      "0011" when "01110000001010", -- t[7178] = 3
      "0011" when "01110000001011", -- t[7179] = 3
      "0011" when "01110000001100", -- t[7180] = 3
      "0011" when "01110000001101", -- t[7181] = 3
      "0011" when "01110000001110", -- t[7182] = 3
      "0011" when "01110000001111", -- t[7183] = 3
      "0011" when "01110000010000", -- t[7184] = 3
      "0011" when "01110000010001", -- t[7185] = 3
      "0011" when "01110000010010", -- t[7186] = 3
      "0011" when "01110000010011", -- t[7187] = 3
      "0011" when "01110000010100", -- t[7188] = 3
      "0011" when "01110000010101", -- t[7189] = 3
      "0011" when "01110000010110", -- t[7190] = 3
      "0011" when "01110000010111", -- t[7191] = 3
      "0011" when "01110000011000", -- t[7192] = 3
      "0011" when "01110000011001", -- t[7193] = 3
      "0011" when "01110000011010", -- t[7194] = 3
      "0011" when "01110000011011", -- t[7195] = 3
      "0011" when "01110000011100", -- t[7196] = 3
      "0011" when "01110000011101", -- t[7197] = 3
      "0011" when "01110000011110", -- t[7198] = 3
      "0011" when "01110000011111", -- t[7199] = 3
      "0011" when "01110000100000", -- t[7200] = 3
      "0011" when "01110000100001", -- t[7201] = 3
      "0011" when "01110000100010", -- t[7202] = 3
      "0011" when "01110000100011", -- t[7203] = 3
      "0011" when "01110000100100", -- t[7204] = 3
      "0011" when "01110000100101", -- t[7205] = 3
      "0011" when "01110000100110", -- t[7206] = 3
      "0011" when "01110000100111", -- t[7207] = 3
      "0011" when "01110000101000", -- t[7208] = 3
      "0011" when "01110000101001", -- t[7209] = 3
      "0011" when "01110000101010", -- t[7210] = 3
      "0011" when "01110000101011", -- t[7211] = 3
      "0011" when "01110000101100", -- t[7212] = 3
      "0011" when "01110000101101", -- t[7213] = 3
      "0011" when "01110000101110", -- t[7214] = 3
      "0011" when "01110000101111", -- t[7215] = 3
      "0011" when "01110000110000", -- t[7216] = 3
      "0011" when "01110000110001", -- t[7217] = 3
      "0011" when "01110000110010", -- t[7218] = 3
      "0011" when "01110000110011", -- t[7219] = 3
      "0011" when "01110000110100", -- t[7220] = 3
      "0011" when "01110000110101", -- t[7221] = 3
      "0011" when "01110000110110", -- t[7222] = 3
      "0011" when "01110000110111", -- t[7223] = 3
      "0011" when "01110000111000", -- t[7224] = 3
      "0011" when "01110000111001", -- t[7225] = 3
      "0011" when "01110000111010", -- t[7226] = 3
      "0011" when "01110000111011", -- t[7227] = 3
      "0011" when "01110000111100", -- t[7228] = 3
      "0011" when "01110000111101", -- t[7229] = 3
      "0011" when "01110000111110", -- t[7230] = 3
      "0011" when "01110000111111", -- t[7231] = 3
      "0011" when "01110001000000", -- t[7232] = 3
      "0011" when "01110001000001", -- t[7233] = 3
      "0011" when "01110001000010", -- t[7234] = 3
      "0011" when "01110001000011", -- t[7235] = 3
      "0011" when "01110001000100", -- t[7236] = 3
      "0011" when "01110001000101", -- t[7237] = 3
      "0011" when "01110001000110", -- t[7238] = 3
      "0011" when "01110001000111", -- t[7239] = 3
      "0011" when "01110001001000", -- t[7240] = 3
      "0011" when "01110001001001", -- t[7241] = 3
      "0011" when "01110001001010", -- t[7242] = 3
      "0011" when "01110001001011", -- t[7243] = 3
      "0011" when "01110001001100", -- t[7244] = 3
      "0011" when "01110001001101", -- t[7245] = 3
      "0011" when "01110001001110", -- t[7246] = 3
      "0011" when "01110001001111", -- t[7247] = 3
      "0011" when "01110001010000", -- t[7248] = 3
      "0011" when "01110001010001", -- t[7249] = 3
      "0011" when "01110001010010", -- t[7250] = 3
      "0011" when "01110001010011", -- t[7251] = 3
      "0011" when "01110001010100", -- t[7252] = 3
      "0011" when "01110001010101", -- t[7253] = 3
      "0011" when "01110001010110", -- t[7254] = 3
      "0011" when "01110001010111", -- t[7255] = 3
      "0011" when "01110001011000", -- t[7256] = 3
      "0011" when "01110001011001", -- t[7257] = 3
      "0011" when "01110001011010", -- t[7258] = 3
      "0011" when "01110001011011", -- t[7259] = 3
      "0011" when "01110001011100", -- t[7260] = 3
      "0011" when "01110001011101", -- t[7261] = 3
      "0011" when "01110001011110", -- t[7262] = 3
      "0011" when "01110001011111", -- t[7263] = 3
      "0011" when "01110001100000", -- t[7264] = 3
      "0011" when "01110001100001", -- t[7265] = 3
      "0011" when "01110001100010", -- t[7266] = 3
      "0011" when "01110001100011", -- t[7267] = 3
      "0011" when "01110001100100", -- t[7268] = 3
      "0011" when "01110001100101", -- t[7269] = 3
      "0011" when "01110001100110", -- t[7270] = 3
      "0011" when "01110001100111", -- t[7271] = 3
      "0011" when "01110001101000", -- t[7272] = 3
      "0011" when "01110001101001", -- t[7273] = 3
      "0011" when "01110001101010", -- t[7274] = 3
      "0011" when "01110001101011", -- t[7275] = 3
      "0011" when "01110001101100", -- t[7276] = 3
      "0011" when "01110001101101", -- t[7277] = 3
      "0011" when "01110001101110", -- t[7278] = 3
      "0011" when "01110001101111", -- t[7279] = 3
      "0011" when "01110001110000", -- t[7280] = 3
      "0011" when "01110001110001", -- t[7281] = 3
      "0011" when "01110001110010", -- t[7282] = 3
      "0011" when "01110001110011", -- t[7283] = 3
      "0011" when "01110001110100", -- t[7284] = 3
      "0011" when "01110001110101", -- t[7285] = 3
      "0011" when "01110001110110", -- t[7286] = 3
      "0011" when "01110001110111", -- t[7287] = 3
      "0011" when "01110001111000", -- t[7288] = 3
      "0011" when "01110001111001", -- t[7289] = 3
      "0011" when "01110001111010", -- t[7290] = 3
      "0011" when "01110001111011", -- t[7291] = 3
      "0011" when "01110001111100", -- t[7292] = 3
      "0011" when "01110001111101", -- t[7293] = 3
      "0011" when "01110001111110", -- t[7294] = 3
      "0011" when "01110001111111", -- t[7295] = 3
      "0011" when "01110010000000", -- t[7296] = 3
      "0011" when "01110010000001", -- t[7297] = 3
      "0011" when "01110010000010", -- t[7298] = 3
      "0011" when "01110010000011", -- t[7299] = 3
      "0011" when "01110010000100", -- t[7300] = 3
      "0011" when "01110010000101", -- t[7301] = 3
      "0011" when "01110010000110", -- t[7302] = 3
      "0011" when "01110010000111", -- t[7303] = 3
      "0011" when "01110010001000", -- t[7304] = 3
      "0011" when "01110010001001", -- t[7305] = 3
      "0011" when "01110010001010", -- t[7306] = 3
      "0011" when "01110010001011", -- t[7307] = 3
      "0011" when "01110010001100", -- t[7308] = 3
      "0011" when "01110010001101", -- t[7309] = 3
      "0011" when "01110010001110", -- t[7310] = 3
      "0011" when "01110010001111", -- t[7311] = 3
      "0011" when "01110010010000", -- t[7312] = 3
      "0011" when "01110010010001", -- t[7313] = 3
      "0011" when "01110010010010", -- t[7314] = 3
      "0011" when "01110010010011", -- t[7315] = 3
      "0011" when "01110010010100", -- t[7316] = 3
      "0011" when "01110010010101", -- t[7317] = 3
      "0011" when "01110010010110", -- t[7318] = 3
      "0011" when "01110010010111", -- t[7319] = 3
      "0011" when "01110010011000", -- t[7320] = 3
      "0011" when "01110010011001", -- t[7321] = 3
      "0011" when "01110010011010", -- t[7322] = 3
      "0011" when "01110010011011", -- t[7323] = 3
      "0011" when "01110010011100", -- t[7324] = 3
      "0011" when "01110010011101", -- t[7325] = 3
      "0011" when "01110010011110", -- t[7326] = 3
      "0011" when "01110010011111", -- t[7327] = 3
      "0011" when "01110010100000", -- t[7328] = 3
      "0011" when "01110010100001", -- t[7329] = 3
      "0011" when "01110010100010", -- t[7330] = 3
      "0011" when "01110010100011", -- t[7331] = 3
      "0011" when "01110010100100", -- t[7332] = 3
      "0011" when "01110010100101", -- t[7333] = 3
      "0011" when "01110010100110", -- t[7334] = 3
      "0011" when "01110010100111", -- t[7335] = 3
      "0011" when "01110010101000", -- t[7336] = 3
      "0011" when "01110010101001", -- t[7337] = 3
      "0011" when "01110010101010", -- t[7338] = 3
      "0011" when "01110010101011", -- t[7339] = 3
      "0011" when "01110010101100", -- t[7340] = 3
      "0011" when "01110010101101", -- t[7341] = 3
      "0011" when "01110010101110", -- t[7342] = 3
      "0011" when "01110010101111", -- t[7343] = 3
      "0011" when "01110010110000", -- t[7344] = 3
      "0011" when "01110010110001", -- t[7345] = 3
      "0011" when "01110010110010", -- t[7346] = 3
      "0011" when "01110010110011", -- t[7347] = 3
      "0011" when "01110010110100", -- t[7348] = 3
      "0011" when "01110010110101", -- t[7349] = 3
      "0011" when "01110010110110", -- t[7350] = 3
      "0011" when "01110010110111", -- t[7351] = 3
      "0011" when "01110010111000", -- t[7352] = 3
      "0011" when "01110010111001", -- t[7353] = 3
      "0011" when "01110010111010", -- t[7354] = 3
      "0011" when "01110010111011", -- t[7355] = 3
      "0011" when "01110010111100", -- t[7356] = 3
      "0011" when "01110010111101", -- t[7357] = 3
      "0011" when "01110010111110", -- t[7358] = 3
      "0011" when "01110010111111", -- t[7359] = 3
      "0011" when "01110011000000", -- t[7360] = 3
      "0011" when "01110011000001", -- t[7361] = 3
      "0011" when "01110011000010", -- t[7362] = 3
      "0011" when "01110011000011", -- t[7363] = 3
      "0011" when "01110011000100", -- t[7364] = 3
      "0011" when "01110011000101", -- t[7365] = 3
      "0011" when "01110011000110", -- t[7366] = 3
      "0011" when "01110011000111", -- t[7367] = 3
      "0011" when "01110011001000", -- t[7368] = 3
      "0011" when "01110011001001", -- t[7369] = 3
      "0011" when "01110011001010", -- t[7370] = 3
      "0011" when "01110011001011", -- t[7371] = 3
      "0011" when "01110011001100", -- t[7372] = 3
      "0011" when "01110011001101", -- t[7373] = 3
      "0011" when "01110011001110", -- t[7374] = 3
      "0011" when "01110011001111", -- t[7375] = 3
      "0011" when "01110011010000", -- t[7376] = 3
      "0011" when "01110011010001", -- t[7377] = 3
      "0011" when "01110011010010", -- t[7378] = 3
      "0011" when "01110011010011", -- t[7379] = 3
      "0011" when "01110011010100", -- t[7380] = 3
      "0011" when "01110011010101", -- t[7381] = 3
      "0011" when "01110011010110", -- t[7382] = 3
      "0011" when "01110011010111", -- t[7383] = 3
      "0011" when "01110011011000", -- t[7384] = 3
      "0011" when "01110011011001", -- t[7385] = 3
      "0011" when "01110011011010", -- t[7386] = 3
      "0011" when "01110011011011", -- t[7387] = 3
      "0011" when "01110011011100", -- t[7388] = 3
      "0011" when "01110011011101", -- t[7389] = 3
      "0011" when "01110011011110", -- t[7390] = 3
      "0011" when "01110011011111", -- t[7391] = 3
      "0011" when "01110011100000", -- t[7392] = 3
      "0011" when "01110011100001", -- t[7393] = 3
      "0011" when "01110011100010", -- t[7394] = 3
      "0011" when "01110011100011", -- t[7395] = 3
      "0011" when "01110011100100", -- t[7396] = 3
      "0011" when "01110011100101", -- t[7397] = 3
      "0011" when "01110011100110", -- t[7398] = 3
      "0011" when "01110011100111", -- t[7399] = 3
      "0011" when "01110011101000", -- t[7400] = 3
      "0011" when "01110011101001", -- t[7401] = 3
      "0011" when "01110011101010", -- t[7402] = 3
      "0011" when "01110011101011", -- t[7403] = 3
      "0011" when "01110011101100", -- t[7404] = 3
      "0011" when "01110011101101", -- t[7405] = 3
      "0011" when "01110011101110", -- t[7406] = 3
      "0011" when "01110011101111", -- t[7407] = 3
      "0011" when "01110011110000", -- t[7408] = 3
      "0011" when "01110011110001", -- t[7409] = 3
      "0011" when "01110011110010", -- t[7410] = 3
      "0011" when "01110011110011", -- t[7411] = 3
      "0011" when "01110011110100", -- t[7412] = 3
      "0011" when "01110011110101", -- t[7413] = 3
      "0011" when "01110011110110", -- t[7414] = 3
      "0011" when "01110011110111", -- t[7415] = 3
      "0011" when "01110011111000", -- t[7416] = 3
      "0011" when "01110011111001", -- t[7417] = 3
      "0011" when "01110011111010", -- t[7418] = 3
      "0011" when "01110011111011", -- t[7419] = 3
      "0011" when "01110011111100", -- t[7420] = 3
      "0011" when "01110011111101", -- t[7421] = 3
      "0011" when "01110011111110", -- t[7422] = 3
      "0011" when "01110011111111", -- t[7423] = 3
      "0011" when "01110100000000", -- t[7424] = 3
      "0011" when "01110100000001", -- t[7425] = 3
      "0011" when "01110100000010", -- t[7426] = 3
      "0011" when "01110100000011", -- t[7427] = 3
      "0011" when "01110100000100", -- t[7428] = 3
      "0011" when "01110100000101", -- t[7429] = 3
      "0011" when "01110100000110", -- t[7430] = 3
      "0011" when "01110100000111", -- t[7431] = 3
      "0011" when "01110100001000", -- t[7432] = 3
      "0011" when "01110100001001", -- t[7433] = 3
      "0011" when "01110100001010", -- t[7434] = 3
      "0011" when "01110100001011", -- t[7435] = 3
      "0011" when "01110100001100", -- t[7436] = 3
      "0011" when "01110100001101", -- t[7437] = 3
      "0011" when "01110100001110", -- t[7438] = 3
      "0011" when "01110100001111", -- t[7439] = 3
      "0011" when "01110100010000", -- t[7440] = 3
      "0011" when "01110100010001", -- t[7441] = 3
      "0011" when "01110100010010", -- t[7442] = 3
      "0011" when "01110100010011", -- t[7443] = 3
      "0011" when "01110100010100", -- t[7444] = 3
      "0011" when "01110100010101", -- t[7445] = 3
      "0011" when "01110100010110", -- t[7446] = 3
      "0011" when "01110100010111", -- t[7447] = 3
      "0011" when "01110100011000", -- t[7448] = 3
      "0011" when "01110100011001", -- t[7449] = 3
      "0011" when "01110100011010", -- t[7450] = 3
      "0011" when "01110100011011", -- t[7451] = 3
      "0100" when "01110100011100", -- t[7452] = 4
      "0100" when "01110100011101", -- t[7453] = 4
      "0100" when "01110100011110", -- t[7454] = 4
      "0100" when "01110100011111", -- t[7455] = 4
      "0100" when "01110100100000", -- t[7456] = 4
      "0100" when "01110100100001", -- t[7457] = 4
      "0100" when "01110100100010", -- t[7458] = 4
      "0100" when "01110100100011", -- t[7459] = 4
      "0100" when "01110100100100", -- t[7460] = 4
      "0100" when "01110100100101", -- t[7461] = 4
      "0100" when "01110100100110", -- t[7462] = 4
      "0100" when "01110100100111", -- t[7463] = 4
      "0100" when "01110100101000", -- t[7464] = 4
      "0100" when "01110100101001", -- t[7465] = 4
      "0100" when "01110100101010", -- t[7466] = 4
      "0100" when "01110100101011", -- t[7467] = 4
      "0100" when "01110100101100", -- t[7468] = 4
      "0100" when "01110100101101", -- t[7469] = 4
      "0100" when "01110100101110", -- t[7470] = 4
      "0100" when "01110100101111", -- t[7471] = 4
      "0100" when "01110100110000", -- t[7472] = 4
      "0100" when "01110100110001", -- t[7473] = 4
      "0100" when "01110100110010", -- t[7474] = 4
      "0100" when "01110100110011", -- t[7475] = 4
      "0100" when "01110100110100", -- t[7476] = 4
      "0100" when "01110100110101", -- t[7477] = 4
      "0100" when "01110100110110", -- t[7478] = 4
      "0100" when "01110100110111", -- t[7479] = 4
      "0100" when "01110100111000", -- t[7480] = 4
      "0100" when "01110100111001", -- t[7481] = 4
      "0100" when "01110100111010", -- t[7482] = 4
      "0100" when "01110100111011", -- t[7483] = 4
      "0100" when "01110100111100", -- t[7484] = 4
      "0100" when "01110100111101", -- t[7485] = 4
      "0100" when "01110100111110", -- t[7486] = 4
      "0100" when "01110100111111", -- t[7487] = 4
      "0100" when "01110101000000", -- t[7488] = 4
      "0100" when "01110101000001", -- t[7489] = 4
      "0100" when "01110101000010", -- t[7490] = 4
      "0100" when "01110101000011", -- t[7491] = 4
      "0100" when "01110101000100", -- t[7492] = 4
      "0100" when "01110101000101", -- t[7493] = 4
      "0100" when "01110101000110", -- t[7494] = 4
      "0100" when "01110101000111", -- t[7495] = 4
      "0100" when "01110101001000", -- t[7496] = 4
      "0100" when "01110101001001", -- t[7497] = 4
      "0100" when "01110101001010", -- t[7498] = 4
      "0100" when "01110101001011", -- t[7499] = 4
      "0100" when "01110101001100", -- t[7500] = 4
      "0100" when "01110101001101", -- t[7501] = 4
      "0100" when "01110101001110", -- t[7502] = 4
      "0100" when "01110101001111", -- t[7503] = 4
      "0100" when "01110101010000", -- t[7504] = 4
      "0100" when "01110101010001", -- t[7505] = 4
      "0100" when "01110101010010", -- t[7506] = 4
      "0100" when "01110101010011", -- t[7507] = 4
      "0100" when "01110101010100", -- t[7508] = 4
      "0100" when "01110101010101", -- t[7509] = 4
      "0100" when "01110101010110", -- t[7510] = 4
      "0100" when "01110101010111", -- t[7511] = 4
      "0100" when "01110101011000", -- t[7512] = 4
      "0100" when "01110101011001", -- t[7513] = 4
      "0100" when "01110101011010", -- t[7514] = 4
      "0100" when "01110101011011", -- t[7515] = 4
      "0100" when "01110101011100", -- t[7516] = 4
      "0100" when "01110101011101", -- t[7517] = 4
      "0100" when "01110101011110", -- t[7518] = 4
      "0100" when "01110101011111", -- t[7519] = 4
      "0100" when "01110101100000", -- t[7520] = 4
      "0100" when "01110101100001", -- t[7521] = 4
      "0100" when "01110101100010", -- t[7522] = 4
      "0100" when "01110101100011", -- t[7523] = 4
      "0100" when "01110101100100", -- t[7524] = 4
      "0100" when "01110101100101", -- t[7525] = 4
      "0100" when "01110101100110", -- t[7526] = 4
      "0100" when "01110101100111", -- t[7527] = 4
      "0100" when "01110101101000", -- t[7528] = 4
      "0100" when "01110101101001", -- t[7529] = 4
      "0100" when "01110101101010", -- t[7530] = 4
      "0100" when "01110101101011", -- t[7531] = 4
      "0100" when "01110101101100", -- t[7532] = 4
      "0100" when "01110101101101", -- t[7533] = 4
      "0100" when "01110101101110", -- t[7534] = 4
      "0100" when "01110101101111", -- t[7535] = 4
      "0100" when "01110101110000", -- t[7536] = 4
      "0100" when "01110101110001", -- t[7537] = 4
      "0100" when "01110101110010", -- t[7538] = 4
      "0100" when "01110101110011", -- t[7539] = 4
      "0100" when "01110101110100", -- t[7540] = 4
      "0100" when "01110101110101", -- t[7541] = 4
      "0100" when "01110101110110", -- t[7542] = 4
      "0100" when "01110101110111", -- t[7543] = 4
      "0100" when "01110101111000", -- t[7544] = 4
      "0100" when "01110101111001", -- t[7545] = 4
      "0100" when "01110101111010", -- t[7546] = 4
      "0100" when "01110101111011", -- t[7547] = 4
      "0100" when "01110101111100", -- t[7548] = 4
      "0100" when "01110101111101", -- t[7549] = 4
      "0100" when "01110101111110", -- t[7550] = 4
      "0100" when "01110101111111", -- t[7551] = 4
      "0100" when "01110110000000", -- t[7552] = 4
      "0100" when "01110110000001", -- t[7553] = 4
      "0100" when "01110110000010", -- t[7554] = 4
      "0100" when "01110110000011", -- t[7555] = 4
      "0100" when "01110110000100", -- t[7556] = 4
      "0100" when "01110110000101", -- t[7557] = 4
      "0100" when "01110110000110", -- t[7558] = 4
      "0100" when "01110110000111", -- t[7559] = 4
      "0100" when "01110110001000", -- t[7560] = 4
      "0100" when "01110110001001", -- t[7561] = 4
      "0100" when "01110110001010", -- t[7562] = 4
      "0100" when "01110110001011", -- t[7563] = 4
      "0100" when "01110110001100", -- t[7564] = 4
      "0100" when "01110110001101", -- t[7565] = 4
      "0100" when "01110110001110", -- t[7566] = 4
      "0100" when "01110110001111", -- t[7567] = 4
      "0100" when "01110110010000", -- t[7568] = 4
      "0100" when "01110110010001", -- t[7569] = 4
      "0100" when "01110110010010", -- t[7570] = 4
      "0100" when "01110110010011", -- t[7571] = 4
      "0100" when "01110110010100", -- t[7572] = 4
      "0100" when "01110110010101", -- t[7573] = 4
      "0100" when "01110110010110", -- t[7574] = 4
      "0100" when "01110110010111", -- t[7575] = 4
      "0100" when "01110110011000", -- t[7576] = 4
      "0100" when "01110110011001", -- t[7577] = 4
      "0100" when "01110110011010", -- t[7578] = 4
      "0100" when "01110110011011", -- t[7579] = 4
      "0100" when "01110110011100", -- t[7580] = 4
      "0100" when "01110110011101", -- t[7581] = 4
      "0100" when "01110110011110", -- t[7582] = 4
      "0100" when "01110110011111", -- t[7583] = 4
      "0100" when "01110110100000", -- t[7584] = 4
      "0100" when "01110110100001", -- t[7585] = 4
      "0100" when "01110110100010", -- t[7586] = 4
      "0100" when "01110110100011", -- t[7587] = 4
      "0100" when "01110110100100", -- t[7588] = 4
      "0100" when "01110110100101", -- t[7589] = 4
      "0100" when "01110110100110", -- t[7590] = 4
      "0100" when "01110110100111", -- t[7591] = 4
      "0100" when "01110110101000", -- t[7592] = 4
      "0100" when "01110110101001", -- t[7593] = 4
      "0100" when "01110110101010", -- t[7594] = 4
      "0100" when "01110110101011", -- t[7595] = 4
      "0100" when "01110110101100", -- t[7596] = 4
      "0100" when "01110110101101", -- t[7597] = 4
      "0100" when "01110110101110", -- t[7598] = 4
      "0100" when "01110110101111", -- t[7599] = 4
      "0100" when "01110110110000", -- t[7600] = 4
      "0100" when "01110110110001", -- t[7601] = 4
      "0100" when "01110110110010", -- t[7602] = 4
      "0100" when "01110110110011", -- t[7603] = 4
      "0100" when "01110110110100", -- t[7604] = 4
      "0100" when "01110110110101", -- t[7605] = 4
      "0100" when "01110110110110", -- t[7606] = 4
      "0100" when "01110110110111", -- t[7607] = 4
      "0100" when "01110110111000", -- t[7608] = 4
      "0100" when "01110110111001", -- t[7609] = 4
      "0100" when "01110110111010", -- t[7610] = 4
      "0100" when "01110110111011", -- t[7611] = 4
      "0100" when "01110110111100", -- t[7612] = 4
      "0100" when "01110110111101", -- t[7613] = 4
      "0100" when "01110110111110", -- t[7614] = 4
      "0100" when "01110110111111", -- t[7615] = 4
      "0100" when "01110111000000", -- t[7616] = 4
      "0100" when "01110111000001", -- t[7617] = 4
      "0100" when "01110111000010", -- t[7618] = 4
      "0100" when "01110111000011", -- t[7619] = 4
      "0100" when "01110111000100", -- t[7620] = 4
      "0100" when "01110111000101", -- t[7621] = 4
      "0100" when "01110111000110", -- t[7622] = 4
      "0100" when "01110111000111", -- t[7623] = 4
      "0100" when "01110111001000", -- t[7624] = 4
      "0100" when "01110111001001", -- t[7625] = 4
      "0100" when "01110111001010", -- t[7626] = 4
      "0100" when "01110111001011", -- t[7627] = 4
      "0100" when "01110111001100", -- t[7628] = 4
      "0100" when "01110111001101", -- t[7629] = 4
      "0100" when "01110111001110", -- t[7630] = 4
      "0100" when "01110111001111", -- t[7631] = 4
      "0100" when "01110111010000", -- t[7632] = 4
      "0100" when "01110111010001", -- t[7633] = 4
      "0100" when "01110111010010", -- t[7634] = 4
      "0100" when "01110111010011", -- t[7635] = 4
      "0100" when "01110111010100", -- t[7636] = 4
      "0100" when "01110111010101", -- t[7637] = 4
      "0100" when "01110111010110", -- t[7638] = 4
      "0100" when "01110111010111", -- t[7639] = 4
      "0100" when "01110111011000", -- t[7640] = 4
      "0100" when "01110111011001", -- t[7641] = 4
      "0100" when "01110111011010", -- t[7642] = 4
      "0100" when "01110111011011", -- t[7643] = 4
      "0100" when "01110111011100", -- t[7644] = 4
      "0100" when "01110111011101", -- t[7645] = 4
      "0100" when "01110111011110", -- t[7646] = 4
      "0100" when "01110111011111", -- t[7647] = 4
      "0100" when "01110111100000", -- t[7648] = 4
      "0100" when "01110111100001", -- t[7649] = 4
      "0100" when "01110111100010", -- t[7650] = 4
      "0100" when "01110111100011", -- t[7651] = 4
      "0100" when "01110111100100", -- t[7652] = 4
      "0100" when "01110111100101", -- t[7653] = 4
      "0100" when "01110111100110", -- t[7654] = 4
      "0100" when "01110111100111", -- t[7655] = 4
      "0100" when "01110111101000", -- t[7656] = 4
      "0100" when "01110111101001", -- t[7657] = 4
      "0100" when "01110111101010", -- t[7658] = 4
      "0100" when "01110111101011", -- t[7659] = 4
      "0100" when "01110111101100", -- t[7660] = 4
      "0100" when "01110111101101", -- t[7661] = 4
      "0100" when "01110111101110", -- t[7662] = 4
      "0100" when "01110111101111", -- t[7663] = 4
      "0100" when "01110111110000", -- t[7664] = 4
      "0100" when "01110111110001", -- t[7665] = 4
      "0100" when "01110111110010", -- t[7666] = 4
      "0100" when "01110111110011", -- t[7667] = 4
      "0100" when "01110111110100", -- t[7668] = 4
      "0100" when "01110111110101", -- t[7669] = 4
      "0100" when "01110111110110", -- t[7670] = 4
      "0100" when "01110111110111", -- t[7671] = 4
      "0100" when "01110111111000", -- t[7672] = 4
      "0100" when "01110111111001", -- t[7673] = 4
      "0100" when "01110111111010", -- t[7674] = 4
      "0100" when "01110111111011", -- t[7675] = 4
      "0100" when "01110111111100", -- t[7676] = 4
      "0100" when "01110111111101", -- t[7677] = 4
      "0100" when "01110111111110", -- t[7678] = 4
      "0100" when "01110111111111", -- t[7679] = 4
      "0100" when "01111000000000", -- t[7680] = 4
      "0100" when "01111000000001", -- t[7681] = 4
      "0100" when "01111000000010", -- t[7682] = 4
      "0100" when "01111000000011", -- t[7683] = 4
      "0100" when "01111000000100", -- t[7684] = 4
      "0100" when "01111000000101", -- t[7685] = 4
      "0100" when "01111000000110", -- t[7686] = 4
      "0100" when "01111000000111", -- t[7687] = 4
      "0100" when "01111000001000", -- t[7688] = 4
      "0100" when "01111000001001", -- t[7689] = 4
      "0100" when "01111000001010", -- t[7690] = 4
      "0100" when "01111000001011", -- t[7691] = 4
      "0100" when "01111000001100", -- t[7692] = 4
      "0100" when "01111000001101", -- t[7693] = 4
      "0100" when "01111000001110", -- t[7694] = 4
      "0100" when "01111000001111", -- t[7695] = 4
      "0100" when "01111000010000", -- t[7696] = 4
      "0100" when "01111000010001", -- t[7697] = 4
      "0100" when "01111000010010", -- t[7698] = 4
      "0100" when "01111000010011", -- t[7699] = 4
      "0100" when "01111000010100", -- t[7700] = 4
      "0100" when "01111000010101", -- t[7701] = 4
      "0100" when "01111000010110", -- t[7702] = 4
      "0100" when "01111000010111", -- t[7703] = 4
      "0100" when "01111000011000", -- t[7704] = 4
      "0100" when "01111000011001", -- t[7705] = 4
      "0100" when "01111000011010", -- t[7706] = 4
      "0100" when "01111000011011", -- t[7707] = 4
      "0100" when "01111000011100", -- t[7708] = 4
      "0100" when "01111000011101", -- t[7709] = 4
      "0100" when "01111000011110", -- t[7710] = 4
      "0100" when "01111000011111", -- t[7711] = 4
      "0100" when "01111000100000", -- t[7712] = 4
      "0100" when "01111000100001", -- t[7713] = 4
      "0100" when "01111000100010", -- t[7714] = 4
      "0100" when "01111000100011", -- t[7715] = 4
      "0100" when "01111000100100", -- t[7716] = 4
      "0100" when "01111000100101", -- t[7717] = 4
      "0100" when "01111000100110", -- t[7718] = 4
      "0100" when "01111000100111", -- t[7719] = 4
      "0100" when "01111000101000", -- t[7720] = 4
      "0100" when "01111000101001", -- t[7721] = 4
      "0100" when "01111000101010", -- t[7722] = 4
      "0100" when "01111000101011", -- t[7723] = 4
      "0100" when "01111000101100", -- t[7724] = 4
      "0100" when "01111000101101", -- t[7725] = 4
      "0100" when "01111000101110", -- t[7726] = 4
      "0100" when "01111000101111", -- t[7727] = 4
      "0100" when "01111000110000", -- t[7728] = 4
      "0100" when "01111000110001", -- t[7729] = 4
      "0100" when "01111000110010", -- t[7730] = 4
      "0100" when "01111000110011", -- t[7731] = 4
      "0100" when "01111000110100", -- t[7732] = 4
      "0100" when "01111000110101", -- t[7733] = 4
      "0100" when "01111000110110", -- t[7734] = 4
      "0100" when "01111000110111", -- t[7735] = 4
      "0100" when "01111000111000", -- t[7736] = 4
      "0100" when "01111000111001", -- t[7737] = 4
      "0100" when "01111000111010", -- t[7738] = 4
      "0100" when "01111000111011", -- t[7739] = 4
      "0100" when "01111000111100", -- t[7740] = 4
      "0100" when "01111000111101", -- t[7741] = 4
      "0100" when "01111000111110", -- t[7742] = 4
      "0100" when "01111000111111", -- t[7743] = 4
      "0100" when "01111001000000", -- t[7744] = 4
      "0100" when "01111001000001", -- t[7745] = 4
      "0100" when "01111001000010", -- t[7746] = 4
      "0100" when "01111001000011", -- t[7747] = 4
      "0100" when "01111001000100", -- t[7748] = 4
      "0100" when "01111001000101", -- t[7749] = 4
      "0100" when "01111001000110", -- t[7750] = 4
      "0100" when "01111001000111", -- t[7751] = 4
      "0100" when "01111001001000", -- t[7752] = 4
      "0100" when "01111001001001", -- t[7753] = 4
      "0100" when "01111001001010", -- t[7754] = 4
      "0100" when "01111001001011", -- t[7755] = 4
      "0100" when "01111001001100", -- t[7756] = 4
      "0100" when "01111001001101", -- t[7757] = 4
      "0100" when "01111001001110", -- t[7758] = 4
      "0100" when "01111001001111", -- t[7759] = 4
      "0100" when "01111001010000", -- t[7760] = 4
      "0100" when "01111001010001", -- t[7761] = 4
      "0100" when "01111001010010", -- t[7762] = 4
      "0100" when "01111001010011", -- t[7763] = 4
      "0100" when "01111001010100", -- t[7764] = 4
      "0100" when "01111001010101", -- t[7765] = 4
      "0100" when "01111001010110", -- t[7766] = 4
      "0100" when "01111001010111", -- t[7767] = 4
      "0100" when "01111001011000", -- t[7768] = 4
      "0100" when "01111001011001", -- t[7769] = 4
      "0100" when "01111001011010", -- t[7770] = 4
      "0100" when "01111001011011", -- t[7771] = 4
      "0100" when "01111001011100", -- t[7772] = 4
      "0100" when "01111001011101", -- t[7773] = 4
      "0100" when "01111001011110", -- t[7774] = 4
      "0100" when "01111001011111", -- t[7775] = 4
      "0100" when "01111001100000", -- t[7776] = 4
      "0100" when "01111001100001", -- t[7777] = 4
      "0100" when "01111001100010", -- t[7778] = 4
      "0100" when "01111001100011", -- t[7779] = 4
      "0100" when "01111001100100", -- t[7780] = 4
      "0100" when "01111001100101", -- t[7781] = 4
      "0100" when "01111001100110", -- t[7782] = 4
      "0100" when "01111001100111", -- t[7783] = 4
      "0100" when "01111001101000", -- t[7784] = 4
      "0100" when "01111001101001", -- t[7785] = 4
      "0100" when "01111001101010", -- t[7786] = 4
      "0100" when "01111001101011", -- t[7787] = 4
      "0100" when "01111001101100", -- t[7788] = 4
      "0100" when "01111001101101", -- t[7789] = 4
      "0100" when "01111001101110", -- t[7790] = 4
      "0100" when "01111001101111", -- t[7791] = 4
      "0100" when "01111001110000", -- t[7792] = 4
      "0100" when "01111001110001", -- t[7793] = 4
      "0100" when "01111001110010", -- t[7794] = 4
      "0100" when "01111001110011", -- t[7795] = 4
      "0100" when "01111001110100", -- t[7796] = 4
      "0100" when "01111001110101", -- t[7797] = 4
      "0100" when "01111001110110", -- t[7798] = 4
      "0100" when "01111001110111", -- t[7799] = 4
      "0100" when "01111001111000", -- t[7800] = 4
      "0100" when "01111001111001", -- t[7801] = 4
      "0100" when "01111001111010", -- t[7802] = 4
      "0100" when "01111001111011", -- t[7803] = 4
      "0100" when "01111001111100", -- t[7804] = 4
      "0100" when "01111001111101", -- t[7805] = 4
      "0100" when "01111001111110", -- t[7806] = 4
      "0100" when "01111001111111", -- t[7807] = 4
      "0100" when "01111010000000", -- t[7808] = 4
      "0100" when "01111010000001", -- t[7809] = 4
      "0100" when "01111010000010", -- t[7810] = 4
      "0100" when "01111010000011", -- t[7811] = 4
      "0100" when "01111010000100", -- t[7812] = 4
      "0100" when "01111010000101", -- t[7813] = 4
      "0100" when "01111010000110", -- t[7814] = 4
      "0100" when "01111010000111", -- t[7815] = 4
      "0100" when "01111010001000", -- t[7816] = 4
      "0100" when "01111010001001", -- t[7817] = 4
      "0100" when "01111010001010", -- t[7818] = 4
      "0100" when "01111010001011", -- t[7819] = 4
      "0100" when "01111010001100", -- t[7820] = 4
      "0100" when "01111010001101", -- t[7821] = 4
      "0100" when "01111010001110", -- t[7822] = 4
      "0101" when "01111010001111", -- t[7823] = 5
      "0101" when "01111010010000", -- t[7824] = 5
      "0101" when "01111010010001", -- t[7825] = 5
      "0101" when "01111010010010", -- t[7826] = 5
      "0101" when "01111010010011", -- t[7827] = 5
      "0101" when "01111010010100", -- t[7828] = 5
      "0101" when "01111010010101", -- t[7829] = 5
      "0101" when "01111010010110", -- t[7830] = 5
      "0101" when "01111010010111", -- t[7831] = 5
      "0101" when "01111010011000", -- t[7832] = 5
      "0101" when "01111010011001", -- t[7833] = 5
      "0101" when "01111010011010", -- t[7834] = 5
      "0101" when "01111010011011", -- t[7835] = 5
      "0101" when "01111010011100", -- t[7836] = 5
      "0101" when "01111010011101", -- t[7837] = 5
      "0101" when "01111010011110", -- t[7838] = 5
      "0101" when "01111010011111", -- t[7839] = 5
      "0101" when "01111010100000", -- t[7840] = 5
      "0101" when "01111010100001", -- t[7841] = 5
      "0101" when "01111010100010", -- t[7842] = 5
      "0101" when "01111010100011", -- t[7843] = 5
      "0101" when "01111010100100", -- t[7844] = 5
      "0101" when "01111010100101", -- t[7845] = 5
      "0101" when "01111010100110", -- t[7846] = 5
      "0101" when "01111010100111", -- t[7847] = 5
      "0101" when "01111010101000", -- t[7848] = 5
      "0101" when "01111010101001", -- t[7849] = 5
      "0101" when "01111010101010", -- t[7850] = 5
      "0101" when "01111010101011", -- t[7851] = 5
      "0101" when "01111010101100", -- t[7852] = 5
      "0101" when "01111010101101", -- t[7853] = 5
      "0101" when "01111010101110", -- t[7854] = 5
      "0101" when "01111010101111", -- t[7855] = 5
      "0101" when "01111010110000", -- t[7856] = 5
      "0101" when "01111010110001", -- t[7857] = 5
      "0101" when "01111010110010", -- t[7858] = 5
      "0101" when "01111010110011", -- t[7859] = 5
      "0101" when "01111010110100", -- t[7860] = 5
      "0101" when "01111010110101", -- t[7861] = 5
      "0101" when "01111010110110", -- t[7862] = 5
      "0101" when "01111010110111", -- t[7863] = 5
      "0101" when "01111010111000", -- t[7864] = 5
      "0101" when "01111010111001", -- t[7865] = 5
      "0101" when "01111010111010", -- t[7866] = 5
      "0101" when "01111010111011", -- t[7867] = 5
      "0101" when "01111010111100", -- t[7868] = 5
      "0101" when "01111010111101", -- t[7869] = 5
      "0101" when "01111010111110", -- t[7870] = 5
      "0101" when "01111010111111", -- t[7871] = 5
      "0101" when "01111011000000", -- t[7872] = 5
      "0101" when "01111011000001", -- t[7873] = 5
      "0101" when "01111011000010", -- t[7874] = 5
      "0101" when "01111011000011", -- t[7875] = 5
      "0101" when "01111011000100", -- t[7876] = 5
      "0101" when "01111011000101", -- t[7877] = 5
      "0101" when "01111011000110", -- t[7878] = 5
      "0101" when "01111011000111", -- t[7879] = 5
      "0101" when "01111011001000", -- t[7880] = 5
      "0101" when "01111011001001", -- t[7881] = 5
      "0101" when "01111011001010", -- t[7882] = 5
      "0101" when "01111011001011", -- t[7883] = 5
      "0101" when "01111011001100", -- t[7884] = 5
      "0101" when "01111011001101", -- t[7885] = 5
      "0101" when "01111011001110", -- t[7886] = 5
      "0101" when "01111011001111", -- t[7887] = 5
      "0101" when "01111011010000", -- t[7888] = 5
      "0101" when "01111011010001", -- t[7889] = 5
      "0101" when "01111011010010", -- t[7890] = 5
      "0101" when "01111011010011", -- t[7891] = 5
      "0101" when "01111011010100", -- t[7892] = 5
      "0101" when "01111011010101", -- t[7893] = 5
      "0101" when "01111011010110", -- t[7894] = 5
      "0101" when "01111011010111", -- t[7895] = 5
      "0101" when "01111011011000", -- t[7896] = 5
      "0101" when "01111011011001", -- t[7897] = 5
      "0101" when "01111011011010", -- t[7898] = 5
      "0101" when "01111011011011", -- t[7899] = 5
      "0101" when "01111011011100", -- t[7900] = 5
      "0101" when "01111011011101", -- t[7901] = 5
      "0101" when "01111011011110", -- t[7902] = 5
      "0101" when "01111011011111", -- t[7903] = 5
      "0101" when "01111011100000", -- t[7904] = 5
      "0101" when "01111011100001", -- t[7905] = 5
      "0101" when "01111011100010", -- t[7906] = 5
      "0101" when "01111011100011", -- t[7907] = 5
      "0101" when "01111011100100", -- t[7908] = 5
      "0101" when "01111011100101", -- t[7909] = 5
      "0101" when "01111011100110", -- t[7910] = 5
      "0101" when "01111011100111", -- t[7911] = 5
      "0101" when "01111011101000", -- t[7912] = 5
      "0101" when "01111011101001", -- t[7913] = 5
      "0101" when "01111011101010", -- t[7914] = 5
      "0101" when "01111011101011", -- t[7915] = 5
      "0101" when "01111011101100", -- t[7916] = 5
      "0101" when "01111011101101", -- t[7917] = 5
      "0101" when "01111011101110", -- t[7918] = 5
      "0101" when "01111011101111", -- t[7919] = 5
      "0101" when "01111011110000", -- t[7920] = 5
      "0101" when "01111011110001", -- t[7921] = 5
      "0101" when "01111011110010", -- t[7922] = 5
      "0101" when "01111011110011", -- t[7923] = 5
      "0101" when "01111011110100", -- t[7924] = 5
      "0101" when "01111011110101", -- t[7925] = 5
      "0101" when "01111011110110", -- t[7926] = 5
      "0101" when "01111011110111", -- t[7927] = 5
      "0101" when "01111011111000", -- t[7928] = 5
      "0101" when "01111011111001", -- t[7929] = 5
      "0101" when "01111011111010", -- t[7930] = 5
      "0101" when "01111011111011", -- t[7931] = 5
      "0101" when "01111011111100", -- t[7932] = 5
      "0101" when "01111011111101", -- t[7933] = 5
      "0101" when "01111011111110", -- t[7934] = 5
      "0101" when "01111011111111", -- t[7935] = 5
      "0101" when "01111100000000", -- t[7936] = 5
      "0101" when "01111100000001", -- t[7937] = 5
      "0101" when "01111100000010", -- t[7938] = 5
      "0101" when "01111100000011", -- t[7939] = 5
      "0101" when "01111100000100", -- t[7940] = 5
      "0101" when "01111100000101", -- t[7941] = 5
      "0101" when "01111100000110", -- t[7942] = 5
      "0101" when "01111100000111", -- t[7943] = 5
      "0101" when "01111100001000", -- t[7944] = 5
      "0101" when "01111100001001", -- t[7945] = 5
      "0101" when "01111100001010", -- t[7946] = 5
      "0101" when "01111100001011", -- t[7947] = 5
      "0101" when "01111100001100", -- t[7948] = 5
      "0101" when "01111100001101", -- t[7949] = 5
      "0101" when "01111100001110", -- t[7950] = 5
      "0101" when "01111100001111", -- t[7951] = 5
      "0101" when "01111100010000", -- t[7952] = 5
      "0101" when "01111100010001", -- t[7953] = 5
      "0101" when "01111100010010", -- t[7954] = 5
      "0101" when "01111100010011", -- t[7955] = 5
      "0101" when "01111100010100", -- t[7956] = 5
      "0101" when "01111100010101", -- t[7957] = 5
      "0101" when "01111100010110", -- t[7958] = 5
      "0101" when "01111100010111", -- t[7959] = 5
      "0101" when "01111100011000", -- t[7960] = 5
      "0101" when "01111100011001", -- t[7961] = 5
      "0101" when "01111100011010", -- t[7962] = 5
      "0101" when "01111100011011", -- t[7963] = 5
      "0101" when "01111100011100", -- t[7964] = 5
      "0101" when "01111100011101", -- t[7965] = 5
      "0101" when "01111100011110", -- t[7966] = 5
      "0101" when "01111100011111", -- t[7967] = 5
      "0101" when "01111100100000", -- t[7968] = 5
      "0101" when "01111100100001", -- t[7969] = 5
      "0101" when "01111100100010", -- t[7970] = 5
      "0101" when "01111100100011", -- t[7971] = 5
      "0101" when "01111100100100", -- t[7972] = 5
      "0101" when "01111100100101", -- t[7973] = 5
      "0101" when "01111100100110", -- t[7974] = 5
      "0101" when "01111100100111", -- t[7975] = 5
      "0101" when "01111100101000", -- t[7976] = 5
      "0101" when "01111100101001", -- t[7977] = 5
      "0101" when "01111100101010", -- t[7978] = 5
      "0101" when "01111100101011", -- t[7979] = 5
      "0101" when "01111100101100", -- t[7980] = 5
      "0101" when "01111100101101", -- t[7981] = 5
      "0101" when "01111100101110", -- t[7982] = 5
      "0101" when "01111100101111", -- t[7983] = 5
      "0101" when "01111100110000", -- t[7984] = 5
      "0101" when "01111100110001", -- t[7985] = 5
      "0101" when "01111100110010", -- t[7986] = 5
      "0101" when "01111100110011", -- t[7987] = 5
      "0101" when "01111100110100", -- t[7988] = 5
      "0101" when "01111100110101", -- t[7989] = 5
      "0101" when "01111100110110", -- t[7990] = 5
      "0101" when "01111100110111", -- t[7991] = 5
      "0101" when "01111100111000", -- t[7992] = 5
      "0101" when "01111100111001", -- t[7993] = 5
      "0101" when "01111100111010", -- t[7994] = 5
      "0101" when "01111100111011", -- t[7995] = 5
      "0101" when "01111100111100", -- t[7996] = 5
      "0101" when "01111100111101", -- t[7997] = 5
      "0101" when "01111100111110", -- t[7998] = 5
      "0101" when "01111100111111", -- t[7999] = 5
      "0101" when "01111101000000", -- t[8000] = 5
      "0101" when "01111101000001", -- t[8001] = 5
      "0101" when "01111101000010", -- t[8002] = 5
      "0101" when "01111101000011", -- t[8003] = 5
      "0101" when "01111101000100", -- t[8004] = 5
      "0101" when "01111101000101", -- t[8005] = 5
      "0101" when "01111101000110", -- t[8006] = 5
      "0101" when "01111101000111", -- t[8007] = 5
      "0101" when "01111101001000", -- t[8008] = 5
      "0101" when "01111101001001", -- t[8009] = 5
      "0101" when "01111101001010", -- t[8010] = 5
      "0101" when "01111101001011", -- t[8011] = 5
      "0101" when "01111101001100", -- t[8012] = 5
      "0101" when "01111101001101", -- t[8013] = 5
      "0101" when "01111101001110", -- t[8014] = 5
      "0101" when "01111101001111", -- t[8015] = 5
      "0101" when "01111101010000", -- t[8016] = 5
      "0101" when "01111101010001", -- t[8017] = 5
      "0101" when "01111101010010", -- t[8018] = 5
      "0101" when "01111101010011", -- t[8019] = 5
      "0101" when "01111101010100", -- t[8020] = 5
      "0101" when "01111101010101", -- t[8021] = 5
      "0101" when "01111101010110", -- t[8022] = 5
      "0101" when "01111101010111", -- t[8023] = 5
      "0101" when "01111101011000", -- t[8024] = 5
      "0101" when "01111101011001", -- t[8025] = 5
      "0101" when "01111101011010", -- t[8026] = 5
      "0101" when "01111101011011", -- t[8027] = 5
      "0101" when "01111101011100", -- t[8028] = 5
      "0101" when "01111101011101", -- t[8029] = 5
      "0101" when "01111101011110", -- t[8030] = 5
      "0101" when "01111101011111", -- t[8031] = 5
      "0101" when "01111101100000", -- t[8032] = 5
      "0101" when "01111101100001", -- t[8033] = 5
      "0101" when "01111101100010", -- t[8034] = 5
      "0101" when "01111101100011", -- t[8035] = 5
      "0101" when "01111101100100", -- t[8036] = 5
      "0101" when "01111101100101", -- t[8037] = 5
      "0101" when "01111101100110", -- t[8038] = 5
      "0101" when "01111101100111", -- t[8039] = 5
      "0101" when "01111101101000", -- t[8040] = 5
      "0101" when "01111101101001", -- t[8041] = 5
      "0101" when "01111101101010", -- t[8042] = 5
      "0101" when "01111101101011", -- t[8043] = 5
      "0101" when "01111101101100", -- t[8044] = 5
      "0101" when "01111101101101", -- t[8045] = 5
      "0101" when "01111101101110", -- t[8046] = 5
      "0101" when "01111101101111", -- t[8047] = 5
      "0101" when "01111101110000", -- t[8048] = 5
      "0101" when "01111101110001", -- t[8049] = 5
      "0101" when "01111101110010", -- t[8050] = 5
      "0101" when "01111101110011", -- t[8051] = 5
      "0101" when "01111101110100", -- t[8052] = 5
      "0101" when "01111101110101", -- t[8053] = 5
      "0101" when "01111101110110", -- t[8054] = 5
      "0101" when "01111101110111", -- t[8055] = 5
      "0101" when "01111101111000", -- t[8056] = 5
      "0101" when "01111101111001", -- t[8057] = 5
      "0101" when "01111101111010", -- t[8058] = 5
      "0101" when "01111101111011", -- t[8059] = 5
      "0101" when "01111101111100", -- t[8060] = 5
      "0101" when "01111101111101", -- t[8061] = 5
      "0101" when "01111101111110", -- t[8062] = 5
      "0101" when "01111101111111", -- t[8063] = 5
      "0101" when "01111110000000", -- t[8064] = 5
      "0101" when "01111110000001", -- t[8065] = 5
      "0101" when "01111110000010", -- t[8066] = 5
      "0101" when "01111110000011", -- t[8067] = 5
      "0101" when "01111110000100", -- t[8068] = 5
      "0101" when "01111110000101", -- t[8069] = 5
      "0101" when "01111110000110", -- t[8070] = 5
      "0101" when "01111110000111", -- t[8071] = 5
      "0101" when "01111110001000", -- t[8072] = 5
      "0101" when "01111110001001", -- t[8073] = 5
      "0101" when "01111110001010", -- t[8074] = 5
      "0101" when "01111110001011", -- t[8075] = 5
      "0101" when "01111110001100", -- t[8076] = 5
      "0101" when "01111110001101", -- t[8077] = 5
      "0101" when "01111110001110", -- t[8078] = 5
      "0101" when "01111110001111", -- t[8079] = 5
      "0101" when "01111110010000", -- t[8080] = 5
      "0101" when "01111110010001", -- t[8081] = 5
      "0101" when "01111110010010", -- t[8082] = 5
      "0101" when "01111110010011", -- t[8083] = 5
      "0101" when "01111110010100", -- t[8084] = 5
      "0101" when "01111110010101", -- t[8085] = 5
      "0101" when "01111110010110", -- t[8086] = 5
      "0101" when "01111110010111", -- t[8087] = 5
      "0101" when "01111110011000", -- t[8088] = 5
      "0101" when "01111110011001", -- t[8089] = 5
      "0101" when "01111110011010", -- t[8090] = 5
      "0101" when "01111110011011", -- t[8091] = 5
      "0101" when "01111110011100", -- t[8092] = 5
      "0101" when "01111110011101", -- t[8093] = 5
      "0101" when "01111110011110", -- t[8094] = 5
      "0101" when "01111110011111", -- t[8095] = 5
      "0101" when "01111110100000", -- t[8096] = 5
      "0101" when "01111110100001", -- t[8097] = 5
      "0101" when "01111110100010", -- t[8098] = 5
      "0101" when "01111110100011", -- t[8099] = 5
      "0101" when "01111110100100", -- t[8100] = 5
      "0101" when "01111110100101", -- t[8101] = 5
      "0101" when "01111110100110", -- t[8102] = 5
      "0101" when "01111110100111", -- t[8103] = 5
      "0101" when "01111110101000", -- t[8104] = 5
      "0101" when "01111110101001", -- t[8105] = 5
      "0101" when "01111110101010", -- t[8106] = 5
      "0101" when "01111110101011", -- t[8107] = 5
      "0101" when "01111110101100", -- t[8108] = 5
      "0101" when "01111110101101", -- t[8109] = 5
      "0101" when "01111110101110", -- t[8110] = 5
      "0101" when "01111110101111", -- t[8111] = 5
      "0101" when "01111110110000", -- t[8112] = 5
      "0101" when "01111110110001", -- t[8113] = 5
      "0101" when "01111110110010", -- t[8114] = 5
      "0101" when "01111110110011", -- t[8115] = 5
      "0101" when "01111110110100", -- t[8116] = 5
      "0101" when "01111110110101", -- t[8117] = 5
      "0101" when "01111110110110", -- t[8118] = 5
      "0110" when "01111110110111", -- t[8119] = 6
      "0110" when "01111110111000", -- t[8120] = 6
      "0110" when "01111110111001", -- t[8121] = 6
      "0110" when "01111110111010", -- t[8122] = 6
      "0110" when "01111110111011", -- t[8123] = 6
      "0110" when "01111110111100", -- t[8124] = 6
      "0110" when "01111110111101", -- t[8125] = 6
      "0110" when "01111110111110", -- t[8126] = 6
      "0110" when "01111110111111", -- t[8127] = 6
      "0110" when "01111111000000", -- t[8128] = 6
      "0110" when "01111111000001", -- t[8129] = 6
      "0110" when "01111111000010", -- t[8130] = 6
      "0110" when "01111111000011", -- t[8131] = 6
      "0110" when "01111111000100", -- t[8132] = 6
      "0110" when "01111111000101", -- t[8133] = 6
      "0110" when "01111111000110", -- t[8134] = 6
      "0110" when "01111111000111", -- t[8135] = 6
      "0110" when "01111111001000", -- t[8136] = 6
      "0110" when "01111111001001", -- t[8137] = 6
      "0110" when "01111111001010", -- t[8138] = 6
      "0110" when "01111111001011", -- t[8139] = 6
      "0110" when "01111111001100", -- t[8140] = 6
      "0110" when "01111111001101", -- t[8141] = 6
      "0110" when "01111111001110", -- t[8142] = 6
      "0110" when "01111111001111", -- t[8143] = 6
      "0110" when "01111111010000", -- t[8144] = 6
      "0110" when "01111111010001", -- t[8145] = 6
      "0110" when "01111111010010", -- t[8146] = 6
      "0110" when "01111111010011", -- t[8147] = 6
      "0110" when "01111111010100", -- t[8148] = 6
      "0110" when "01111111010101", -- t[8149] = 6
      "0110" when "01111111010110", -- t[8150] = 6
      "0110" when "01111111010111", -- t[8151] = 6
      "0110" when "01111111011000", -- t[8152] = 6
      "0110" when "01111111011001", -- t[8153] = 6
      "0110" when "01111111011010", -- t[8154] = 6
      "0110" when "01111111011011", -- t[8155] = 6
      "0110" when "01111111011100", -- t[8156] = 6
      "0110" when "01111111011101", -- t[8157] = 6
      "0110" when "01111111011110", -- t[8158] = 6
      "0110" when "01111111011111", -- t[8159] = 6
      "0110" when "01111111100000", -- t[8160] = 6
      "0110" when "01111111100001", -- t[8161] = 6
      "0110" when "01111111100010", -- t[8162] = 6
      "0110" when "01111111100011", -- t[8163] = 6
      "0110" when "01111111100100", -- t[8164] = 6
      "0110" when "01111111100101", -- t[8165] = 6
      "0110" when "01111111100110", -- t[8166] = 6
      "0110" when "01111111100111", -- t[8167] = 6
      "0110" when "01111111101000", -- t[8168] = 6
      "0110" when "01111111101001", -- t[8169] = 6
      "0110" when "01111111101010", -- t[8170] = 6
      "0110" when "01111111101011", -- t[8171] = 6
      "0110" when "01111111101100", -- t[8172] = 6
      "0110" when "01111111101101", -- t[8173] = 6
      "0110" when "01111111101110", -- t[8174] = 6
      "0110" when "01111111101111", -- t[8175] = 6
      "0110" when "01111111110000", -- t[8176] = 6
      "0110" when "01111111110001", -- t[8177] = 6
      "0110" when "01111111110010", -- t[8178] = 6
      "0110" when "01111111110011", -- t[8179] = 6
      "0110" when "01111111110100", -- t[8180] = 6
      "0110" when "01111111110101", -- t[8181] = 6
      "0110" when "01111111110110", -- t[8182] = 6
      "0110" when "01111111110111", -- t[8183] = 6
      "0110" when "01111111111000", -- t[8184] = 6
      "0110" when "01111111111001", -- t[8185] = 6
      "0110" when "01111111111010", -- t[8186] = 6
      "0110" when "01111111111011", -- t[8187] = 6
      "0110" when "01111111111100", -- t[8188] = 6
      "0110" when "01111111111101", -- t[8189] = 6
      "0110" when "01111111111110", -- t[8190] = 6
      "0110" when "01111111111111", -- t[8191] = 6
      "----" when others;
end architecture;


-- Minimax-Defour: LNS subtraction function [ -8.000000, -4.000000 [ -> [ 0.000000, 0.125000 [
-- Input:  wE =   2, wF =  10, w =  12
-- Output: wE =  -3, wF =  10, w =   7
-- Decomposition: a  =  5, b  =  7
--                a0 =  5, b0 =  5, p0 =  5
--                a1 =  3, b1 =  2, p1 = 10
--                a2 =  3, b2 =  2, p2 =  5
--                g0 =  3, g1 =  -2
-- ROMs: 2^ 5 x 10  +  2^ 5 x  5  +  2^ 5 x  0  +  2^ 5 x  0  =     480 bits
-- Mult: 5 x 5 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T1_10 is
  component LNSSub_MNMX_T1_10_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_t2 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_t3 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T1_10_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_10_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_t0 is
begin
  with x select
    r <=
      "0000110011" when "00000", -- t[0] = 51
      "0000110110" when "00001", -- t[1] = 54
      "0000111100" when "00010", -- t[2] = 60
      "0001000010" when "00011", -- t[3] = 66
      "0001000110" when "00100", -- t[4] = 70
      "0001001100" when "00101", -- t[5] = 76
      "0001010010" when "00110", -- t[6] = 82
      "0001011001" when "00111", -- t[7] = 89
      "0001100001" when "01000", -- t[8] = 97
      "0001101010" when "01001", -- t[9] = 106
      "0001110010" when "01010", -- t[10] = 114
      "0001111100" when "01011", -- t[11] = 124
      "0010001000" when "01100", -- t[12] = 136
      "0010010100" when "01101", -- t[13] = 148
      "0010100000" when "01110", -- t[14] = 160
      "0010101111" when "01111", -- t[15] = 175
      "0010111111" when "10000", -- t[16] = 191
      "0011001111" when "10001", -- t[17] = 207
      "0011100010" when "10010", -- t[18] = 226
      "0011110101" when "10011", -- t[19] = 245
      "0100001101" when "10100", -- t[20] = 269
      "0100100100" when "10101", -- t[21] = 292
      "0100111111" when "10110", -- t[22] = 319
      "0101011100" when "10111", -- t[23] = 348
      "0101111011" when "11000", -- t[24] = 379
      "0110011111" when "11001", -- t[25] = 415
      "0111000101" when "11010", -- t[26] = 453
      "0111101110" when "11011", -- t[27] = 494
      "1000011011" when "11100", -- t[28] = 539
      "1001001100" when "11101", -- t[29] = 588
      "1010000011" when "11110", -- t[30] = 643
      "1010111111" when "11111", -- t[31] = 703
      "----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_10_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_t1 is
begin
  with x select
    r <=
      "00001" when "00000", -- t[0] = 1
      "00001" when "00001", -- t[1] = 1
      "00001" when "00010", -- t[2] = 1
      "00001" when "00011", -- t[3] = 1
      "00001" when "00100", -- t[4] = 1
      "00010" when "00101", -- t[5] = 2
      "00010" when "00110", -- t[6] = 2
      "00010" when "00111", -- t[7] = 2
      "00010" when "01000", -- t[8] = 2
      "00010" when "01001", -- t[9] = 2
      "00011" when "01010", -- t[10] = 3
      "00011" when "01011", -- t[11] = 3
      "00011" when "01100", -- t[12] = 3
      "00011" when "01101", -- t[13] = 3
      "00100" when "01110", -- t[14] = 4
      "00100" when "01111", -- t[15] = 4
      "00100" when "10000", -- t[16] = 4
      "00101" when "10001", -- t[17] = 5
      "00101" when "10010", -- t[18] = 5
      "00110" when "10011", -- t[19] = 6
      "00110" when "10100", -- t[20] = 6
      "00111" when "10101", -- t[21] = 7
      "00111" when "10110", -- t[22] = 7
      "01000" when "10111", -- t[23] = 8
      "01001" when "11000", -- t[24] = 9
      "01001" when "11001", -- t[25] = 9
      "01010" when "11010", -- t[26] = 10
      "01011" when "11011", -- t[27] = 11
      "01100" when "11100", -- t[28] = 12
      "01110" when "11101", -- t[29] = 14
      "01111" when "11110", -- t[30] = 15
      "10000" when "11111", -- t[31] = 16
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_10_t2 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_t2 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "0" when "1101", -- t[13] = 0
      "0" when "1110", -- t[14] = 0
      "0" when "1111", -- t[15] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T1_10_t3 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_t3 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "0" when "1101", -- t[13] = 0
      "0" when "1110", -- t[14] = 0
      "0" when "1111", -- t[15] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_10.all;

entity LNSSub_MNMX_T1_10_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_mult is
  signal out_t : std_logic_vector(4 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T1_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_10.all;

entity LNSSub_MNMX_T1_10_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T1_10_t2
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_10.all;

entity LNSSub_MNMX_T1_10_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T1_10_t3
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T1_10.all;

entity LNSSub_MNMX_T1_10 is
  port ( x : in  std_logic_vector(11 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T1_10 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(9 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(4 downto 0);
  signal r1  : std_logic_vector(9 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(9 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(9 downto 0);
  signal sum : std_logic_vector(9 downto 0);
begin
  a0 <= x(11 downto 7);
  inst_t0 : LNSSub_MNMX_T1_10_t0
    port map ( x => a0,
               r => r0(9 downto 0) );

  a1 <= x(11 downto 7);
  b1 <= x(6 downto 2);
  inst_mult : LNSSub_MNMX_T1_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(6 downto 0) );
  r1(9 downto 7) <= (9 downto 7 => '0');

  a2 <= x(11 downto 9);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T1_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(9 downto 0) );

  a3 <= x(11 downto 9);
  b3 <= x(6 downto 5);
  inst_xor3 : LNSSub_MNMX_T1_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(9 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(9 downto 3);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -4.000000, -2.000000 [ -> [ 0.000000, 0.500000 [
-- Input:  wE =   1, wF =  10, w =  11
-- Output: wE =  -1, wF =  10, w =   9
-- Decomposition: a  =  5, b  =  6
--                a0 =  5, b0 =  4, p0 =  5
--                a1 =  3, b1 =  2, p1 =  9
--                a2 =  3, b2 =  2, p2 =  5
--                g0 =  3, g1 =  -3
-- ROMs: 2^ 5 x 12  +  2^ 5 x  6  +  2^ 5 x  2  +  2^ 5 x  0  =     640 bits
-- Mult: 4 x 6 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T2_10 is
  component LNSSub_MNMX_T2_10_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_t2 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_t3 is
    port ( x : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MNMX_T2_10_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_10_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_t0 is
begin
  with x select
    r <=
      "001011111111" when "00000", -- t[0] = 767
      "001100100011" when "00001", -- t[1] = 803
      "001101000110" when "00010", -- t[2] = 838
      "001101101110" when "00011", -- t[3] = 878
      "001110010101" when "00100", -- t[4] = 917
      "001111000000" when "00101", -- t[5] = 960
      "001111101011" when "00110", -- t[6] = 1003
      "010000011010" when "00111", -- t[7] = 1050
      "010001001011" when "01000", -- t[8] = 1099
      "010001111110" when "01001", -- t[9] = 1150
      "010010110011" when "01010", -- t[10] = 1203
      "010011101011" when "01011", -- t[11] = 1259
      "010100100111" when "01100", -- t[12] = 1319
      "010101100100" when "01101", -- t[13] = 1380
      "010110100101" when "01110", -- t[14] = 1445
      "010111101000" when "01111", -- t[15] = 1512
      "011000110000" when "10000", -- t[16] = 1584
      "011001111010" when "10001", -- t[17] = 1658
      "011011001001" when "10010", -- t[18] = 1737
      "011100011101" when "10011", -- t[19] = 1821
      "011101110100" when "10100", -- t[20] = 1908
      "011111010000" when "10101", -- t[21] = 2000
      "100000110010" when "10110", -- t[22] = 2098
      "100010010110" when "10111", -- t[23] = 2198
      "100100000010" when "11000", -- t[24] = 2306
      "100101110010" when "11001", -- t[25] = 2418
      "100111101010" when "11010", -- t[26] = 2538
      "101001101000" when "11011", -- t[27] = 2664
      "101011101100" when "11100", -- t[28] = 2796
      "101101111000" when "11101", -- t[29] = 2936
      "110000001101" when "11110", -- t[30] = 3085
      "110010101010" when "11111", -- t[31] = 3242
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_10_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_t1 is
begin
  with x select
    r <=
      "001001" when "00000", -- t[0] = 9
      "001001" when "00001", -- t[1] = 9
      "001010" when "00010", -- t[2] = 10
      "001010" when "00011", -- t[3] = 10
      "001011" when "00100", -- t[4] = 11
      "001011" when "00101", -- t[5] = 11
      "001100" when "00110", -- t[6] = 12
      "001100" when "00111", -- t[7] = 12
      "001101" when "01000", -- t[8] = 13
      "001101" when "01001", -- t[9] = 13
      "001110" when "01010", -- t[10] = 14
      "001111" when "01011", -- t[11] = 15
      "001111" when "01100", -- t[12] = 15
      "010000" when "01101", -- t[13] = 16
      "010001" when "01110", -- t[14] = 17
      "010010" when "01111", -- t[15] = 18
      "010011" when "10000", -- t[16] = 19
      "010100" when "10001", -- t[17] = 20
      "010101" when "10010", -- t[18] = 21
      "010110" when "10011", -- t[19] = 22
      "010111" when "10100", -- t[20] = 23
      "011000" when "10101", -- t[21] = 24
      "011001" when "10110", -- t[22] = 25
      "011011" when "10111", -- t[23] = 27
      "011100" when "11000", -- t[24] = 28
      "011110" when "11001", -- t[25] = 30
      "011111" when "11010", -- t[26] = 31
      "100001" when "11011", -- t[27] = 33
      "100011" when "11100", -- t[28] = 35
      "100101" when "11101", -- t[29] = 37
      "100111" when "11110", -- t[30] = 39
      "101001" when "11111", -- t[31] = 41
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_10_t2 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_t2 is
begin
  with x select
    r <=
      "00" when "0000", -- t[0] = 0
      "00" when "0001", -- t[1] = 0
      "00" when "0010", -- t[2] = 0
      "01" when "0011", -- t[3] = 1
      "00" when "0100", -- t[4] = 0
      "01" when "0101", -- t[5] = 1
      "00" when "0110", -- t[6] = 0
      "01" when "0111", -- t[7] = 1
      "00" when "1000", -- t[8] = 0
      "01" when "1001", -- t[9] = 1
      "00" when "1010", -- t[10] = 0
      "10" when "1011", -- t[11] = 2
      "00" when "1100", -- t[12] = 0
      "10" when "1101", -- t[13] = 2
      "01" when "1110", -- t[14] = 1
      "11" when "1111", -- t[15] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T2_10_t3 is
  port ( x : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_t3 is
begin
  with x select
    r <=
      "0" when "0000", -- t[0] = 0
      "0" when "0001", -- t[1] = 0
      "0" when "0010", -- t[2] = 0
      "0" when "0011", -- t[3] = 0
      "0" when "0100", -- t[4] = 0
      "0" when "0101", -- t[5] = 0
      "0" when "0110", -- t[6] = 0
      "0" when "0111", -- t[7] = 0
      "0" when "1000", -- t[8] = 0
      "0" when "1001", -- t[9] = 0
      "0" when "1010", -- t[10] = 0
      "0" when "1011", -- t[11] = 0
      "0" when "1100", -- t[12] = 0
      "0" when "1101", -- t[13] = 0
      "0" when "1110", -- t[14] = 0
      "0" when "1111", -- t[15] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_10.all;

entity LNSSub_MNMX_T2_10_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_mult is
  signal out_t : std_logic_vector(5 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T2_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_10.all;

entity LNSSub_MNMX_T2_10_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T2_10_t2
    port map ( x => in_t,
               r => out_t );

  r(11 downto 2) <= (11 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_10.all;

entity LNSSub_MNMX_T2_10_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T2_10_t3
    port map ( x => in_t,
               r => out_t );

  r(11 downto 1) <= (11 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T2_10.all;

entity LNSSub_MNMX_T2_10 is
  port ( x : in  std_logic_vector(10 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T2_10 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(11 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(11 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(11 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(11 downto 0);
  signal sum : std_logic_vector(11 downto 0);
begin
  a0 <= x(10 downto 6);
  inst_t0 : LNSSub_MNMX_T2_10_t0
    port map ( x => a0,
               r => r0(11 downto 0) );

  a1 <= x(10 downto 6);
  b1 <= x(5 downto 2);
  inst_mult : LNSSub_MNMX_T2_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(11 downto 8) <= (11 downto 8 => '0');

  a2 <= x(10 downto 8);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T2_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(11 downto 0) );

  a3 <= x(10 downto 8);
  b3 <= x(5 downto 4);
  inst_xor3 : LNSSub_MNMX_T2_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(11 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(11 downto 3);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -2.000000, -1.000000 [ -> [ 0.000000, 1.000000 [
-- Input:  wE =   0, wF =  10, w =  10
-- Output: wE =   0, wF =  10, w =  10
-- Decomposition: a  =  5, b  =  5
--                a0 =  5, b0 =  4, p0 =  5
--                a1 =  3, b1 =  1, p1 =  9
--                a2 =  3, b2 =  1, p2 =  5
--                g0 =  3, g1 =  -4
-- ROMs: 2^ 5 x 13  +  2^ 5 x  6  +  2^ 4 x  2  +  2^ 4 x  0  =     640 bits
-- Mult: 4 x 6 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T3_10 is
  component LNSSub_MNMX_T3_10_t0 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_t1 is
    port ( x : in  std_logic_vector(4 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_t2 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_t3 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_mult is
    port ( a : in  std_logic_vector(4 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_xor2 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MNMX_T3_10_xor3 is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_10_t0 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_t0 is
begin
  with x select
    r <=
      "0110101001100" when "00000", -- t[0] = 3404
      "0110110100100" when "00001", -- t[1] = 3492
      "0110111111101" when "00010", -- t[2] = 3581
      "0111001011000" when "00011", -- t[3] = 3672
      "0111010111000" when "00100", -- t[4] = 3768
      "0111100011001" when "00101", -- t[5] = 3865
      "0111101111101" when "00110", -- t[6] = 3965
      "0111111100100" when "00111", -- t[7] = 4068
      "1000001010000" when "01000", -- t[8] = 4176
      "1000010111110" when "01001", -- t[9] = 4286
      "1000100110000" when "01010", -- t[10] = 4400
      "1000110100101" when "01011", -- t[11] = 4517
      "1001000011110" when "01100", -- t[12] = 4638
      "1001010011001" when "01101", -- t[13] = 4761
      "1001100011100" when "01110", -- t[14] = 4892
      "1001110100001" when "01111", -- t[15] = 5025
      "1010000101001" when "10000", -- t[16] = 5161
      "1010010111000" when "10001", -- t[17] = 5304
      "1010101001100" when "10010", -- t[18] = 5452
      "1010111100101" when "10011", -- t[19] = 5605
      "1011010000010" when "10100", -- t[20] = 5762
      "1011100100110" when "10101", -- t[21] = 5926
      "1011111001111" when "10110", -- t[22] = 6095
      "1100001111111" when "10111", -- t[23] = 6271
      "1100100110110" when "11000", -- t[24] = 6454
      "1100111110011" when "11001", -- t[25] = 6643
      "1101010111000" when "11010", -- t[26] = 6840
      "1101110000100" when "11011", -- t[27] = 7044
      "1110001011001" when "11100", -- t[28] = 7257
      "1110100110101" when "11101", -- t[29] = 7477
      "1111000011100" when "11110", -- t[30] = 7708
      "1111100001100" when "11111", -- t[31] = 7948
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_10_t1 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_t1 is
begin
  with x select
    r <=
      "010110" when "00000", -- t[0] = 22
      "010110" when "00001", -- t[1] = 22
      "010111" when "00010", -- t[2] = 23
      "011000" when "00011", -- t[3] = 24
      "011000" when "00100", -- t[4] = 24
      "011001" when "00101", -- t[5] = 25
      "011010" when "00110", -- t[6] = 26
      "011011" when "00111", -- t[7] = 27
      "011011" when "01000", -- t[8] = 27
      "011100" when "01001", -- t[9] = 28
      "011101" when "01010", -- t[10] = 29
      "011110" when "01011", -- t[11] = 30
      "011111" when "01100", -- t[12] = 31
      "100000" when "01101", -- t[13] = 32
      "100001" when "01110", -- t[14] = 33
      "100010" when "01111", -- t[15] = 34
      "100100" when "10000", -- t[16] = 36
      "100101" when "10001", -- t[17] = 37
      "100110" when "10010", -- t[18] = 38
      "100111" when "10011", -- t[19] = 39
      "101001" when "10100", -- t[20] = 41
      "101010" when "10101", -- t[21] = 42
      "101100" when "10110", -- t[22] = 44
      "101110" when "10111", -- t[23] = 46
      "101111" when "11000", -- t[24] = 47
      "110001" when "11001", -- t[25] = 49
      "110011" when "11010", -- t[26] = 51
      "110101" when "11011", -- t[27] = 53
      "110111" when "11100", -- t[28] = 55
      "111010" when "11101", -- t[29] = 58
      "111100" when "11110", -- t[30] = 60
      "111111" when "11111", -- t[31] = 63
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_10_t2 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_t2 is
begin
  with x select
    r <=
      "01" when "000", -- t[0] = 1
      "01" when "001", -- t[1] = 1
      "01" when "010", -- t[2] = 1
      "10" when "011", -- t[3] = 2
      "10" when "100", -- t[4] = 2
      "10" when "101", -- t[5] = 2
      "11" when "110", -- t[6] = 3
      "11" when "111", -- t[7] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T3_10_t3 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_t3 is
begin
  with x select
    r <=
      "0" when "000", -- t[0] = 0
      "0" when "001", -- t[1] = 0
      "0" when "010", -- t[2] = 0
      "0" when "011", -- t[3] = 0
      "0" when "100", -- t[4] = 0
      "0" when "101", -- t[5] = 0
      "0" when "110", -- t[6] = 0
      "0" when "111", -- t[7] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_10.all;

entity LNSSub_MNMX_T3_10_mult is
  port ( a : in  std_logic_vector(4 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_mult is
  signal out_t : std_logic_vector(5 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T3_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_10.all;

entity LNSSub_MNMX_T3_10_xor2 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(0);
  in_t(2 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T3_10_t2
    port map ( x => in_t,
               r => out_t );

  r(12 downto 2) <= (12 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_10.all;

entity LNSSub_MNMX_T3_10_xor3 is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(2 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T3_10_t3
    port map ( x => in_t,
               r => out_t );

  r(12 downto 1) <= (12 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T3_10.all;

entity LNSSub_MNMX_T3_10 is
  port ( x : in  std_logic_vector(9 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T3_10 is
  signal a0  : std_logic_vector(4 downto 0);
  signal r0  : std_logic_vector(12 downto 0);
  signal a1  : std_logic_vector(4 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(12 downto 0);
  signal a2  : std_logic_vector(2 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(12 downto 0);
  signal a3  : std_logic_vector(2 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(12 downto 0);
  signal sum : std_logic_vector(12 downto 0);
begin
  a0 <= x(9 downto 5);
  inst_t0 : LNSSub_MNMX_T3_10_t0
    port map ( x => a0,
               r => r0(12 downto 0) );

  a1 <= x(9 downto 5);
  b1 <= x(4 downto 1);
  inst_mult : LNSSub_MNMX_T3_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(12 downto 8) <= (12 downto 8 => '0');

  a2 <= x(9 downto 7);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T3_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(12 downto 0) );

  a3 <= x(9 downto 7);
  b3 <= x(4 downto 4);
  inst_xor3 : LNSSub_MNMX_T3_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(12 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(12 downto 3);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -1.000000, -0.500000 [ -> [ 0.000000, 2.000000 [
-- Input:  wE =  -1, wF =  10, w =   9
-- Output: wE =   1, wF =  10, w =  11
-- Decomposition: a  =  3, b  =  6
--                a0 =  3, b0 =  4, p0 =  3
--                a1 =  2, b1 =  2, p1 =  7
--                a2 =  2, b2 =  2, p2 =  3
--                g0 =  0, g1 =  -4
-- ROMs: 2^ 3 x 11  +  2^ 3 x  8  +  2^ 4 x  2  +  2^ 4 x  1  =     200 bits
-- Mult: 4 x 8 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T4_10 is
  component LNSSub_MNMX_T4_10_t0 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_t1 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_t2 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_t3 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_mult is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T4_10_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_10_t0 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_t0 is
begin
  with x select
    r <=
      "10000000010" when "000", -- t[0] = 1026
      "10001000101" when "001", -- t[1] = 1093
      "10010001110" when "010", -- t[2] = 1166
      "10011011111" when "011", -- t[3] = 1247
      "10100111001" when "100", -- t[4] = 1337
      "10110011100" when "101", -- t[5] = 1436
      "11000001010" when "110", -- t[6] = 1546
      "11010001000" when "111", -- t[7] = 1672
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_10_t1 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_t1 is
begin
  with x select
    r <=
      "01000011" when "000", -- t[0] = 67
      "01001001" when "001", -- t[1] = 73
      "01010001" when "010", -- t[2] = 81
      "01011001" when "011", -- t[3] = 89
      "01100011" when "100", -- t[4] = 99
      "01101111" when "101", -- t[5] = 111
      "01111110" when "110", -- t[6] = 126
      "10010000" when "111", -- t[7] = 144
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_10_t2 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_t2 is
begin
  with x select
    r <=
      "00" when "000", -- t[0] = 0
      "01" when "001", -- t[1] = 1
      "00" when "010", -- t[2] = 0
      "01" when "011", -- t[3] = 1
      "00" when "100", -- t[4] = 0
      "10" when "101", -- t[5] = 2
      "01" when "110", -- t[6] = 1
      "11" when "111", -- t[7] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T4_10_t3 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_t3 is
begin
  with x select
    r <=
      "0" when "000", -- t[0] = 0
      "0" when "001", -- t[1] = 0
      "0" when "010", -- t[2] = 0
      "0" when "011", -- t[3] = 0
      "0" when "100", -- t[4] = 0
      "0" when "101", -- t[5] = 0
      "0" when "110", -- t[6] = 0
      "1" when "111", -- t[7] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_10.all;

entity LNSSub_MNMX_T4_10_mult is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_mult is
  signal out_t : std_logic_vector(7 downto 0);
  signal r0    : std_logic_vector(11 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T4_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(11 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_10.all;

entity LNSSub_MNMX_T4_10_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T4_10_t2
    port map ( x => in_t,
               r => out_t );

  r(10 downto 2) <= (10 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_10.all;

entity LNSSub_MNMX_T4_10_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t3 : LNSSub_MNMX_T4_10_t3
    port map ( x => in_t,
               r => out_t );

  r(10 downto 1) <= (10 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T4_10.all;

entity LNSSub_MNMX_T4_10 is
  port ( x : in  std_logic_vector(8 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T4_10 is
  signal a0  : std_logic_vector(2 downto 0);
  signal r0  : std_logic_vector(10 downto 0);
  signal a1  : std_logic_vector(2 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(10 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(10 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(1 downto 0);
  signal r3  : std_logic_vector(10 downto 0);
  signal sum : std_logic_vector(10 downto 0);
begin
  a0 <= x(8 downto 6);
  inst_t0 : LNSSub_MNMX_T4_10_t0
    port map ( x => a0,
               r => r0(10 downto 0) );

  a1 <= x(8 downto 6);
  b1 <= x(5 downto 2);
  inst_mult : LNSSub_MNMX_T4_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(7 downto 0) );
  r1(10 downto 8) <= (10 downto 8 => '0');

  a2 <= x(8 downto 7);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T4_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(10 downto 0) );

  a3 <= x(8 downto 7);
  b3 <= x(5 downto 4);
  inst_xor3 : LNSSub_MNMX_T4_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(10 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(10 downto 0);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.500000, -0.250000 [ -> [ 0.000000, 4.000000 [
-- Input:  wE =  -2, wF =  10, w =   8
-- Output: wE =   2, wF =   8, w =  10
-- Decomposition: a  =  3, b  =  5
--                a0 =  3, b0 =  4, p0 =  3
--                a1 =  2, b1 =  1, p1 =  7
--                a2 =  2, b2 =  1, p2 =  3
--                g0 =  1, g1 =  -5
-- ROMs: 2^ 3 x 11  +  2^ 3 x  6  +  2^ 3 x  1  +  2^ 3 x  0  =     144 bits
-- Mult: 4 x 6 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T5_10 is
  component LNSSub_MNMX_T5_10_t0 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_t1 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_t2 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_t3 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_mult is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(3 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MNMX_T5_10_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_10_t0 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_t0 is
begin
  with x select
    r <=
      "01110001101" when "000", -- t[0] = 909
      "01110110101" when "001", -- t[1] = 949
      "01111100000" when "010", -- t[2] = 992
      "10000001111" when "011", -- t[3] = 1039
      "10001000011" when "100", -- t[4] = 1091
      "10001111100" when "101", -- t[5] = 1148
      "10010111010" when "110", -- t[6] = 1210
      "10100000000" when "111", -- t[7] = 1280
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_10_t1 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_t1 is
begin
  with x select
    r <=
      "010100" when "000", -- t[0] = 20
      "010110" when "001", -- t[1] = 22
      "011000" when "010", -- t[2] = 24
      "011010" when "011", -- t[3] = 26
      "011100" when "100", -- t[4] = 28
      "011111" when "101", -- t[5] = 31
      "100011" when "110", -- t[6] = 35
      "101000" when "111", -- t[7] = 40
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_10_t2 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_t2 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "0" when "01", -- t[1] = 0
      "0" when "10", -- t[2] = 0
      "1" when "11", -- t[3] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T5_10_t3 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_t3 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "0" when "01", -- t[1] = 0
      "0" when "10", -- t[2] = 0
      "0" when "11", -- t[3] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_10.all;

entity LNSSub_MNMX_T5_10_mult is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(3 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_mult is
  signal out_t : std_logic_vector(5 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T5_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_10.all;

entity LNSSub_MNMX_T5_10_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T5_10_t2
    port map ( x => in_t,
               r => out_t );

  r(10 downto 1) <= (10 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_10.all;

entity LNSSub_MNMX_T5_10_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T5_10_t3
    port map ( x => in_t,
               r => out_t );

  r(10 downto 1) <= (10 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T5_10.all;

entity LNSSub_MNMX_T5_10 is
  port ( x : in  std_logic_vector(7 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T5_10 is
  signal a0  : std_logic_vector(2 downto 0);
  signal r0  : std_logic_vector(10 downto 0);
  signal a1  : std_logic_vector(2 downto 0);
  signal b1  : std_logic_vector(3 downto 0);
  signal r1  : std_logic_vector(10 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(10 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(10 downto 0);
  signal sum : std_logic_vector(10 downto 0);
begin
  a0 <= x(7 downto 5);
  inst_t0 : LNSSub_MNMX_T5_10_t0
    port map ( x => a0,
               r => r0(10 downto 0) );

  a1 <= x(7 downto 5);
  b1 <= x(4 downto 1);
  inst_mult : LNSSub_MNMX_T5_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(6 downto 0) );
  r1(10 downto 7) <= (10 downto 7 => '0');

  a2 <= x(7 downto 6);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T5_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(10 downto 0) );

  a3 <= x(7 downto 6);
  b3 <= x(4 downto 4);
  inst_xor3 : LNSSub_MNMX_T5_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(10 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(10 downto 1);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.250000, -0.125000 [ -> [ 0.000000, 4.000000 [
-- Input:  wE =  -3, wF =  10, w =   7
-- Output: wE =   2, wF =   7, w =   9
-- Decomposition: a  =  3, b  =  4
--                a0 =  3, b0 =  3, p0 =  3
--                a1 =  2, b1 =  1, p1 =  6
--                a2 =  2, b2 =  1, p2 =  3
--                g0 =  1, g1 =  -4
-- ROMs: 2^ 3 x 10  +  2^ 3 x  7  +  2^ 3 x  1  +  2^ 3 x  0  =     144 bits
-- Mult: 3 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T6_10 is
  component LNSSub_MNMX_T6_10_t0 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_t1 is
    port ( x : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_t2 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_t3 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_mult is
    port ( a : in  std_logic_vector(2 downto 0);
           b : in  std_logic_vector(2 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_xor2 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T6_10_xor3 is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_10_t0 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_t0 is
begin
  with x select
    r <=
      "1010101001" when "000", -- t[0] = 681
      "1010111111" when "001", -- t[1] = 703
      "1011010110" when "010", -- t[2] = 726
      "1011110000" when "011", -- t[3] = 752
      "1100001100" when "100", -- t[4] = 780
      "1100101010" when "101", -- t[5] = 810
      "1101001011" when "110", -- t[6] = 843
      "1101110000" when "111", -- t[7] = 880
      "----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_10_t1 is
  port ( x : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_t1 is
begin
  with x select
    r <=
      "0101100" when "000", -- t[0] = 44
      "0101111" when "001", -- t[1] = 47
      "0110011" when "010", -- t[2] = 51
      "0110111" when "011", -- t[3] = 55
      "0111100" when "100", -- t[4] = 60
      "1000010" when "101", -- t[5] = 66
      "1001010" when "110", -- t[6] = 74
      "1010011" when "111", -- t[7] = 83
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_10_t2 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_t2 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "0" when "01", -- t[1] = 0
      "0" when "10", -- t[2] = 0
      "1" when "11", -- t[3] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T6_10_t3 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_t3 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "0" when "01", -- t[1] = 0
      "0" when "10", -- t[2] = 0
      "0" when "11", -- t[3] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_10.all;

entity LNSSub_MNMX_T6_10_mult is
  port ( a : in  std_logic_vector(2 downto 0);
         b : in  std_logic_vector(2 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(9 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T6_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(9 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_10.all;

entity LNSSub_MNMX_T6_10_xor2 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T6_10_t2
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_10.all;

entity LNSSub_MNMX_T6_10_xor3 is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(1 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T6_10_t3
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T6_10.all;

entity LNSSub_MNMX_T6_10 is
  port ( x : in  std_logic_vector(6 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T6_10 is
  signal a0  : std_logic_vector(2 downto 0);
  signal r0  : std_logic_vector(9 downto 0);
  signal a1  : std_logic_vector(2 downto 0);
  signal b1  : std_logic_vector(2 downto 0);
  signal r1  : std_logic_vector(9 downto 0);
  signal a2  : std_logic_vector(1 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(9 downto 0);
  signal a3  : std_logic_vector(1 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(9 downto 0);
  signal sum : std_logic_vector(9 downto 0);
begin
  a0 <= x(6 downto 4);
  inst_t0 : LNSSub_MNMX_T6_10_t0
    port map ( x => a0,
               r => r0(9 downto 0) );

  a1 <= x(6 downto 4);
  b1 <= x(3 downto 1);
  inst_mult : LNSSub_MNMX_T6_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(5 downto 0) );
  r1(9 downto 6) <= (9 downto 6 => '0');

  a2 <= x(6 downto 5);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T6_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(9 downto 0) );

  a3 <= x(6 downto 5);
  b3 <= x(3 downto 3);
  inst_xor3 : LNSSub_MNMX_T6_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(9 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(9 downto 1);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.125000, -0.062500 [ -> [ 0.000000, 8.000000 [
-- Input:  wE =  -4, wF =  10, w =   6
-- Output: wE =   3, wF =   6, w =   9
-- Decomposition: a  =  2, b  =  4
--                a0 =  2, b0 =  2, p0 =  2
--                a1 =  1, b1 =  2, p1 =  4
--                a2 =  1, b2 =  1, p2 =  2
--                g0 =  1, g1 =  -4
-- ROMs: 2^ 2 x 10  +  2^ 2 x  7  +  2^ 3 x  2  +  2^ 2 x  0  =      84 bits
-- Mult: 2 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T7_10 is
  component LNSSub_MNMX_T7_10_t0 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_t1 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_t2 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_t3 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_mult is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_xor2 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MNMX_T7_10_xor3 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(9 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_10_t0 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_t0 is
begin
  with x select
    r <=
      "0111001111" when "00", -- t[0] = 463
      "0111100111" when "01", -- t[1] = 487
      "1000000011" when "10", -- t[2] = 515
      "1000100100" when "11", -- t[3] = 548
      "----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_10_t1 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_t1 is
begin
  with x select
    r <=
      "0101111" when "00", -- t[0] = 47
      "0110111" when "01", -- t[1] = 55
      "1000001" when "10", -- t[2] = 65
      "1010000" when "11", -- t[3] = 80
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_10_t2 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_t2 is
begin
  with x select
    r <=
      "00" when "00", -- t[0] = 0
      "10" when "01", -- t[1] = 2
      "01" when "10", -- t[2] = 1
      "11" when "11", -- t[3] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T7_10_t3 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_t3 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_10.all;

entity LNSSub_MNMX_T7_10_mult is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T7_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(8 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_10.all;

entity LNSSub_MNMX_T7_10_xor2 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a;
  in_t(0) <= b(0) xor sign;

  inst_t2 : LNSSub_MNMX_T7_10_t2
    port map ( x => in_t,
               r => out_t );

  r(9 downto 2) <= (9 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_10.all;

entity LNSSub_MNMX_T7_10_xor3 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T7_10_t3
    port map ( x => in_t,
               r => out_t );

  r(9 downto 1) <= (9 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T7_10.all;

entity LNSSub_MNMX_T7_10 is
  port ( x : in  std_logic_vector(5 downto 0);
         r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T7_10 is
  signal a0  : std_logic_vector(1 downto 0);
  signal r0  : std_logic_vector(9 downto 0);
  signal a1  : std_logic_vector(1 downto 0);
  signal b1  : std_logic_vector(1 downto 0);
  signal r1  : std_logic_vector(9 downto 0);
  signal a2  : std_logic_vector(0 downto 0);
  signal b2  : std_logic_vector(1 downto 0);
  signal r2  : std_logic_vector(9 downto 0);
  signal a3  : std_logic_vector(0 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(9 downto 0);
  signal sum : std_logic_vector(9 downto 0);
begin
  a0 <= x(5 downto 4);
  inst_t0 : LNSSub_MNMX_T7_10_t0
    port map ( x => a0,
               r => r0(9 downto 0) );

  a1 <= x(5 downto 4);
  b1 <= x(3 downto 2);
  inst_mult : LNSSub_MNMX_T7_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(5 downto 0) );
  r1(9 downto 6) <= (9 downto 6 => '0');

  a2 <= x(5 downto 5);
  b2 <= x(1 downto 0);
  inst_xor2 : LNSSub_MNMX_T7_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(9 downto 0) );

  a3 <= x(5 downto 5);
  b3 <= x(3 downto 3);
  inst_xor3 : LNSSub_MNMX_T7_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(9 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(9 downto 1);
end architecture;


-- Minimax-Defour: LNS subtraction function [ -0.062500, -0.031250 [ -> [ 0.000000, 8.000000 [
-- Input:  wE =  -5, wF =  10, w =   5
-- Output: wE =   3, wF =   5, w =   8
-- Decomposition: a  =  2, b  =  3
--                a0 =  2, b0 =  2, p0 =  2
--                a1 =  1, b1 =  1, p1 =  4
--                a2 =  1, b2 =  1, p2 =  2
--                g0 =  0, g1 =  -4
-- ROMs: 2^ 2 x  8  +  2^ 2 x  7  +  2^ 2 x  0  +  2^ 2 x  0  =      60 bits
-- Mult: 2 x 7 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MNMX_T8_10 is
  component LNSSub_MNMX_T8_10_t0 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_t1 is
    port ( x : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_t2 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_t3 is
    port ( x : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_mult is
    port ( a : in  std_logic_vector(1 downto 0);
           b : in  std_logic_vector(1 downto 0);
           r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_xor2 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MNMX_T8_10_xor3 is
    port ( a : in  std_logic_vector(0 downto 0);
           b : in  std_logic_vector(0 downto 0);
           r : out std_logic_vector(7 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_10_t0 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_t0 is
begin
  with x select
    r <=
      "10010011" when "00", -- t[0] = 147
      "10011001" when "01", -- t[1] = 153
      "10100000" when "10", -- t[2] = 160
      "10101001" when "11", -- t[3] = 169
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_10_t1 is
  port ( x : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_t1 is
begin
  with x select
    r <=
      "0110000" when "00", -- t[0] = 48
      "0110111" when "01", -- t[1] = 55
      "1000010" when "10", -- t[2] = 66
      "1010000" when "11", -- t[3] = 80
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_10_t2 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_t2 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T8_10_t3 is
  port ( x : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_t3 is
begin
  with x select
    r <=
      "0" when "0", -- t[0] = 0
      "0" when "1", -- t[1] = 0
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_10.all;

entity LNSSub_MNMX_T8_10_mult is
  port ( a : in  std_logic_vector(1 downto 0);
         b : in  std_logic_vector(1 downto 0);
         r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_mult is
  signal out_t : std_logic_vector(6 downto 0);
  signal r0    : std_logic_vector(8 downto 0);
begin
  inst_t1 : LNSSub_MNMX_T8_10_t1
    port map ( x => a,
               r => out_t );
  r0 <= out_t * b;
  r <= r0(8 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_10.all;

entity LNSSub_MNMX_T8_10_xor2 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_xor2 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t2 : LNSSub_MNMX_T8_10_t2
    port map ( x => in_t,
               r => out_t );

  r(7 downto 1) <= (7 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_10.all;

entity LNSSub_MNMX_T8_10_xor3 is
  port ( a : in  std_logic_vector(0 downto 0);
         b : in  std_logic_vector(0 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10_xor3 is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(0 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(0);
  in_t(0 downto 0) <= a;

  inst_t3 : LNSSub_MNMX_T8_10_t3
    port map ( x => in_t,
               r => out_t );

  r(7 downto 1) <= (7 downto 1 => '0');
  r(0) <= out_t(0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MNMX_T8_10.all;

entity LNSSub_MNMX_T8_10 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T8_10 is
  signal a0  : std_logic_vector(1 downto 0);
  signal r0  : std_logic_vector(7 downto 0);
  signal a1  : std_logic_vector(1 downto 0);
  signal b1  : std_logic_vector(1 downto 0);
  signal r1  : std_logic_vector(7 downto 0);
  signal a2  : std_logic_vector(0 downto 0);
  signal b2  : std_logic_vector(0 downto 0);
  signal r2  : std_logic_vector(7 downto 0);
  signal a3  : std_logic_vector(0 downto 0);
  signal b3  : std_logic_vector(0 downto 0);
  signal r3  : std_logic_vector(7 downto 0);
  signal sum : std_logic_vector(7 downto 0);
begin
  a0 <= x(4 downto 3);
  inst_t0 : LNSSub_MNMX_T8_10_t0
    port map ( x => a0,
               r => r0(7 downto 0) );

  a1 <= x(4 downto 3);
  b1 <= x(2 downto 1);
  inst_mult : LNSSub_MNMX_T8_10_mult
    port map ( a => a1,
               b => b1,
               r => r1(3 downto 0) );
  r1(7 downto 4) <= (7 downto 4 => '0');

  a2 <= x(4 downto 4);
  b2 <= x(0 downto 0);
  inst_xor2 : LNSSub_MNMX_T8_10_xor2
    port map ( a => a2,
               b => b2,
               r => r2(7 downto 0) );

  a3 <= x(4 downto 4);
  b3 <= x(2 downto 2);
  inst_xor3 : LNSSub_MNMX_T8_10_xor3
    port map ( a => a3,
               b => b3,
               r => r3(7 downto 0) );

  sum <= r0 + r1 + r2 + r3;
  r <= sum(7 downto 0);
end architecture;


-- Simple table: LNS subtraction function [ -0.031250, 0.000000 [ -> [ 0.000000, 16.000000 [
-- Input:  wE =  -5, wF =  10, w =   5
-- Output: wE =   4, wF =   4, w =   8

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MNMX_T9_10 is
  port ( x : in  std_logic_vector(4 downto 0);
         r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_T9_10 is
begin
  with x select
    r <=
      "01011001" when "00000", -- t[0] = 89
      "01011001" when "00001", -- t[1] = 89
      "01011010" when "00010", -- t[2] = 90
      "01011011" when "00011", -- t[3] = 91
      "01011100" when "00100", -- t[4] = 92
      "01011101" when "00101", -- t[5] = 93
      "01011101" when "00110", -- t[6] = 93
      "01011110" when "00111", -- t[7] = 94
      "01011111" when "01000", -- t[8] = 95
      "01100000" when "01001", -- t[9] = 96
      "01100001" when "01010", -- t[10] = 97
      "01100010" when "01011", -- t[11] = 98
      "01100011" when "01100", -- t[12] = 99
      "01100101" when "01101", -- t[13] = 101
      "01100110" when "01110", -- t[14] = 102
      "01100111" when "01111", -- t[15] = 103
      "01101001" when "10000", -- t[16] = 105
      "01101010" when "10001", -- t[17] = 106
      "01101100" when "10010", -- t[18] = 108
      "01101101" when "10011", -- t[19] = 109
      "01101111" when "10100", -- t[20] = 111
      "01110001" when "10101", -- t[21] = 113
      "01110011" when "10110", -- t[22] = 115
      "01110110" when "10111", -- t[23] = 118
      "01111001" when "11000", -- t[24] = 121
      "01111100" when "11001", -- t[25] = 124
      "01111111" when "11010", -- t[26] = 127
      "10000011" when "11011", -- t[27] = 131
      "10001000" when "11100", -- t[28] = 136
      "10001111" when "11101", -- t[29] = 143
      "10011000" when "11110", -- t[30] = 152
      "10101000" when "11111", -- t[31] = 168
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_lnssub_mnmx_10.all;

entity LNSSub_MNMX_10 is
  port ( x : in  std_logic_vector(13 downto 0);
         r : out std_logic_vector(13 downto 0) );
end entity;

architecture arch of LNSSub_MNMX_10 is
  signal out_t0 : std_logic_vector(3 downto 0);
  signal out_t1 : std_logic_vector(6 downto 0);
  signal out_t2 : std_logic_vector(8 downto 0);
  signal out_t3 : std_logic_vector(9 downto 0);
  signal out_t4 : std_logic_vector(10 downto 0);
  signal out_t5 : std_logic_vector(9 downto 0);
  signal out_t6 : std_logic_vector(8 downto 0);
  signal out_t7 : std_logic_vector(8 downto 0);
  signal out_t8 : std_logic_vector(7 downto 0);
  signal out_t9 : std_logic_vector(7 downto 0);
begin
  inst_t0 : LNSSub_MNMX_T0_10
    port map ( x => x(13 downto 0),
               r => out_t0 );

  inst_t1 : LNSSub_MNMX_T1_10
    port map ( x => x(11 downto 0),
               r => out_t1 );

  inst_t2 : LNSSub_MNMX_T2_10
    port map ( x => x(10 downto 0),
               r => out_t2 );

  inst_t3 : LNSSub_MNMX_T3_10
    port map ( x => x(9 downto 0),
               r => out_t3 );

  inst_t4 : LNSSub_MNMX_T4_10
    port map ( x => x(8 downto 0),
               r => out_t4 );

  inst_t5 : LNSSub_MNMX_T5_10
    port map ( x => x(7 downto 0),
               r => out_t5 );

  inst_t6 : LNSSub_MNMX_T6_10
    port map ( x => x(6 downto 0),
               r => out_t6 );

  inst_t7 : LNSSub_MNMX_T7_10
    port map ( x => x(5 downto 0),
               r => out_t7 );

  inst_t8 : LNSSub_MNMX_T8_10
    port map ( x => x(4 downto 0),
               r => out_t8 );

  inst_t9 : LNSSub_MNMX_T9_10
    port map ( x => x(4 downto 0),
               r => out_t9 );

  r <= (13 downto 4 => '0') & out_t0
         when x(13 downto 13) /= (13 downto 13 => '1') else
       (13 downto 7 => '0') & out_t1
         when x(12) /= '1' else
       (13 downto 9 => '0') & out_t2
         when x(11) /= '1' else
       (13 downto 10 => '0') & out_t3
         when x(10) /= '1' else
       (13 downto 11 => '0') & out_t4
         when x(9) /= '1' else
       (13 downto 12 => '0') & out_t5 & (1 downto 0 => '0')
         when x(8) /= '1' else
       (13 downto 12 => '0') & out_t6 & (2 downto 0 => '0')
         when x(7) /= '1' else
       (13 downto 13 => '0') & out_t7 & (3 downto 0 => '0')
         when x(6) /= '1' else
       (13 downto 13 => '0') & out_t8 & (4 downto 0 => '0')
         when x(5) /= '1' else
       out_t9 & (5 downto 0 => '0');
end architecture;
