-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


-- Implementation of MultiPartiteSubtracter object for LNS arithmetic in base 2.0 with 8-bit integer part and 12-bit fractional part
-- wI = 16 bits
-- wO = 16 bits

library ieee;
use ieee.std_logic_1164.all;

package pkg_lnssub_mpt_12 is
  component LNSSub_MPT_T0_12 is
    port( x : in  std_logic_vector(15 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T1_12 is
    port( x : in  std_logic_vector(13 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T1_12_Clk is
    port( x   : in  std_logic_vector(13 downto 0);
          r   : out std_logic_vector(8 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T2_12 is
    port( x : in  std_logic_vector(12 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_Clk is
    port( x   : in  std_logic_vector(12 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T3_12 is
    port( x : in  std_logic_vector(11 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_Clk is
    port( x   : in  std_logic_vector(11 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T4_12 is
    port( x : in  std_logic_vector(10 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_Clk is
    port( x   : in  std_logic_vector(10 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T5_12 is
    port( x : in  std_logic_vector(9 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T5_12_Clk is
    port( x   : in  std_logic_vector(9 downto 0);
          r   : out std_logic_vector(10 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T6_12 is
    port( x : in  std_logic_vector(8 downto 0);
          r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MPT_T6_12_Clk is
    port( x   : in  std_logic_vector(8 downto 0);
          r   : out std_logic_vector(9 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T7_12 is
    port( x : in  std_logic_vector(7 downto 0);
          r : out std_logic_vector(9 downto 0) );
  end component;

  component LNSSub_MPT_T7_12_Clk is
    port( x   : in  std_logic_vector(7 downto 0);
          r   : out std_logic_vector(9 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T8_12 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T8_12_Clk is
    port( x   : in  std_logic_vector(6 downto 0);
          r   : out std_logic_vector(8 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T9_12 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T9_12_Clk is
    port( x   : in  std_logic_vector(5 downto 0);
          r   : out std_logic_vector(7 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T10_12 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T10_12_Clk is
    port( x   : in  std_logic_vector(4 downto 0);
          r   : out std_logic_vector(6 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T11_12 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T11_12_Clk is
    port( x   : in  std_logic_vector(3 downto 0);
          r   : out std_logic_vector(6 downto 0);
          clk : in  std_logic );
  end component;

  component LNSSub_MPT_T12_12 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T12_12_Clk is
    port( x   : in  std_logic_vector(3 downto 0);
          r   : out std_logic_vector(6 downto 0);
          clk : in  std_logic );
  end component;
end package;


-- SimpleTable: LNS subtraction function: [-16.0 0.0[ -> [0.0 1.0[
-- (bounded to [-16.0; -8.0[)
-- wI = 16 bits
-- wO = 6 bits

library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T0_12 is
  port( x : in  std_logic_vector(15 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T0_12 is
begin
  with x select
    r <=
      "000000" when "0000000000000000", -- t[0] = 0
      "000000" when "0000000000000001", -- t[1] = 0
      "000000" when "0000000000000010", -- t[2] = 0
      "000000" when "0000000000000011", -- t[3] = 0
      "000000" when "0000000000000100", -- t[4] = 0
      "000000" when "0000000000000101", -- t[5] = 0
      "000000" when "0000000000000110", -- t[6] = 0
      "000000" when "0000000000000111", -- t[7] = 0
      "000000" when "0000000000001000", -- t[8] = 0
      "000000" when "0000000000001001", -- t[9] = 0
      "000000" when "0000000000001010", -- t[10] = 0
      "000000" when "0000000000001011", -- t[11] = 0
      "000000" when "0000000000001100", -- t[12] = 0
      "000000" when "0000000000001101", -- t[13] = 0
      "000000" when "0000000000001110", -- t[14] = 0
      "000000" when "0000000000001111", -- t[15] = 0
      "000000" when "0000000000010000", -- t[16] = 0
      "000000" when "0000000000010001", -- t[17] = 0
      "000000" when "0000000000010010", -- t[18] = 0
      "000000" when "0000000000010011", -- t[19] = 0
      "000000" when "0000000000010100", -- t[20] = 0
      "000000" when "0000000000010101", -- t[21] = 0
      "000000" when "0000000000010110", -- t[22] = 0
      "000000" when "0000000000010111", -- t[23] = 0
      "000000" when "0000000000011000", -- t[24] = 0
      "000000" when "0000000000011001", -- t[25] = 0
      "000000" when "0000000000011010", -- t[26] = 0
      "000000" when "0000000000011011", -- t[27] = 0
      "000000" when "0000000000011100", -- t[28] = 0
      "000000" when "0000000000011101", -- t[29] = 0
      "000000" when "0000000000011110", -- t[30] = 0
      "000000" when "0000000000011111", -- t[31] = 0
      "000000" when "0000000000100000", -- t[32] = 0
      "000000" when "0000000000100001", -- t[33] = 0
      "000000" when "0000000000100010", -- t[34] = 0
      "000000" when "0000000000100011", -- t[35] = 0
      "000000" when "0000000000100100", -- t[36] = 0
      "000000" when "0000000000100101", -- t[37] = 0
      "000000" when "0000000000100110", -- t[38] = 0
      "000000" when "0000000000100111", -- t[39] = 0
      "000000" when "0000000000101000", -- t[40] = 0
      "000000" when "0000000000101001", -- t[41] = 0
      "000000" when "0000000000101010", -- t[42] = 0
      "000000" when "0000000000101011", -- t[43] = 0
      "000000" when "0000000000101100", -- t[44] = 0
      "000000" when "0000000000101101", -- t[45] = 0
      "000000" when "0000000000101110", -- t[46] = 0
      "000000" when "0000000000101111", -- t[47] = 0
      "000000" when "0000000000110000", -- t[48] = 0
      "000000" when "0000000000110001", -- t[49] = 0
      "000000" when "0000000000110010", -- t[50] = 0
      "000000" when "0000000000110011", -- t[51] = 0
      "000000" when "0000000000110100", -- t[52] = 0
      "000000" when "0000000000110101", -- t[53] = 0
      "000000" when "0000000000110110", -- t[54] = 0
      "000000" when "0000000000110111", -- t[55] = 0
      "000000" when "0000000000111000", -- t[56] = 0
      "000000" when "0000000000111001", -- t[57] = 0
      "000000" when "0000000000111010", -- t[58] = 0
      "000000" when "0000000000111011", -- t[59] = 0
      "000000" when "0000000000111100", -- t[60] = 0
      "000000" when "0000000000111101", -- t[61] = 0
      "000000" when "0000000000111110", -- t[62] = 0
      "000000" when "0000000000111111", -- t[63] = 0
      "000000" when "0000000001000000", -- t[64] = 0
      "000000" when "0000000001000001", -- t[65] = 0
      "000000" when "0000000001000010", -- t[66] = 0
      "000000" when "0000000001000011", -- t[67] = 0
      "000000" when "0000000001000100", -- t[68] = 0
      "000000" when "0000000001000101", -- t[69] = 0
      "000000" when "0000000001000110", -- t[70] = 0
      "000000" when "0000000001000111", -- t[71] = 0
      "000000" when "0000000001001000", -- t[72] = 0
      "000000" when "0000000001001001", -- t[73] = 0
      "000000" when "0000000001001010", -- t[74] = 0
      "000000" when "0000000001001011", -- t[75] = 0
      "000000" when "0000000001001100", -- t[76] = 0
      "000000" when "0000000001001101", -- t[77] = 0
      "000000" when "0000000001001110", -- t[78] = 0
      "000000" when "0000000001001111", -- t[79] = 0
      "000000" when "0000000001010000", -- t[80] = 0
      "000000" when "0000000001010001", -- t[81] = 0
      "000000" when "0000000001010010", -- t[82] = 0
      "000000" when "0000000001010011", -- t[83] = 0
      "000000" when "0000000001010100", -- t[84] = 0
      "000000" when "0000000001010101", -- t[85] = 0
      "000000" when "0000000001010110", -- t[86] = 0
      "000000" when "0000000001010111", -- t[87] = 0
      "000000" when "0000000001011000", -- t[88] = 0
      "000000" when "0000000001011001", -- t[89] = 0
      "000000" when "0000000001011010", -- t[90] = 0
      "000000" when "0000000001011011", -- t[91] = 0
      "000000" when "0000000001011100", -- t[92] = 0
      "000000" when "0000000001011101", -- t[93] = 0
      "000000" when "0000000001011110", -- t[94] = 0
      "000000" when "0000000001011111", -- t[95] = 0
      "000000" when "0000000001100000", -- t[96] = 0
      "000000" when "0000000001100001", -- t[97] = 0
      "000000" when "0000000001100010", -- t[98] = 0
      "000000" when "0000000001100011", -- t[99] = 0
      "000000" when "0000000001100100", -- t[100] = 0
      "000000" when "0000000001100101", -- t[101] = 0
      "000000" when "0000000001100110", -- t[102] = 0
      "000000" when "0000000001100111", -- t[103] = 0
      "000000" when "0000000001101000", -- t[104] = 0
      "000000" when "0000000001101001", -- t[105] = 0
      "000000" when "0000000001101010", -- t[106] = 0
      "000000" when "0000000001101011", -- t[107] = 0
      "000000" when "0000000001101100", -- t[108] = 0
      "000000" when "0000000001101101", -- t[109] = 0
      "000000" when "0000000001101110", -- t[110] = 0
      "000000" when "0000000001101111", -- t[111] = 0
      "000000" when "0000000001110000", -- t[112] = 0
      "000000" when "0000000001110001", -- t[113] = 0
      "000000" when "0000000001110010", -- t[114] = 0
      "000000" when "0000000001110011", -- t[115] = 0
      "000000" when "0000000001110100", -- t[116] = 0
      "000000" when "0000000001110101", -- t[117] = 0
      "000000" when "0000000001110110", -- t[118] = 0
      "000000" when "0000000001110111", -- t[119] = 0
      "000000" when "0000000001111000", -- t[120] = 0
      "000000" when "0000000001111001", -- t[121] = 0
      "000000" when "0000000001111010", -- t[122] = 0
      "000000" when "0000000001111011", -- t[123] = 0
      "000000" when "0000000001111100", -- t[124] = 0
      "000000" when "0000000001111101", -- t[125] = 0
      "000000" when "0000000001111110", -- t[126] = 0
      "000000" when "0000000001111111", -- t[127] = 0
      "000000" when "0000000010000000", -- t[128] = 0
      "000000" when "0000000010000001", -- t[129] = 0
      "000000" when "0000000010000010", -- t[130] = 0
      "000000" when "0000000010000011", -- t[131] = 0
      "000000" when "0000000010000100", -- t[132] = 0
      "000000" when "0000000010000101", -- t[133] = 0
      "000000" when "0000000010000110", -- t[134] = 0
      "000000" when "0000000010000111", -- t[135] = 0
      "000000" when "0000000010001000", -- t[136] = 0
      "000000" when "0000000010001001", -- t[137] = 0
      "000000" when "0000000010001010", -- t[138] = 0
      "000000" when "0000000010001011", -- t[139] = 0
      "000000" when "0000000010001100", -- t[140] = 0
      "000000" when "0000000010001101", -- t[141] = 0
      "000000" when "0000000010001110", -- t[142] = 0
      "000000" when "0000000010001111", -- t[143] = 0
      "000000" when "0000000010010000", -- t[144] = 0
      "000000" when "0000000010010001", -- t[145] = 0
      "000000" when "0000000010010010", -- t[146] = 0
      "000000" when "0000000010010011", -- t[147] = 0
      "000000" when "0000000010010100", -- t[148] = 0
      "000000" when "0000000010010101", -- t[149] = 0
      "000000" when "0000000010010110", -- t[150] = 0
      "000000" when "0000000010010111", -- t[151] = 0
      "000000" when "0000000010011000", -- t[152] = 0
      "000000" when "0000000010011001", -- t[153] = 0
      "000000" when "0000000010011010", -- t[154] = 0
      "000000" when "0000000010011011", -- t[155] = 0
      "000000" when "0000000010011100", -- t[156] = 0
      "000000" when "0000000010011101", -- t[157] = 0
      "000000" when "0000000010011110", -- t[158] = 0
      "000000" when "0000000010011111", -- t[159] = 0
      "000000" when "0000000010100000", -- t[160] = 0
      "000000" when "0000000010100001", -- t[161] = 0
      "000000" when "0000000010100010", -- t[162] = 0
      "000000" when "0000000010100011", -- t[163] = 0
      "000000" when "0000000010100100", -- t[164] = 0
      "000000" when "0000000010100101", -- t[165] = 0
      "000000" when "0000000010100110", -- t[166] = 0
      "000000" when "0000000010100111", -- t[167] = 0
      "000000" when "0000000010101000", -- t[168] = 0
      "000000" when "0000000010101001", -- t[169] = 0
      "000000" when "0000000010101010", -- t[170] = 0
      "000000" when "0000000010101011", -- t[171] = 0
      "000000" when "0000000010101100", -- t[172] = 0
      "000000" when "0000000010101101", -- t[173] = 0
      "000000" when "0000000010101110", -- t[174] = 0
      "000000" when "0000000010101111", -- t[175] = 0
      "000000" when "0000000010110000", -- t[176] = 0
      "000000" when "0000000010110001", -- t[177] = 0
      "000000" when "0000000010110010", -- t[178] = 0
      "000000" when "0000000010110011", -- t[179] = 0
      "000000" when "0000000010110100", -- t[180] = 0
      "000000" when "0000000010110101", -- t[181] = 0
      "000000" when "0000000010110110", -- t[182] = 0
      "000000" when "0000000010110111", -- t[183] = 0
      "000000" when "0000000010111000", -- t[184] = 0
      "000000" when "0000000010111001", -- t[185] = 0
      "000000" when "0000000010111010", -- t[186] = 0
      "000000" when "0000000010111011", -- t[187] = 0
      "000000" when "0000000010111100", -- t[188] = 0
      "000000" when "0000000010111101", -- t[189] = 0
      "000000" when "0000000010111110", -- t[190] = 0
      "000000" when "0000000010111111", -- t[191] = 0
      "000000" when "0000000011000000", -- t[192] = 0
      "000000" when "0000000011000001", -- t[193] = 0
      "000000" when "0000000011000010", -- t[194] = 0
      "000000" when "0000000011000011", -- t[195] = 0
      "000000" when "0000000011000100", -- t[196] = 0
      "000000" when "0000000011000101", -- t[197] = 0
      "000000" when "0000000011000110", -- t[198] = 0
      "000000" when "0000000011000111", -- t[199] = 0
      "000000" when "0000000011001000", -- t[200] = 0
      "000000" when "0000000011001001", -- t[201] = 0
      "000000" when "0000000011001010", -- t[202] = 0
      "000000" when "0000000011001011", -- t[203] = 0
      "000000" when "0000000011001100", -- t[204] = 0
      "000000" when "0000000011001101", -- t[205] = 0
      "000000" when "0000000011001110", -- t[206] = 0
      "000000" when "0000000011001111", -- t[207] = 0
      "000000" when "0000000011010000", -- t[208] = 0
      "000000" when "0000000011010001", -- t[209] = 0
      "000000" when "0000000011010010", -- t[210] = 0
      "000000" when "0000000011010011", -- t[211] = 0
      "000000" when "0000000011010100", -- t[212] = 0
      "000000" when "0000000011010101", -- t[213] = 0
      "000000" when "0000000011010110", -- t[214] = 0
      "000000" when "0000000011010111", -- t[215] = 0
      "000000" when "0000000011011000", -- t[216] = 0
      "000000" when "0000000011011001", -- t[217] = 0
      "000000" when "0000000011011010", -- t[218] = 0
      "000000" when "0000000011011011", -- t[219] = 0
      "000000" when "0000000011011100", -- t[220] = 0
      "000000" when "0000000011011101", -- t[221] = 0
      "000000" when "0000000011011110", -- t[222] = 0
      "000000" when "0000000011011111", -- t[223] = 0
      "000000" when "0000000011100000", -- t[224] = 0
      "000000" when "0000000011100001", -- t[225] = 0
      "000000" when "0000000011100010", -- t[226] = 0
      "000000" when "0000000011100011", -- t[227] = 0
      "000000" when "0000000011100100", -- t[228] = 0
      "000000" when "0000000011100101", -- t[229] = 0
      "000000" when "0000000011100110", -- t[230] = 0
      "000000" when "0000000011100111", -- t[231] = 0
      "000000" when "0000000011101000", -- t[232] = 0
      "000000" when "0000000011101001", -- t[233] = 0
      "000000" when "0000000011101010", -- t[234] = 0
      "000000" when "0000000011101011", -- t[235] = 0
      "000000" when "0000000011101100", -- t[236] = 0
      "000000" when "0000000011101101", -- t[237] = 0
      "000000" when "0000000011101110", -- t[238] = 0
      "000000" when "0000000011101111", -- t[239] = 0
      "000000" when "0000000011110000", -- t[240] = 0
      "000000" when "0000000011110001", -- t[241] = 0
      "000000" when "0000000011110010", -- t[242] = 0
      "000000" when "0000000011110011", -- t[243] = 0
      "000000" when "0000000011110100", -- t[244] = 0
      "000000" when "0000000011110101", -- t[245] = 0
      "000000" when "0000000011110110", -- t[246] = 0
      "000000" when "0000000011110111", -- t[247] = 0
      "000000" when "0000000011111000", -- t[248] = 0
      "000000" when "0000000011111001", -- t[249] = 0
      "000000" when "0000000011111010", -- t[250] = 0
      "000000" when "0000000011111011", -- t[251] = 0
      "000000" when "0000000011111100", -- t[252] = 0
      "000000" when "0000000011111101", -- t[253] = 0
      "000000" when "0000000011111110", -- t[254] = 0
      "000000" when "0000000011111111", -- t[255] = 0
      "000000" when "0000000100000000", -- t[256] = 0
      "000000" when "0000000100000001", -- t[257] = 0
      "000000" when "0000000100000010", -- t[258] = 0
      "000000" when "0000000100000011", -- t[259] = 0
      "000000" when "0000000100000100", -- t[260] = 0
      "000000" when "0000000100000101", -- t[261] = 0
      "000000" when "0000000100000110", -- t[262] = 0
      "000000" when "0000000100000111", -- t[263] = 0
      "000000" when "0000000100001000", -- t[264] = 0
      "000000" when "0000000100001001", -- t[265] = 0
      "000000" when "0000000100001010", -- t[266] = 0
      "000000" when "0000000100001011", -- t[267] = 0
      "000000" when "0000000100001100", -- t[268] = 0
      "000000" when "0000000100001101", -- t[269] = 0
      "000000" when "0000000100001110", -- t[270] = 0
      "000000" when "0000000100001111", -- t[271] = 0
      "000000" when "0000000100010000", -- t[272] = 0
      "000000" when "0000000100010001", -- t[273] = 0
      "000000" when "0000000100010010", -- t[274] = 0
      "000000" when "0000000100010011", -- t[275] = 0
      "000000" when "0000000100010100", -- t[276] = 0
      "000000" when "0000000100010101", -- t[277] = 0
      "000000" when "0000000100010110", -- t[278] = 0
      "000000" when "0000000100010111", -- t[279] = 0
      "000000" when "0000000100011000", -- t[280] = 0
      "000000" when "0000000100011001", -- t[281] = 0
      "000000" when "0000000100011010", -- t[282] = 0
      "000000" when "0000000100011011", -- t[283] = 0
      "000000" when "0000000100011100", -- t[284] = 0
      "000000" when "0000000100011101", -- t[285] = 0
      "000000" when "0000000100011110", -- t[286] = 0
      "000000" when "0000000100011111", -- t[287] = 0
      "000000" when "0000000100100000", -- t[288] = 0
      "000000" when "0000000100100001", -- t[289] = 0
      "000000" when "0000000100100010", -- t[290] = 0
      "000000" when "0000000100100011", -- t[291] = 0
      "000000" when "0000000100100100", -- t[292] = 0
      "000000" when "0000000100100101", -- t[293] = 0
      "000000" when "0000000100100110", -- t[294] = 0
      "000000" when "0000000100100111", -- t[295] = 0
      "000000" when "0000000100101000", -- t[296] = 0
      "000000" when "0000000100101001", -- t[297] = 0
      "000000" when "0000000100101010", -- t[298] = 0
      "000000" when "0000000100101011", -- t[299] = 0
      "000000" when "0000000100101100", -- t[300] = 0
      "000000" when "0000000100101101", -- t[301] = 0
      "000000" when "0000000100101110", -- t[302] = 0
      "000000" when "0000000100101111", -- t[303] = 0
      "000000" when "0000000100110000", -- t[304] = 0
      "000000" when "0000000100110001", -- t[305] = 0
      "000000" when "0000000100110010", -- t[306] = 0
      "000000" when "0000000100110011", -- t[307] = 0
      "000000" when "0000000100110100", -- t[308] = 0
      "000000" when "0000000100110101", -- t[309] = 0
      "000000" when "0000000100110110", -- t[310] = 0
      "000000" when "0000000100110111", -- t[311] = 0
      "000000" when "0000000100111000", -- t[312] = 0
      "000000" when "0000000100111001", -- t[313] = 0
      "000000" when "0000000100111010", -- t[314] = 0
      "000000" when "0000000100111011", -- t[315] = 0
      "000000" when "0000000100111100", -- t[316] = 0
      "000000" when "0000000100111101", -- t[317] = 0
      "000000" when "0000000100111110", -- t[318] = 0
      "000000" when "0000000100111111", -- t[319] = 0
      "000000" when "0000000101000000", -- t[320] = 0
      "000000" when "0000000101000001", -- t[321] = 0
      "000000" when "0000000101000010", -- t[322] = 0
      "000000" when "0000000101000011", -- t[323] = 0
      "000000" when "0000000101000100", -- t[324] = 0
      "000000" when "0000000101000101", -- t[325] = 0
      "000000" when "0000000101000110", -- t[326] = 0
      "000000" when "0000000101000111", -- t[327] = 0
      "000000" when "0000000101001000", -- t[328] = 0
      "000000" when "0000000101001001", -- t[329] = 0
      "000000" when "0000000101001010", -- t[330] = 0
      "000000" when "0000000101001011", -- t[331] = 0
      "000000" when "0000000101001100", -- t[332] = 0
      "000000" when "0000000101001101", -- t[333] = 0
      "000000" when "0000000101001110", -- t[334] = 0
      "000000" when "0000000101001111", -- t[335] = 0
      "000000" when "0000000101010000", -- t[336] = 0
      "000000" when "0000000101010001", -- t[337] = 0
      "000000" when "0000000101010010", -- t[338] = 0
      "000000" when "0000000101010011", -- t[339] = 0
      "000000" when "0000000101010100", -- t[340] = 0
      "000000" when "0000000101010101", -- t[341] = 0
      "000000" when "0000000101010110", -- t[342] = 0
      "000000" when "0000000101010111", -- t[343] = 0
      "000000" when "0000000101011000", -- t[344] = 0
      "000000" when "0000000101011001", -- t[345] = 0
      "000000" when "0000000101011010", -- t[346] = 0
      "000000" when "0000000101011011", -- t[347] = 0
      "000000" when "0000000101011100", -- t[348] = 0
      "000000" when "0000000101011101", -- t[349] = 0
      "000000" when "0000000101011110", -- t[350] = 0
      "000000" when "0000000101011111", -- t[351] = 0
      "000000" when "0000000101100000", -- t[352] = 0
      "000000" when "0000000101100001", -- t[353] = 0
      "000000" when "0000000101100010", -- t[354] = 0
      "000000" when "0000000101100011", -- t[355] = 0
      "000000" when "0000000101100100", -- t[356] = 0
      "000000" when "0000000101100101", -- t[357] = 0
      "000000" when "0000000101100110", -- t[358] = 0
      "000000" when "0000000101100111", -- t[359] = 0
      "000000" when "0000000101101000", -- t[360] = 0
      "000000" when "0000000101101001", -- t[361] = 0
      "000000" when "0000000101101010", -- t[362] = 0
      "000000" when "0000000101101011", -- t[363] = 0
      "000000" when "0000000101101100", -- t[364] = 0
      "000000" when "0000000101101101", -- t[365] = 0
      "000000" when "0000000101101110", -- t[366] = 0
      "000000" when "0000000101101111", -- t[367] = 0
      "000000" when "0000000101110000", -- t[368] = 0
      "000000" when "0000000101110001", -- t[369] = 0
      "000000" when "0000000101110010", -- t[370] = 0
      "000000" when "0000000101110011", -- t[371] = 0
      "000000" when "0000000101110100", -- t[372] = 0
      "000000" when "0000000101110101", -- t[373] = 0
      "000000" when "0000000101110110", -- t[374] = 0
      "000000" when "0000000101110111", -- t[375] = 0
      "000000" when "0000000101111000", -- t[376] = 0
      "000000" when "0000000101111001", -- t[377] = 0
      "000000" when "0000000101111010", -- t[378] = 0
      "000000" when "0000000101111011", -- t[379] = 0
      "000000" when "0000000101111100", -- t[380] = 0
      "000000" when "0000000101111101", -- t[381] = 0
      "000000" when "0000000101111110", -- t[382] = 0
      "000000" when "0000000101111111", -- t[383] = 0
      "000000" when "0000000110000000", -- t[384] = 0
      "000000" when "0000000110000001", -- t[385] = 0
      "000000" when "0000000110000010", -- t[386] = 0
      "000000" when "0000000110000011", -- t[387] = 0
      "000000" when "0000000110000100", -- t[388] = 0
      "000000" when "0000000110000101", -- t[389] = 0
      "000000" when "0000000110000110", -- t[390] = 0
      "000000" when "0000000110000111", -- t[391] = 0
      "000000" when "0000000110001000", -- t[392] = 0
      "000000" when "0000000110001001", -- t[393] = 0
      "000000" when "0000000110001010", -- t[394] = 0
      "000000" when "0000000110001011", -- t[395] = 0
      "000000" when "0000000110001100", -- t[396] = 0
      "000000" when "0000000110001101", -- t[397] = 0
      "000000" when "0000000110001110", -- t[398] = 0
      "000000" when "0000000110001111", -- t[399] = 0
      "000000" when "0000000110010000", -- t[400] = 0
      "000000" when "0000000110010001", -- t[401] = 0
      "000000" when "0000000110010010", -- t[402] = 0
      "000000" when "0000000110010011", -- t[403] = 0
      "000000" when "0000000110010100", -- t[404] = 0
      "000000" when "0000000110010101", -- t[405] = 0
      "000000" when "0000000110010110", -- t[406] = 0
      "000000" when "0000000110010111", -- t[407] = 0
      "000000" when "0000000110011000", -- t[408] = 0
      "000000" when "0000000110011001", -- t[409] = 0
      "000000" when "0000000110011010", -- t[410] = 0
      "000000" when "0000000110011011", -- t[411] = 0
      "000000" when "0000000110011100", -- t[412] = 0
      "000000" when "0000000110011101", -- t[413] = 0
      "000000" when "0000000110011110", -- t[414] = 0
      "000000" when "0000000110011111", -- t[415] = 0
      "000000" when "0000000110100000", -- t[416] = 0
      "000000" when "0000000110100001", -- t[417] = 0
      "000000" when "0000000110100010", -- t[418] = 0
      "000000" when "0000000110100011", -- t[419] = 0
      "000000" when "0000000110100100", -- t[420] = 0
      "000000" when "0000000110100101", -- t[421] = 0
      "000000" when "0000000110100110", -- t[422] = 0
      "000000" when "0000000110100111", -- t[423] = 0
      "000000" when "0000000110101000", -- t[424] = 0
      "000000" when "0000000110101001", -- t[425] = 0
      "000000" when "0000000110101010", -- t[426] = 0
      "000000" when "0000000110101011", -- t[427] = 0
      "000000" when "0000000110101100", -- t[428] = 0
      "000000" when "0000000110101101", -- t[429] = 0
      "000000" when "0000000110101110", -- t[430] = 0
      "000000" when "0000000110101111", -- t[431] = 0
      "000000" when "0000000110110000", -- t[432] = 0
      "000000" when "0000000110110001", -- t[433] = 0
      "000000" when "0000000110110010", -- t[434] = 0
      "000000" when "0000000110110011", -- t[435] = 0
      "000000" when "0000000110110100", -- t[436] = 0
      "000000" when "0000000110110101", -- t[437] = 0
      "000000" when "0000000110110110", -- t[438] = 0
      "000000" when "0000000110110111", -- t[439] = 0
      "000000" when "0000000110111000", -- t[440] = 0
      "000000" when "0000000110111001", -- t[441] = 0
      "000000" when "0000000110111010", -- t[442] = 0
      "000000" when "0000000110111011", -- t[443] = 0
      "000000" when "0000000110111100", -- t[444] = 0
      "000000" when "0000000110111101", -- t[445] = 0
      "000000" when "0000000110111110", -- t[446] = 0
      "000000" when "0000000110111111", -- t[447] = 0
      "000000" when "0000000111000000", -- t[448] = 0
      "000000" when "0000000111000001", -- t[449] = 0
      "000000" when "0000000111000010", -- t[450] = 0
      "000000" when "0000000111000011", -- t[451] = 0
      "000000" when "0000000111000100", -- t[452] = 0
      "000000" when "0000000111000101", -- t[453] = 0
      "000000" when "0000000111000110", -- t[454] = 0
      "000000" when "0000000111000111", -- t[455] = 0
      "000000" when "0000000111001000", -- t[456] = 0
      "000000" when "0000000111001001", -- t[457] = 0
      "000000" when "0000000111001010", -- t[458] = 0
      "000000" when "0000000111001011", -- t[459] = 0
      "000000" when "0000000111001100", -- t[460] = 0
      "000000" when "0000000111001101", -- t[461] = 0
      "000000" when "0000000111001110", -- t[462] = 0
      "000000" when "0000000111001111", -- t[463] = 0
      "000000" when "0000000111010000", -- t[464] = 0
      "000000" when "0000000111010001", -- t[465] = 0
      "000000" when "0000000111010010", -- t[466] = 0
      "000000" when "0000000111010011", -- t[467] = 0
      "000000" when "0000000111010100", -- t[468] = 0
      "000000" when "0000000111010101", -- t[469] = 0
      "000000" when "0000000111010110", -- t[470] = 0
      "000000" when "0000000111010111", -- t[471] = 0
      "000000" when "0000000111011000", -- t[472] = 0
      "000000" when "0000000111011001", -- t[473] = 0
      "000000" when "0000000111011010", -- t[474] = 0
      "000000" when "0000000111011011", -- t[475] = 0
      "000000" when "0000000111011100", -- t[476] = 0
      "000000" when "0000000111011101", -- t[477] = 0
      "000000" when "0000000111011110", -- t[478] = 0
      "000000" when "0000000111011111", -- t[479] = 0
      "000000" when "0000000111100000", -- t[480] = 0
      "000000" when "0000000111100001", -- t[481] = 0
      "000000" when "0000000111100010", -- t[482] = 0
      "000000" when "0000000111100011", -- t[483] = 0
      "000000" when "0000000111100100", -- t[484] = 0
      "000000" when "0000000111100101", -- t[485] = 0
      "000000" when "0000000111100110", -- t[486] = 0
      "000000" when "0000000111100111", -- t[487] = 0
      "000000" when "0000000111101000", -- t[488] = 0
      "000000" when "0000000111101001", -- t[489] = 0
      "000000" when "0000000111101010", -- t[490] = 0
      "000000" when "0000000111101011", -- t[491] = 0
      "000000" when "0000000111101100", -- t[492] = 0
      "000000" when "0000000111101101", -- t[493] = 0
      "000000" when "0000000111101110", -- t[494] = 0
      "000000" when "0000000111101111", -- t[495] = 0
      "000000" when "0000000111110000", -- t[496] = 0
      "000000" when "0000000111110001", -- t[497] = 0
      "000000" when "0000000111110010", -- t[498] = 0
      "000000" when "0000000111110011", -- t[499] = 0
      "000000" when "0000000111110100", -- t[500] = 0
      "000000" when "0000000111110101", -- t[501] = 0
      "000000" when "0000000111110110", -- t[502] = 0
      "000000" when "0000000111110111", -- t[503] = 0
      "000000" when "0000000111111000", -- t[504] = 0
      "000000" when "0000000111111001", -- t[505] = 0
      "000000" when "0000000111111010", -- t[506] = 0
      "000000" when "0000000111111011", -- t[507] = 0
      "000000" when "0000000111111100", -- t[508] = 0
      "000000" when "0000000111111101", -- t[509] = 0
      "000000" when "0000000111111110", -- t[510] = 0
      "000000" when "0000000111111111", -- t[511] = 0
      "000000" when "0000001000000000", -- t[512] = 0
      "000000" when "0000001000000001", -- t[513] = 0
      "000000" when "0000001000000010", -- t[514] = 0
      "000000" when "0000001000000011", -- t[515] = 0
      "000000" when "0000001000000100", -- t[516] = 0
      "000000" when "0000001000000101", -- t[517] = 0
      "000000" when "0000001000000110", -- t[518] = 0
      "000000" when "0000001000000111", -- t[519] = 0
      "000000" when "0000001000001000", -- t[520] = 0
      "000000" when "0000001000001001", -- t[521] = 0
      "000000" when "0000001000001010", -- t[522] = 0
      "000000" when "0000001000001011", -- t[523] = 0
      "000000" when "0000001000001100", -- t[524] = 0
      "000000" when "0000001000001101", -- t[525] = 0
      "000000" when "0000001000001110", -- t[526] = 0
      "000000" when "0000001000001111", -- t[527] = 0
      "000000" when "0000001000010000", -- t[528] = 0
      "000000" when "0000001000010001", -- t[529] = 0
      "000000" when "0000001000010010", -- t[530] = 0
      "000000" when "0000001000010011", -- t[531] = 0
      "000000" when "0000001000010100", -- t[532] = 0
      "000000" when "0000001000010101", -- t[533] = 0
      "000000" when "0000001000010110", -- t[534] = 0
      "000000" when "0000001000010111", -- t[535] = 0
      "000000" when "0000001000011000", -- t[536] = 0
      "000000" when "0000001000011001", -- t[537] = 0
      "000000" when "0000001000011010", -- t[538] = 0
      "000000" when "0000001000011011", -- t[539] = 0
      "000000" when "0000001000011100", -- t[540] = 0
      "000000" when "0000001000011101", -- t[541] = 0
      "000000" when "0000001000011110", -- t[542] = 0
      "000000" when "0000001000011111", -- t[543] = 0
      "000000" when "0000001000100000", -- t[544] = 0
      "000000" when "0000001000100001", -- t[545] = 0
      "000000" when "0000001000100010", -- t[546] = 0
      "000000" when "0000001000100011", -- t[547] = 0
      "000000" when "0000001000100100", -- t[548] = 0
      "000000" when "0000001000100101", -- t[549] = 0
      "000000" when "0000001000100110", -- t[550] = 0
      "000000" when "0000001000100111", -- t[551] = 0
      "000000" when "0000001000101000", -- t[552] = 0
      "000000" when "0000001000101001", -- t[553] = 0
      "000000" when "0000001000101010", -- t[554] = 0
      "000000" when "0000001000101011", -- t[555] = 0
      "000000" when "0000001000101100", -- t[556] = 0
      "000000" when "0000001000101101", -- t[557] = 0
      "000000" when "0000001000101110", -- t[558] = 0
      "000000" when "0000001000101111", -- t[559] = 0
      "000000" when "0000001000110000", -- t[560] = 0
      "000000" when "0000001000110001", -- t[561] = 0
      "000000" when "0000001000110010", -- t[562] = 0
      "000000" when "0000001000110011", -- t[563] = 0
      "000000" when "0000001000110100", -- t[564] = 0
      "000000" when "0000001000110101", -- t[565] = 0
      "000000" when "0000001000110110", -- t[566] = 0
      "000000" when "0000001000110111", -- t[567] = 0
      "000000" when "0000001000111000", -- t[568] = 0
      "000000" when "0000001000111001", -- t[569] = 0
      "000000" when "0000001000111010", -- t[570] = 0
      "000000" when "0000001000111011", -- t[571] = 0
      "000000" when "0000001000111100", -- t[572] = 0
      "000000" when "0000001000111101", -- t[573] = 0
      "000000" when "0000001000111110", -- t[574] = 0
      "000000" when "0000001000111111", -- t[575] = 0
      "000000" when "0000001001000000", -- t[576] = 0
      "000000" when "0000001001000001", -- t[577] = 0
      "000000" when "0000001001000010", -- t[578] = 0
      "000000" when "0000001001000011", -- t[579] = 0
      "000000" when "0000001001000100", -- t[580] = 0
      "000000" when "0000001001000101", -- t[581] = 0
      "000000" when "0000001001000110", -- t[582] = 0
      "000000" when "0000001001000111", -- t[583] = 0
      "000000" when "0000001001001000", -- t[584] = 0
      "000000" when "0000001001001001", -- t[585] = 0
      "000000" when "0000001001001010", -- t[586] = 0
      "000000" when "0000001001001011", -- t[587] = 0
      "000000" when "0000001001001100", -- t[588] = 0
      "000000" when "0000001001001101", -- t[589] = 0
      "000000" when "0000001001001110", -- t[590] = 0
      "000000" when "0000001001001111", -- t[591] = 0
      "000000" when "0000001001010000", -- t[592] = 0
      "000000" when "0000001001010001", -- t[593] = 0
      "000000" when "0000001001010010", -- t[594] = 0
      "000000" when "0000001001010011", -- t[595] = 0
      "000000" when "0000001001010100", -- t[596] = 0
      "000000" when "0000001001010101", -- t[597] = 0
      "000000" when "0000001001010110", -- t[598] = 0
      "000000" when "0000001001010111", -- t[599] = 0
      "000000" when "0000001001011000", -- t[600] = 0
      "000000" when "0000001001011001", -- t[601] = 0
      "000000" when "0000001001011010", -- t[602] = 0
      "000000" when "0000001001011011", -- t[603] = 0
      "000000" when "0000001001011100", -- t[604] = 0
      "000000" when "0000001001011101", -- t[605] = 0
      "000000" when "0000001001011110", -- t[606] = 0
      "000000" when "0000001001011111", -- t[607] = 0
      "000000" when "0000001001100000", -- t[608] = 0
      "000000" when "0000001001100001", -- t[609] = 0
      "000000" when "0000001001100010", -- t[610] = 0
      "000000" when "0000001001100011", -- t[611] = 0
      "000000" when "0000001001100100", -- t[612] = 0
      "000000" when "0000001001100101", -- t[613] = 0
      "000000" when "0000001001100110", -- t[614] = 0
      "000000" when "0000001001100111", -- t[615] = 0
      "000000" when "0000001001101000", -- t[616] = 0
      "000000" when "0000001001101001", -- t[617] = 0
      "000000" when "0000001001101010", -- t[618] = 0
      "000000" when "0000001001101011", -- t[619] = 0
      "000000" when "0000001001101100", -- t[620] = 0
      "000000" when "0000001001101101", -- t[621] = 0
      "000000" when "0000001001101110", -- t[622] = 0
      "000000" when "0000001001101111", -- t[623] = 0
      "000000" when "0000001001110000", -- t[624] = 0
      "000000" when "0000001001110001", -- t[625] = 0
      "000000" when "0000001001110010", -- t[626] = 0
      "000000" when "0000001001110011", -- t[627] = 0
      "000000" when "0000001001110100", -- t[628] = 0
      "000000" when "0000001001110101", -- t[629] = 0
      "000000" when "0000001001110110", -- t[630] = 0
      "000000" when "0000001001110111", -- t[631] = 0
      "000000" when "0000001001111000", -- t[632] = 0
      "000000" when "0000001001111001", -- t[633] = 0
      "000000" when "0000001001111010", -- t[634] = 0
      "000000" when "0000001001111011", -- t[635] = 0
      "000000" when "0000001001111100", -- t[636] = 0
      "000000" when "0000001001111101", -- t[637] = 0
      "000000" when "0000001001111110", -- t[638] = 0
      "000000" when "0000001001111111", -- t[639] = 0
      "000000" when "0000001010000000", -- t[640] = 0
      "000000" when "0000001010000001", -- t[641] = 0
      "000000" when "0000001010000010", -- t[642] = 0
      "000000" when "0000001010000011", -- t[643] = 0
      "000000" when "0000001010000100", -- t[644] = 0
      "000000" when "0000001010000101", -- t[645] = 0
      "000000" when "0000001010000110", -- t[646] = 0
      "000000" when "0000001010000111", -- t[647] = 0
      "000000" when "0000001010001000", -- t[648] = 0
      "000000" when "0000001010001001", -- t[649] = 0
      "000000" when "0000001010001010", -- t[650] = 0
      "000000" when "0000001010001011", -- t[651] = 0
      "000000" when "0000001010001100", -- t[652] = 0
      "000000" when "0000001010001101", -- t[653] = 0
      "000000" when "0000001010001110", -- t[654] = 0
      "000000" when "0000001010001111", -- t[655] = 0
      "000000" when "0000001010010000", -- t[656] = 0
      "000000" when "0000001010010001", -- t[657] = 0
      "000000" when "0000001010010010", -- t[658] = 0
      "000000" when "0000001010010011", -- t[659] = 0
      "000000" when "0000001010010100", -- t[660] = 0
      "000000" when "0000001010010101", -- t[661] = 0
      "000000" when "0000001010010110", -- t[662] = 0
      "000000" when "0000001010010111", -- t[663] = 0
      "000000" when "0000001010011000", -- t[664] = 0
      "000000" when "0000001010011001", -- t[665] = 0
      "000000" when "0000001010011010", -- t[666] = 0
      "000000" when "0000001010011011", -- t[667] = 0
      "000000" when "0000001010011100", -- t[668] = 0
      "000000" when "0000001010011101", -- t[669] = 0
      "000000" when "0000001010011110", -- t[670] = 0
      "000000" when "0000001010011111", -- t[671] = 0
      "000000" when "0000001010100000", -- t[672] = 0
      "000000" when "0000001010100001", -- t[673] = 0
      "000000" when "0000001010100010", -- t[674] = 0
      "000000" when "0000001010100011", -- t[675] = 0
      "000000" when "0000001010100100", -- t[676] = 0
      "000000" when "0000001010100101", -- t[677] = 0
      "000000" when "0000001010100110", -- t[678] = 0
      "000000" when "0000001010100111", -- t[679] = 0
      "000000" when "0000001010101000", -- t[680] = 0
      "000000" when "0000001010101001", -- t[681] = 0
      "000000" when "0000001010101010", -- t[682] = 0
      "000000" when "0000001010101011", -- t[683] = 0
      "000000" when "0000001010101100", -- t[684] = 0
      "000000" when "0000001010101101", -- t[685] = 0
      "000000" when "0000001010101110", -- t[686] = 0
      "000000" when "0000001010101111", -- t[687] = 0
      "000000" when "0000001010110000", -- t[688] = 0
      "000000" when "0000001010110001", -- t[689] = 0
      "000000" when "0000001010110010", -- t[690] = 0
      "000000" when "0000001010110011", -- t[691] = 0
      "000000" when "0000001010110100", -- t[692] = 0
      "000000" when "0000001010110101", -- t[693] = 0
      "000000" when "0000001010110110", -- t[694] = 0
      "000000" when "0000001010110111", -- t[695] = 0
      "000000" when "0000001010111000", -- t[696] = 0
      "000000" when "0000001010111001", -- t[697] = 0
      "000000" when "0000001010111010", -- t[698] = 0
      "000000" when "0000001010111011", -- t[699] = 0
      "000000" when "0000001010111100", -- t[700] = 0
      "000000" when "0000001010111101", -- t[701] = 0
      "000000" when "0000001010111110", -- t[702] = 0
      "000000" when "0000001010111111", -- t[703] = 0
      "000000" when "0000001011000000", -- t[704] = 0
      "000000" when "0000001011000001", -- t[705] = 0
      "000000" when "0000001011000010", -- t[706] = 0
      "000000" when "0000001011000011", -- t[707] = 0
      "000000" when "0000001011000100", -- t[708] = 0
      "000000" when "0000001011000101", -- t[709] = 0
      "000000" when "0000001011000110", -- t[710] = 0
      "000000" when "0000001011000111", -- t[711] = 0
      "000000" when "0000001011001000", -- t[712] = 0
      "000000" when "0000001011001001", -- t[713] = 0
      "000000" when "0000001011001010", -- t[714] = 0
      "000000" when "0000001011001011", -- t[715] = 0
      "000000" when "0000001011001100", -- t[716] = 0
      "000000" when "0000001011001101", -- t[717] = 0
      "000000" when "0000001011001110", -- t[718] = 0
      "000000" when "0000001011001111", -- t[719] = 0
      "000000" when "0000001011010000", -- t[720] = 0
      "000000" when "0000001011010001", -- t[721] = 0
      "000000" when "0000001011010010", -- t[722] = 0
      "000000" when "0000001011010011", -- t[723] = 0
      "000000" when "0000001011010100", -- t[724] = 0
      "000000" when "0000001011010101", -- t[725] = 0
      "000000" when "0000001011010110", -- t[726] = 0
      "000000" when "0000001011010111", -- t[727] = 0
      "000000" when "0000001011011000", -- t[728] = 0
      "000000" when "0000001011011001", -- t[729] = 0
      "000000" when "0000001011011010", -- t[730] = 0
      "000000" when "0000001011011011", -- t[731] = 0
      "000000" when "0000001011011100", -- t[732] = 0
      "000000" when "0000001011011101", -- t[733] = 0
      "000000" when "0000001011011110", -- t[734] = 0
      "000000" when "0000001011011111", -- t[735] = 0
      "000000" when "0000001011100000", -- t[736] = 0
      "000000" when "0000001011100001", -- t[737] = 0
      "000000" when "0000001011100010", -- t[738] = 0
      "000000" when "0000001011100011", -- t[739] = 0
      "000000" when "0000001011100100", -- t[740] = 0
      "000000" when "0000001011100101", -- t[741] = 0
      "000000" when "0000001011100110", -- t[742] = 0
      "000000" when "0000001011100111", -- t[743] = 0
      "000000" when "0000001011101000", -- t[744] = 0
      "000000" when "0000001011101001", -- t[745] = 0
      "000000" when "0000001011101010", -- t[746] = 0
      "000000" when "0000001011101011", -- t[747] = 0
      "000000" when "0000001011101100", -- t[748] = 0
      "000000" when "0000001011101101", -- t[749] = 0
      "000000" when "0000001011101110", -- t[750] = 0
      "000000" when "0000001011101111", -- t[751] = 0
      "000000" when "0000001011110000", -- t[752] = 0
      "000000" when "0000001011110001", -- t[753] = 0
      "000000" when "0000001011110010", -- t[754] = 0
      "000000" when "0000001011110011", -- t[755] = 0
      "000000" when "0000001011110100", -- t[756] = 0
      "000000" when "0000001011110101", -- t[757] = 0
      "000000" when "0000001011110110", -- t[758] = 0
      "000000" when "0000001011110111", -- t[759] = 0
      "000000" when "0000001011111000", -- t[760] = 0
      "000000" when "0000001011111001", -- t[761] = 0
      "000000" when "0000001011111010", -- t[762] = 0
      "000000" when "0000001011111011", -- t[763] = 0
      "000000" when "0000001011111100", -- t[764] = 0
      "000000" when "0000001011111101", -- t[765] = 0
      "000000" when "0000001011111110", -- t[766] = 0
      "000000" when "0000001011111111", -- t[767] = 0
      "000000" when "0000001100000000", -- t[768] = 0
      "000000" when "0000001100000001", -- t[769] = 0
      "000000" when "0000001100000010", -- t[770] = 0
      "000000" when "0000001100000011", -- t[771] = 0
      "000000" when "0000001100000100", -- t[772] = 0
      "000000" when "0000001100000101", -- t[773] = 0
      "000000" when "0000001100000110", -- t[774] = 0
      "000000" when "0000001100000111", -- t[775] = 0
      "000000" when "0000001100001000", -- t[776] = 0
      "000000" when "0000001100001001", -- t[777] = 0
      "000000" when "0000001100001010", -- t[778] = 0
      "000000" when "0000001100001011", -- t[779] = 0
      "000000" when "0000001100001100", -- t[780] = 0
      "000000" when "0000001100001101", -- t[781] = 0
      "000000" when "0000001100001110", -- t[782] = 0
      "000000" when "0000001100001111", -- t[783] = 0
      "000000" when "0000001100010000", -- t[784] = 0
      "000000" when "0000001100010001", -- t[785] = 0
      "000000" when "0000001100010010", -- t[786] = 0
      "000000" when "0000001100010011", -- t[787] = 0
      "000000" when "0000001100010100", -- t[788] = 0
      "000000" when "0000001100010101", -- t[789] = 0
      "000000" when "0000001100010110", -- t[790] = 0
      "000000" when "0000001100010111", -- t[791] = 0
      "000000" when "0000001100011000", -- t[792] = 0
      "000000" when "0000001100011001", -- t[793] = 0
      "000000" when "0000001100011010", -- t[794] = 0
      "000000" when "0000001100011011", -- t[795] = 0
      "000000" when "0000001100011100", -- t[796] = 0
      "000000" when "0000001100011101", -- t[797] = 0
      "000000" when "0000001100011110", -- t[798] = 0
      "000000" when "0000001100011111", -- t[799] = 0
      "000000" when "0000001100100000", -- t[800] = 0
      "000000" when "0000001100100001", -- t[801] = 0
      "000000" when "0000001100100010", -- t[802] = 0
      "000000" when "0000001100100011", -- t[803] = 0
      "000000" when "0000001100100100", -- t[804] = 0
      "000000" when "0000001100100101", -- t[805] = 0
      "000000" when "0000001100100110", -- t[806] = 0
      "000000" when "0000001100100111", -- t[807] = 0
      "000000" when "0000001100101000", -- t[808] = 0
      "000000" when "0000001100101001", -- t[809] = 0
      "000000" when "0000001100101010", -- t[810] = 0
      "000000" when "0000001100101011", -- t[811] = 0
      "000000" when "0000001100101100", -- t[812] = 0
      "000000" when "0000001100101101", -- t[813] = 0
      "000000" when "0000001100101110", -- t[814] = 0
      "000000" when "0000001100101111", -- t[815] = 0
      "000000" when "0000001100110000", -- t[816] = 0
      "000000" when "0000001100110001", -- t[817] = 0
      "000000" when "0000001100110010", -- t[818] = 0
      "000000" when "0000001100110011", -- t[819] = 0
      "000000" when "0000001100110100", -- t[820] = 0
      "000000" when "0000001100110101", -- t[821] = 0
      "000000" when "0000001100110110", -- t[822] = 0
      "000000" when "0000001100110111", -- t[823] = 0
      "000000" when "0000001100111000", -- t[824] = 0
      "000000" when "0000001100111001", -- t[825] = 0
      "000000" when "0000001100111010", -- t[826] = 0
      "000000" when "0000001100111011", -- t[827] = 0
      "000000" when "0000001100111100", -- t[828] = 0
      "000000" when "0000001100111101", -- t[829] = 0
      "000000" when "0000001100111110", -- t[830] = 0
      "000000" when "0000001100111111", -- t[831] = 0
      "000000" when "0000001101000000", -- t[832] = 0
      "000000" when "0000001101000001", -- t[833] = 0
      "000000" when "0000001101000010", -- t[834] = 0
      "000000" when "0000001101000011", -- t[835] = 0
      "000000" when "0000001101000100", -- t[836] = 0
      "000000" when "0000001101000101", -- t[837] = 0
      "000000" when "0000001101000110", -- t[838] = 0
      "000000" when "0000001101000111", -- t[839] = 0
      "000000" when "0000001101001000", -- t[840] = 0
      "000000" when "0000001101001001", -- t[841] = 0
      "000000" when "0000001101001010", -- t[842] = 0
      "000000" when "0000001101001011", -- t[843] = 0
      "000000" when "0000001101001100", -- t[844] = 0
      "000000" when "0000001101001101", -- t[845] = 0
      "000000" when "0000001101001110", -- t[846] = 0
      "000000" when "0000001101001111", -- t[847] = 0
      "000000" when "0000001101010000", -- t[848] = 0
      "000000" when "0000001101010001", -- t[849] = 0
      "000000" when "0000001101010010", -- t[850] = 0
      "000000" when "0000001101010011", -- t[851] = 0
      "000000" when "0000001101010100", -- t[852] = 0
      "000000" when "0000001101010101", -- t[853] = 0
      "000000" when "0000001101010110", -- t[854] = 0
      "000000" when "0000001101010111", -- t[855] = 0
      "000000" when "0000001101011000", -- t[856] = 0
      "000000" when "0000001101011001", -- t[857] = 0
      "000000" when "0000001101011010", -- t[858] = 0
      "000000" when "0000001101011011", -- t[859] = 0
      "000000" when "0000001101011100", -- t[860] = 0
      "000000" when "0000001101011101", -- t[861] = 0
      "000000" when "0000001101011110", -- t[862] = 0
      "000000" when "0000001101011111", -- t[863] = 0
      "000000" when "0000001101100000", -- t[864] = 0
      "000000" when "0000001101100001", -- t[865] = 0
      "000000" when "0000001101100010", -- t[866] = 0
      "000000" when "0000001101100011", -- t[867] = 0
      "000000" when "0000001101100100", -- t[868] = 0
      "000000" when "0000001101100101", -- t[869] = 0
      "000000" when "0000001101100110", -- t[870] = 0
      "000000" when "0000001101100111", -- t[871] = 0
      "000000" when "0000001101101000", -- t[872] = 0
      "000000" when "0000001101101001", -- t[873] = 0
      "000000" when "0000001101101010", -- t[874] = 0
      "000000" when "0000001101101011", -- t[875] = 0
      "000000" when "0000001101101100", -- t[876] = 0
      "000000" when "0000001101101101", -- t[877] = 0
      "000000" when "0000001101101110", -- t[878] = 0
      "000000" when "0000001101101111", -- t[879] = 0
      "000000" when "0000001101110000", -- t[880] = 0
      "000000" when "0000001101110001", -- t[881] = 0
      "000000" when "0000001101110010", -- t[882] = 0
      "000000" when "0000001101110011", -- t[883] = 0
      "000000" when "0000001101110100", -- t[884] = 0
      "000000" when "0000001101110101", -- t[885] = 0
      "000000" when "0000001101110110", -- t[886] = 0
      "000000" when "0000001101110111", -- t[887] = 0
      "000000" when "0000001101111000", -- t[888] = 0
      "000000" when "0000001101111001", -- t[889] = 0
      "000000" when "0000001101111010", -- t[890] = 0
      "000000" when "0000001101111011", -- t[891] = 0
      "000000" when "0000001101111100", -- t[892] = 0
      "000000" when "0000001101111101", -- t[893] = 0
      "000000" when "0000001101111110", -- t[894] = 0
      "000000" when "0000001101111111", -- t[895] = 0
      "000000" when "0000001110000000", -- t[896] = 0
      "000000" when "0000001110000001", -- t[897] = 0
      "000000" when "0000001110000010", -- t[898] = 0
      "000000" when "0000001110000011", -- t[899] = 0
      "000000" when "0000001110000100", -- t[900] = 0
      "000000" when "0000001110000101", -- t[901] = 0
      "000000" when "0000001110000110", -- t[902] = 0
      "000000" when "0000001110000111", -- t[903] = 0
      "000000" when "0000001110001000", -- t[904] = 0
      "000000" when "0000001110001001", -- t[905] = 0
      "000000" when "0000001110001010", -- t[906] = 0
      "000000" when "0000001110001011", -- t[907] = 0
      "000000" when "0000001110001100", -- t[908] = 0
      "000000" when "0000001110001101", -- t[909] = 0
      "000000" when "0000001110001110", -- t[910] = 0
      "000000" when "0000001110001111", -- t[911] = 0
      "000000" when "0000001110010000", -- t[912] = 0
      "000000" when "0000001110010001", -- t[913] = 0
      "000000" when "0000001110010010", -- t[914] = 0
      "000000" when "0000001110010011", -- t[915] = 0
      "000000" when "0000001110010100", -- t[916] = 0
      "000000" when "0000001110010101", -- t[917] = 0
      "000000" when "0000001110010110", -- t[918] = 0
      "000000" when "0000001110010111", -- t[919] = 0
      "000000" when "0000001110011000", -- t[920] = 0
      "000000" when "0000001110011001", -- t[921] = 0
      "000000" when "0000001110011010", -- t[922] = 0
      "000000" when "0000001110011011", -- t[923] = 0
      "000000" when "0000001110011100", -- t[924] = 0
      "000000" when "0000001110011101", -- t[925] = 0
      "000000" when "0000001110011110", -- t[926] = 0
      "000000" when "0000001110011111", -- t[927] = 0
      "000000" when "0000001110100000", -- t[928] = 0
      "000000" when "0000001110100001", -- t[929] = 0
      "000000" when "0000001110100010", -- t[930] = 0
      "000000" when "0000001110100011", -- t[931] = 0
      "000000" when "0000001110100100", -- t[932] = 0
      "000000" when "0000001110100101", -- t[933] = 0
      "000000" when "0000001110100110", -- t[934] = 0
      "000000" when "0000001110100111", -- t[935] = 0
      "000000" when "0000001110101000", -- t[936] = 0
      "000000" when "0000001110101001", -- t[937] = 0
      "000000" when "0000001110101010", -- t[938] = 0
      "000000" when "0000001110101011", -- t[939] = 0
      "000000" when "0000001110101100", -- t[940] = 0
      "000000" when "0000001110101101", -- t[941] = 0
      "000000" when "0000001110101110", -- t[942] = 0
      "000000" when "0000001110101111", -- t[943] = 0
      "000000" when "0000001110110000", -- t[944] = 0
      "000000" when "0000001110110001", -- t[945] = 0
      "000000" when "0000001110110010", -- t[946] = 0
      "000000" when "0000001110110011", -- t[947] = 0
      "000000" when "0000001110110100", -- t[948] = 0
      "000000" when "0000001110110101", -- t[949] = 0
      "000000" when "0000001110110110", -- t[950] = 0
      "000000" when "0000001110110111", -- t[951] = 0
      "000000" when "0000001110111000", -- t[952] = 0
      "000000" when "0000001110111001", -- t[953] = 0
      "000000" when "0000001110111010", -- t[954] = 0
      "000000" when "0000001110111011", -- t[955] = 0
      "000000" when "0000001110111100", -- t[956] = 0
      "000000" when "0000001110111101", -- t[957] = 0
      "000000" when "0000001110111110", -- t[958] = 0
      "000000" when "0000001110111111", -- t[959] = 0
      "000000" when "0000001111000000", -- t[960] = 0
      "000000" when "0000001111000001", -- t[961] = 0
      "000000" when "0000001111000010", -- t[962] = 0
      "000000" when "0000001111000011", -- t[963] = 0
      "000000" when "0000001111000100", -- t[964] = 0
      "000000" when "0000001111000101", -- t[965] = 0
      "000000" when "0000001111000110", -- t[966] = 0
      "000000" when "0000001111000111", -- t[967] = 0
      "000000" when "0000001111001000", -- t[968] = 0
      "000000" when "0000001111001001", -- t[969] = 0
      "000000" when "0000001111001010", -- t[970] = 0
      "000000" when "0000001111001011", -- t[971] = 0
      "000000" when "0000001111001100", -- t[972] = 0
      "000000" when "0000001111001101", -- t[973] = 0
      "000000" when "0000001111001110", -- t[974] = 0
      "000000" when "0000001111001111", -- t[975] = 0
      "000000" when "0000001111010000", -- t[976] = 0
      "000000" when "0000001111010001", -- t[977] = 0
      "000000" when "0000001111010010", -- t[978] = 0
      "000000" when "0000001111010011", -- t[979] = 0
      "000000" when "0000001111010100", -- t[980] = 0
      "000000" when "0000001111010101", -- t[981] = 0
      "000000" when "0000001111010110", -- t[982] = 0
      "000000" when "0000001111010111", -- t[983] = 0
      "000000" when "0000001111011000", -- t[984] = 0
      "000000" when "0000001111011001", -- t[985] = 0
      "000000" when "0000001111011010", -- t[986] = 0
      "000000" when "0000001111011011", -- t[987] = 0
      "000000" when "0000001111011100", -- t[988] = 0
      "000000" when "0000001111011101", -- t[989] = 0
      "000000" when "0000001111011110", -- t[990] = 0
      "000000" when "0000001111011111", -- t[991] = 0
      "000000" when "0000001111100000", -- t[992] = 0
      "000000" when "0000001111100001", -- t[993] = 0
      "000000" when "0000001111100010", -- t[994] = 0
      "000000" when "0000001111100011", -- t[995] = 0
      "000000" when "0000001111100100", -- t[996] = 0
      "000000" when "0000001111100101", -- t[997] = 0
      "000000" when "0000001111100110", -- t[998] = 0
      "000000" when "0000001111100111", -- t[999] = 0
      "000000" when "0000001111101000", -- t[1000] = 0
      "000000" when "0000001111101001", -- t[1001] = 0
      "000000" when "0000001111101010", -- t[1002] = 0
      "000000" when "0000001111101011", -- t[1003] = 0
      "000000" when "0000001111101100", -- t[1004] = 0
      "000000" when "0000001111101101", -- t[1005] = 0
      "000000" when "0000001111101110", -- t[1006] = 0
      "000000" when "0000001111101111", -- t[1007] = 0
      "000000" when "0000001111110000", -- t[1008] = 0
      "000000" when "0000001111110001", -- t[1009] = 0
      "000000" when "0000001111110010", -- t[1010] = 0
      "000000" when "0000001111110011", -- t[1011] = 0
      "000000" when "0000001111110100", -- t[1012] = 0
      "000000" when "0000001111110101", -- t[1013] = 0
      "000000" when "0000001111110110", -- t[1014] = 0
      "000000" when "0000001111110111", -- t[1015] = 0
      "000000" when "0000001111111000", -- t[1016] = 0
      "000000" when "0000001111111001", -- t[1017] = 0
      "000000" when "0000001111111010", -- t[1018] = 0
      "000000" when "0000001111111011", -- t[1019] = 0
      "000000" when "0000001111111100", -- t[1020] = 0
      "000000" when "0000001111111101", -- t[1021] = 0
      "000000" when "0000001111111110", -- t[1022] = 0
      "000000" when "0000001111111111", -- t[1023] = 0
      "000000" when "0000010000000000", -- t[1024] = 0
      "000000" when "0000010000000001", -- t[1025] = 0
      "000000" when "0000010000000010", -- t[1026] = 0
      "000000" when "0000010000000011", -- t[1027] = 0
      "000000" when "0000010000000100", -- t[1028] = 0
      "000000" when "0000010000000101", -- t[1029] = 0
      "000000" when "0000010000000110", -- t[1030] = 0
      "000000" when "0000010000000111", -- t[1031] = 0
      "000000" when "0000010000001000", -- t[1032] = 0
      "000000" when "0000010000001001", -- t[1033] = 0
      "000000" when "0000010000001010", -- t[1034] = 0
      "000000" when "0000010000001011", -- t[1035] = 0
      "000000" when "0000010000001100", -- t[1036] = 0
      "000000" when "0000010000001101", -- t[1037] = 0
      "000000" when "0000010000001110", -- t[1038] = 0
      "000000" when "0000010000001111", -- t[1039] = 0
      "000000" when "0000010000010000", -- t[1040] = 0
      "000000" when "0000010000010001", -- t[1041] = 0
      "000000" when "0000010000010010", -- t[1042] = 0
      "000000" when "0000010000010011", -- t[1043] = 0
      "000000" when "0000010000010100", -- t[1044] = 0
      "000000" when "0000010000010101", -- t[1045] = 0
      "000000" when "0000010000010110", -- t[1046] = 0
      "000000" when "0000010000010111", -- t[1047] = 0
      "000000" when "0000010000011000", -- t[1048] = 0
      "000000" when "0000010000011001", -- t[1049] = 0
      "000000" when "0000010000011010", -- t[1050] = 0
      "000000" when "0000010000011011", -- t[1051] = 0
      "000000" when "0000010000011100", -- t[1052] = 0
      "000000" when "0000010000011101", -- t[1053] = 0
      "000000" when "0000010000011110", -- t[1054] = 0
      "000000" when "0000010000011111", -- t[1055] = 0
      "000000" when "0000010000100000", -- t[1056] = 0
      "000000" when "0000010000100001", -- t[1057] = 0
      "000000" when "0000010000100010", -- t[1058] = 0
      "000000" when "0000010000100011", -- t[1059] = 0
      "000000" when "0000010000100100", -- t[1060] = 0
      "000000" when "0000010000100101", -- t[1061] = 0
      "000000" when "0000010000100110", -- t[1062] = 0
      "000000" when "0000010000100111", -- t[1063] = 0
      "000000" when "0000010000101000", -- t[1064] = 0
      "000000" when "0000010000101001", -- t[1065] = 0
      "000000" when "0000010000101010", -- t[1066] = 0
      "000000" when "0000010000101011", -- t[1067] = 0
      "000000" when "0000010000101100", -- t[1068] = 0
      "000000" when "0000010000101101", -- t[1069] = 0
      "000000" when "0000010000101110", -- t[1070] = 0
      "000000" when "0000010000101111", -- t[1071] = 0
      "000000" when "0000010000110000", -- t[1072] = 0
      "000000" when "0000010000110001", -- t[1073] = 0
      "000000" when "0000010000110010", -- t[1074] = 0
      "000000" when "0000010000110011", -- t[1075] = 0
      "000000" when "0000010000110100", -- t[1076] = 0
      "000000" when "0000010000110101", -- t[1077] = 0
      "000000" when "0000010000110110", -- t[1078] = 0
      "000000" when "0000010000110111", -- t[1079] = 0
      "000000" when "0000010000111000", -- t[1080] = 0
      "000000" when "0000010000111001", -- t[1081] = 0
      "000000" when "0000010000111010", -- t[1082] = 0
      "000000" when "0000010000111011", -- t[1083] = 0
      "000000" when "0000010000111100", -- t[1084] = 0
      "000000" when "0000010000111101", -- t[1085] = 0
      "000000" when "0000010000111110", -- t[1086] = 0
      "000000" when "0000010000111111", -- t[1087] = 0
      "000000" when "0000010001000000", -- t[1088] = 0
      "000000" when "0000010001000001", -- t[1089] = 0
      "000000" when "0000010001000010", -- t[1090] = 0
      "000000" when "0000010001000011", -- t[1091] = 0
      "000000" when "0000010001000100", -- t[1092] = 0
      "000000" when "0000010001000101", -- t[1093] = 0
      "000000" when "0000010001000110", -- t[1094] = 0
      "000000" when "0000010001000111", -- t[1095] = 0
      "000000" when "0000010001001000", -- t[1096] = 0
      "000000" when "0000010001001001", -- t[1097] = 0
      "000000" when "0000010001001010", -- t[1098] = 0
      "000000" when "0000010001001011", -- t[1099] = 0
      "000000" when "0000010001001100", -- t[1100] = 0
      "000000" when "0000010001001101", -- t[1101] = 0
      "000000" when "0000010001001110", -- t[1102] = 0
      "000000" when "0000010001001111", -- t[1103] = 0
      "000000" when "0000010001010000", -- t[1104] = 0
      "000000" when "0000010001010001", -- t[1105] = 0
      "000000" when "0000010001010010", -- t[1106] = 0
      "000000" when "0000010001010011", -- t[1107] = 0
      "000000" when "0000010001010100", -- t[1108] = 0
      "000000" when "0000010001010101", -- t[1109] = 0
      "000000" when "0000010001010110", -- t[1110] = 0
      "000000" when "0000010001010111", -- t[1111] = 0
      "000000" when "0000010001011000", -- t[1112] = 0
      "000000" when "0000010001011001", -- t[1113] = 0
      "000000" when "0000010001011010", -- t[1114] = 0
      "000000" when "0000010001011011", -- t[1115] = 0
      "000000" when "0000010001011100", -- t[1116] = 0
      "000000" when "0000010001011101", -- t[1117] = 0
      "000000" when "0000010001011110", -- t[1118] = 0
      "000000" when "0000010001011111", -- t[1119] = 0
      "000000" when "0000010001100000", -- t[1120] = 0
      "000000" when "0000010001100001", -- t[1121] = 0
      "000000" when "0000010001100010", -- t[1122] = 0
      "000000" when "0000010001100011", -- t[1123] = 0
      "000000" when "0000010001100100", -- t[1124] = 0
      "000000" when "0000010001100101", -- t[1125] = 0
      "000000" when "0000010001100110", -- t[1126] = 0
      "000000" when "0000010001100111", -- t[1127] = 0
      "000000" when "0000010001101000", -- t[1128] = 0
      "000000" when "0000010001101001", -- t[1129] = 0
      "000000" when "0000010001101010", -- t[1130] = 0
      "000000" when "0000010001101011", -- t[1131] = 0
      "000000" when "0000010001101100", -- t[1132] = 0
      "000000" when "0000010001101101", -- t[1133] = 0
      "000000" when "0000010001101110", -- t[1134] = 0
      "000000" when "0000010001101111", -- t[1135] = 0
      "000000" when "0000010001110000", -- t[1136] = 0
      "000000" when "0000010001110001", -- t[1137] = 0
      "000000" when "0000010001110010", -- t[1138] = 0
      "000000" when "0000010001110011", -- t[1139] = 0
      "000000" when "0000010001110100", -- t[1140] = 0
      "000000" when "0000010001110101", -- t[1141] = 0
      "000000" when "0000010001110110", -- t[1142] = 0
      "000000" when "0000010001110111", -- t[1143] = 0
      "000000" when "0000010001111000", -- t[1144] = 0
      "000000" when "0000010001111001", -- t[1145] = 0
      "000000" when "0000010001111010", -- t[1146] = 0
      "000000" when "0000010001111011", -- t[1147] = 0
      "000000" when "0000010001111100", -- t[1148] = 0
      "000000" when "0000010001111101", -- t[1149] = 0
      "000000" when "0000010001111110", -- t[1150] = 0
      "000000" when "0000010001111111", -- t[1151] = 0
      "000000" when "0000010010000000", -- t[1152] = 0
      "000000" when "0000010010000001", -- t[1153] = 0
      "000000" when "0000010010000010", -- t[1154] = 0
      "000000" when "0000010010000011", -- t[1155] = 0
      "000000" when "0000010010000100", -- t[1156] = 0
      "000000" when "0000010010000101", -- t[1157] = 0
      "000000" when "0000010010000110", -- t[1158] = 0
      "000000" when "0000010010000111", -- t[1159] = 0
      "000000" when "0000010010001000", -- t[1160] = 0
      "000000" when "0000010010001001", -- t[1161] = 0
      "000000" when "0000010010001010", -- t[1162] = 0
      "000000" when "0000010010001011", -- t[1163] = 0
      "000000" when "0000010010001100", -- t[1164] = 0
      "000000" when "0000010010001101", -- t[1165] = 0
      "000000" when "0000010010001110", -- t[1166] = 0
      "000000" when "0000010010001111", -- t[1167] = 0
      "000000" when "0000010010010000", -- t[1168] = 0
      "000000" when "0000010010010001", -- t[1169] = 0
      "000000" when "0000010010010010", -- t[1170] = 0
      "000000" when "0000010010010011", -- t[1171] = 0
      "000000" when "0000010010010100", -- t[1172] = 0
      "000000" when "0000010010010101", -- t[1173] = 0
      "000000" when "0000010010010110", -- t[1174] = 0
      "000000" when "0000010010010111", -- t[1175] = 0
      "000000" when "0000010010011000", -- t[1176] = 0
      "000000" when "0000010010011001", -- t[1177] = 0
      "000000" when "0000010010011010", -- t[1178] = 0
      "000000" when "0000010010011011", -- t[1179] = 0
      "000000" when "0000010010011100", -- t[1180] = 0
      "000000" when "0000010010011101", -- t[1181] = 0
      "000000" when "0000010010011110", -- t[1182] = 0
      "000000" when "0000010010011111", -- t[1183] = 0
      "000000" when "0000010010100000", -- t[1184] = 0
      "000000" when "0000010010100001", -- t[1185] = 0
      "000000" when "0000010010100010", -- t[1186] = 0
      "000000" when "0000010010100011", -- t[1187] = 0
      "000000" when "0000010010100100", -- t[1188] = 0
      "000000" when "0000010010100101", -- t[1189] = 0
      "000000" when "0000010010100110", -- t[1190] = 0
      "000000" when "0000010010100111", -- t[1191] = 0
      "000000" when "0000010010101000", -- t[1192] = 0
      "000000" when "0000010010101001", -- t[1193] = 0
      "000000" when "0000010010101010", -- t[1194] = 0
      "000000" when "0000010010101011", -- t[1195] = 0
      "000000" when "0000010010101100", -- t[1196] = 0
      "000000" when "0000010010101101", -- t[1197] = 0
      "000000" when "0000010010101110", -- t[1198] = 0
      "000000" when "0000010010101111", -- t[1199] = 0
      "000000" when "0000010010110000", -- t[1200] = 0
      "000000" when "0000010010110001", -- t[1201] = 0
      "000000" when "0000010010110010", -- t[1202] = 0
      "000000" when "0000010010110011", -- t[1203] = 0
      "000000" when "0000010010110100", -- t[1204] = 0
      "000000" when "0000010010110101", -- t[1205] = 0
      "000000" when "0000010010110110", -- t[1206] = 0
      "000000" when "0000010010110111", -- t[1207] = 0
      "000000" when "0000010010111000", -- t[1208] = 0
      "000000" when "0000010010111001", -- t[1209] = 0
      "000000" when "0000010010111010", -- t[1210] = 0
      "000000" when "0000010010111011", -- t[1211] = 0
      "000000" when "0000010010111100", -- t[1212] = 0
      "000000" when "0000010010111101", -- t[1213] = 0
      "000000" when "0000010010111110", -- t[1214] = 0
      "000000" when "0000010010111111", -- t[1215] = 0
      "000000" when "0000010011000000", -- t[1216] = 0
      "000000" when "0000010011000001", -- t[1217] = 0
      "000000" when "0000010011000010", -- t[1218] = 0
      "000000" when "0000010011000011", -- t[1219] = 0
      "000000" when "0000010011000100", -- t[1220] = 0
      "000000" when "0000010011000101", -- t[1221] = 0
      "000000" when "0000010011000110", -- t[1222] = 0
      "000000" when "0000010011000111", -- t[1223] = 0
      "000000" when "0000010011001000", -- t[1224] = 0
      "000000" when "0000010011001001", -- t[1225] = 0
      "000000" when "0000010011001010", -- t[1226] = 0
      "000000" when "0000010011001011", -- t[1227] = 0
      "000000" when "0000010011001100", -- t[1228] = 0
      "000000" when "0000010011001101", -- t[1229] = 0
      "000000" when "0000010011001110", -- t[1230] = 0
      "000000" when "0000010011001111", -- t[1231] = 0
      "000000" when "0000010011010000", -- t[1232] = 0
      "000000" when "0000010011010001", -- t[1233] = 0
      "000000" when "0000010011010010", -- t[1234] = 0
      "000000" when "0000010011010011", -- t[1235] = 0
      "000000" when "0000010011010100", -- t[1236] = 0
      "000000" when "0000010011010101", -- t[1237] = 0
      "000000" when "0000010011010110", -- t[1238] = 0
      "000000" when "0000010011010111", -- t[1239] = 0
      "000000" when "0000010011011000", -- t[1240] = 0
      "000000" when "0000010011011001", -- t[1241] = 0
      "000000" when "0000010011011010", -- t[1242] = 0
      "000000" when "0000010011011011", -- t[1243] = 0
      "000000" when "0000010011011100", -- t[1244] = 0
      "000000" when "0000010011011101", -- t[1245] = 0
      "000000" when "0000010011011110", -- t[1246] = 0
      "000000" when "0000010011011111", -- t[1247] = 0
      "000000" when "0000010011100000", -- t[1248] = 0
      "000000" when "0000010011100001", -- t[1249] = 0
      "000000" when "0000010011100010", -- t[1250] = 0
      "000000" when "0000010011100011", -- t[1251] = 0
      "000000" when "0000010011100100", -- t[1252] = 0
      "000000" when "0000010011100101", -- t[1253] = 0
      "000000" when "0000010011100110", -- t[1254] = 0
      "000000" when "0000010011100111", -- t[1255] = 0
      "000000" when "0000010011101000", -- t[1256] = 0
      "000000" when "0000010011101001", -- t[1257] = 0
      "000000" when "0000010011101010", -- t[1258] = 0
      "000000" when "0000010011101011", -- t[1259] = 0
      "000000" when "0000010011101100", -- t[1260] = 0
      "000000" when "0000010011101101", -- t[1261] = 0
      "000000" when "0000010011101110", -- t[1262] = 0
      "000000" when "0000010011101111", -- t[1263] = 0
      "000000" when "0000010011110000", -- t[1264] = 0
      "000000" when "0000010011110001", -- t[1265] = 0
      "000000" when "0000010011110010", -- t[1266] = 0
      "000000" when "0000010011110011", -- t[1267] = 0
      "000000" when "0000010011110100", -- t[1268] = 0
      "000000" when "0000010011110101", -- t[1269] = 0
      "000000" when "0000010011110110", -- t[1270] = 0
      "000000" when "0000010011110111", -- t[1271] = 0
      "000000" when "0000010011111000", -- t[1272] = 0
      "000000" when "0000010011111001", -- t[1273] = 0
      "000000" when "0000010011111010", -- t[1274] = 0
      "000000" when "0000010011111011", -- t[1275] = 0
      "000000" when "0000010011111100", -- t[1276] = 0
      "000000" when "0000010011111101", -- t[1277] = 0
      "000000" when "0000010011111110", -- t[1278] = 0
      "000000" when "0000010011111111", -- t[1279] = 0
      "000000" when "0000010100000000", -- t[1280] = 0
      "000000" when "0000010100000001", -- t[1281] = 0
      "000000" when "0000010100000010", -- t[1282] = 0
      "000000" when "0000010100000011", -- t[1283] = 0
      "000000" when "0000010100000100", -- t[1284] = 0
      "000000" when "0000010100000101", -- t[1285] = 0
      "000000" when "0000010100000110", -- t[1286] = 0
      "000000" when "0000010100000111", -- t[1287] = 0
      "000000" when "0000010100001000", -- t[1288] = 0
      "000000" when "0000010100001001", -- t[1289] = 0
      "000000" when "0000010100001010", -- t[1290] = 0
      "000000" when "0000010100001011", -- t[1291] = 0
      "000000" when "0000010100001100", -- t[1292] = 0
      "000000" when "0000010100001101", -- t[1293] = 0
      "000000" when "0000010100001110", -- t[1294] = 0
      "000000" when "0000010100001111", -- t[1295] = 0
      "000000" when "0000010100010000", -- t[1296] = 0
      "000000" when "0000010100010001", -- t[1297] = 0
      "000000" when "0000010100010010", -- t[1298] = 0
      "000000" when "0000010100010011", -- t[1299] = 0
      "000000" when "0000010100010100", -- t[1300] = 0
      "000000" when "0000010100010101", -- t[1301] = 0
      "000000" when "0000010100010110", -- t[1302] = 0
      "000000" when "0000010100010111", -- t[1303] = 0
      "000000" when "0000010100011000", -- t[1304] = 0
      "000000" when "0000010100011001", -- t[1305] = 0
      "000000" when "0000010100011010", -- t[1306] = 0
      "000000" when "0000010100011011", -- t[1307] = 0
      "000000" when "0000010100011100", -- t[1308] = 0
      "000000" when "0000010100011101", -- t[1309] = 0
      "000000" when "0000010100011110", -- t[1310] = 0
      "000000" when "0000010100011111", -- t[1311] = 0
      "000000" when "0000010100100000", -- t[1312] = 0
      "000000" when "0000010100100001", -- t[1313] = 0
      "000000" when "0000010100100010", -- t[1314] = 0
      "000000" when "0000010100100011", -- t[1315] = 0
      "000000" when "0000010100100100", -- t[1316] = 0
      "000000" when "0000010100100101", -- t[1317] = 0
      "000000" when "0000010100100110", -- t[1318] = 0
      "000000" when "0000010100100111", -- t[1319] = 0
      "000000" when "0000010100101000", -- t[1320] = 0
      "000000" when "0000010100101001", -- t[1321] = 0
      "000000" when "0000010100101010", -- t[1322] = 0
      "000000" when "0000010100101011", -- t[1323] = 0
      "000000" when "0000010100101100", -- t[1324] = 0
      "000000" when "0000010100101101", -- t[1325] = 0
      "000000" when "0000010100101110", -- t[1326] = 0
      "000000" when "0000010100101111", -- t[1327] = 0
      "000000" when "0000010100110000", -- t[1328] = 0
      "000000" when "0000010100110001", -- t[1329] = 0
      "000000" when "0000010100110010", -- t[1330] = 0
      "000000" when "0000010100110011", -- t[1331] = 0
      "000000" when "0000010100110100", -- t[1332] = 0
      "000000" when "0000010100110101", -- t[1333] = 0
      "000000" when "0000010100110110", -- t[1334] = 0
      "000000" when "0000010100110111", -- t[1335] = 0
      "000000" when "0000010100111000", -- t[1336] = 0
      "000000" when "0000010100111001", -- t[1337] = 0
      "000000" when "0000010100111010", -- t[1338] = 0
      "000000" when "0000010100111011", -- t[1339] = 0
      "000000" when "0000010100111100", -- t[1340] = 0
      "000000" when "0000010100111101", -- t[1341] = 0
      "000000" when "0000010100111110", -- t[1342] = 0
      "000000" when "0000010100111111", -- t[1343] = 0
      "000000" when "0000010101000000", -- t[1344] = 0
      "000000" when "0000010101000001", -- t[1345] = 0
      "000000" when "0000010101000010", -- t[1346] = 0
      "000000" when "0000010101000011", -- t[1347] = 0
      "000000" when "0000010101000100", -- t[1348] = 0
      "000000" when "0000010101000101", -- t[1349] = 0
      "000000" when "0000010101000110", -- t[1350] = 0
      "000000" when "0000010101000111", -- t[1351] = 0
      "000000" when "0000010101001000", -- t[1352] = 0
      "000000" when "0000010101001001", -- t[1353] = 0
      "000000" when "0000010101001010", -- t[1354] = 0
      "000000" when "0000010101001011", -- t[1355] = 0
      "000000" when "0000010101001100", -- t[1356] = 0
      "000000" when "0000010101001101", -- t[1357] = 0
      "000000" when "0000010101001110", -- t[1358] = 0
      "000000" when "0000010101001111", -- t[1359] = 0
      "000000" when "0000010101010000", -- t[1360] = 0
      "000000" when "0000010101010001", -- t[1361] = 0
      "000000" when "0000010101010010", -- t[1362] = 0
      "000000" when "0000010101010011", -- t[1363] = 0
      "000000" when "0000010101010100", -- t[1364] = 0
      "000000" when "0000010101010101", -- t[1365] = 0
      "000000" when "0000010101010110", -- t[1366] = 0
      "000000" when "0000010101010111", -- t[1367] = 0
      "000000" when "0000010101011000", -- t[1368] = 0
      "000000" when "0000010101011001", -- t[1369] = 0
      "000000" when "0000010101011010", -- t[1370] = 0
      "000000" when "0000010101011011", -- t[1371] = 0
      "000000" when "0000010101011100", -- t[1372] = 0
      "000000" when "0000010101011101", -- t[1373] = 0
      "000000" when "0000010101011110", -- t[1374] = 0
      "000000" when "0000010101011111", -- t[1375] = 0
      "000000" when "0000010101100000", -- t[1376] = 0
      "000000" when "0000010101100001", -- t[1377] = 0
      "000000" when "0000010101100010", -- t[1378] = 0
      "000000" when "0000010101100011", -- t[1379] = 0
      "000000" when "0000010101100100", -- t[1380] = 0
      "000000" when "0000010101100101", -- t[1381] = 0
      "000000" when "0000010101100110", -- t[1382] = 0
      "000000" when "0000010101100111", -- t[1383] = 0
      "000000" when "0000010101101000", -- t[1384] = 0
      "000000" when "0000010101101001", -- t[1385] = 0
      "000000" when "0000010101101010", -- t[1386] = 0
      "000000" when "0000010101101011", -- t[1387] = 0
      "000000" when "0000010101101100", -- t[1388] = 0
      "000000" when "0000010101101101", -- t[1389] = 0
      "000000" when "0000010101101110", -- t[1390] = 0
      "000000" when "0000010101101111", -- t[1391] = 0
      "000000" when "0000010101110000", -- t[1392] = 0
      "000000" when "0000010101110001", -- t[1393] = 0
      "000000" when "0000010101110010", -- t[1394] = 0
      "000000" when "0000010101110011", -- t[1395] = 0
      "000000" when "0000010101110100", -- t[1396] = 0
      "000000" when "0000010101110101", -- t[1397] = 0
      "000000" when "0000010101110110", -- t[1398] = 0
      "000000" when "0000010101110111", -- t[1399] = 0
      "000000" when "0000010101111000", -- t[1400] = 0
      "000000" when "0000010101111001", -- t[1401] = 0
      "000000" when "0000010101111010", -- t[1402] = 0
      "000000" when "0000010101111011", -- t[1403] = 0
      "000000" when "0000010101111100", -- t[1404] = 0
      "000000" when "0000010101111101", -- t[1405] = 0
      "000000" when "0000010101111110", -- t[1406] = 0
      "000000" when "0000010101111111", -- t[1407] = 0
      "000000" when "0000010110000000", -- t[1408] = 0
      "000000" when "0000010110000001", -- t[1409] = 0
      "000000" when "0000010110000010", -- t[1410] = 0
      "000000" when "0000010110000011", -- t[1411] = 0
      "000000" when "0000010110000100", -- t[1412] = 0
      "000000" when "0000010110000101", -- t[1413] = 0
      "000000" when "0000010110000110", -- t[1414] = 0
      "000000" when "0000010110000111", -- t[1415] = 0
      "000000" when "0000010110001000", -- t[1416] = 0
      "000000" when "0000010110001001", -- t[1417] = 0
      "000000" when "0000010110001010", -- t[1418] = 0
      "000000" when "0000010110001011", -- t[1419] = 0
      "000000" when "0000010110001100", -- t[1420] = 0
      "000000" when "0000010110001101", -- t[1421] = 0
      "000000" when "0000010110001110", -- t[1422] = 0
      "000000" when "0000010110001111", -- t[1423] = 0
      "000000" when "0000010110010000", -- t[1424] = 0
      "000000" when "0000010110010001", -- t[1425] = 0
      "000000" when "0000010110010010", -- t[1426] = 0
      "000000" when "0000010110010011", -- t[1427] = 0
      "000000" when "0000010110010100", -- t[1428] = 0
      "000000" when "0000010110010101", -- t[1429] = 0
      "000000" when "0000010110010110", -- t[1430] = 0
      "000000" when "0000010110010111", -- t[1431] = 0
      "000000" when "0000010110011000", -- t[1432] = 0
      "000000" when "0000010110011001", -- t[1433] = 0
      "000000" when "0000010110011010", -- t[1434] = 0
      "000000" when "0000010110011011", -- t[1435] = 0
      "000000" when "0000010110011100", -- t[1436] = 0
      "000000" when "0000010110011101", -- t[1437] = 0
      "000000" when "0000010110011110", -- t[1438] = 0
      "000000" when "0000010110011111", -- t[1439] = 0
      "000000" when "0000010110100000", -- t[1440] = 0
      "000000" when "0000010110100001", -- t[1441] = 0
      "000000" when "0000010110100010", -- t[1442] = 0
      "000000" when "0000010110100011", -- t[1443] = 0
      "000000" when "0000010110100100", -- t[1444] = 0
      "000000" when "0000010110100101", -- t[1445] = 0
      "000000" when "0000010110100110", -- t[1446] = 0
      "000000" when "0000010110100111", -- t[1447] = 0
      "000000" when "0000010110101000", -- t[1448] = 0
      "000000" when "0000010110101001", -- t[1449] = 0
      "000000" when "0000010110101010", -- t[1450] = 0
      "000000" when "0000010110101011", -- t[1451] = 0
      "000000" when "0000010110101100", -- t[1452] = 0
      "000000" when "0000010110101101", -- t[1453] = 0
      "000000" when "0000010110101110", -- t[1454] = 0
      "000000" when "0000010110101111", -- t[1455] = 0
      "000000" when "0000010110110000", -- t[1456] = 0
      "000000" when "0000010110110001", -- t[1457] = 0
      "000000" when "0000010110110010", -- t[1458] = 0
      "000000" when "0000010110110011", -- t[1459] = 0
      "000000" when "0000010110110100", -- t[1460] = 0
      "000000" when "0000010110110101", -- t[1461] = 0
      "000000" when "0000010110110110", -- t[1462] = 0
      "000000" when "0000010110110111", -- t[1463] = 0
      "000000" when "0000010110111000", -- t[1464] = 0
      "000000" when "0000010110111001", -- t[1465] = 0
      "000000" when "0000010110111010", -- t[1466] = 0
      "000000" when "0000010110111011", -- t[1467] = 0
      "000000" when "0000010110111100", -- t[1468] = 0
      "000000" when "0000010110111101", -- t[1469] = 0
      "000000" when "0000010110111110", -- t[1470] = 0
      "000000" when "0000010110111111", -- t[1471] = 0
      "000000" when "0000010111000000", -- t[1472] = 0
      "000000" when "0000010111000001", -- t[1473] = 0
      "000000" when "0000010111000010", -- t[1474] = 0
      "000000" when "0000010111000011", -- t[1475] = 0
      "000000" when "0000010111000100", -- t[1476] = 0
      "000000" when "0000010111000101", -- t[1477] = 0
      "000000" when "0000010111000110", -- t[1478] = 0
      "000000" when "0000010111000111", -- t[1479] = 0
      "000000" when "0000010111001000", -- t[1480] = 0
      "000000" when "0000010111001001", -- t[1481] = 0
      "000000" when "0000010111001010", -- t[1482] = 0
      "000000" when "0000010111001011", -- t[1483] = 0
      "000000" when "0000010111001100", -- t[1484] = 0
      "000000" when "0000010111001101", -- t[1485] = 0
      "000000" when "0000010111001110", -- t[1486] = 0
      "000000" when "0000010111001111", -- t[1487] = 0
      "000000" when "0000010111010000", -- t[1488] = 0
      "000000" when "0000010111010001", -- t[1489] = 0
      "000000" when "0000010111010010", -- t[1490] = 0
      "000000" when "0000010111010011", -- t[1491] = 0
      "000000" when "0000010111010100", -- t[1492] = 0
      "000000" when "0000010111010101", -- t[1493] = 0
      "000000" when "0000010111010110", -- t[1494] = 0
      "000000" when "0000010111010111", -- t[1495] = 0
      "000000" when "0000010111011000", -- t[1496] = 0
      "000000" when "0000010111011001", -- t[1497] = 0
      "000000" when "0000010111011010", -- t[1498] = 0
      "000000" when "0000010111011011", -- t[1499] = 0
      "000000" when "0000010111011100", -- t[1500] = 0
      "000000" when "0000010111011101", -- t[1501] = 0
      "000000" when "0000010111011110", -- t[1502] = 0
      "000000" when "0000010111011111", -- t[1503] = 0
      "000000" when "0000010111100000", -- t[1504] = 0
      "000000" when "0000010111100001", -- t[1505] = 0
      "000000" when "0000010111100010", -- t[1506] = 0
      "000000" when "0000010111100011", -- t[1507] = 0
      "000000" when "0000010111100100", -- t[1508] = 0
      "000000" when "0000010111100101", -- t[1509] = 0
      "000000" when "0000010111100110", -- t[1510] = 0
      "000000" when "0000010111100111", -- t[1511] = 0
      "000000" when "0000010111101000", -- t[1512] = 0
      "000000" when "0000010111101001", -- t[1513] = 0
      "000000" when "0000010111101010", -- t[1514] = 0
      "000000" when "0000010111101011", -- t[1515] = 0
      "000000" when "0000010111101100", -- t[1516] = 0
      "000000" when "0000010111101101", -- t[1517] = 0
      "000000" when "0000010111101110", -- t[1518] = 0
      "000000" when "0000010111101111", -- t[1519] = 0
      "000000" when "0000010111110000", -- t[1520] = 0
      "000000" when "0000010111110001", -- t[1521] = 0
      "000000" when "0000010111110010", -- t[1522] = 0
      "000000" when "0000010111110011", -- t[1523] = 0
      "000000" when "0000010111110100", -- t[1524] = 0
      "000000" when "0000010111110101", -- t[1525] = 0
      "000000" when "0000010111110110", -- t[1526] = 0
      "000000" when "0000010111110111", -- t[1527] = 0
      "000000" when "0000010111111000", -- t[1528] = 0
      "000000" when "0000010111111001", -- t[1529] = 0
      "000000" when "0000010111111010", -- t[1530] = 0
      "000000" when "0000010111111011", -- t[1531] = 0
      "000000" when "0000010111111100", -- t[1532] = 0
      "000000" when "0000010111111101", -- t[1533] = 0
      "000000" when "0000010111111110", -- t[1534] = 0
      "000000" when "0000010111111111", -- t[1535] = 0
      "000000" when "0000011000000000", -- t[1536] = 0
      "000000" when "0000011000000001", -- t[1537] = 0
      "000000" when "0000011000000010", -- t[1538] = 0
      "000000" when "0000011000000011", -- t[1539] = 0
      "000000" when "0000011000000100", -- t[1540] = 0
      "000000" when "0000011000000101", -- t[1541] = 0
      "000000" when "0000011000000110", -- t[1542] = 0
      "000000" when "0000011000000111", -- t[1543] = 0
      "000000" when "0000011000001000", -- t[1544] = 0
      "000000" when "0000011000001001", -- t[1545] = 0
      "000000" when "0000011000001010", -- t[1546] = 0
      "000000" when "0000011000001011", -- t[1547] = 0
      "000000" when "0000011000001100", -- t[1548] = 0
      "000000" when "0000011000001101", -- t[1549] = 0
      "000000" when "0000011000001110", -- t[1550] = 0
      "000000" when "0000011000001111", -- t[1551] = 0
      "000000" when "0000011000010000", -- t[1552] = 0
      "000000" when "0000011000010001", -- t[1553] = 0
      "000000" when "0000011000010010", -- t[1554] = 0
      "000000" when "0000011000010011", -- t[1555] = 0
      "000000" when "0000011000010100", -- t[1556] = 0
      "000000" when "0000011000010101", -- t[1557] = 0
      "000000" when "0000011000010110", -- t[1558] = 0
      "000000" when "0000011000010111", -- t[1559] = 0
      "000000" when "0000011000011000", -- t[1560] = 0
      "000000" when "0000011000011001", -- t[1561] = 0
      "000000" when "0000011000011010", -- t[1562] = 0
      "000000" when "0000011000011011", -- t[1563] = 0
      "000000" when "0000011000011100", -- t[1564] = 0
      "000000" when "0000011000011101", -- t[1565] = 0
      "000000" when "0000011000011110", -- t[1566] = 0
      "000000" when "0000011000011111", -- t[1567] = 0
      "000000" when "0000011000100000", -- t[1568] = 0
      "000000" when "0000011000100001", -- t[1569] = 0
      "000000" when "0000011000100010", -- t[1570] = 0
      "000000" when "0000011000100011", -- t[1571] = 0
      "000000" when "0000011000100100", -- t[1572] = 0
      "000000" when "0000011000100101", -- t[1573] = 0
      "000000" when "0000011000100110", -- t[1574] = 0
      "000000" when "0000011000100111", -- t[1575] = 0
      "000000" when "0000011000101000", -- t[1576] = 0
      "000000" when "0000011000101001", -- t[1577] = 0
      "000000" when "0000011000101010", -- t[1578] = 0
      "000000" when "0000011000101011", -- t[1579] = 0
      "000000" when "0000011000101100", -- t[1580] = 0
      "000000" when "0000011000101101", -- t[1581] = 0
      "000000" when "0000011000101110", -- t[1582] = 0
      "000000" when "0000011000101111", -- t[1583] = 0
      "000000" when "0000011000110000", -- t[1584] = 0
      "000000" when "0000011000110001", -- t[1585] = 0
      "000000" when "0000011000110010", -- t[1586] = 0
      "000000" when "0000011000110011", -- t[1587] = 0
      "000000" when "0000011000110100", -- t[1588] = 0
      "000000" when "0000011000110101", -- t[1589] = 0
      "000000" when "0000011000110110", -- t[1590] = 0
      "000000" when "0000011000110111", -- t[1591] = 0
      "000000" when "0000011000111000", -- t[1592] = 0
      "000000" when "0000011000111001", -- t[1593] = 0
      "000000" when "0000011000111010", -- t[1594] = 0
      "000000" when "0000011000111011", -- t[1595] = 0
      "000000" when "0000011000111100", -- t[1596] = 0
      "000000" when "0000011000111101", -- t[1597] = 0
      "000000" when "0000011000111110", -- t[1598] = 0
      "000000" when "0000011000111111", -- t[1599] = 0
      "000000" when "0000011001000000", -- t[1600] = 0
      "000000" when "0000011001000001", -- t[1601] = 0
      "000000" when "0000011001000010", -- t[1602] = 0
      "000000" when "0000011001000011", -- t[1603] = 0
      "000000" when "0000011001000100", -- t[1604] = 0
      "000000" when "0000011001000101", -- t[1605] = 0
      "000000" when "0000011001000110", -- t[1606] = 0
      "000000" when "0000011001000111", -- t[1607] = 0
      "000000" when "0000011001001000", -- t[1608] = 0
      "000000" when "0000011001001001", -- t[1609] = 0
      "000000" when "0000011001001010", -- t[1610] = 0
      "000000" when "0000011001001011", -- t[1611] = 0
      "000000" when "0000011001001100", -- t[1612] = 0
      "000000" when "0000011001001101", -- t[1613] = 0
      "000000" when "0000011001001110", -- t[1614] = 0
      "000000" when "0000011001001111", -- t[1615] = 0
      "000000" when "0000011001010000", -- t[1616] = 0
      "000000" when "0000011001010001", -- t[1617] = 0
      "000000" when "0000011001010010", -- t[1618] = 0
      "000000" when "0000011001010011", -- t[1619] = 0
      "000000" when "0000011001010100", -- t[1620] = 0
      "000000" when "0000011001010101", -- t[1621] = 0
      "000000" when "0000011001010110", -- t[1622] = 0
      "000000" when "0000011001010111", -- t[1623] = 0
      "000000" when "0000011001011000", -- t[1624] = 0
      "000000" when "0000011001011001", -- t[1625] = 0
      "000000" when "0000011001011010", -- t[1626] = 0
      "000000" when "0000011001011011", -- t[1627] = 0
      "000000" when "0000011001011100", -- t[1628] = 0
      "000000" when "0000011001011101", -- t[1629] = 0
      "000000" when "0000011001011110", -- t[1630] = 0
      "000000" when "0000011001011111", -- t[1631] = 0
      "000000" when "0000011001100000", -- t[1632] = 0
      "000000" when "0000011001100001", -- t[1633] = 0
      "000000" when "0000011001100010", -- t[1634] = 0
      "000000" when "0000011001100011", -- t[1635] = 0
      "000000" when "0000011001100100", -- t[1636] = 0
      "000000" when "0000011001100101", -- t[1637] = 0
      "000000" when "0000011001100110", -- t[1638] = 0
      "000000" when "0000011001100111", -- t[1639] = 0
      "000000" when "0000011001101000", -- t[1640] = 0
      "000000" when "0000011001101001", -- t[1641] = 0
      "000000" when "0000011001101010", -- t[1642] = 0
      "000000" when "0000011001101011", -- t[1643] = 0
      "000000" when "0000011001101100", -- t[1644] = 0
      "000000" when "0000011001101101", -- t[1645] = 0
      "000000" when "0000011001101110", -- t[1646] = 0
      "000000" when "0000011001101111", -- t[1647] = 0
      "000000" when "0000011001110000", -- t[1648] = 0
      "000000" when "0000011001110001", -- t[1649] = 0
      "000000" when "0000011001110010", -- t[1650] = 0
      "000000" when "0000011001110011", -- t[1651] = 0
      "000000" when "0000011001110100", -- t[1652] = 0
      "000000" when "0000011001110101", -- t[1653] = 0
      "000000" when "0000011001110110", -- t[1654] = 0
      "000000" when "0000011001110111", -- t[1655] = 0
      "000000" when "0000011001111000", -- t[1656] = 0
      "000000" when "0000011001111001", -- t[1657] = 0
      "000000" when "0000011001111010", -- t[1658] = 0
      "000000" when "0000011001111011", -- t[1659] = 0
      "000000" when "0000011001111100", -- t[1660] = 0
      "000000" when "0000011001111101", -- t[1661] = 0
      "000000" when "0000011001111110", -- t[1662] = 0
      "000000" when "0000011001111111", -- t[1663] = 0
      "000000" when "0000011010000000", -- t[1664] = 0
      "000000" when "0000011010000001", -- t[1665] = 0
      "000000" when "0000011010000010", -- t[1666] = 0
      "000000" when "0000011010000011", -- t[1667] = 0
      "000000" when "0000011010000100", -- t[1668] = 0
      "000000" when "0000011010000101", -- t[1669] = 0
      "000000" when "0000011010000110", -- t[1670] = 0
      "000000" when "0000011010000111", -- t[1671] = 0
      "000000" when "0000011010001000", -- t[1672] = 0
      "000000" when "0000011010001001", -- t[1673] = 0
      "000000" when "0000011010001010", -- t[1674] = 0
      "000000" when "0000011010001011", -- t[1675] = 0
      "000000" when "0000011010001100", -- t[1676] = 0
      "000000" when "0000011010001101", -- t[1677] = 0
      "000000" when "0000011010001110", -- t[1678] = 0
      "000000" when "0000011010001111", -- t[1679] = 0
      "000000" when "0000011010010000", -- t[1680] = 0
      "000000" when "0000011010010001", -- t[1681] = 0
      "000000" when "0000011010010010", -- t[1682] = 0
      "000000" when "0000011010010011", -- t[1683] = 0
      "000000" when "0000011010010100", -- t[1684] = 0
      "000000" when "0000011010010101", -- t[1685] = 0
      "000000" when "0000011010010110", -- t[1686] = 0
      "000000" when "0000011010010111", -- t[1687] = 0
      "000000" when "0000011010011000", -- t[1688] = 0
      "000000" when "0000011010011001", -- t[1689] = 0
      "000000" when "0000011010011010", -- t[1690] = 0
      "000000" when "0000011010011011", -- t[1691] = 0
      "000000" when "0000011010011100", -- t[1692] = 0
      "000000" when "0000011010011101", -- t[1693] = 0
      "000000" when "0000011010011110", -- t[1694] = 0
      "000000" when "0000011010011111", -- t[1695] = 0
      "000000" when "0000011010100000", -- t[1696] = 0
      "000000" when "0000011010100001", -- t[1697] = 0
      "000000" when "0000011010100010", -- t[1698] = 0
      "000000" when "0000011010100011", -- t[1699] = 0
      "000000" when "0000011010100100", -- t[1700] = 0
      "000000" when "0000011010100101", -- t[1701] = 0
      "000000" when "0000011010100110", -- t[1702] = 0
      "000000" when "0000011010100111", -- t[1703] = 0
      "000000" when "0000011010101000", -- t[1704] = 0
      "000000" when "0000011010101001", -- t[1705] = 0
      "000000" when "0000011010101010", -- t[1706] = 0
      "000000" when "0000011010101011", -- t[1707] = 0
      "000000" when "0000011010101100", -- t[1708] = 0
      "000000" when "0000011010101101", -- t[1709] = 0
      "000000" when "0000011010101110", -- t[1710] = 0
      "000000" when "0000011010101111", -- t[1711] = 0
      "000000" when "0000011010110000", -- t[1712] = 0
      "000000" when "0000011010110001", -- t[1713] = 0
      "000000" when "0000011010110010", -- t[1714] = 0
      "000000" when "0000011010110011", -- t[1715] = 0
      "000000" when "0000011010110100", -- t[1716] = 0
      "000000" when "0000011010110101", -- t[1717] = 0
      "000000" when "0000011010110110", -- t[1718] = 0
      "000000" when "0000011010110111", -- t[1719] = 0
      "000000" when "0000011010111000", -- t[1720] = 0
      "000000" when "0000011010111001", -- t[1721] = 0
      "000000" when "0000011010111010", -- t[1722] = 0
      "000000" when "0000011010111011", -- t[1723] = 0
      "000000" when "0000011010111100", -- t[1724] = 0
      "000000" when "0000011010111101", -- t[1725] = 0
      "000000" when "0000011010111110", -- t[1726] = 0
      "000000" when "0000011010111111", -- t[1727] = 0
      "000000" when "0000011011000000", -- t[1728] = 0
      "000000" when "0000011011000001", -- t[1729] = 0
      "000000" when "0000011011000010", -- t[1730] = 0
      "000000" when "0000011011000011", -- t[1731] = 0
      "000000" when "0000011011000100", -- t[1732] = 0
      "000000" when "0000011011000101", -- t[1733] = 0
      "000000" when "0000011011000110", -- t[1734] = 0
      "000000" when "0000011011000111", -- t[1735] = 0
      "000000" when "0000011011001000", -- t[1736] = 0
      "000000" when "0000011011001001", -- t[1737] = 0
      "000000" when "0000011011001010", -- t[1738] = 0
      "000000" when "0000011011001011", -- t[1739] = 0
      "000000" when "0000011011001100", -- t[1740] = 0
      "000000" when "0000011011001101", -- t[1741] = 0
      "000000" when "0000011011001110", -- t[1742] = 0
      "000000" when "0000011011001111", -- t[1743] = 0
      "000000" when "0000011011010000", -- t[1744] = 0
      "000000" when "0000011011010001", -- t[1745] = 0
      "000000" when "0000011011010010", -- t[1746] = 0
      "000000" when "0000011011010011", -- t[1747] = 0
      "000000" when "0000011011010100", -- t[1748] = 0
      "000000" when "0000011011010101", -- t[1749] = 0
      "000000" when "0000011011010110", -- t[1750] = 0
      "000000" when "0000011011010111", -- t[1751] = 0
      "000000" when "0000011011011000", -- t[1752] = 0
      "000000" when "0000011011011001", -- t[1753] = 0
      "000000" when "0000011011011010", -- t[1754] = 0
      "000000" when "0000011011011011", -- t[1755] = 0
      "000000" when "0000011011011100", -- t[1756] = 0
      "000000" when "0000011011011101", -- t[1757] = 0
      "000000" when "0000011011011110", -- t[1758] = 0
      "000000" when "0000011011011111", -- t[1759] = 0
      "000000" when "0000011011100000", -- t[1760] = 0
      "000000" when "0000011011100001", -- t[1761] = 0
      "000000" when "0000011011100010", -- t[1762] = 0
      "000000" when "0000011011100011", -- t[1763] = 0
      "000000" when "0000011011100100", -- t[1764] = 0
      "000000" when "0000011011100101", -- t[1765] = 0
      "000000" when "0000011011100110", -- t[1766] = 0
      "000000" when "0000011011100111", -- t[1767] = 0
      "000000" when "0000011011101000", -- t[1768] = 0
      "000000" when "0000011011101001", -- t[1769] = 0
      "000000" when "0000011011101010", -- t[1770] = 0
      "000000" when "0000011011101011", -- t[1771] = 0
      "000000" when "0000011011101100", -- t[1772] = 0
      "000000" when "0000011011101101", -- t[1773] = 0
      "000000" when "0000011011101110", -- t[1774] = 0
      "000000" when "0000011011101111", -- t[1775] = 0
      "000000" when "0000011011110000", -- t[1776] = 0
      "000000" when "0000011011110001", -- t[1777] = 0
      "000000" when "0000011011110010", -- t[1778] = 0
      "000000" when "0000011011110011", -- t[1779] = 0
      "000000" when "0000011011110100", -- t[1780] = 0
      "000000" when "0000011011110101", -- t[1781] = 0
      "000000" when "0000011011110110", -- t[1782] = 0
      "000000" when "0000011011110111", -- t[1783] = 0
      "000000" when "0000011011111000", -- t[1784] = 0
      "000000" when "0000011011111001", -- t[1785] = 0
      "000000" when "0000011011111010", -- t[1786] = 0
      "000000" when "0000011011111011", -- t[1787] = 0
      "000000" when "0000011011111100", -- t[1788] = 0
      "000000" when "0000011011111101", -- t[1789] = 0
      "000000" when "0000011011111110", -- t[1790] = 0
      "000000" when "0000011011111111", -- t[1791] = 0
      "000000" when "0000011100000000", -- t[1792] = 0
      "000000" when "0000011100000001", -- t[1793] = 0
      "000000" when "0000011100000010", -- t[1794] = 0
      "000000" when "0000011100000011", -- t[1795] = 0
      "000000" when "0000011100000100", -- t[1796] = 0
      "000000" when "0000011100000101", -- t[1797] = 0
      "000000" when "0000011100000110", -- t[1798] = 0
      "000000" when "0000011100000111", -- t[1799] = 0
      "000000" when "0000011100001000", -- t[1800] = 0
      "000000" when "0000011100001001", -- t[1801] = 0
      "000000" when "0000011100001010", -- t[1802] = 0
      "000000" when "0000011100001011", -- t[1803] = 0
      "000000" when "0000011100001100", -- t[1804] = 0
      "000000" when "0000011100001101", -- t[1805] = 0
      "000000" when "0000011100001110", -- t[1806] = 0
      "000000" when "0000011100001111", -- t[1807] = 0
      "000000" when "0000011100010000", -- t[1808] = 0
      "000000" when "0000011100010001", -- t[1809] = 0
      "000000" when "0000011100010010", -- t[1810] = 0
      "000000" when "0000011100010011", -- t[1811] = 0
      "000000" when "0000011100010100", -- t[1812] = 0
      "000000" when "0000011100010101", -- t[1813] = 0
      "000000" when "0000011100010110", -- t[1814] = 0
      "000000" when "0000011100010111", -- t[1815] = 0
      "000000" when "0000011100011000", -- t[1816] = 0
      "000000" when "0000011100011001", -- t[1817] = 0
      "000000" when "0000011100011010", -- t[1818] = 0
      "000000" when "0000011100011011", -- t[1819] = 0
      "000000" when "0000011100011100", -- t[1820] = 0
      "000000" when "0000011100011101", -- t[1821] = 0
      "000000" when "0000011100011110", -- t[1822] = 0
      "000000" when "0000011100011111", -- t[1823] = 0
      "000000" when "0000011100100000", -- t[1824] = 0
      "000000" when "0000011100100001", -- t[1825] = 0
      "000000" when "0000011100100010", -- t[1826] = 0
      "000000" when "0000011100100011", -- t[1827] = 0
      "000000" when "0000011100100100", -- t[1828] = 0
      "000000" when "0000011100100101", -- t[1829] = 0
      "000000" when "0000011100100110", -- t[1830] = 0
      "000000" when "0000011100100111", -- t[1831] = 0
      "000000" when "0000011100101000", -- t[1832] = 0
      "000000" when "0000011100101001", -- t[1833] = 0
      "000000" when "0000011100101010", -- t[1834] = 0
      "000000" when "0000011100101011", -- t[1835] = 0
      "000000" when "0000011100101100", -- t[1836] = 0
      "000000" when "0000011100101101", -- t[1837] = 0
      "000000" when "0000011100101110", -- t[1838] = 0
      "000000" when "0000011100101111", -- t[1839] = 0
      "000000" when "0000011100110000", -- t[1840] = 0
      "000000" when "0000011100110001", -- t[1841] = 0
      "000000" when "0000011100110010", -- t[1842] = 0
      "000000" when "0000011100110011", -- t[1843] = 0
      "000000" when "0000011100110100", -- t[1844] = 0
      "000000" when "0000011100110101", -- t[1845] = 0
      "000000" when "0000011100110110", -- t[1846] = 0
      "000000" when "0000011100110111", -- t[1847] = 0
      "000000" when "0000011100111000", -- t[1848] = 0
      "000000" when "0000011100111001", -- t[1849] = 0
      "000000" when "0000011100111010", -- t[1850] = 0
      "000000" when "0000011100111011", -- t[1851] = 0
      "000000" when "0000011100111100", -- t[1852] = 0
      "000000" when "0000011100111101", -- t[1853] = 0
      "000000" when "0000011100111110", -- t[1854] = 0
      "000000" when "0000011100111111", -- t[1855] = 0
      "000000" when "0000011101000000", -- t[1856] = 0
      "000000" when "0000011101000001", -- t[1857] = 0
      "000000" when "0000011101000010", -- t[1858] = 0
      "000000" when "0000011101000011", -- t[1859] = 0
      "000000" when "0000011101000100", -- t[1860] = 0
      "000000" when "0000011101000101", -- t[1861] = 0
      "000000" when "0000011101000110", -- t[1862] = 0
      "000000" when "0000011101000111", -- t[1863] = 0
      "000000" when "0000011101001000", -- t[1864] = 0
      "000000" when "0000011101001001", -- t[1865] = 0
      "000000" when "0000011101001010", -- t[1866] = 0
      "000000" when "0000011101001011", -- t[1867] = 0
      "000000" when "0000011101001100", -- t[1868] = 0
      "000000" when "0000011101001101", -- t[1869] = 0
      "000000" when "0000011101001110", -- t[1870] = 0
      "000000" when "0000011101001111", -- t[1871] = 0
      "000000" when "0000011101010000", -- t[1872] = 0
      "000000" when "0000011101010001", -- t[1873] = 0
      "000000" when "0000011101010010", -- t[1874] = 0
      "000000" when "0000011101010011", -- t[1875] = 0
      "000000" when "0000011101010100", -- t[1876] = 0
      "000000" when "0000011101010101", -- t[1877] = 0
      "000000" when "0000011101010110", -- t[1878] = 0
      "000000" when "0000011101010111", -- t[1879] = 0
      "000000" when "0000011101011000", -- t[1880] = 0
      "000000" when "0000011101011001", -- t[1881] = 0
      "000000" when "0000011101011010", -- t[1882] = 0
      "000000" when "0000011101011011", -- t[1883] = 0
      "000000" when "0000011101011100", -- t[1884] = 0
      "000000" when "0000011101011101", -- t[1885] = 0
      "000000" when "0000011101011110", -- t[1886] = 0
      "000000" when "0000011101011111", -- t[1887] = 0
      "000000" when "0000011101100000", -- t[1888] = 0
      "000000" when "0000011101100001", -- t[1889] = 0
      "000000" when "0000011101100010", -- t[1890] = 0
      "000000" when "0000011101100011", -- t[1891] = 0
      "000000" when "0000011101100100", -- t[1892] = 0
      "000000" when "0000011101100101", -- t[1893] = 0
      "000000" when "0000011101100110", -- t[1894] = 0
      "000000" when "0000011101100111", -- t[1895] = 0
      "000000" when "0000011101101000", -- t[1896] = 0
      "000000" when "0000011101101001", -- t[1897] = 0
      "000000" when "0000011101101010", -- t[1898] = 0
      "000000" when "0000011101101011", -- t[1899] = 0
      "000000" when "0000011101101100", -- t[1900] = 0
      "000000" when "0000011101101101", -- t[1901] = 0
      "000000" when "0000011101101110", -- t[1902] = 0
      "000000" when "0000011101101111", -- t[1903] = 0
      "000000" when "0000011101110000", -- t[1904] = 0
      "000000" when "0000011101110001", -- t[1905] = 0
      "000000" when "0000011101110010", -- t[1906] = 0
      "000000" when "0000011101110011", -- t[1907] = 0
      "000000" when "0000011101110100", -- t[1908] = 0
      "000000" when "0000011101110101", -- t[1909] = 0
      "000000" when "0000011101110110", -- t[1910] = 0
      "000000" when "0000011101110111", -- t[1911] = 0
      "000000" when "0000011101111000", -- t[1912] = 0
      "000000" when "0000011101111001", -- t[1913] = 0
      "000000" when "0000011101111010", -- t[1914] = 0
      "000000" when "0000011101111011", -- t[1915] = 0
      "000000" when "0000011101111100", -- t[1916] = 0
      "000000" when "0000011101111101", -- t[1917] = 0
      "000000" when "0000011101111110", -- t[1918] = 0
      "000000" when "0000011101111111", -- t[1919] = 0
      "000000" when "0000011110000000", -- t[1920] = 0
      "000000" when "0000011110000001", -- t[1921] = 0
      "000000" when "0000011110000010", -- t[1922] = 0
      "000000" when "0000011110000011", -- t[1923] = 0
      "000000" when "0000011110000100", -- t[1924] = 0
      "000000" when "0000011110000101", -- t[1925] = 0
      "000000" when "0000011110000110", -- t[1926] = 0
      "000000" when "0000011110000111", -- t[1927] = 0
      "000000" when "0000011110001000", -- t[1928] = 0
      "000000" when "0000011110001001", -- t[1929] = 0
      "000000" when "0000011110001010", -- t[1930] = 0
      "000000" when "0000011110001011", -- t[1931] = 0
      "000000" when "0000011110001100", -- t[1932] = 0
      "000000" when "0000011110001101", -- t[1933] = 0
      "000000" when "0000011110001110", -- t[1934] = 0
      "000000" when "0000011110001111", -- t[1935] = 0
      "000000" when "0000011110010000", -- t[1936] = 0
      "000000" when "0000011110010001", -- t[1937] = 0
      "000000" when "0000011110010010", -- t[1938] = 0
      "000000" when "0000011110010011", -- t[1939] = 0
      "000000" when "0000011110010100", -- t[1940] = 0
      "000000" when "0000011110010101", -- t[1941] = 0
      "000000" when "0000011110010110", -- t[1942] = 0
      "000000" when "0000011110010111", -- t[1943] = 0
      "000000" when "0000011110011000", -- t[1944] = 0
      "000000" when "0000011110011001", -- t[1945] = 0
      "000000" when "0000011110011010", -- t[1946] = 0
      "000000" when "0000011110011011", -- t[1947] = 0
      "000000" when "0000011110011100", -- t[1948] = 0
      "000000" when "0000011110011101", -- t[1949] = 0
      "000000" when "0000011110011110", -- t[1950] = 0
      "000000" when "0000011110011111", -- t[1951] = 0
      "000000" when "0000011110100000", -- t[1952] = 0
      "000000" when "0000011110100001", -- t[1953] = 0
      "000000" when "0000011110100010", -- t[1954] = 0
      "000000" when "0000011110100011", -- t[1955] = 0
      "000000" when "0000011110100100", -- t[1956] = 0
      "000000" when "0000011110100101", -- t[1957] = 0
      "000000" when "0000011110100110", -- t[1958] = 0
      "000000" when "0000011110100111", -- t[1959] = 0
      "000000" when "0000011110101000", -- t[1960] = 0
      "000000" when "0000011110101001", -- t[1961] = 0
      "000000" when "0000011110101010", -- t[1962] = 0
      "000000" when "0000011110101011", -- t[1963] = 0
      "000000" when "0000011110101100", -- t[1964] = 0
      "000000" when "0000011110101101", -- t[1965] = 0
      "000000" when "0000011110101110", -- t[1966] = 0
      "000000" when "0000011110101111", -- t[1967] = 0
      "000000" when "0000011110110000", -- t[1968] = 0
      "000000" when "0000011110110001", -- t[1969] = 0
      "000000" when "0000011110110010", -- t[1970] = 0
      "000000" when "0000011110110011", -- t[1971] = 0
      "000000" when "0000011110110100", -- t[1972] = 0
      "000000" when "0000011110110101", -- t[1973] = 0
      "000000" when "0000011110110110", -- t[1974] = 0
      "000000" when "0000011110110111", -- t[1975] = 0
      "000000" when "0000011110111000", -- t[1976] = 0
      "000000" when "0000011110111001", -- t[1977] = 0
      "000000" when "0000011110111010", -- t[1978] = 0
      "000000" when "0000011110111011", -- t[1979] = 0
      "000000" when "0000011110111100", -- t[1980] = 0
      "000000" when "0000011110111101", -- t[1981] = 0
      "000000" when "0000011110111110", -- t[1982] = 0
      "000000" when "0000011110111111", -- t[1983] = 0
      "000000" when "0000011111000000", -- t[1984] = 0
      "000000" when "0000011111000001", -- t[1985] = 0
      "000000" when "0000011111000010", -- t[1986] = 0
      "000000" when "0000011111000011", -- t[1987] = 0
      "000000" when "0000011111000100", -- t[1988] = 0
      "000000" when "0000011111000101", -- t[1989] = 0
      "000000" when "0000011111000110", -- t[1990] = 0
      "000000" when "0000011111000111", -- t[1991] = 0
      "000000" when "0000011111001000", -- t[1992] = 0
      "000000" when "0000011111001001", -- t[1993] = 0
      "000000" when "0000011111001010", -- t[1994] = 0
      "000000" when "0000011111001011", -- t[1995] = 0
      "000000" when "0000011111001100", -- t[1996] = 0
      "000000" when "0000011111001101", -- t[1997] = 0
      "000000" when "0000011111001110", -- t[1998] = 0
      "000000" when "0000011111001111", -- t[1999] = 0
      "000000" when "0000011111010000", -- t[2000] = 0
      "000000" when "0000011111010001", -- t[2001] = 0
      "000000" when "0000011111010010", -- t[2002] = 0
      "000000" when "0000011111010011", -- t[2003] = 0
      "000000" when "0000011111010100", -- t[2004] = 0
      "000000" when "0000011111010101", -- t[2005] = 0
      "000000" when "0000011111010110", -- t[2006] = 0
      "000000" when "0000011111010111", -- t[2007] = 0
      "000000" when "0000011111011000", -- t[2008] = 0
      "000000" when "0000011111011001", -- t[2009] = 0
      "000000" when "0000011111011010", -- t[2010] = 0
      "000000" when "0000011111011011", -- t[2011] = 0
      "000000" when "0000011111011100", -- t[2012] = 0
      "000000" when "0000011111011101", -- t[2013] = 0
      "000000" when "0000011111011110", -- t[2014] = 0
      "000000" when "0000011111011111", -- t[2015] = 0
      "000000" when "0000011111100000", -- t[2016] = 0
      "000000" when "0000011111100001", -- t[2017] = 0
      "000000" when "0000011111100010", -- t[2018] = 0
      "000000" when "0000011111100011", -- t[2019] = 0
      "000000" when "0000011111100100", -- t[2020] = 0
      "000000" when "0000011111100101", -- t[2021] = 0
      "000000" when "0000011111100110", -- t[2022] = 0
      "000000" when "0000011111100111", -- t[2023] = 0
      "000000" when "0000011111101000", -- t[2024] = 0
      "000000" when "0000011111101001", -- t[2025] = 0
      "000000" when "0000011111101010", -- t[2026] = 0
      "000000" when "0000011111101011", -- t[2027] = 0
      "000000" when "0000011111101100", -- t[2028] = 0
      "000000" when "0000011111101101", -- t[2029] = 0
      "000000" when "0000011111101110", -- t[2030] = 0
      "000000" when "0000011111101111", -- t[2031] = 0
      "000000" when "0000011111110000", -- t[2032] = 0
      "000000" when "0000011111110001", -- t[2033] = 0
      "000000" when "0000011111110010", -- t[2034] = 0
      "000000" when "0000011111110011", -- t[2035] = 0
      "000000" when "0000011111110100", -- t[2036] = 0
      "000000" when "0000011111110101", -- t[2037] = 0
      "000000" when "0000011111110110", -- t[2038] = 0
      "000000" when "0000011111110111", -- t[2039] = 0
      "000000" when "0000011111111000", -- t[2040] = 0
      "000000" when "0000011111111001", -- t[2041] = 0
      "000000" when "0000011111111010", -- t[2042] = 0
      "000000" when "0000011111111011", -- t[2043] = 0
      "000000" when "0000011111111100", -- t[2044] = 0
      "000000" when "0000011111111101", -- t[2045] = 0
      "000000" when "0000011111111110", -- t[2046] = 0
      "000000" when "0000011111111111", -- t[2047] = 0
      "000000" when "0000100000000000", -- t[2048] = 0
      "000000" when "0000100000000001", -- t[2049] = 0
      "000000" when "0000100000000010", -- t[2050] = 0
      "000000" when "0000100000000011", -- t[2051] = 0
      "000000" when "0000100000000100", -- t[2052] = 0
      "000000" when "0000100000000101", -- t[2053] = 0
      "000000" when "0000100000000110", -- t[2054] = 0
      "000000" when "0000100000000111", -- t[2055] = 0
      "000000" when "0000100000001000", -- t[2056] = 0
      "000000" when "0000100000001001", -- t[2057] = 0
      "000000" when "0000100000001010", -- t[2058] = 0
      "000000" when "0000100000001011", -- t[2059] = 0
      "000000" when "0000100000001100", -- t[2060] = 0
      "000000" when "0000100000001101", -- t[2061] = 0
      "000000" when "0000100000001110", -- t[2062] = 0
      "000000" when "0000100000001111", -- t[2063] = 0
      "000000" when "0000100000010000", -- t[2064] = 0
      "000000" when "0000100000010001", -- t[2065] = 0
      "000000" when "0000100000010010", -- t[2066] = 0
      "000000" when "0000100000010011", -- t[2067] = 0
      "000000" when "0000100000010100", -- t[2068] = 0
      "000000" when "0000100000010101", -- t[2069] = 0
      "000000" when "0000100000010110", -- t[2070] = 0
      "000000" when "0000100000010111", -- t[2071] = 0
      "000000" when "0000100000011000", -- t[2072] = 0
      "000000" when "0000100000011001", -- t[2073] = 0
      "000000" when "0000100000011010", -- t[2074] = 0
      "000000" when "0000100000011011", -- t[2075] = 0
      "000000" when "0000100000011100", -- t[2076] = 0
      "000000" when "0000100000011101", -- t[2077] = 0
      "000000" when "0000100000011110", -- t[2078] = 0
      "000000" when "0000100000011111", -- t[2079] = 0
      "000000" when "0000100000100000", -- t[2080] = 0
      "000000" when "0000100000100001", -- t[2081] = 0
      "000000" when "0000100000100010", -- t[2082] = 0
      "000000" when "0000100000100011", -- t[2083] = 0
      "000000" when "0000100000100100", -- t[2084] = 0
      "000000" when "0000100000100101", -- t[2085] = 0
      "000000" when "0000100000100110", -- t[2086] = 0
      "000000" when "0000100000100111", -- t[2087] = 0
      "000000" when "0000100000101000", -- t[2088] = 0
      "000000" when "0000100000101001", -- t[2089] = 0
      "000000" when "0000100000101010", -- t[2090] = 0
      "000000" when "0000100000101011", -- t[2091] = 0
      "000000" when "0000100000101100", -- t[2092] = 0
      "000000" when "0000100000101101", -- t[2093] = 0
      "000000" when "0000100000101110", -- t[2094] = 0
      "000000" when "0000100000101111", -- t[2095] = 0
      "000000" when "0000100000110000", -- t[2096] = 0
      "000000" when "0000100000110001", -- t[2097] = 0
      "000000" when "0000100000110010", -- t[2098] = 0
      "000000" when "0000100000110011", -- t[2099] = 0
      "000000" when "0000100000110100", -- t[2100] = 0
      "000000" when "0000100000110101", -- t[2101] = 0
      "000000" when "0000100000110110", -- t[2102] = 0
      "000000" when "0000100000110111", -- t[2103] = 0
      "000000" when "0000100000111000", -- t[2104] = 0
      "000000" when "0000100000111001", -- t[2105] = 0
      "000000" when "0000100000111010", -- t[2106] = 0
      "000000" when "0000100000111011", -- t[2107] = 0
      "000000" when "0000100000111100", -- t[2108] = 0
      "000000" when "0000100000111101", -- t[2109] = 0
      "000000" when "0000100000111110", -- t[2110] = 0
      "000000" when "0000100000111111", -- t[2111] = 0
      "000000" when "0000100001000000", -- t[2112] = 0
      "000000" when "0000100001000001", -- t[2113] = 0
      "000000" when "0000100001000010", -- t[2114] = 0
      "000000" when "0000100001000011", -- t[2115] = 0
      "000000" when "0000100001000100", -- t[2116] = 0
      "000000" when "0000100001000101", -- t[2117] = 0
      "000000" when "0000100001000110", -- t[2118] = 0
      "000000" when "0000100001000111", -- t[2119] = 0
      "000000" when "0000100001001000", -- t[2120] = 0
      "000000" when "0000100001001001", -- t[2121] = 0
      "000000" when "0000100001001010", -- t[2122] = 0
      "000000" when "0000100001001011", -- t[2123] = 0
      "000000" when "0000100001001100", -- t[2124] = 0
      "000000" when "0000100001001101", -- t[2125] = 0
      "000000" when "0000100001001110", -- t[2126] = 0
      "000000" when "0000100001001111", -- t[2127] = 0
      "000000" when "0000100001010000", -- t[2128] = 0
      "000000" when "0000100001010001", -- t[2129] = 0
      "000000" when "0000100001010010", -- t[2130] = 0
      "000000" when "0000100001010011", -- t[2131] = 0
      "000000" when "0000100001010100", -- t[2132] = 0
      "000000" when "0000100001010101", -- t[2133] = 0
      "000000" when "0000100001010110", -- t[2134] = 0
      "000000" when "0000100001010111", -- t[2135] = 0
      "000000" when "0000100001011000", -- t[2136] = 0
      "000000" when "0000100001011001", -- t[2137] = 0
      "000000" when "0000100001011010", -- t[2138] = 0
      "000000" when "0000100001011011", -- t[2139] = 0
      "000000" when "0000100001011100", -- t[2140] = 0
      "000000" when "0000100001011101", -- t[2141] = 0
      "000000" when "0000100001011110", -- t[2142] = 0
      "000000" when "0000100001011111", -- t[2143] = 0
      "000000" when "0000100001100000", -- t[2144] = 0
      "000000" when "0000100001100001", -- t[2145] = 0
      "000000" when "0000100001100010", -- t[2146] = 0
      "000000" when "0000100001100011", -- t[2147] = 0
      "000000" when "0000100001100100", -- t[2148] = 0
      "000000" when "0000100001100101", -- t[2149] = 0
      "000000" when "0000100001100110", -- t[2150] = 0
      "000000" when "0000100001100111", -- t[2151] = 0
      "000000" when "0000100001101000", -- t[2152] = 0
      "000000" when "0000100001101001", -- t[2153] = 0
      "000000" when "0000100001101010", -- t[2154] = 0
      "000000" when "0000100001101011", -- t[2155] = 0
      "000000" when "0000100001101100", -- t[2156] = 0
      "000000" when "0000100001101101", -- t[2157] = 0
      "000000" when "0000100001101110", -- t[2158] = 0
      "000000" when "0000100001101111", -- t[2159] = 0
      "000000" when "0000100001110000", -- t[2160] = 0
      "000000" when "0000100001110001", -- t[2161] = 0
      "000000" when "0000100001110010", -- t[2162] = 0
      "000000" when "0000100001110011", -- t[2163] = 0
      "000000" when "0000100001110100", -- t[2164] = 0
      "000000" when "0000100001110101", -- t[2165] = 0
      "000000" when "0000100001110110", -- t[2166] = 0
      "000000" when "0000100001110111", -- t[2167] = 0
      "000000" when "0000100001111000", -- t[2168] = 0
      "000000" when "0000100001111001", -- t[2169] = 0
      "000000" when "0000100001111010", -- t[2170] = 0
      "000000" when "0000100001111011", -- t[2171] = 0
      "000000" when "0000100001111100", -- t[2172] = 0
      "000000" when "0000100001111101", -- t[2173] = 0
      "000000" when "0000100001111110", -- t[2174] = 0
      "000000" when "0000100001111111", -- t[2175] = 0
      "000000" when "0000100010000000", -- t[2176] = 0
      "000000" when "0000100010000001", -- t[2177] = 0
      "000000" when "0000100010000010", -- t[2178] = 0
      "000000" when "0000100010000011", -- t[2179] = 0
      "000000" when "0000100010000100", -- t[2180] = 0
      "000000" when "0000100010000101", -- t[2181] = 0
      "000000" when "0000100010000110", -- t[2182] = 0
      "000000" when "0000100010000111", -- t[2183] = 0
      "000000" when "0000100010001000", -- t[2184] = 0
      "000000" when "0000100010001001", -- t[2185] = 0
      "000000" when "0000100010001010", -- t[2186] = 0
      "000000" when "0000100010001011", -- t[2187] = 0
      "000000" when "0000100010001100", -- t[2188] = 0
      "000000" when "0000100010001101", -- t[2189] = 0
      "000000" when "0000100010001110", -- t[2190] = 0
      "000000" when "0000100010001111", -- t[2191] = 0
      "000000" when "0000100010010000", -- t[2192] = 0
      "000000" when "0000100010010001", -- t[2193] = 0
      "000000" when "0000100010010010", -- t[2194] = 0
      "000000" when "0000100010010011", -- t[2195] = 0
      "000000" when "0000100010010100", -- t[2196] = 0
      "000000" when "0000100010010101", -- t[2197] = 0
      "000000" when "0000100010010110", -- t[2198] = 0
      "000000" when "0000100010010111", -- t[2199] = 0
      "000000" when "0000100010011000", -- t[2200] = 0
      "000000" when "0000100010011001", -- t[2201] = 0
      "000000" when "0000100010011010", -- t[2202] = 0
      "000000" when "0000100010011011", -- t[2203] = 0
      "000000" when "0000100010011100", -- t[2204] = 0
      "000000" when "0000100010011101", -- t[2205] = 0
      "000000" when "0000100010011110", -- t[2206] = 0
      "000000" when "0000100010011111", -- t[2207] = 0
      "000000" when "0000100010100000", -- t[2208] = 0
      "000000" when "0000100010100001", -- t[2209] = 0
      "000000" when "0000100010100010", -- t[2210] = 0
      "000000" when "0000100010100011", -- t[2211] = 0
      "000000" when "0000100010100100", -- t[2212] = 0
      "000000" when "0000100010100101", -- t[2213] = 0
      "000000" when "0000100010100110", -- t[2214] = 0
      "000000" when "0000100010100111", -- t[2215] = 0
      "000000" when "0000100010101000", -- t[2216] = 0
      "000000" when "0000100010101001", -- t[2217] = 0
      "000000" when "0000100010101010", -- t[2218] = 0
      "000000" when "0000100010101011", -- t[2219] = 0
      "000000" when "0000100010101100", -- t[2220] = 0
      "000000" when "0000100010101101", -- t[2221] = 0
      "000000" when "0000100010101110", -- t[2222] = 0
      "000000" when "0000100010101111", -- t[2223] = 0
      "000000" when "0000100010110000", -- t[2224] = 0
      "000000" when "0000100010110001", -- t[2225] = 0
      "000000" when "0000100010110010", -- t[2226] = 0
      "000000" when "0000100010110011", -- t[2227] = 0
      "000000" when "0000100010110100", -- t[2228] = 0
      "000000" when "0000100010110101", -- t[2229] = 0
      "000000" when "0000100010110110", -- t[2230] = 0
      "000000" when "0000100010110111", -- t[2231] = 0
      "000000" when "0000100010111000", -- t[2232] = 0
      "000000" when "0000100010111001", -- t[2233] = 0
      "000000" when "0000100010111010", -- t[2234] = 0
      "000000" when "0000100010111011", -- t[2235] = 0
      "000000" when "0000100010111100", -- t[2236] = 0
      "000000" when "0000100010111101", -- t[2237] = 0
      "000000" when "0000100010111110", -- t[2238] = 0
      "000000" when "0000100010111111", -- t[2239] = 0
      "000000" when "0000100011000000", -- t[2240] = 0
      "000000" when "0000100011000001", -- t[2241] = 0
      "000000" when "0000100011000010", -- t[2242] = 0
      "000000" when "0000100011000011", -- t[2243] = 0
      "000000" when "0000100011000100", -- t[2244] = 0
      "000000" when "0000100011000101", -- t[2245] = 0
      "000000" when "0000100011000110", -- t[2246] = 0
      "000000" when "0000100011000111", -- t[2247] = 0
      "000000" when "0000100011001000", -- t[2248] = 0
      "000000" when "0000100011001001", -- t[2249] = 0
      "000000" when "0000100011001010", -- t[2250] = 0
      "000000" when "0000100011001011", -- t[2251] = 0
      "000000" when "0000100011001100", -- t[2252] = 0
      "000000" when "0000100011001101", -- t[2253] = 0
      "000000" when "0000100011001110", -- t[2254] = 0
      "000000" when "0000100011001111", -- t[2255] = 0
      "000000" when "0000100011010000", -- t[2256] = 0
      "000000" when "0000100011010001", -- t[2257] = 0
      "000000" when "0000100011010010", -- t[2258] = 0
      "000000" when "0000100011010011", -- t[2259] = 0
      "000000" when "0000100011010100", -- t[2260] = 0
      "000000" when "0000100011010101", -- t[2261] = 0
      "000000" when "0000100011010110", -- t[2262] = 0
      "000000" when "0000100011010111", -- t[2263] = 0
      "000000" when "0000100011011000", -- t[2264] = 0
      "000000" when "0000100011011001", -- t[2265] = 0
      "000000" when "0000100011011010", -- t[2266] = 0
      "000000" when "0000100011011011", -- t[2267] = 0
      "000000" when "0000100011011100", -- t[2268] = 0
      "000000" when "0000100011011101", -- t[2269] = 0
      "000000" when "0000100011011110", -- t[2270] = 0
      "000000" when "0000100011011111", -- t[2271] = 0
      "000000" when "0000100011100000", -- t[2272] = 0
      "000000" when "0000100011100001", -- t[2273] = 0
      "000000" when "0000100011100010", -- t[2274] = 0
      "000000" when "0000100011100011", -- t[2275] = 0
      "000000" when "0000100011100100", -- t[2276] = 0
      "000000" when "0000100011100101", -- t[2277] = 0
      "000000" when "0000100011100110", -- t[2278] = 0
      "000000" when "0000100011100111", -- t[2279] = 0
      "000000" when "0000100011101000", -- t[2280] = 0
      "000000" when "0000100011101001", -- t[2281] = 0
      "000000" when "0000100011101010", -- t[2282] = 0
      "000000" when "0000100011101011", -- t[2283] = 0
      "000000" when "0000100011101100", -- t[2284] = 0
      "000000" when "0000100011101101", -- t[2285] = 0
      "000000" when "0000100011101110", -- t[2286] = 0
      "000000" when "0000100011101111", -- t[2287] = 0
      "000000" when "0000100011110000", -- t[2288] = 0
      "000000" when "0000100011110001", -- t[2289] = 0
      "000000" when "0000100011110010", -- t[2290] = 0
      "000000" when "0000100011110011", -- t[2291] = 0
      "000000" when "0000100011110100", -- t[2292] = 0
      "000000" when "0000100011110101", -- t[2293] = 0
      "000000" when "0000100011110110", -- t[2294] = 0
      "000000" when "0000100011110111", -- t[2295] = 0
      "000000" when "0000100011111000", -- t[2296] = 0
      "000000" when "0000100011111001", -- t[2297] = 0
      "000000" when "0000100011111010", -- t[2298] = 0
      "000000" when "0000100011111011", -- t[2299] = 0
      "000000" when "0000100011111100", -- t[2300] = 0
      "000000" when "0000100011111101", -- t[2301] = 0
      "000000" when "0000100011111110", -- t[2302] = 0
      "000000" when "0000100011111111", -- t[2303] = 0
      "000000" when "0000100100000000", -- t[2304] = 0
      "000000" when "0000100100000001", -- t[2305] = 0
      "000000" when "0000100100000010", -- t[2306] = 0
      "000000" when "0000100100000011", -- t[2307] = 0
      "000000" when "0000100100000100", -- t[2308] = 0
      "000000" when "0000100100000101", -- t[2309] = 0
      "000000" when "0000100100000110", -- t[2310] = 0
      "000000" when "0000100100000111", -- t[2311] = 0
      "000000" when "0000100100001000", -- t[2312] = 0
      "000000" when "0000100100001001", -- t[2313] = 0
      "000000" when "0000100100001010", -- t[2314] = 0
      "000000" when "0000100100001011", -- t[2315] = 0
      "000000" when "0000100100001100", -- t[2316] = 0
      "000000" when "0000100100001101", -- t[2317] = 0
      "000000" when "0000100100001110", -- t[2318] = 0
      "000000" when "0000100100001111", -- t[2319] = 0
      "000000" when "0000100100010000", -- t[2320] = 0
      "000000" when "0000100100010001", -- t[2321] = 0
      "000000" when "0000100100010010", -- t[2322] = 0
      "000000" when "0000100100010011", -- t[2323] = 0
      "000000" when "0000100100010100", -- t[2324] = 0
      "000000" when "0000100100010101", -- t[2325] = 0
      "000000" when "0000100100010110", -- t[2326] = 0
      "000000" when "0000100100010111", -- t[2327] = 0
      "000000" when "0000100100011000", -- t[2328] = 0
      "000000" when "0000100100011001", -- t[2329] = 0
      "000000" when "0000100100011010", -- t[2330] = 0
      "000000" when "0000100100011011", -- t[2331] = 0
      "000000" when "0000100100011100", -- t[2332] = 0
      "000000" when "0000100100011101", -- t[2333] = 0
      "000000" when "0000100100011110", -- t[2334] = 0
      "000000" when "0000100100011111", -- t[2335] = 0
      "000000" when "0000100100100000", -- t[2336] = 0
      "000000" when "0000100100100001", -- t[2337] = 0
      "000000" when "0000100100100010", -- t[2338] = 0
      "000000" when "0000100100100011", -- t[2339] = 0
      "000000" when "0000100100100100", -- t[2340] = 0
      "000000" when "0000100100100101", -- t[2341] = 0
      "000000" when "0000100100100110", -- t[2342] = 0
      "000000" when "0000100100100111", -- t[2343] = 0
      "000000" when "0000100100101000", -- t[2344] = 0
      "000000" when "0000100100101001", -- t[2345] = 0
      "000000" when "0000100100101010", -- t[2346] = 0
      "000000" when "0000100100101011", -- t[2347] = 0
      "000000" when "0000100100101100", -- t[2348] = 0
      "000000" when "0000100100101101", -- t[2349] = 0
      "000000" when "0000100100101110", -- t[2350] = 0
      "000000" when "0000100100101111", -- t[2351] = 0
      "000000" when "0000100100110000", -- t[2352] = 0
      "000000" when "0000100100110001", -- t[2353] = 0
      "000000" when "0000100100110010", -- t[2354] = 0
      "000000" when "0000100100110011", -- t[2355] = 0
      "000000" when "0000100100110100", -- t[2356] = 0
      "000000" when "0000100100110101", -- t[2357] = 0
      "000000" when "0000100100110110", -- t[2358] = 0
      "000000" when "0000100100110111", -- t[2359] = 0
      "000000" when "0000100100111000", -- t[2360] = 0
      "000000" when "0000100100111001", -- t[2361] = 0
      "000000" when "0000100100111010", -- t[2362] = 0
      "000000" when "0000100100111011", -- t[2363] = 0
      "000000" when "0000100100111100", -- t[2364] = 0
      "000000" when "0000100100111101", -- t[2365] = 0
      "000000" when "0000100100111110", -- t[2366] = 0
      "000000" when "0000100100111111", -- t[2367] = 0
      "000000" when "0000100101000000", -- t[2368] = 0
      "000000" when "0000100101000001", -- t[2369] = 0
      "000000" when "0000100101000010", -- t[2370] = 0
      "000000" when "0000100101000011", -- t[2371] = 0
      "000000" when "0000100101000100", -- t[2372] = 0
      "000000" when "0000100101000101", -- t[2373] = 0
      "000000" when "0000100101000110", -- t[2374] = 0
      "000000" when "0000100101000111", -- t[2375] = 0
      "000000" when "0000100101001000", -- t[2376] = 0
      "000000" when "0000100101001001", -- t[2377] = 0
      "000000" when "0000100101001010", -- t[2378] = 0
      "000000" when "0000100101001011", -- t[2379] = 0
      "000000" when "0000100101001100", -- t[2380] = 0
      "000000" when "0000100101001101", -- t[2381] = 0
      "000000" when "0000100101001110", -- t[2382] = 0
      "000000" when "0000100101001111", -- t[2383] = 0
      "000000" when "0000100101010000", -- t[2384] = 0
      "000000" when "0000100101010001", -- t[2385] = 0
      "000000" when "0000100101010010", -- t[2386] = 0
      "000000" when "0000100101010011", -- t[2387] = 0
      "000000" when "0000100101010100", -- t[2388] = 0
      "000000" when "0000100101010101", -- t[2389] = 0
      "000000" when "0000100101010110", -- t[2390] = 0
      "000000" when "0000100101010111", -- t[2391] = 0
      "000000" when "0000100101011000", -- t[2392] = 0
      "000000" when "0000100101011001", -- t[2393] = 0
      "000000" when "0000100101011010", -- t[2394] = 0
      "000000" when "0000100101011011", -- t[2395] = 0
      "000000" when "0000100101011100", -- t[2396] = 0
      "000000" when "0000100101011101", -- t[2397] = 0
      "000000" when "0000100101011110", -- t[2398] = 0
      "000000" when "0000100101011111", -- t[2399] = 0
      "000000" when "0000100101100000", -- t[2400] = 0
      "000000" when "0000100101100001", -- t[2401] = 0
      "000000" when "0000100101100010", -- t[2402] = 0
      "000000" when "0000100101100011", -- t[2403] = 0
      "000000" when "0000100101100100", -- t[2404] = 0
      "000000" when "0000100101100101", -- t[2405] = 0
      "000000" when "0000100101100110", -- t[2406] = 0
      "000000" when "0000100101100111", -- t[2407] = 0
      "000000" when "0000100101101000", -- t[2408] = 0
      "000000" when "0000100101101001", -- t[2409] = 0
      "000000" when "0000100101101010", -- t[2410] = 0
      "000000" when "0000100101101011", -- t[2411] = 0
      "000000" when "0000100101101100", -- t[2412] = 0
      "000000" when "0000100101101101", -- t[2413] = 0
      "000000" when "0000100101101110", -- t[2414] = 0
      "000000" when "0000100101101111", -- t[2415] = 0
      "000000" when "0000100101110000", -- t[2416] = 0
      "000000" when "0000100101110001", -- t[2417] = 0
      "000000" when "0000100101110010", -- t[2418] = 0
      "000000" when "0000100101110011", -- t[2419] = 0
      "000000" when "0000100101110100", -- t[2420] = 0
      "000000" when "0000100101110101", -- t[2421] = 0
      "000000" when "0000100101110110", -- t[2422] = 0
      "000000" when "0000100101110111", -- t[2423] = 0
      "000000" when "0000100101111000", -- t[2424] = 0
      "000000" when "0000100101111001", -- t[2425] = 0
      "000000" when "0000100101111010", -- t[2426] = 0
      "000000" when "0000100101111011", -- t[2427] = 0
      "000000" when "0000100101111100", -- t[2428] = 0
      "000000" when "0000100101111101", -- t[2429] = 0
      "000000" when "0000100101111110", -- t[2430] = 0
      "000000" when "0000100101111111", -- t[2431] = 0
      "000000" when "0000100110000000", -- t[2432] = 0
      "000000" when "0000100110000001", -- t[2433] = 0
      "000000" when "0000100110000010", -- t[2434] = 0
      "000000" when "0000100110000011", -- t[2435] = 0
      "000000" when "0000100110000100", -- t[2436] = 0
      "000000" when "0000100110000101", -- t[2437] = 0
      "000000" when "0000100110000110", -- t[2438] = 0
      "000000" when "0000100110000111", -- t[2439] = 0
      "000000" when "0000100110001000", -- t[2440] = 0
      "000000" when "0000100110001001", -- t[2441] = 0
      "000000" when "0000100110001010", -- t[2442] = 0
      "000000" when "0000100110001011", -- t[2443] = 0
      "000000" when "0000100110001100", -- t[2444] = 0
      "000000" when "0000100110001101", -- t[2445] = 0
      "000000" when "0000100110001110", -- t[2446] = 0
      "000000" when "0000100110001111", -- t[2447] = 0
      "000000" when "0000100110010000", -- t[2448] = 0
      "000000" when "0000100110010001", -- t[2449] = 0
      "000000" when "0000100110010010", -- t[2450] = 0
      "000000" when "0000100110010011", -- t[2451] = 0
      "000000" when "0000100110010100", -- t[2452] = 0
      "000000" when "0000100110010101", -- t[2453] = 0
      "000000" when "0000100110010110", -- t[2454] = 0
      "000000" when "0000100110010111", -- t[2455] = 0
      "000000" when "0000100110011000", -- t[2456] = 0
      "000000" when "0000100110011001", -- t[2457] = 0
      "000000" when "0000100110011010", -- t[2458] = 0
      "000000" when "0000100110011011", -- t[2459] = 0
      "000000" when "0000100110011100", -- t[2460] = 0
      "000000" when "0000100110011101", -- t[2461] = 0
      "000000" when "0000100110011110", -- t[2462] = 0
      "000000" when "0000100110011111", -- t[2463] = 0
      "000000" when "0000100110100000", -- t[2464] = 0
      "000000" when "0000100110100001", -- t[2465] = 0
      "000000" when "0000100110100010", -- t[2466] = 0
      "000000" when "0000100110100011", -- t[2467] = 0
      "000000" when "0000100110100100", -- t[2468] = 0
      "000000" when "0000100110100101", -- t[2469] = 0
      "000000" when "0000100110100110", -- t[2470] = 0
      "000000" when "0000100110100111", -- t[2471] = 0
      "000000" when "0000100110101000", -- t[2472] = 0
      "000000" when "0000100110101001", -- t[2473] = 0
      "000000" when "0000100110101010", -- t[2474] = 0
      "000000" when "0000100110101011", -- t[2475] = 0
      "000000" when "0000100110101100", -- t[2476] = 0
      "000000" when "0000100110101101", -- t[2477] = 0
      "000000" when "0000100110101110", -- t[2478] = 0
      "000000" when "0000100110101111", -- t[2479] = 0
      "000000" when "0000100110110000", -- t[2480] = 0
      "000000" when "0000100110110001", -- t[2481] = 0
      "000000" when "0000100110110010", -- t[2482] = 0
      "000000" when "0000100110110011", -- t[2483] = 0
      "000000" when "0000100110110100", -- t[2484] = 0
      "000000" when "0000100110110101", -- t[2485] = 0
      "000000" when "0000100110110110", -- t[2486] = 0
      "000000" when "0000100110110111", -- t[2487] = 0
      "000000" when "0000100110111000", -- t[2488] = 0
      "000000" when "0000100110111001", -- t[2489] = 0
      "000000" when "0000100110111010", -- t[2490] = 0
      "000000" when "0000100110111011", -- t[2491] = 0
      "000000" when "0000100110111100", -- t[2492] = 0
      "000000" when "0000100110111101", -- t[2493] = 0
      "000000" when "0000100110111110", -- t[2494] = 0
      "000000" when "0000100110111111", -- t[2495] = 0
      "000000" when "0000100111000000", -- t[2496] = 0
      "000000" when "0000100111000001", -- t[2497] = 0
      "000000" when "0000100111000010", -- t[2498] = 0
      "000000" when "0000100111000011", -- t[2499] = 0
      "000000" when "0000100111000100", -- t[2500] = 0
      "000000" when "0000100111000101", -- t[2501] = 0
      "000000" when "0000100111000110", -- t[2502] = 0
      "000000" when "0000100111000111", -- t[2503] = 0
      "000000" when "0000100111001000", -- t[2504] = 0
      "000000" when "0000100111001001", -- t[2505] = 0
      "000000" when "0000100111001010", -- t[2506] = 0
      "000000" when "0000100111001011", -- t[2507] = 0
      "000000" when "0000100111001100", -- t[2508] = 0
      "000000" when "0000100111001101", -- t[2509] = 0
      "000000" when "0000100111001110", -- t[2510] = 0
      "000000" when "0000100111001111", -- t[2511] = 0
      "000000" when "0000100111010000", -- t[2512] = 0
      "000000" when "0000100111010001", -- t[2513] = 0
      "000000" when "0000100111010010", -- t[2514] = 0
      "000000" when "0000100111010011", -- t[2515] = 0
      "000000" when "0000100111010100", -- t[2516] = 0
      "000000" when "0000100111010101", -- t[2517] = 0
      "000000" when "0000100111010110", -- t[2518] = 0
      "000000" when "0000100111010111", -- t[2519] = 0
      "000000" when "0000100111011000", -- t[2520] = 0
      "000000" when "0000100111011001", -- t[2521] = 0
      "000000" when "0000100111011010", -- t[2522] = 0
      "000000" when "0000100111011011", -- t[2523] = 0
      "000000" when "0000100111011100", -- t[2524] = 0
      "000000" when "0000100111011101", -- t[2525] = 0
      "000000" when "0000100111011110", -- t[2526] = 0
      "000000" when "0000100111011111", -- t[2527] = 0
      "000000" when "0000100111100000", -- t[2528] = 0
      "000000" when "0000100111100001", -- t[2529] = 0
      "000000" when "0000100111100010", -- t[2530] = 0
      "000000" when "0000100111100011", -- t[2531] = 0
      "000000" when "0000100111100100", -- t[2532] = 0
      "000000" when "0000100111100101", -- t[2533] = 0
      "000000" when "0000100111100110", -- t[2534] = 0
      "000000" when "0000100111100111", -- t[2535] = 0
      "000000" when "0000100111101000", -- t[2536] = 0
      "000000" when "0000100111101001", -- t[2537] = 0
      "000000" when "0000100111101010", -- t[2538] = 0
      "000000" when "0000100111101011", -- t[2539] = 0
      "000000" when "0000100111101100", -- t[2540] = 0
      "000000" when "0000100111101101", -- t[2541] = 0
      "000000" when "0000100111101110", -- t[2542] = 0
      "000000" when "0000100111101111", -- t[2543] = 0
      "000000" when "0000100111110000", -- t[2544] = 0
      "000000" when "0000100111110001", -- t[2545] = 0
      "000000" when "0000100111110010", -- t[2546] = 0
      "000000" when "0000100111110011", -- t[2547] = 0
      "000000" when "0000100111110100", -- t[2548] = 0
      "000000" when "0000100111110101", -- t[2549] = 0
      "000000" when "0000100111110110", -- t[2550] = 0
      "000000" when "0000100111110111", -- t[2551] = 0
      "000000" when "0000100111111000", -- t[2552] = 0
      "000000" when "0000100111111001", -- t[2553] = 0
      "000000" when "0000100111111010", -- t[2554] = 0
      "000000" when "0000100111111011", -- t[2555] = 0
      "000000" when "0000100111111100", -- t[2556] = 0
      "000000" when "0000100111111101", -- t[2557] = 0
      "000000" when "0000100111111110", -- t[2558] = 0
      "000000" when "0000100111111111", -- t[2559] = 0
      "000000" when "0000101000000000", -- t[2560] = 0
      "000000" when "0000101000000001", -- t[2561] = 0
      "000000" when "0000101000000010", -- t[2562] = 0
      "000000" when "0000101000000011", -- t[2563] = 0
      "000000" when "0000101000000100", -- t[2564] = 0
      "000000" when "0000101000000101", -- t[2565] = 0
      "000000" when "0000101000000110", -- t[2566] = 0
      "000000" when "0000101000000111", -- t[2567] = 0
      "000000" when "0000101000001000", -- t[2568] = 0
      "000000" when "0000101000001001", -- t[2569] = 0
      "000000" when "0000101000001010", -- t[2570] = 0
      "000000" when "0000101000001011", -- t[2571] = 0
      "000000" when "0000101000001100", -- t[2572] = 0
      "000000" when "0000101000001101", -- t[2573] = 0
      "000000" when "0000101000001110", -- t[2574] = 0
      "000000" when "0000101000001111", -- t[2575] = 0
      "000000" when "0000101000010000", -- t[2576] = 0
      "000000" when "0000101000010001", -- t[2577] = 0
      "000000" when "0000101000010010", -- t[2578] = 0
      "000000" when "0000101000010011", -- t[2579] = 0
      "000000" when "0000101000010100", -- t[2580] = 0
      "000000" when "0000101000010101", -- t[2581] = 0
      "000000" when "0000101000010110", -- t[2582] = 0
      "000000" when "0000101000010111", -- t[2583] = 0
      "000000" when "0000101000011000", -- t[2584] = 0
      "000000" when "0000101000011001", -- t[2585] = 0
      "000000" when "0000101000011010", -- t[2586] = 0
      "000000" when "0000101000011011", -- t[2587] = 0
      "000000" when "0000101000011100", -- t[2588] = 0
      "000000" when "0000101000011101", -- t[2589] = 0
      "000000" when "0000101000011110", -- t[2590] = 0
      "000000" when "0000101000011111", -- t[2591] = 0
      "000000" when "0000101000100000", -- t[2592] = 0
      "000000" when "0000101000100001", -- t[2593] = 0
      "000000" when "0000101000100010", -- t[2594] = 0
      "000000" when "0000101000100011", -- t[2595] = 0
      "000000" when "0000101000100100", -- t[2596] = 0
      "000000" when "0000101000100101", -- t[2597] = 0
      "000000" when "0000101000100110", -- t[2598] = 0
      "000000" when "0000101000100111", -- t[2599] = 0
      "000000" when "0000101000101000", -- t[2600] = 0
      "000000" when "0000101000101001", -- t[2601] = 0
      "000000" when "0000101000101010", -- t[2602] = 0
      "000000" when "0000101000101011", -- t[2603] = 0
      "000000" when "0000101000101100", -- t[2604] = 0
      "000000" when "0000101000101101", -- t[2605] = 0
      "000000" when "0000101000101110", -- t[2606] = 0
      "000000" when "0000101000101111", -- t[2607] = 0
      "000000" when "0000101000110000", -- t[2608] = 0
      "000000" when "0000101000110001", -- t[2609] = 0
      "000000" when "0000101000110010", -- t[2610] = 0
      "000000" when "0000101000110011", -- t[2611] = 0
      "000000" when "0000101000110100", -- t[2612] = 0
      "000000" when "0000101000110101", -- t[2613] = 0
      "000000" when "0000101000110110", -- t[2614] = 0
      "000000" when "0000101000110111", -- t[2615] = 0
      "000000" when "0000101000111000", -- t[2616] = 0
      "000000" when "0000101000111001", -- t[2617] = 0
      "000000" when "0000101000111010", -- t[2618] = 0
      "000000" when "0000101000111011", -- t[2619] = 0
      "000000" when "0000101000111100", -- t[2620] = 0
      "000000" when "0000101000111101", -- t[2621] = 0
      "000000" when "0000101000111110", -- t[2622] = 0
      "000000" when "0000101000111111", -- t[2623] = 0
      "000000" when "0000101001000000", -- t[2624] = 0
      "000000" when "0000101001000001", -- t[2625] = 0
      "000000" when "0000101001000010", -- t[2626] = 0
      "000000" when "0000101001000011", -- t[2627] = 0
      "000000" when "0000101001000100", -- t[2628] = 0
      "000000" when "0000101001000101", -- t[2629] = 0
      "000000" when "0000101001000110", -- t[2630] = 0
      "000000" when "0000101001000111", -- t[2631] = 0
      "000000" when "0000101001001000", -- t[2632] = 0
      "000000" when "0000101001001001", -- t[2633] = 0
      "000000" when "0000101001001010", -- t[2634] = 0
      "000000" when "0000101001001011", -- t[2635] = 0
      "000000" when "0000101001001100", -- t[2636] = 0
      "000000" when "0000101001001101", -- t[2637] = 0
      "000000" when "0000101001001110", -- t[2638] = 0
      "000000" when "0000101001001111", -- t[2639] = 0
      "000000" when "0000101001010000", -- t[2640] = 0
      "000000" when "0000101001010001", -- t[2641] = 0
      "000000" when "0000101001010010", -- t[2642] = 0
      "000000" when "0000101001010011", -- t[2643] = 0
      "000000" when "0000101001010100", -- t[2644] = 0
      "000000" when "0000101001010101", -- t[2645] = 0
      "000000" when "0000101001010110", -- t[2646] = 0
      "000000" when "0000101001010111", -- t[2647] = 0
      "000000" when "0000101001011000", -- t[2648] = 0
      "000000" when "0000101001011001", -- t[2649] = 0
      "000000" when "0000101001011010", -- t[2650] = 0
      "000000" when "0000101001011011", -- t[2651] = 0
      "000000" when "0000101001011100", -- t[2652] = 0
      "000000" when "0000101001011101", -- t[2653] = 0
      "000000" when "0000101001011110", -- t[2654] = 0
      "000000" when "0000101001011111", -- t[2655] = 0
      "000000" when "0000101001100000", -- t[2656] = 0
      "000000" when "0000101001100001", -- t[2657] = 0
      "000000" when "0000101001100010", -- t[2658] = 0
      "000000" when "0000101001100011", -- t[2659] = 0
      "000000" when "0000101001100100", -- t[2660] = 0
      "000000" when "0000101001100101", -- t[2661] = 0
      "000000" when "0000101001100110", -- t[2662] = 0
      "000000" when "0000101001100111", -- t[2663] = 0
      "000000" when "0000101001101000", -- t[2664] = 0
      "000000" when "0000101001101001", -- t[2665] = 0
      "000000" when "0000101001101010", -- t[2666] = 0
      "000000" when "0000101001101011", -- t[2667] = 0
      "000000" when "0000101001101100", -- t[2668] = 0
      "000000" when "0000101001101101", -- t[2669] = 0
      "000000" when "0000101001101110", -- t[2670] = 0
      "000000" when "0000101001101111", -- t[2671] = 0
      "000000" when "0000101001110000", -- t[2672] = 0
      "000000" when "0000101001110001", -- t[2673] = 0
      "000000" when "0000101001110010", -- t[2674] = 0
      "000000" when "0000101001110011", -- t[2675] = 0
      "000000" when "0000101001110100", -- t[2676] = 0
      "000000" when "0000101001110101", -- t[2677] = 0
      "000000" when "0000101001110110", -- t[2678] = 0
      "000000" when "0000101001110111", -- t[2679] = 0
      "000000" when "0000101001111000", -- t[2680] = 0
      "000000" when "0000101001111001", -- t[2681] = 0
      "000000" when "0000101001111010", -- t[2682] = 0
      "000000" when "0000101001111011", -- t[2683] = 0
      "000000" when "0000101001111100", -- t[2684] = 0
      "000000" when "0000101001111101", -- t[2685] = 0
      "000000" when "0000101001111110", -- t[2686] = 0
      "000000" when "0000101001111111", -- t[2687] = 0
      "000000" when "0000101010000000", -- t[2688] = 0
      "000000" when "0000101010000001", -- t[2689] = 0
      "000000" when "0000101010000010", -- t[2690] = 0
      "000000" when "0000101010000011", -- t[2691] = 0
      "000000" when "0000101010000100", -- t[2692] = 0
      "000000" when "0000101010000101", -- t[2693] = 0
      "000000" when "0000101010000110", -- t[2694] = 0
      "000000" when "0000101010000111", -- t[2695] = 0
      "000000" when "0000101010001000", -- t[2696] = 0
      "000000" when "0000101010001001", -- t[2697] = 0
      "000000" when "0000101010001010", -- t[2698] = 0
      "000000" when "0000101010001011", -- t[2699] = 0
      "000000" when "0000101010001100", -- t[2700] = 0
      "000000" when "0000101010001101", -- t[2701] = 0
      "000000" when "0000101010001110", -- t[2702] = 0
      "000000" when "0000101010001111", -- t[2703] = 0
      "000000" when "0000101010010000", -- t[2704] = 0
      "000000" when "0000101010010001", -- t[2705] = 0
      "000000" when "0000101010010010", -- t[2706] = 0
      "000000" when "0000101010010011", -- t[2707] = 0
      "000000" when "0000101010010100", -- t[2708] = 0
      "000000" when "0000101010010101", -- t[2709] = 0
      "000000" when "0000101010010110", -- t[2710] = 0
      "000000" when "0000101010010111", -- t[2711] = 0
      "000000" when "0000101010011000", -- t[2712] = 0
      "000000" when "0000101010011001", -- t[2713] = 0
      "000000" when "0000101010011010", -- t[2714] = 0
      "000000" when "0000101010011011", -- t[2715] = 0
      "000000" when "0000101010011100", -- t[2716] = 0
      "000000" when "0000101010011101", -- t[2717] = 0
      "000000" when "0000101010011110", -- t[2718] = 0
      "000000" when "0000101010011111", -- t[2719] = 0
      "000000" when "0000101010100000", -- t[2720] = 0
      "000000" when "0000101010100001", -- t[2721] = 0
      "000000" when "0000101010100010", -- t[2722] = 0
      "000000" when "0000101010100011", -- t[2723] = 0
      "000000" when "0000101010100100", -- t[2724] = 0
      "000000" when "0000101010100101", -- t[2725] = 0
      "000000" when "0000101010100110", -- t[2726] = 0
      "000000" when "0000101010100111", -- t[2727] = 0
      "000000" when "0000101010101000", -- t[2728] = 0
      "000000" when "0000101010101001", -- t[2729] = 0
      "000000" when "0000101010101010", -- t[2730] = 0
      "000000" when "0000101010101011", -- t[2731] = 0
      "000000" when "0000101010101100", -- t[2732] = 0
      "000000" when "0000101010101101", -- t[2733] = 0
      "000000" when "0000101010101110", -- t[2734] = 0
      "000000" when "0000101010101111", -- t[2735] = 0
      "000000" when "0000101010110000", -- t[2736] = 0
      "000000" when "0000101010110001", -- t[2737] = 0
      "000000" when "0000101010110010", -- t[2738] = 0
      "000000" when "0000101010110011", -- t[2739] = 0
      "000000" when "0000101010110100", -- t[2740] = 0
      "000000" when "0000101010110101", -- t[2741] = 0
      "000000" when "0000101010110110", -- t[2742] = 0
      "000000" when "0000101010110111", -- t[2743] = 0
      "000000" when "0000101010111000", -- t[2744] = 0
      "000000" when "0000101010111001", -- t[2745] = 0
      "000000" when "0000101010111010", -- t[2746] = 0
      "000000" when "0000101010111011", -- t[2747] = 0
      "000000" when "0000101010111100", -- t[2748] = 0
      "000000" when "0000101010111101", -- t[2749] = 0
      "000000" when "0000101010111110", -- t[2750] = 0
      "000000" when "0000101010111111", -- t[2751] = 0
      "000000" when "0000101011000000", -- t[2752] = 0
      "000000" when "0000101011000001", -- t[2753] = 0
      "000000" when "0000101011000010", -- t[2754] = 0
      "000000" when "0000101011000011", -- t[2755] = 0
      "000000" when "0000101011000100", -- t[2756] = 0
      "000000" when "0000101011000101", -- t[2757] = 0
      "000000" when "0000101011000110", -- t[2758] = 0
      "000000" when "0000101011000111", -- t[2759] = 0
      "000000" when "0000101011001000", -- t[2760] = 0
      "000000" when "0000101011001001", -- t[2761] = 0
      "000000" when "0000101011001010", -- t[2762] = 0
      "000000" when "0000101011001011", -- t[2763] = 0
      "000000" when "0000101011001100", -- t[2764] = 0
      "000000" when "0000101011001101", -- t[2765] = 0
      "000000" when "0000101011001110", -- t[2766] = 0
      "000000" when "0000101011001111", -- t[2767] = 0
      "000000" when "0000101011010000", -- t[2768] = 0
      "000000" when "0000101011010001", -- t[2769] = 0
      "000000" when "0000101011010010", -- t[2770] = 0
      "000000" when "0000101011010011", -- t[2771] = 0
      "000000" when "0000101011010100", -- t[2772] = 0
      "000000" when "0000101011010101", -- t[2773] = 0
      "000000" when "0000101011010110", -- t[2774] = 0
      "000000" when "0000101011010111", -- t[2775] = 0
      "000000" when "0000101011011000", -- t[2776] = 0
      "000000" when "0000101011011001", -- t[2777] = 0
      "000000" when "0000101011011010", -- t[2778] = 0
      "000000" when "0000101011011011", -- t[2779] = 0
      "000000" when "0000101011011100", -- t[2780] = 0
      "000000" when "0000101011011101", -- t[2781] = 0
      "000000" when "0000101011011110", -- t[2782] = 0
      "000000" when "0000101011011111", -- t[2783] = 0
      "000000" when "0000101011100000", -- t[2784] = 0
      "000000" when "0000101011100001", -- t[2785] = 0
      "000000" when "0000101011100010", -- t[2786] = 0
      "000000" when "0000101011100011", -- t[2787] = 0
      "000000" when "0000101011100100", -- t[2788] = 0
      "000000" when "0000101011100101", -- t[2789] = 0
      "000000" when "0000101011100110", -- t[2790] = 0
      "000000" when "0000101011100111", -- t[2791] = 0
      "000000" when "0000101011101000", -- t[2792] = 0
      "000000" when "0000101011101001", -- t[2793] = 0
      "000000" when "0000101011101010", -- t[2794] = 0
      "000000" when "0000101011101011", -- t[2795] = 0
      "000000" when "0000101011101100", -- t[2796] = 0
      "000000" when "0000101011101101", -- t[2797] = 0
      "000000" when "0000101011101110", -- t[2798] = 0
      "000000" when "0000101011101111", -- t[2799] = 0
      "000000" when "0000101011110000", -- t[2800] = 0
      "000000" when "0000101011110001", -- t[2801] = 0
      "000000" when "0000101011110010", -- t[2802] = 0
      "000000" when "0000101011110011", -- t[2803] = 0
      "000000" when "0000101011110100", -- t[2804] = 0
      "000000" when "0000101011110101", -- t[2805] = 0
      "000000" when "0000101011110110", -- t[2806] = 0
      "000000" when "0000101011110111", -- t[2807] = 0
      "000000" when "0000101011111000", -- t[2808] = 0
      "000000" when "0000101011111001", -- t[2809] = 0
      "000000" when "0000101011111010", -- t[2810] = 0
      "000000" when "0000101011111011", -- t[2811] = 0
      "000000" when "0000101011111100", -- t[2812] = 0
      "000000" when "0000101011111101", -- t[2813] = 0
      "000000" when "0000101011111110", -- t[2814] = 0
      "000000" when "0000101011111111", -- t[2815] = 0
      "000000" when "0000101100000000", -- t[2816] = 0
      "000000" when "0000101100000001", -- t[2817] = 0
      "000000" when "0000101100000010", -- t[2818] = 0
      "000000" when "0000101100000011", -- t[2819] = 0
      "000000" when "0000101100000100", -- t[2820] = 0
      "000000" when "0000101100000101", -- t[2821] = 0
      "000000" when "0000101100000110", -- t[2822] = 0
      "000000" when "0000101100000111", -- t[2823] = 0
      "000000" when "0000101100001000", -- t[2824] = 0
      "000000" when "0000101100001001", -- t[2825] = 0
      "000000" when "0000101100001010", -- t[2826] = 0
      "000000" when "0000101100001011", -- t[2827] = 0
      "000000" when "0000101100001100", -- t[2828] = 0
      "000000" when "0000101100001101", -- t[2829] = 0
      "000000" when "0000101100001110", -- t[2830] = 0
      "000000" when "0000101100001111", -- t[2831] = 0
      "000000" when "0000101100010000", -- t[2832] = 0
      "000000" when "0000101100010001", -- t[2833] = 0
      "000000" when "0000101100010010", -- t[2834] = 0
      "000000" when "0000101100010011", -- t[2835] = 0
      "000000" when "0000101100010100", -- t[2836] = 0
      "000000" when "0000101100010101", -- t[2837] = 0
      "000000" when "0000101100010110", -- t[2838] = 0
      "000000" when "0000101100010111", -- t[2839] = 0
      "000000" when "0000101100011000", -- t[2840] = 0
      "000000" when "0000101100011001", -- t[2841] = 0
      "000000" when "0000101100011010", -- t[2842] = 0
      "000000" when "0000101100011011", -- t[2843] = 0
      "000000" when "0000101100011100", -- t[2844] = 0
      "000000" when "0000101100011101", -- t[2845] = 0
      "000000" when "0000101100011110", -- t[2846] = 0
      "000000" when "0000101100011111", -- t[2847] = 0
      "000000" when "0000101100100000", -- t[2848] = 0
      "000000" when "0000101100100001", -- t[2849] = 0
      "000000" when "0000101100100010", -- t[2850] = 0
      "000000" when "0000101100100011", -- t[2851] = 0
      "000000" when "0000101100100100", -- t[2852] = 0
      "000000" when "0000101100100101", -- t[2853] = 0
      "000000" when "0000101100100110", -- t[2854] = 0
      "000000" when "0000101100100111", -- t[2855] = 0
      "000000" when "0000101100101000", -- t[2856] = 0
      "000000" when "0000101100101001", -- t[2857] = 0
      "000000" when "0000101100101010", -- t[2858] = 0
      "000000" when "0000101100101011", -- t[2859] = 0
      "000000" when "0000101100101100", -- t[2860] = 0
      "000000" when "0000101100101101", -- t[2861] = 0
      "000000" when "0000101100101110", -- t[2862] = 0
      "000000" when "0000101100101111", -- t[2863] = 0
      "000000" when "0000101100110000", -- t[2864] = 0
      "000000" when "0000101100110001", -- t[2865] = 0
      "000000" when "0000101100110010", -- t[2866] = 0
      "000000" when "0000101100110011", -- t[2867] = 0
      "000000" when "0000101100110100", -- t[2868] = 0
      "000000" when "0000101100110101", -- t[2869] = 0
      "000000" when "0000101100110110", -- t[2870] = 0
      "000000" when "0000101100110111", -- t[2871] = 0
      "000000" when "0000101100111000", -- t[2872] = 0
      "000000" when "0000101100111001", -- t[2873] = 0
      "000000" when "0000101100111010", -- t[2874] = 0
      "000000" when "0000101100111011", -- t[2875] = 0
      "000000" when "0000101100111100", -- t[2876] = 0
      "000000" when "0000101100111101", -- t[2877] = 0
      "000000" when "0000101100111110", -- t[2878] = 0
      "000000" when "0000101100111111", -- t[2879] = 0
      "000000" when "0000101101000000", -- t[2880] = 0
      "000000" when "0000101101000001", -- t[2881] = 0
      "000000" when "0000101101000010", -- t[2882] = 0
      "000000" when "0000101101000011", -- t[2883] = 0
      "000000" when "0000101101000100", -- t[2884] = 0
      "000000" when "0000101101000101", -- t[2885] = 0
      "000000" when "0000101101000110", -- t[2886] = 0
      "000000" when "0000101101000111", -- t[2887] = 0
      "000000" when "0000101101001000", -- t[2888] = 0
      "000000" when "0000101101001001", -- t[2889] = 0
      "000000" when "0000101101001010", -- t[2890] = 0
      "000000" when "0000101101001011", -- t[2891] = 0
      "000000" when "0000101101001100", -- t[2892] = 0
      "000000" when "0000101101001101", -- t[2893] = 0
      "000000" when "0000101101001110", -- t[2894] = 0
      "000000" when "0000101101001111", -- t[2895] = 0
      "000000" when "0000101101010000", -- t[2896] = 0
      "000000" when "0000101101010001", -- t[2897] = 0
      "000000" when "0000101101010010", -- t[2898] = 0
      "000000" when "0000101101010011", -- t[2899] = 0
      "000000" when "0000101101010100", -- t[2900] = 0
      "000000" when "0000101101010101", -- t[2901] = 0
      "000000" when "0000101101010110", -- t[2902] = 0
      "000000" when "0000101101010111", -- t[2903] = 0
      "000000" when "0000101101011000", -- t[2904] = 0
      "000000" when "0000101101011001", -- t[2905] = 0
      "000000" when "0000101101011010", -- t[2906] = 0
      "000000" when "0000101101011011", -- t[2907] = 0
      "000000" when "0000101101011100", -- t[2908] = 0
      "000000" when "0000101101011101", -- t[2909] = 0
      "000000" when "0000101101011110", -- t[2910] = 0
      "000000" when "0000101101011111", -- t[2911] = 0
      "000000" when "0000101101100000", -- t[2912] = 0
      "000000" when "0000101101100001", -- t[2913] = 0
      "000000" when "0000101101100010", -- t[2914] = 0
      "000000" when "0000101101100011", -- t[2915] = 0
      "000000" when "0000101101100100", -- t[2916] = 0
      "000000" when "0000101101100101", -- t[2917] = 0
      "000000" when "0000101101100110", -- t[2918] = 0
      "000000" when "0000101101100111", -- t[2919] = 0
      "000000" when "0000101101101000", -- t[2920] = 0
      "000000" when "0000101101101001", -- t[2921] = 0
      "000000" when "0000101101101010", -- t[2922] = 0
      "000000" when "0000101101101011", -- t[2923] = 0
      "000000" when "0000101101101100", -- t[2924] = 0
      "000000" when "0000101101101101", -- t[2925] = 0
      "000000" when "0000101101101110", -- t[2926] = 0
      "000000" when "0000101101101111", -- t[2927] = 0
      "000000" when "0000101101110000", -- t[2928] = 0
      "000000" when "0000101101110001", -- t[2929] = 0
      "000000" when "0000101101110010", -- t[2930] = 0
      "000000" when "0000101101110011", -- t[2931] = 0
      "000000" when "0000101101110100", -- t[2932] = 0
      "000000" when "0000101101110101", -- t[2933] = 0
      "000000" when "0000101101110110", -- t[2934] = 0
      "000000" when "0000101101110111", -- t[2935] = 0
      "000000" when "0000101101111000", -- t[2936] = 0
      "000000" when "0000101101111001", -- t[2937] = 0
      "000000" when "0000101101111010", -- t[2938] = 0
      "000000" when "0000101101111011", -- t[2939] = 0
      "000000" when "0000101101111100", -- t[2940] = 0
      "000000" when "0000101101111101", -- t[2941] = 0
      "000000" when "0000101101111110", -- t[2942] = 0
      "000000" when "0000101101111111", -- t[2943] = 0
      "000000" when "0000101110000000", -- t[2944] = 0
      "000000" when "0000101110000001", -- t[2945] = 0
      "000000" when "0000101110000010", -- t[2946] = 0
      "000000" when "0000101110000011", -- t[2947] = 0
      "000000" when "0000101110000100", -- t[2948] = 0
      "000000" when "0000101110000101", -- t[2949] = 0
      "000000" when "0000101110000110", -- t[2950] = 0
      "000000" when "0000101110000111", -- t[2951] = 0
      "000000" when "0000101110001000", -- t[2952] = 0
      "000000" when "0000101110001001", -- t[2953] = 0
      "000000" when "0000101110001010", -- t[2954] = 0
      "000000" when "0000101110001011", -- t[2955] = 0
      "000000" when "0000101110001100", -- t[2956] = 0
      "000000" when "0000101110001101", -- t[2957] = 0
      "000000" when "0000101110001110", -- t[2958] = 0
      "000000" when "0000101110001111", -- t[2959] = 0
      "000000" when "0000101110010000", -- t[2960] = 0
      "000000" when "0000101110010001", -- t[2961] = 0
      "000000" when "0000101110010010", -- t[2962] = 0
      "000000" when "0000101110010011", -- t[2963] = 0
      "000000" when "0000101110010100", -- t[2964] = 0
      "000000" when "0000101110010101", -- t[2965] = 0
      "000000" when "0000101110010110", -- t[2966] = 0
      "000000" when "0000101110010111", -- t[2967] = 0
      "000000" when "0000101110011000", -- t[2968] = 0
      "000000" when "0000101110011001", -- t[2969] = 0
      "000000" when "0000101110011010", -- t[2970] = 0
      "000000" when "0000101110011011", -- t[2971] = 0
      "000000" when "0000101110011100", -- t[2972] = 0
      "000000" when "0000101110011101", -- t[2973] = 0
      "000000" when "0000101110011110", -- t[2974] = 0
      "000000" when "0000101110011111", -- t[2975] = 0
      "000000" when "0000101110100000", -- t[2976] = 0
      "000000" when "0000101110100001", -- t[2977] = 0
      "000000" when "0000101110100010", -- t[2978] = 0
      "000000" when "0000101110100011", -- t[2979] = 0
      "000000" when "0000101110100100", -- t[2980] = 0
      "000000" when "0000101110100101", -- t[2981] = 0
      "000000" when "0000101110100110", -- t[2982] = 0
      "000000" when "0000101110100111", -- t[2983] = 0
      "000000" when "0000101110101000", -- t[2984] = 0
      "000000" when "0000101110101001", -- t[2985] = 0
      "000000" when "0000101110101010", -- t[2986] = 0
      "000000" when "0000101110101011", -- t[2987] = 0
      "000000" when "0000101110101100", -- t[2988] = 0
      "000000" when "0000101110101101", -- t[2989] = 0
      "000000" when "0000101110101110", -- t[2990] = 0
      "000000" when "0000101110101111", -- t[2991] = 0
      "000000" when "0000101110110000", -- t[2992] = 0
      "000000" when "0000101110110001", -- t[2993] = 0
      "000000" when "0000101110110010", -- t[2994] = 0
      "000000" when "0000101110110011", -- t[2995] = 0
      "000000" when "0000101110110100", -- t[2996] = 0
      "000000" when "0000101110110101", -- t[2997] = 0
      "000000" when "0000101110110110", -- t[2998] = 0
      "000000" when "0000101110110111", -- t[2999] = 0
      "000000" when "0000101110111000", -- t[3000] = 0
      "000000" when "0000101110111001", -- t[3001] = 0
      "000000" when "0000101110111010", -- t[3002] = 0
      "000000" when "0000101110111011", -- t[3003] = 0
      "000000" when "0000101110111100", -- t[3004] = 0
      "000000" when "0000101110111101", -- t[3005] = 0
      "000000" when "0000101110111110", -- t[3006] = 0
      "000000" when "0000101110111111", -- t[3007] = 0
      "000000" when "0000101111000000", -- t[3008] = 0
      "000000" when "0000101111000001", -- t[3009] = 0
      "000000" when "0000101111000010", -- t[3010] = 0
      "000000" when "0000101111000011", -- t[3011] = 0
      "000000" when "0000101111000100", -- t[3012] = 0
      "000000" when "0000101111000101", -- t[3013] = 0
      "000000" when "0000101111000110", -- t[3014] = 0
      "000000" when "0000101111000111", -- t[3015] = 0
      "000000" when "0000101111001000", -- t[3016] = 0
      "000000" when "0000101111001001", -- t[3017] = 0
      "000000" when "0000101111001010", -- t[3018] = 0
      "000000" when "0000101111001011", -- t[3019] = 0
      "000000" when "0000101111001100", -- t[3020] = 0
      "000000" when "0000101111001101", -- t[3021] = 0
      "000000" when "0000101111001110", -- t[3022] = 0
      "000000" when "0000101111001111", -- t[3023] = 0
      "000000" when "0000101111010000", -- t[3024] = 0
      "000000" when "0000101111010001", -- t[3025] = 0
      "000000" when "0000101111010010", -- t[3026] = 0
      "000000" when "0000101111010011", -- t[3027] = 0
      "000000" when "0000101111010100", -- t[3028] = 0
      "000000" when "0000101111010101", -- t[3029] = 0
      "000000" when "0000101111010110", -- t[3030] = 0
      "000000" when "0000101111010111", -- t[3031] = 0
      "000000" when "0000101111011000", -- t[3032] = 0
      "000000" when "0000101111011001", -- t[3033] = 0
      "000000" when "0000101111011010", -- t[3034] = 0
      "000000" when "0000101111011011", -- t[3035] = 0
      "000000" when "0000101111011100", -- t[3036] = 0
      "000000" when "0000101111011101", -- t[3037] = 0
      "000000" when "0000101111011110", -- t[3038] = 0
      "000000" when "0000101111011111", -- t[3039] = 0
      "000000" when "0000101111100000", -- t[3040] = 0
      "000000" when "0000101111100001", -- t[3041] = 0
      "000000" when "0000101111100010", -- t[3042] = 0
      "000000" when "0000101111100011", -- t[3043] = 0
      "000000" when "0000101111100100", -- t[3044] = 0
      "000000" when "0000101111100101", -- t[3045] = 0
      "000000" when "0000101111100110", -- t[3046] = 0
      "000000" when "0000101111100111", -- t[3047] = 0
      "000000" when "0000101111101000", -- t[3048] = 0
      "000000" when "0000101111101001", -- t[3049] = 0
      "000000" when "0000101111101010", -- t[3050] = 0
      "000000" when "0000101111101011", -- t[3051] = 0
      "000000" when "0000101111101100", -- t[3052] = 0
      "000000" when "0000101111101101", -- t[3053] = 0
      "000000" when "0000101111101110", -- t[3054] = 0
      "000000" when "0000101111101111", -- t[3055] = 0
      "000000" when "0000101111110000", -- t[3056] = 0
      "000000" when "0000101111110001", -- t[3057] = 0
      "000000" when "0000101111110010", -- t[3058] = 0
      "000000" when "0000101111110011", -- t[3059] = 0
      "000000" when "0000101111110100", -- t[3060] = 0
      "000000" when "0000101111110101", -- t[3061] = 0
      "000000" when "0000101111110110", -- t[3062] = 0
      "000000" when "0000101111110111", -- t[3063] = 0
      "000000" when "0000101111111000", -- t[3064] = 0
      "000000" when "0000101111111001", -- t[3065] = 0
      "000000" when "0000101111111010", -- t[3066] = 0
      "000000" when "0000101111111011", -- t[3067] = 0
      "000000" when "0000101111111100", -- t[3068] = 0
      "000000" when "0000101111111101", -- t[3069] = 0
      "000000" when "0000101111111110", -- t[3070] = 0
      "000000" when "0000101111111111", -- t[3071] = 0
      "000000" when "0000110000000000", -- t[3072] = 0
      "000000" when "0000110000000001", -- t[3073] = 0
      "000000" when "0000110000000010", -- t[3074] = 0
      "000000" when "0000110000000011", -- t[3075] = 0
      "000000" when "0000110000000100", -- t[3076] = 0
      "000000" when "0000110000000101", -- t[3077] = 0
      "000000" when "0000110000000110", -- t[3078] = 0
      "000000" when "0000110000000111", -- t[3079] = 0
      "000000" when "0000110000001000", -- t[3080] = 0
      "000000" when "0000110000001001", -- t[3081] = 0
      "000000" when "0000110000001010", -- t[3082] = 0
      "000000" when "0000110000001011", -- t[3083] = 0
      "000000" when "0000110000001100", -- t[3084] = 0
      "000000" when "0000110000001101", -- t[3085] = 0
      "000000" when "0000110000001110", -- t[3086] = 0
      "000000" when "0000110000001111", -- t[3087] = 0
      "000000" when "0000110000010000", -- t[3088] = 0
      "000000" when "0000110000010001", -- t[3089] = 0
      "000000" when "0000110000010010", -- t[3090] = 0
      "000000" when "0000110000010011", -- t[3091] = 0
      "000000" when "0000110000010100", -- t[3092] = 0
      "000000" when "0000110000010101", -- t[3093] = 0
      "000000" when "0000110000010110", -- t[3094] = 0
      "000000" when "0000110000010111", -- t[3095] = 0
      "000000" when "0000110000011000", -- t[3096] = 0
      "000000" when "0000110000011001", -- t[3097] = 0
      "000000" when "0000110000011010", -- t[3098] = 0
      "000000" when "0000110000011011", -- t[3099] = 0
      "000000" when "0000110000011100", -- t[3100] = 0
      "000000" when "0000110000011101", -- t[3101] = 0
      "000000" when "0000110000011110", -- t[3102] = 0
      "000000" when "0000110000011111", -- t[3103] = 0
      "000000" when "0000110000100000", -- t[3104] = 0
      "000000" when "0000110000100001", -- t[3105] = 0
      "000000" when "0000110000100010", -- t[3106] = 0
      "000000" when "0000110000100011", -- t[3107] = 0
      "000000" when "0000110000100100", -- t[3108] = 0
      "000000" when "0000110000100101", -- t[3109] = 0
      "000000" when "0000110000100110", -- t[3110] = 0
      "000000" when "0000110000100111", -- t[3111] = 0
      "000000" when "0000110000101000", -- t[3112] = 0
      "000000" when "0000110000101001", -- t[3113] = 0
      "000000" when "0000110000101010", -- t[3114] = 0
      "000000" when "0000110000101011", -- t[3115] = 0
      "000000" when "0000110000101100", -- t[3116] = 0
      "000000" when "0000110000101101", -- t[3117] = 0
      "000000" when "0000110000101110", -- t[3118] = 0
      "000000" when "0000110000101111", -- t[3119] = 0
      "000000" when "0000110000110000", -- t[3120] = 0
      "000000" when "0000110000110001", -- t[3121] = 0
      "000000" when "0000110000110010", -- t[3122] = 0
      "000000" when "0000110000110011", -- t[3123] = 0
      "000000" when "0000110000110100", -- t[3124] = 0
      "000000" when "0000110000110101", -- t[3125] = 0
      "000000" when "0000110000110110", -- t[3126] = 0
      "000000" when "0000110000110111", -- t[3127] = 0
      "000000" when "0000110000111000", -- t[3128] = 0
      "000000" when "0000110000111001", -- t[3129] = 0
      "000000" when "0000110000111010", -- t[3130] = 0
      "000000" when "0000110000111011", -- t[3131] = 0
      "000000" when "0000110000111100", -- t[3132] = 0
      "000000" when "0000110000111101", -- t[3133] = 0
      "000000" when "0000110000111110", -- t[3134] = 0
      "000000" when "0000110000111111", -- t[3135] = 0
      "000000" when "0000110001000000", -- t[3136] = 0
      "000000" when "0000110001000001", -- t[3137] = 0
      "000000" when "0000110001000010", -- t[3138] = 0
      "000000" when "0000110001000011", -- t[3139] = 0
      "000000" when "0000110001000100", -- t[3140] = 0
      "000000" when "0000110001000101", -- t[3141] = 0
      "000000" when "0000110001000110", -- t[3142] = 0
      "000000" when "0000110001000111", -- t[3143] = 0
      "000000" when "0000110001001000", -- t[3144] = 0
      "000000" when "0000110001001001", -- t[3145] = 0
      "000000" when "0000110001001010", -- t[3146] = 0
      "000000" when "0000110001001011", -- t[3147] = 0
      "000000" when "0000110001001100", -- t[3148] = 0
      "000000" when "0000110001001101", -- t[3149] = 0
      "000000" when "0000110001001110", -- t[3150] = 0
      "000000" when "0000110001001111", -- t[3151] = 0
      "000000" when "0000110001010000", -- t[3152] = 0
      "000000" when "0000110001010001", -- t[3153] = 0
      "000000" when "0000110001010010", -- t[3154] = 0
      "000000" when "0000110001010011", -- t[3155] = 0
      "000000" when "0000110001010100", -- t[3156] = 0
      "000000" when "0000110001010101", -- t[3157] = 0
      "000000" when "0000110001010110", -- t[3158] = 0
      "000000" when "0000110001010111", -- t[3159] = 0
      "000000" when "0000110001011000", -- t[3160] = 0
      "000000" when "0000110001011001", -- t[3161] = 0
      "000000" when "0000110001011010", -- t[3162] = 0
      "000000" when "0000110001011011", -- t[3163] = 0
      "000000" when "0000110001011100", -- t[3164] = 0
      "000000" when "0000110001011101", -- t[3165] = 0
      "000000" when "0000110001011110", -- t[3166] = 0
      "000000" when "0000110001011111", -- t[3167] = 0
      "000000" when "0000110001100000", -- t[3168] = 0
      "000000" when "0000110001100001", -- t[3169] = 0
      "000000" when "0000110001100010", -- t[3170] = 0
      "000000" when "0000110001100011", -- t[3171] = 0
      "000000" when "0000110001100100", -- t[3172] = 0
      "000000" when "0000110001100101", -- t[3173] = 0
      "000000" when "0000110001100110", -- t[3174] = 0
      "000000" when "0000110001100111", -- t[3175] = 0
      "000000" when "0000110001101000", -- t[3176] = 0
      "000000" when "0000110001101001", -- t[3177] = 0
      "000000" when "0000110001101010", -- t[3178] = 0
      "000000" when "0000110001101011", -- t[3179] = 0
      "000000" when "0000110001101100", -- t[3180] = 0
      "000000" when "0000110001101101", -- t[3181] = 0
      "000000" when "0000110001101110", -- t[3182] = 0
      "000000" when "0000110001101111", -- t[3183] = 0
      "000000" when "0000110001110000", -- t[3184] = 0
      "000000" when "0000110001110001", -- t[3185] = 0
      "000000" when "0000110001110010", -- t[3186] = 0
      "000000" when "0000110001110011", -- t[3187] = 0
      "000000" when "0000110001110100", -- t[3188] = 0
      "000000" when "0000110001110101", -- t[3189] = 0
      "000000" when "0000110001110110", -- t[3190] = 0
      "000000" when "0000110001110111", -- t[3191] = 0
      "000000" when "0000110001111000", -- t[3192] = 0
      "000000" when "0000110001111001", -- t[3193] = 0
      "000000" when "0000110001111010", -- t[3194] = 0
      "000000" when "0000110001111011", -- t[3195] = 0
      "000000" when "0000110001111100", -- t[3196] = 0
      "000000" when "0000110001111101", -- t[3197] = 0
      "000000" when "0000110001111110", -- t[3198] = 0
      "000000" when "0000110001111111", -- t[3199] = 0
      "000000" when "0000110010000000", -- t[3200] = 0
      "000000" when "0000110010000001", -- t[3201] = 0
      "000000" when "0000110010000010", -- t[3202] = 0
      "000000" when "0000110010000011", -- t[3203] = 0
      "000000" when "0000110010000100", -- t[3204] = 0
      "000000" when "0000110010000101", -- t[3205] = 0
      "000000" when "0000110010000110", -- t[3206] = 0
      "000000" when "0000110010000111", -- t[3207] = 0
      "000000" when "0000110010001000", -- t[3208] = 0
      "000000" when "0000110010001001", -- t[3209] = 0
      "000000" when "0000110010001010", -- t[3210] = 0
      "000000" when "0000110010001011", -- t[3211] = 0
      "000000" when "0000110010001100", -- t[3212] = 0
      "000000" when "0000110010001101", -- t[3213] = 0
      "000000" when "0000110010001110", -- t[3214] = 0
      "000000" when "0000110010001111", -- t[3215] = 0
      "000000" when "0000110010010000", -- t[3216] = 0
      "000000" when "0000110010010001", -- t[3217] = 0
      "000000" when "0000110010010010", -- t[3218] = 0
      "000000" when "0000110010010011", -- t[3219] = 0
      "000000" when "0000110010010100", -- t[3220] = 0
      "000000" when "0000110010010101", -- t[3221] = 0
      "000000" when "0000110010010110", -- t[3222] = 0
      "000000" when "0000110010010111", -- t[3223] = 0
      "000000" when "0000110010011000", -- t[3224] = 0
      "000000" when "0000110010011001", -- t[3225] = 0
      "000000" when "0000110010011010", -- t[3226] = 0
      "000000" when "0000110010011011", -- t[3227] = 0
      "000000" when "0000110010011100", -- t[3228] = 0
      "000000" when "0000110010011101", -- t[3229] = 0
      "000000" when "0000110010011110", -- t[3230] = 0
      "000000" when "0000110010011111", -- t[3231] = 0
      "000000" when "0000110010100000", -- t[3232] = 0
      "000000" when "0000110010100001", -- t[3233] = 0
      "000000" when "0000110010100010", -- t[3234] = 0
      "000000" when "0000110010100011", -- t[3235] = 0
      "000000" when "0000110010100100", -- t[3236] = 0
      "000000" when "0000110010100101", -- t[3237] = 0
      "000000" when "0000110010100110", -- t[3238] = 0
      "000000" when "0000110010100111", -- t[3239] = 0
      "000000" when "0000110010101000", -- t[3240] = 0
      "000000" when "0000110010101001", -- t[3241] = 0
      "000000" when "0000110010101010", -- t[3242] = 0
      "000000" when "0000110010101011", -- t[3243] = 0
      "000000" when "0000110010101100", -- t[3244] = 0
      "000000" when "0000110010101101", -- t[3245] = 0
      "000000" when "0000110010101110", -- t[3246] = 0
      "000000" when "0000110010101111", -- t[3247] = 0
      "000000" when "0000110010110000", -- t[3248] = 0
      "000000" when "0000110010110001", -- t[3249] = 0
      "000000" when "0000110010110010", -- t[3250] = 0
      "000000" when "0000110010110011", -- t[3251] = 0
      "000000" when "0000110010110100", -- t[3252] = 0
      "000000" when "0000110010110101", -- t[3253] = 0
      "000000" when "0000110010110110", -- t[3254] = 0
      "000000" when "0000110010110111", -- t[3255] = 0
      "000000" when "0000110010111000", -- t[3256] = 0
      "000000" when "0000110010111001", -- t[3257] = 0
      "000000" when "0000110010111010", -- t[3258] = 0
      "000000" when "0000110010111011", -- t[3259] = 0
      "000000" when "0000110010111100", -- t[3260] = 0
      "000000" when "0000110010111101", -- t[3261] = 0
      "000000" when "0000110010111110", -- t[3262] = 0
      "000000" when "0000110010111111", -- t[3263] = 0
      "000000" when "0000110011000000", -- t[3264] = 0
      "000000" when "0000110011000001", -- t[3265] = 0
      "000000" when "0000110011000010", -- t[3266] = 0
      "000000" when "0000110011000011", -- t[3267] = 0
      "000000" when "0000110011000100", -- t[3268] = 0
      "000000" when "0000110011000101", -- t[3269] = 0
      "000000" when "0000110011000110", -- t[3270] = 0
      "000000" when "0000110011000111", -- t[3271] = 0
      "000000" when "0000110011001000", -- t[3272] = 0
      "000000" when "0000110011001001", -- t[3273] = 0
      "000000" when "0000110011001010", -- t[3274] = 0
      "000000" when "0000110011001011", -- t[3275] = 0
      "000000" when "0000110011001100", -- t[3276] = 0
      "000000" when "0000110011001101", -- t[3277] = 0
      "000000" when "0000110011001110", -- t[3278] = 0
      "000000" when "0000110011001111", -- t[3279] = 0
      "000000" when "0000110011010000", -- t[3280] = 0
      "000000" when "0000110011010001", -- t[3281] = 0
      "000000" when "0000110011010010", -- t[3282] = 0
      "000000" when "0000110011010011", -- t[3283] = 0
      "000000" when "0000110011010100", -- t[3284] = 0
      "000000" when "0000110011010101", -- t[3285] = 0
      "000000" when "0000110011010110", -- t[3286] = 0
      "000000" when "0000110011010111", -- t[3287] = 0
      "000000" when "0000110011011000", -- t[3288] = 0
      "000000" when "0000110011011001", -- t[3289] = 0
      "000000" when "0000110011011010", -- t[3290] = 0
      "000000" when "0000110011011011", -- t[3291] = 0
      "000000" when "0000110011011100", -- t[3292] = 0
      "000000" when "0000110011011101", -- t[3293] = 0
      "000000" when "0000110011011110", -- t[3294] = 0
      "000000" when "0000110011011111", -- t[3295] = 0
      "000000" when "0000110011100000", -- t[3296] = 0
      "000000" when "0000110011100001", -- t[3297] = 0
      "000000" when "0000110011100010", -- t[3298] = 0
      "000000" when "0000110011100011", -- t[3299] = 0
      "000000" when "0000110011100100", -- t[3300] = 0
      "000000" when "0000110011100101", -- t[3301] = 0
      "000000" when "0000110011100110", -- t[3302] = 0
      "000000" when "0000110011100111", -- t[3303] = 0
      "000000" when "0000110011101000", -- t[3304] = 0
      "000000" when "0000110011101001", -- t[3305] = 0
      "000000" when "0000110011101010", -- t[3306] = 0
      "000000" when "0000110011101011", -- t[3307] = 0
      "000000" when "0000110011101100", -- t[3308] = 0
      "000000" when "0000110011101101", -- t[3309] = 0
      "000000" when "0000110011101110", -- t[3310] = 0
      "000000" when "0000110011101111", -- t[3311] = 0
      "000000" when "0000110011110000", -- t[3312] = 0
      "000000" when "0000110011110001", -- t[3313] = 0
      "000000" when "0000110011110010", -- t[3314] = 0
      "000000" when "0000110011110011", -- t[3315] = 0
      "000000" when "0000110011110100", -- t[3316] = 0
      "000000" when "0000110011110101", -- t[3317] = 0
      "000000" when "0000110011110110", -- t[3318] = 0
      "000000" when "0000110011110111", -- t[3319] = 0
      "000000" when "0000110011111000", -- t[3320] = 0
      "000000" when "0000110011111001", -- t[3321] = 0
      "000000" when "0000110011111010", -- t[3322] = 0
      "000000" when "0000110011111011", -- t[3323] = 0
      "000000" when "0000110011111100", -- t[3324] = 0
      "000000" when "0000110011111101", -- t[3325] = 0
      "000000" when "0000110011111110", -- t[3326] = 0
      "000000" when "0000110011111111", -- t[3327] = 0
      "000000" when "0000110100000000", -- t[3328] = 0
      "000000" when "0000110100000001", -- t[3329] = 0
      "000000" when "0000110100000010", -- t[3330] = 0
      "000000" when "0000110100000011", -- t[3331] = 0
      "000000" when "0000110100000100", -- t[3332] = 0
      "000000" when "0000110100000101", -- t[3333] = 0
      "000000" when "0000110100000110", -- t[3334] = 0
      "000000" when "0000110100000111", -- t[3335] = 0
      "000000" when "0000110100001000", -- t[3336] = 0
      "000000" when "0000110100001001", -- t[3337] = 0
      "000000" when "0000110100001010", -- t[3338] = 0
      "000000" when "0000110100001011", -- t[3339] = 0
      "000000" when "0000110100001100", -- t[3340] = 0
      "000000" when "0000110100001101", -- t[3341] = 0
      "000000" when "0000110100001110", -- t[3342] = 0
      "000000" when "0000110100001111", -- t[3343] = 0
      "000000" when "0000110100010000", -- t[3344] = 0
      "000000" when "0000110100010001", -- t[3345] = 0
      "000000" when "0000110100010010", -- t[3346] = 0
      "000000" when "0000110100010011", -- t[3347] = 0
      "000000" when "0000110100010100", -- t[3348] = 0
      "000000" when "0000110100010101", -- t[3349] = 0
      "000000" when "0000110100010110", -- t[3350] = 0
      "000000" when "0000110100010111", -- t[3351] = 0
      "000000" when "0000110100011000", -- t[3352] = 0
      "000000" when "0000110100011001", -- t[3353] = 0
      "000000" when "0000110100011010", -- t[3354] = 0
      "000000" when "0000110100011011", -- t[3355] = 0
      "000000" when "0000110100011100", -- t[3356] = 0
      "000000" when "0000110100011101", -- t[3357] = 0
      "000000" when "0000110100011110", -- t[3358] = 0
      "000000" when "0000110100011111", -- t[3359] = 0
      "000000" when "0000110100100000", -- t[3360] = 0
      "000000" when "0000110100100001", -- t[3361] = 0
      "000000" when "0000110100100010", -- t[3362] = 0
      "000000" when "0000110100100011", -- t[3363] = 0
      "000000" when "0000110100100100", -- t[3364] = 0
      "000000" when "0000110100100101", -- t[3365] = 0
      "000000" when "0000110100100110", -- t[3366] = 0
      "000000" when "0000110100100111", -- t[3367] = 0
      "000000" when "0000110100101000", -- t[3368] = 0
      "000000" when "0000110100101001", -- t[3369] = 0
      "000000" when "0000110100101010", -- t[3370] = 0
      "000000" when "0000110100101011", -- t[3371] = 0
      "000000" when "0000110100101100", -- t[3372] = 0
      "000000" when "0000110100101101", -- t[3373] = 0
      "000000" when "0000110100101110", -- t[3374] = 0
      "000000" when "0000110100101111", -- t[3375] = 0
      "000000" when "0000110100110000", -- t[3376] = 0
      "000000" when "0000110100110001", -- t[3377] = 0
      "000000" when "0000110100110010", -- t[3378] = 0
      "000000" when "0000110100110011", -- t[3379] = 0
      "000000" when "0000110100110100", -- t[3380] = 0
      "000000" when "0000110100110101", -- t[3381] = 0
      "000000" when "0000110100110110", -- t[3382] = 0
      "000000" when "0000110100110111", -- t[3383] = 0
      "000000" when "0000110100111000", -- t[3384] = 0
      "000000" when "0000110100111001", -- t[3385] = 0
      "000000" when "0000110100111010", -- t[3386] = 0
      "000000" when "0000110100111011", -- t[3387] = 0
      "000000" when "0000110100111100", -- t[3388] = 0
      "000000" when "0000110100111101", -- t[3389] = 0
      "000000" when "0000110100111110", -- t[3390] = 0
      "000000" when "0000110100111111", -- t[3391] = 0
      "000000" when "0000110101000000", -- t[3392] = 0
      "000000" when "0000110101000001", -- t[3393] = 0
      "000000" when "0000110101000010", -- t[3394] = 0
      "000000" when "0000110101000011", -- t[3395] = 0
      "000000" when "0000110101000100", -- t[3396] = 0
      "000000" when "0000110101000101", -- t[3397] = 0
      "000000" when "0000110101000110", -- t[3398] = 0
      "000000" when "0000110101000111", -- t[3399] = 0
      "000000" when "0000110101001000", -- t[3400] = 0
      "000000" when "0000110101001001", -- t[3401] = 0
      "000000" when "0000110101001010", -- t[3402] = 0
      "000000" when "0000110101001011", -- t[3403] = 0
      "000000" when "0000110101001100", -- t[3404] = 0
      "000000" when "0000110101001101", -- t[3405] = 0
      "000000" when "0000110101001110", -- t[3406] = 0
      "000000" when "0000110101001111", -- t[3407] = 0
      "000000" when "0000110101010000", -- t[3408] = 0
      "000000" when "0000110101010001", -- t[3409] = 0
      "000000" when "0000110101010010", -- t[3410] = 0
      "000000" when "0000110101010011", -- t[3411] = 0
      "000000" when "0000110101010100", -- t[3412] = 0
      "000000" when "0000110101010101", -- t[3413] = 0
      "000000" when "0000110101010110", -- t[3414] = 0
      "000000" when "0000110101010111", -- t[3415] = 0
      "000000" when "0000110101011000", -- t[3416] = 0
      "000000" when "0000110101011001", -- t[3417] = 0
      "000000" when "0000110101011010", -- t[3418] = 0
      "000000" when "0000110101011011", -- t[3419] = 0
      "000000" when "0000110101011100", -- t[3420] = 0
      "000000" when "0000110101011101", -- t[3421] = 0
      "000000" when "0000110101011110", -- t[3422] = 0
      "000000" when "0000110101011111", -- t[3423] = 0
      "000000" when "0000110101100000", -- t[3424] = 0
      "000000" when "0000110101100001", -- t[3425] = 0
      "000000" when "0000110101100010", -- t[3426] = 0
      "000000" when "0000110101100011", -- t[3427] = 0
      "000000" when "0000110101100100", -- t[3428] = 0
      "000000" when "0000110101100101", -- t[3429] = 0
      "000000" when "0000110101100110", -- t[3430] = 0
      "000000" when "0000110101100111", -- t[3431] = 0
      "000000" when "0000110101101000", -- t[3432] = 0
      "000000" when "0000110101101001", -- t[3433] = 0
      "000000" when "0000110101101010", -- t[3434] = 0
      "000000" when "0000110101101011", -- t[3435] = 0
      "000000" when "0000110101101100", -- t[3436] = 0
      "000000" when "0000110101101101", -- t[3437] = 0
      "000000" when "0000110101101110", -- t[3438] = 0
      "000000" when "0000110101101111", -- t[3439] = 0
      "000000" when "0000110101110000", -- t[3440] = 0
      "000000" when "0000110101110001", -- t[3441] = 0
      "000000" when "0000110101110010", -- t[3442] = 0
      "000000" when "0000110101110011", -- t[3443] = 0
      "000000" when "0000110101110100", -- t[3444] = 0
      "000000" when "0000110101110101", -- t[3445] = 0
      "000000" when "0000110101110110", -- t[3446] = 0
      "000000" when "0000110101110111", -- t[3447] = 0
      "000000" when "0000110101111000", -- t[3448] = 0
      "000000" when "0000110101111001", -- t[3449] = 0
      "000000" when "0000110101111010", -- t[3450] = 0
      "000000" when "0000110101111011", -- t[3451] = 0
      "000000" when "0000110101111100", -- t[3452] = 0
      "000000" when "0000110101111101", -- t[3453] = 0
      "000000" when "0000110101111110", -- t[3454] = 0
      "000000" when "0000110101111111", -- t[3455] = 0
      "000000" when "0000110110000000", -- t[3456] = 0
      "000000" when "0000110110000001", -- t[3457] = 0
      "000000" when "0000110110000010", -- t[3458] = 0
      "000000" when "0000110110000011", -- t[3459] = 0
      "000000" when "0000110110000100", -- t[3460] = 0
      "000000" when "0000110110000101", -- t[3461] = 0
      "000000" when "0000110110000110", -- t[3462] = 0
      "000000" when "0000110110000111", -- t[3463] = 0
      "000000" when "0000110110001000", -- t[3464] = 0
      "000000" when "0000110110001001", -- t[3465] = 0
      "000000" when "0000110110001010", -- t[3466] = 0
      "000000" when "0000110110001011", -- t[3467] = 0
      "000000" when "0000110110001100", -- t[3468] = 0
      "000000" when "0000110110001101", -- t[3469] = 0
      "000000" when "0000110110001110", -- t[3470] = 0
      "000000" when "0000110110001111", -- t[3471] = 0
      "000000" when "0000110110010000", -- t[3472] = 0
      "000000" when "0000110110010001", -- t[3473] = 0
      "000000" when "0000110110010010", -- t[3474] = 0
      "000000" when "0000110110010011", -- t[3475] = 0
      "000000" when "0000110110010100", -- t[3476] = 0
      "000000" when "0000110110010101", -- t[3477] = 0
      "000000" when "0000110110010110", -- t[3478] = 0
      "000000" when "0000110110010111", -- t[3479] = 0
      "000000" when "0000110110011000", -- t[3480] = 0
      "000000" when "0000110110011001", -- t[3481] = 0
      "000000" when "0000110110011010", -- t[3482] = 0
      "000000" when "0000110110011011", -- t[3483] = 0
      "000000" when "0000110110011100", -- t[3484] = 0
      "000000" when "0000110110011101", -- t[3485] = 0
      "000000" when "0000110110011110", -- t[3486] = 0
      "000000" when "0000110110011111", -- t[3487] = 0
      "000000" when "0000110110100000", -- t[3488] = 0
      "000000" when "0000110110100001", -- t[3489] = 0
      "000000" when "0000110110100010", -- t[3490] = 0
      "000000" when "0000110110100011", -- t[3491] = 0
      "000000" when "0000110110100100", -- t[3492] = 0
      "000000" when "0000110110100101", -- t[3493] = 0
      "000000" when "0000110110100110", -- t[3494] = 0
      "000000" when "0000110110100111", -- t[3495] = 0
      "000000" when "0000110110101000", -- t[3496] = 0
      "000000" when "0000110110101001", -- t[3497] = 0
      "000000" when "0000110110101010", -- t[3498] = 0
      "000000" when "0000110110101011", -- t[3499] = 0
      "000000" when "0000110110101100", -- t[3500] = 0
      "000000" when "0000110110101101", -- t[3501] = 0
      "000000" when "0000110110101110", -- t[3502] = 0
      "000000" when "0000110110101111", -- t[3503] = 0
      "000000" when "0000110110110000", -- t[3504] = 0
      "000000" when "0000110110110001", -- t[3505] = 0
      "000000" when "0000110110110010", -- t[3506] = 0
      "000000" when "0000110110110011", -- t[3507] = 0
      "000000" when "0000110110110100", -- t[3508] = 0
      "000000" when "0000110110110101", -- t[3509] = 0
      "000000" when "0000110110110110", -- t[3510] = 0
      "000000" when "0000110110110111", -- t[3511] = 0
      "000000" when "0000110110111000", -- t[3512] = 0
      "000000" when "0000110110111001", -- t[3513] = 0
      "000000" when "0000110110111010", -- t[3514] = 0
      "000000" when "0000110110111011", -- t[3515] = 0
      "000000" when "0000110110111100", -- t[3516] = 0
      "000000" when "0000110110111101", -- t[3517] = 0
      "000000" when "0000110110111110", -- t[3518] = 0
      "000000" when "0000110110111111", -- t[3519] = 0
      "000000" when "0000110111000000", -- t[3520] = 0
      "000000" when "0000110111000001", -- t[3521] = 0
      "000000" when "0000110111000010", -- t[3522] = 0
      "000000" when "0000110111000011", -- t[3523] = 0
      "000000" when "0000110111000100", -- t[3524] = 0
      "000000" when "0000110111000101", -- t[3525] = 0
      "000000" when "0000110111000110", -- t[3526] = 0
      "000000" when "0000110111000111", -- t[3527] = 0
      "000000" when "0000110111001000", -- t[3528] = 0
      "000000" when "0000110111001001", -- t[3529] = 0
      "000000" when "0000110111001010", -- t[3530] = 0
      "000000" when "0000110111001011", -- t[3531] = 0
      "000000" when "0000110111001100", -- t[3532] = 0
      "000000" when "0000110111001101", -- t[3533] = 0
      "000000" when "0000110111001110", -- t[3534] = 0
      "000000" when "0000110111001111", -- t[3535] = 0
      "000000" when "0000110111010000", -- t[3536] = 0
      "000000" when "0000110111010001", -- t[3537] = 0
      "000000" when "0000110111010010", -- t[3538] = 0
      "000000" when "0000110111010011", -- t[3539] = 0
      "000000" when "0000110111010100", -- t[3540] = 0
      "000000" when "0000110111010101", -- t[3541] = 0
      "000000" when "0000110111010110", -- t[3542] = 0
      "000000" when "0000110111010111", -- t[3543] = 0
      "000000" when "0000110111011000", -- t[3544] = 0
      "000000" when "0000110111011001", -- t[3545] = 0
      "000000" when "0000110111011010", -- t[3546] = 0
      "000000" when "0000110111011011", -- t[3547] = 0
      "000000" when "0000110111011100", -- t[3548] = 0
      "000000" when "0000110111011101", -- t[3549] = 0
      "000000" when "0000110111011110", -- t[3550] = 0
      "000000" when "0000110111011111", -- t[3551] = 0
      "000000" when "0000110111100000", -- t[3552] = 0
      "000000" when "0000110111100001", -- t[3553] = 0
      "000000" when "0000110111100010", -- t[3554] = 0
      "000000" when "0000110111100011", -- t[3555] = 0
      "000000" when "0000110111100100", -- t[3556] = 0
      "000000" when "0000110111100101", -- t[3557] = 0
      "000000" when "0000110111100110", -- t[3558] = 0
      "000000" when "0000110111100111", -- t[3559] = 0
      "000000" when "0000110111101000", -- t[3560] = 0
      "000000" when "0000110111101001", -- t[3561] = 0
      "000000" when "0000110111101010", -- t[3562] = 0
      "000000" when "0000110111101011", -- t[3563] = 0
      "000000" when "0000110111101100", -- t[3564] = 0
      "000000" when "0000110111101101", -- t[3565] = 0
      "000000" when "0000110111101110", -- t[3566] = 0
      "000000" when "0000110111101111", -- t[3567] = 0
      "000000" when "0000110111110000", -- t[3568] = 0
      "000000" when "0000110111110001", -- t[3569] = 0
      "000000" when "0000110111110010", -- t[3570] = 0
      "000000" when "0000110111110011", -- t[3571] = 0
      "000000" when "0000110111110100", -- t[3572] = 0
      "000000" when "0000110111110101", -- t[3573] = 0
      "000000" when "0000110111110110", -- t[3574] = 0
      "000000" when "0000110111110111", -- t[3575] = 0
      "000000" when "0000110111111000", -- t[3576] = 0
      "000000" when "0000110111111001", -- t[3577] = 0
      "000000" when "0000110111111010", -- t[3578] = 0
      "000000" when "0000110111111011", -- t[3579] = 0
      "000000" when "0000110111111100", -- t[3580] = 0
      "000000" when "0000110111111101", -- t[3581] = 0
      "000000" when "0000110111111110", -- t[3582] = 0
      "000000" when "0000110111111111", -- t[3583] = 0
      "000000" when "0000111000000000", -- t[3584] = 0
      "000000" when "0000111000000001", -- t[3585] = 0
      "000000" when "0000111000000010", -- t[3586] = 0
      "000000" when "0000111000000011", -- t[3587] = 0
      "000000" when "0000111000000100", -- t[3588] = 0
      "000000" when "0000111000000101", -- t[3589] = 0
      "000000" when "0000111000000110", -- t[3590] = 0
      "000000" when "0000111000000111", -- t[3591] = 0
      "000000" when "0000111000001000", -- t[3592] = 0
      "000000" when "0000111000001001", -- t[3593] = 0
      "000000" when "0000111000001010", -- t[3594] = 0
      "000000" when "0000111000001011", -- t[3595] = 0
      "000000" when "0000111000001100", -- t[3596] = 0
      "000000" when "0000111000001101", -- t[3597] = 0
      "000000" when "0000111000001110", -- t[3598] = 0
      "000000" when "0000111000001111", -- t[3599] = 0
      "000000" when "0000111000010000", -- t[3600] = 0
      "000000" when "0000111000010001", -- t[3601] = 0
      "000000" when "0000111000010010", -- t[3602] = 0
      "000000" when "0000111000010011", -- t[3603] = 0
      "000000" when "0000111000010100", -- t[3604] = 0
      "000000" when "0000111000010101", -- t[3605] = 0
      "000000" when "0000111000010110", -- t[3606] = 0
      "000000" when "0000111000010111", -- t[3607] = 0
      "000000" when "0000111000011000", -- t[3608] = 0
      "000000" when "0000111000011001", -- t[3609] = 0
      "000000" when "0000111000011010", -- t[3610] = 0
      "000000" when "0000111000011011", -- t[3611] = 0
      "000000" when "0000111000011100", -- t[3612] = 0
      "000000" when "0000111000011101", -- t[3613] = 0
      "000000" when "0000111000011110", -- t[3614] = 0
      "000000" when "0000111000011111", -- t[3615] = 0
      "000000" when "0000111000100000", -- t[3616] = 0
      "000000" when "0000111000100001", -- t[3617] = 0
      "000000" when "0000111000100010", -- t[3618] = 0
      "000000" when "0000111000100011", -- t[3619] = 0
      "000000" when "0000111000100100", -- t[3620] = 0
      "000000" when "0000111000100101", -- t[3621] = 0
      "000000" when "0000111000100110", -- t[3622] = 0
      "000000" when "0000111000100111", -- t[3623] = 0
      "000000" when "0000111000101000", -- t[3624] = 0
      "000000" when "0000111000101001", -- t[3625] = 0
      "000000" when "0000111000101010", -- t[3626] = 0
      "000000" when "0000111000101011", -- t[3627] = 0
      "000000" when "0000111000101100", -- t[3628] = 0
      "000000" when "0000111000101101", -- t[3629] = 0
      "000000" when "0000111000101110", -- t[3630] = 0
      "000000" when "0000111000101111", -- t[3631] = 0
      "000000" when "0000111000110000", -- t[3632] = 0
      "000000" when "0000111000110001", -- t[3633] = 0
      "000000" when "0000111000110010", -- t[3634] = 0
      "000000" when "0000111000110011", -- t[3635] = 0
      "000000" when "0000111000110100", -- t[3636] = 0
      "000000" when "0000111000110101", -- t[3637] = 0
      "000000" when "0000111000110110", -- t[3638] = 0
      "000000" when "0000111000110111", -- t[3639] = 0
      "000000" when "0000111000111000", -- t[3640] = 0
      "000000" when "0000111000111001", -- t[3641] = 0
      "000000" when "0000111000111010", -- t[3642] = 0
      "000000" when "0000111000111011", -- t[3643] = 0
      "000000" when "0000111000111100", -- t[3644] = 0
      "000000" when "0000111000111101", -- t[3645] = 0
      "000000" when "0000111000111110", -- t[3646] = 0
      "000000" when "0000111000111111", -- t[3647] = 0
      "000000" when "0000111001000000", -- t[3648] = 0
      "000000" when "0000111001000001", -- t[3649] = 0
      "000000" when "0000111001000010", -- t[3650] = 0
      "000000" when "0000111001000011", -- t[3651] = 0
      "000000" when "0000111001000100", -- t[3652] = 0
      "000000" when "0000111001000101", -- t[3653] = 0
      "000000" when "0000111001000110", -- t[3654] = 0
      "000000" when "0000111001000111", -- t[3655] = 0
      "000000" when "0000111001001000", -- t[3656] = 0
      "000000" when "0000111001001001", -- t[3657] = 0
      "000000" when "0000111001001010", -- t[3658] = 0
      "000000" when "0000111001001011", -- t[3659] = 0
      "000000" when "0000111001001100", -- t[3660] = 0
      "000000" when "0000111001001101", -- t[3661] = 0
      "000000" when "0000111001001110", -- t[3662] = 0
      "000000" when "0000111001001111", -- t[3663] = 0
      "000000" when "0000111001010000", -- t[3664] = 0
      "000000" when "0000111001010001", -- t[3665] = 0
      "000000" when "0000111001010010", -- t[3666] = 0
      "000000" when "0000111001010011", -- t[3667] = 0
      "000000" when "0000111001010100", -- t[3668] = 0
      "000000" when "0000111001010101", -- t[3669] = 0
      "000000" when "0000111001010110", -- t[3670] = 0
      "000000" when "0000111001010111", -- t[3671] = 0
      "000000" when "0000111001011000", -- t[3672] = 0
      "000000" when "0000111001011001", -- t[3673] = 0
      "000000" when "0000111001011010", -- t[3674] = 0
      "000000" when "0000111001011011", -- t[3675] = 0
      "000000" when "0000111001011100", -- t[3676] = 0
      "000000" when "0000111001011101", -- t[3677] = 0
      "000000" when "0000111001011110", -- t[3678] = 0
      "000000" when "0000111001011111", -- t[3679] = 0
      "000000" when "0000111001100000", -- t[3680] = 0
      "000000" when "0000111001100001", -- t[3681] = 0
      "000000" when "0000111001100010", -- t[3682] = 0
      "000000" when "0000111001100011", -- t[3683] = 0
      "000000" when "0000111001100100", -- t[3684] = 0
      "000000" when "0000111001100101", -- t[3685] = 0
      "000000" when "0000111001100110", -- t[3686] = 0
      "000000" when "0000111001100111", -- t[3687] = 0
      "000000" when "0000111001101000", -- t[3688] = 0
      "000000" when "0000111001101001", -- t[3689] = 0
      "000000" when "0000111001101010", -- t[3690] = 0
      "000000" when "0000111001101011", -- t[3691] = 0
      "000000" when "0000111001101100", -- t[3692] = 0
      "000000" when "0000111001101101", -- t[3693] = 0
      "000000" when "0000111001101110", -- t[3694] = 0
      "000000" when "0000111001101111", -- t[3695] = 0
      "000000" when "0000111001110000", -- t[3696] = 0
      "000000" when "0000111001110001", -- t[3697] = 0
      "000000" when "0000111001110010", -- t[3698] = 0
      "000000" when "0000111001110011", -- t[3699] = 0
      "000000" when "0000111001110100", -- t[3700] = 0
      "000000" when "0000111001110101", -- t[3701] = 0
      "000000" when "0000111001110110", -- t[3702] = 0
      "000000" when "0000111001110111", -- t[3703] = 0
      "000000" when "0000111001111000", -- t[3704] = 0
      "000000" when "0000111001111001", -- t[3705] = 0
      "000000" when "0000111001111010", -- t[3706] = 0
      "000000" when "0000111001111011", -- t[3707] = 0
      "000000" when "0000111001111100", -- t[3708] = 0
      "000000" when "0000111001111101", -- t[3709] = 0
      "000000" when "0000111001111110", -- t[3710] = 0
      "000000" when "0000111001111111", -- t[3711] = 0
      "000000" when "0000111010000000", -- t[3712] = 0
      "000000" when "0000111010000001", -- t[3713] = 0
      "000000" when "0000111010000010", -- t[3714] = 0
      "000000" when "0000111010000011", -- t[3715] = 0
      "000000" when "0000111010000100", -- t[3716] = 0
      "000000" when "0000111010000101", -- t[3717] = 0
      "000000" when "0000111010000110", -- t[3718] = 0
      "000000" when "0000111010000111", -- t[3719] = 0
      "000000" when "0000111010001000", -- t[3720] = 0
      "000000" when "0000111010001001", -- t[3721] = 0
      "000000" when "0000111010001010", -- t[3722] = 0
      "000000" when "0000111010001011", -- t[3723] = 0
      "000000" when "0000111010001100", -- t[3724] = 0
      "000000" when "0000111010001101", -- t[3725] = 0
      "000000" when "0000111010001110", -- t[3726] = 0
      "000000" when "0000111010001111", -- t[3727] = 0
      "000000" when "0000111010010000", -- t[3728] = 0
      "000000" when "0000111010010001", -- t[3729] = 0
      "000000" when "0000111010010010", -- t[3730] = 0
      "000000" when "0000111010010011", -- t[3731] = 0
      "000000" when "0000111010010100", -- t[3732] = 0
      "000000" when "0000111010010101", -- t[3733] = 0
      "000000" when "0000111010010110", -- t[3734] = 0
      "000000" when "0000111010010111", -- t[3735] = 0
      "000000" when "0000111010011000", -- t[3736] = 0
      "000000" when "0000111010011001", -- t[3737] = 0
      "000000" when "0000111010011010", -- t[3738] = 0
      "000000" when "0000111010011011", -- t[3739] = 0
      "000000" when "0000111010011100", -- t[3740] = 0
      "000000" when "0000111010011101", -- t[3741] = 0
      "000000" when "0000111010011110", -- t[3742] = 0
      "000000" when "0000111010011111", -- t[3743] = 0
      "000000" when "0000111010100000", -- t[3744] = 0
      "000000" when "0000111010100001", -- t[3745] = 0
      "000000" when "0000111010100010", -- t[3746] = 0
      "000000" when "0000111010100011", -- t[3747] = 0
      "000000" when "0000111010100100", -- t[3748] = 0
      "000000" when "0000111010100101", -- t[3749] = 0
      "000000" when "0000111010100110", -- t[3750] = 0
      "000000" when "0000111010100111", -- t[3751] = 0
      "000000" when "0000111010101000", -- t[3752] = 0
      "000000" when "0000111010101001", -- t[3753] = 0
      "000000" when "0000111010101010", -- t[3754] = 0
      "000000" when "0000111010101011", -- t[3755] = 0
      "000000" when "0000111010101100", -- t[3756] = 0
      "000000" when "0000111010101101", -- t[3757] = 0
      "000000" when "0000111010101110", -- t[3758] = 0
      "000000" when "0000111010101111", -- t[3759] = 0
      "000000" when "0000111010110000", -- t[3760] = 0
      "000000" when "0000111010110001", -- t[3761] = 0
      "000000" when "0000111010110010", -- t[3762] = 0
      "000000" when "0000111010110011", -- t[3763] = 0
      "000000" when "0000111010110100", -- t[3764] = 0
      "000000" when "0000111010110101", -- t[3765] = 0
      "000000" when "0000111010110110", -- t[3766] = 0
      "000000" when "0000111010110111", -- t[3767] = 0
      "000000" when "0000111010111000", -- t[3768] = 0
      "000000" when "0000111010111001", -- t[3769] = 0
      "000000" when "0000111010111010", -- t[3770] = 0
      "000000" when "0000111010111011", -- t[3771] = 0
      "000000" when "0000111010111100", -- t[3772] = 0
      "000000" when "0000111010111101", -- t[3773] = 0
      "000000" when "0000111010111110", -- t[3774] = 0
      "000000" when "0000111010111111", -- t[3775] = 0
      "000000" when "0000111011000000", -- t[3776] = 0
      "000000" when "0000111011000001", -- t[3777] = 0
      "000000" when "0000111011000010", -- t[3778] = 0
      "000000" when "0000111011000011", -- t[3779] = 0
      "000000" when "0000111011000100", -- t[3780] = 0
      "000000" when "0000111011000101", -- t[3781] = 0
      "000000" when "0000111011000110", -- t[3782] = 0
      "000000" when "0000111011000111", -- t[3783] = 0
      "000000" when "0000111011001000", -- t[3784] = 0
      "000000" when "0000111011001001", -- t[3785] = 0
      "000000" when "0000111011001010", -- t[3786] = 0
      "000000" when "0000111011001011", -- t[3787] = 0
      "000000" when "0000111011001100", -- t[3788] = 0
      "000000" when "0000111011001101", -- t[3789] = 0
      "000000" when "0000111011001110", -- t[3790] = 0
      "000000" when "0000111011001111", -- t[3791] = 0
      "000000" when "0000111011010000", -- t[3792] = 0
      "000000" when "0000111011010001", -- t[3793] = 0
      "000000" when "0000111011010010", -- t[3794] = 0
      "000000" when "0000111011010011", -- t[3795] = 0
      "000000" when "0000111011010100", -- t[3796] = 0
      "000000" when "0000111011010101", -- t[3797] = 0
      "000000" when "0000111011010110", -- t[3798] = 0
      "000000" when "0000111011010111", -- t[3799] = 0
      "000000" when "0000111011011000", -- t[3800] = 0
      "000000" when "0000111011011001", -- t[3801] = 0
      "000000" when "0000111011011010", -- t[3802] = 0
      "000000" when "0000111011011011", -- t[3803] = 0
      "000000" when "0000111011011100", -- t[3804] = 0
      "000000" when "0000111011011101", -- t[3805] = 0
      "000000" when "0000111011011110", -- t[3806] = 0
      "000000" when "0000111011011111", -- t[3807] = 0
      "000000" when "0000111011100000", -- t[3808] = 0
      "000000" when "0000111011100001", -- t[3809] = 0
      "000000" when "0000111011100010", -- t[3810] = 0
      "000000" when "0000111011100011", -- t[3811] = 0
      "000000" when "0000111011100100", -- t[3812] = 0
      "000000" when "0000111011100101", -- t[3813] = 0
      "000000" when "0000111011100110", -- t[3814] = 0
      "000000" when "0000111011100111", -- t[3815] = 0
      "000000" when "0000111011101000", -- t[3816] = 0
      "000000" when "0000111011101001", -- t[3817] = 0
      "000000" when "0000111011101010", -- t[3818] = 0
      "000000" when "0000111011101011", -- t[3819] = 0
      "000000" when "0000111011101100", -- t[3820] = 0
      "000000" when "0000111011101101", -- t[3821] = 0
      "000000" when "0000111011101110", -- t[3822] = 0
      "000000" when "0000111011101111", -- t[3823] = 0
      "000000" when "0000111011110000", -- t[3824] = 0
      "000000" when "0000111011110001", -- t[3825] = 0
      "000000" when "0000111011110010", -- t[3826] = 0
      "000000" when "0000111011110011", -- t[3827] = 0
      "000000" when "0000111011110100", -- t[3828] = 0
      "000000" when "0000111011110101", -- t[3829] = 0
      "000000" when "0000111011110110", -- t[3830] = 0
      "000000" when "0000111011110111", -- t[3831] = 0
      "000000" when "0000111011111000", -- t[3832] = 0
      "000000" when "0000111011111001", -- t[3833] = 0
      "000000" when "0000111011111010", -- t[3834] = 0
      "000000" when "0000111011111011", -- t[3835] = 0
      "000000" when "0000111011111100", -- t[3836] = 0
      "000000" when "0000111011111101", -- t[3837] = 0
      "000000" when "0000111011111110", -- t[3838] = 0
      "000000" when "0000111011111111", -- t[3839] = 0
      "000000" when "0000111100000000", -- t[3840] = 0
      "000000" when "0000111100000001", -- t[3841] = 0
      "000000" when "0000111100000010", -- t[3842] = 0
      "000000" when "0000111100000011", -- t[3843] = 0
      "000000" when "0000111100000100", -- t[3844] = 0
      "000000" when "0000111100000101", -- t[3845] = 0
      "000000" when "0000111100000110", -- t[3846] = 0
      "000000" when "0000111100000111", -- t[3847] = 0
      "000000" when "0000111100001000", -- t[3848] = 0
      "000000" when "0000111100001001", -- t[3849] = 0
      "000000" when "0000111100001010", -- t[3850] = 0
      "000000" when "0000111100001011", -- t[3851] = 0
      "000000" when "0000111100001100", -- t[3852] = 0
      "000000" when "0000111100001101", -- t[3853] = 0
      "000000" when "0000111100001110", -- t[3854] = 0
      "000000" when "0000111100001111", -- t[3855] = 0
      "000000" when "0000111100010000", -- t[3856] = 0
      "000000" when "0000111100010001", -- t[3857] = 0
      "000000" when "0000111100010010", -- t[3858] = 0
      "000000" when "0000111100010011", -- t[3859] = 0
      "000000" when "0000111100010100", -- t[3860] = 0
      "000000" when "0000111100010101", -- t[3861] = 0
      "000000" when "0000111100010110", -- t[3862] = 0
      "000000" when "0000111100010111", -- t[3863] = 0
      "000000" when "0000111100011000", -- t[3864] = 0
      "000000" when "0000111100011001", -- t[3865] = 0
      "000000" when "0000111100011010", -- t[3866] = 0
      "000000" when "0000111100011011", -- t[3867] = 0
      "000000" when "0000111100011100", -- t[3868] = 0
      "000000" when "0000111100011101", -- t[3869] = 0
      "000000" when "0000111100011110", -- t[3870] = 0
      "000000" when "0000111100011111", -- t[3871] = 0
      "000000" when "0000111100100000", -- t[3872] = 0
      "000000" when "0000111100100001", -- t[3873] = 0
      "000000" when "0000111100100010", -- t[3874] = 0
      "000000" when "0000111100100011", -- t[3875] = 0
      "000000" when "0000111100100100", -- t[3876] = 0
      "000000" when "0000111100100101", -- t[3877] = 0
      "000000" when "0000111100100110", -- t[3878] = 0
      "000000" when "0000111100100111", -- t[3879] = 0
      "000000" when "0000111100101000", -- t[3880] = 0
      "000000" when "0000111100101001", -- t[3881] = 0
      "000000" when "0000111100101010", -- t[3882] = 0
      "000000" when "0000111100101011", -- t[3883] = 0
      "000000" when "0000111100101100", -- t[3884] = 0
      "000000" when "0000111100101101", -- t[3885] = 0
      "000000" when "0000111100101110", -- t[3886] = 0
      "000000" when "0000111100101111", -- t[3887] = 0
      "000000" when "0000111100110000", -- t[3888] = 0
      "000000" when "0000111100110001", -- t[3889] = 0
      "000000" when "0000111100110010", -- t[3890] = 0
      "000000" when "0000111100110011", -- t[3891] = 0
      "000000" when "0000111100110100", -- t[3892] = 0
      "000000" when "0000111100110101", -- t[3893] = 0
      "000000" when "0000111100110110", -- t[3894] = 0
      "000000" when "0000111100110111", -- t[3895] = 0
      "000000" when "0000111100111000", -- t[3896] = 0
      "000000" when "0000111100111001", -- t[3897] = 0
      "000000" when "0000111100111010", -- t[3898] = 0
      "000000" when "0000111100111011", -- t[3899] = 0
      "000000" when "0000111100111100", -- t[3900] = 0
      "000000" when "0000111100111101", -- t[3901] = 0
      "000000" when "0000111100111110", -- t[3902] = 0
      "000000" when "0000111100111111", -- t[3903] = 0
      "000000" when "0000111101000000", -- t[3904] = 0
      "000000" when "0000111101000001", -- t[3905] = 0
      "000000" when "0000111101000010", -- t[3906] = 0
      "000000" when "0000111101000011", -- t[3907] = 0
      "000000" when "0000111101000100", -- t[3908] = 0
      "000000" when "0000111101000101", -- t[3909] = 0
      "000000" when "0000111101000110", -- t[3910] = 0
      "000000" when "0000111101000111", -- t[3911] = 0
      "000000" when "0000111101001000", -- t[3912] = 0
      "000000" when "0000111101001001", -- t[3913] = 0
      "000000" when "0000111101001010", -- t[3914] = 0
      "000000" when "0000111101001011", -- t[3915] = 0
      "000000" when "0000111101001100", -- t[3916] = 0
      "000000" when "0000111101001101", -- t[3917] = 0
      "000000" when "0000111101001110", -- t[3918] = 0
      "000000" when "0000111101001111", -- t[3919] = 0
      "000000" when "0000111101010000", -- t[3920] = 0
      "000000" when "0000111101010001", -- t[3921] = 0
      "000000" when "0000111101010010", -- t[3922] = 0
      "000000" when "0000111101010011", -- t[3923] = 0
      "000000" when "0000111101010100", -- t[3924] = 0
      "000000" when "0000111101010101", -- t[3925] = 0
      "000000" when "0000111101010110", -- t[3926] = 0
      "000000" when "0000111101010111", -- t[3927] = 0
      "000000" when "0000111101011000", -- t[3928] = 0
      "000000" when "0000111101011001", -- t[3929] = 0
      "000000" when "0000111101011010", -- t[3930] = 0
      "000000" when "0000111101011011", -- t[3931] = 0
      "000000" when "0000111101011100", -- t[3932] = 0
      "000000" when "0000111101011101", -- t[3933] = 0
      "000000" when "0000111101011110", -- t[3934] = 0
      "000000" when "0000111101011111", -- t[3935] = 0
      "000000" when "0000111101100000", -- t[3936] = 0
      "000000" when "0000111101100001", -- t[3937] = 0
      "000000" when "0000111101100010", -- t[3938] = 0
      "000000" when "0000111101100011", -- t[3939] = 0
      "000000" when "0000111101100100", -- t[3940] = 0
      "000000" when "0000111101100101", -- t[3941] = 0
      "000000" when "0000111101100110", -- t[3942] = 0
      "000000" when "0000111101100111", -- t[3943] = 0
      "000000" when "0000111101101000", -- t[3944] = 0
      "000000" when "0000111101101001", -- t[3945] = 0
      "000000" when "0000111101101010", -- t[3946] = 0
      "000000" when "0000111101101011", -- t[3947] = 0
      "000000" when "0000111101101100", -- t[3948] = 0
      "000000" when "0000111101101101", -- t[3949] = 0
      "000000" when "0000111101101110", -- t[3950] = 0
      "000000" when "0000111101101111", -- t[3951] = 0
      "000000" when "0000111101110000", -- t[3952] = 0
      "000000" when "0000111101110001", -- t[3953] = 0
      "000000" when "0000111101110010", -- t[3954] = 0
      "000000" when "0000111101110011", -- t[3955] = 0
      "000000" when "0000111101110100", -- t[3956] = 0
      "000000" when "0000111101110101", -- t[3957] = 0
      "000000" when "0000111101110110", -- t[3958] = 0
      "000000" when "0000111101110111", -- t[3959] = 0
      "000000" when "0000111101111000", -- t[3960] = 0
      "000000" when "0000111101111001", -- t[3961] = 0
      "000000" when "0000111101111010", -- t[3962] = 0
      "000000" when "0000111101111011", -- t[3963] = 0
      "000000" when "0000111101111100", -- t[3964] = 0
      "000000" when "0000111101111101", -- t[3965] = 0
      "000000" when "0000111101111110", -- t[3966] = 0
      "000000" when "0000111101111111", -- t[3967] = 0
      "000000" when "0000111110000000", -- t[3968] = 0
      "000000" when "0000111110000001", -- t[3969] = 0
      "000000" when "0000111110000010", -- t[3970] = 0
      "000000" when "0000111110000011", -- t[3971] = 0
      "000000" when "0000111110000100", -- t[3972] = 0
      "000000" when "0000111110000101", -- t[3973] = 0
      "000000" when "0000111110000110", -- t[3974] = 0
      "000000" when "0000111110000111", -- t[3975] = 0
      "000000" when "0000111110001000", -- t[3976] = 0
      "000000" when "0000111110001001", -- t[3977] = 0
      "000000" when "0000111110001010", -- t[3978] = 0
      "000000" when "0000111110001011", -- t[3979] = 0
      "000000" when "0000111110001100", -- t[3980] = 0
      "000000" when "0000111110001101", -- t[3981] = 0
      "000000" when "0000111110001110", -- t[3982] = 0
      "000000" when "0000111110001111", -- t[3983] = 0
      "000000" when "0000111110010000", -- t[3984] = 0
      "000000" when "0000111110010001", -- t[3985] = 0
      "000000" when "0000111110010010", -- t[3986] = 0
      "000000" when "0000111110010011", -- t[3987] = 0
      "000000" when "0000111110010100", -- t[3988] = 0
      "000000" when "0000111110010101", -- t[3989] = 0
      "000000" when "0000111110010110", -- t[3990] = 0
      "000000" when "0000111110010111", -- t[3991] = 0
      "000000" when "0000111110011000", -- t[3992] = 0
      "000000" when "0000111110011001", -- t[3993] = 0
      "000000" when "0000111110011010", -- t[3994] = 0
      "000000" when "0000111110011011", -- t[3995] = 0
      "000000" when "0000111110011100", -- t[3996] = 0
      "000000" when "0000111110011101", -- t[3997] = 0
      "000000" when "0000111110011110", -- t[3998] = 0
      "000000" when "0000111110011111", -- t[3999] = 0
      "000000" when "0000111110100000", -- t[4000] = 0
      "000000" when "0000111110100001", -- t[4001] = 0
      "000000" when "0000111110100010", -- t[4002] = 0
      "000000" when "0000111110100011", -- t[4003] = 0
      "000000" when "0000111110100100", -- t[4004] = 0
      "000000" when "0000111110100101", -- t[4005] = 0
      "000000" when "0000111110100110", -- t[4006] = 0
      "000000" when "0000111110100111", -- t[4007] = 0
      "000000" when "0000111110101000", -- t[4008] = 0
      "000000" when "0000111110101001", -- t[4009] = 0
      "000000" when "0000111110101010", -- t[4010] = 0
      "000000" when "0000111110101011", -- t[4011] = 0
      "000000" when "0000111110101100", -- t[4012] = 0
      "000000" when "0000111110101101", -- t[4013] = 0
      "000000" when "0000111110101110", -- t[4014] = 0
      "000000" when "0000111110101111", -- t[4015] = 0
      "000000" when "0000111110110000", -- t[4016] = 0
      "000000" when "0000111110110001", -- t[4017] = 0
      "000000" when "0000111110110010", -- t[4018] = 0
      "000000" when "0000111110110011", -- t[4019] = 0
      "000000" when "0000111110110100", -- t[4020] = 0
      "000000" when "0000111110110101", -- t[4021] = 0
      "000000" when "0000111110110110", -- t[4022] = 0
      "000000" when "0000111110110111", -- t[4023] = 0
      "000000" when "0000111110111000", -- t[4024] = 0
      "000000" when "0000111110111001", -- t[4025] = 0
      "000000" when "0000111110111010", -- t[4026] = 0
      "000000" when "0000111110111011", -- t[4027] = 0
      "000000" when "0000111110111100", -- t[4028] = 0
      "000000" when "0000111110111101", -- t[4029] = 0
      "000000" when "0000111110111110", -- t[4030] = 0
      "000000" when "0000111110111111", -- t[4031] = 0
      "000000" when "0000111111000000", -- t[4032] = 0
      "000000" when "0000111111000001", -- t[4033] = 0
      "000000" when "0000111111000010", -- t[4034] = 0
      "000000" when "0000111111000011", -- t[4035] = 0
      "000000" when "0000111111000100", -- t[4036] = 0
      "000000" when "0000111111000101", -- t[4037] = 0
      "000000" when "0000111111000110", -- t[4038] = 0
      "000000" when "0000111111000111", -- t[4039] = 0
      "000000" when "0000111111001000", -- t[4040] = 0
      "000000" when "0000111111001001", -- t[4041] = 0
      "000000" when "0000111111001010", -- t[4042] = 0
      "000000" when "0000111111001011", -- t[4043] = 0
      "000000" when "0000111111001100", -- t[4044] = 0
      "000000" when "0000111111001101", -- t[4045] = 0
      "000000" when "0000111111001110", -- t[4046] = 0
      "000000" when "0000111111001111", -- t[4047] = 0
      "000000" when "0000111111010000", -- t[4048] = 0
      "000000" when "0000111111010001", -- t[4049] = 0
      "000000" when "0000111111010010", -- t[4050] = 0
      "000000" when "0000111111010011", -- t[4051] = 0
      "000000" when "0000111111010100", -- t[4052] = 0
      "000000" when "0000111111010101", -- t[4053] = 0
      "000000" when "0000111111010110", -- t[4054] = 0
      "000000" when "0000111111010111", -- t[4055] = 0
      "000000" when "0000111111011000", -- t[4056] = 0
      "000000" when "0000111111011001", -- t[4057] = 0
      "000000" when "0000111111011010", -- t[4058] = 0
      "000000" when "0000111111011011", -- t[4059] = 0
      "000000" when "0000111111011100", -- t[4060] = 0
      "000000" when "0000111111011101", -- t[4061] = 0
      "000000" when "0000111111011110", -- t[4062] = 0
      "000000" when "0000111111011111", -- t[4063] = 0
      "000000" when "0000111111100000", -- t[4064] = 0
      "000000" when "0000111111100001", -- t[4065] = 0
      "000000" when "0000111111100010", -- t[4066] = 0
      "000000" when "0000111111100011", -- t[4067] = 0
      "000000" when "0000111111100100", -- t[4068] = 0
      "000000" when "0000111111100101", -- t[4069] = 0
      "000000" when "0000111111100110", -- t[4070] = 0
      "000000" when "0000111111100111", -- t[4071] = 0
      "000000" when "0000111111101000", -- t[4072] = 0
      "000000" when "0000111111101001", -- t[4073] = 0
      "000000" when "0000111111101010", -- t[4074] = 0
      "000000" when "0000111111101011", -- t[4075] = 0
      "000000" when "0000111111101100", -- t[4076] = 0
      "000000" when "0000111111101101", -- t[4077] = 0
      "000000" when "0000111111101110", -- t[4078] = 0
      "000000" when "0000111111101111", -- t[4079] = 0
      "000000" when "0000111111110000", -- t[4080] = 0
      "000000" when "0000111111110001", -- t[4081] = 0
      "000000" when "0000111111110010", -- t[4082] = 0
      "000000" when "0000111111110011", -- t[4083] = 0
      "000000" when "0000111111110100", -- t[4084] = 0
      "000000" when "0000111111110101", -- t[4085] = 0
      "000000" when "0000111111110110", -- t[4086] = 0
      "000000" when "0000111111110111", -- t[4087] = 0
      "000000" when "0000111111111000", -- t[4088] = 0
      "000000" when "0000111111111001", -- t[4089] = 0
      "000000" when "0000111111111010", -- t[4090] = 0
      "000000" when "0000111111111011", -- t[4091] = 0
      "000000" when "0000111111111100", -- t[4092] = 0
      "000000" when "0000111111111101", -- t[4093] = 0
      "000000" when "0000111111111110", -- t[4094] = 0
      "000000" when "0000111111111111", -- t[4095] = 0
      "000000" when "0001000000000000", -- t[4096] = 0
      "000000" when "0001000000000001", -- t[4097] = 0
      "000000" when "0001000000000010", -- t[4098] = 0
      "000000" when "0001000000000011", -- t[4099] = 0
      "000000" when "0001000000000100", -- t[4100] = 0
      "000000" when "0001000000000101", -- t[4101] = 0
      "000000" when "0001000000000110", -- t[4102] = 0
      "000000" when "0001000000000111", -- t[4103] = 0
      "000000" when "0001000000001000", -- t[4104] = 0
      "000000" when "0001000000001001", -- t[4105] = 0
      "000000" when "0001000000001010", -- t[4106] = 0
      "000000" when "0001000000001011", -- t[4107] = 0
      "000000" when "0001000000001100", -- t[4108] = 0
      "000000" when "0001000000001101", -- t[4109] = 0
      "000000" when "0001000000001110", -- t[4110] = 0
      "000000" when "0001000000001111", -- t[4111] = 0
      "000000" when "0001000000010000", -- t[4112] = 0
      "000000" when "0001000000010001", -- t[4113] = 0
      "000000" when "0001000000010010", -- t[4114] = 0
      "000000" when "0001000000010011", -- t[4115] = 0
      "000000" when "0001000000010100", -- t[4116] = 0
      "000000" when "0001000000010101", -- t[4117] = 0
      "000000" when "0001000000010110", -- t[4118] = 0
      "000000" when "0001000000010111", -- t[4119] = 0
      "000000" when "0001000000011000", -- t[4120] = 0
      "000000" when "0001000000011001", -- t[4121] = 0
      "000000" when "0001000000011010", -- t[4122] = 0
      "000000" when "0001000000011011", -- t[4123] = 0
      "000000" when "0001000000011100", -- t[4124] = 0
      "000000" when "0001000000011101", -- t[4125] = 0
      "000000" when "0001000000011110", -- t[4126] = 0
      "000000" when "0001000000011111", -- t[4127] = 0
      "000000" when "0001000000100000", -- t[4128] = 0
      "000000" when "0001000000100001", -- t[4129] = 0
      "000000" when "0001000000100010", -- t[4130] = 0
      "000000" when "0001000000100011", -- t[4131] = 0
      "000000" when "0001000000100100", -- t[4132] = 0
      "000000" when "0001000000100101", -- t[4133] = 0
      "000000" when "0001000000100110", -- t[4134] = 0
      "000000" when "0001000000100111", -- t[4135] = 0
      "000000" when "0001000000101000", -- t[4136] = 0
      "000000" when "0001000000101001", -- t[4137] = 0
      "000000" when "0001000000101010", -- t[4138] = 0
      "000000" when "0001000000101011", -- t[4139] = 0
      "000000" when "0001000000101100", -- t[4140] = 0
      "000000" when "0001000000101101", -- t[4141] = 0
      "000000" when "0001000000101110", -- t[4142] = 0
      "000000" when "0001000000101111", -- t[4143] = 0
      "000000" when "0001000000110000", -- t[4144] = 0
      "000000" when "0001000000110001", -- t[4145] = 0
      "000000" when "0001000000110010", -- t[4146] = 0
      "000000" when "0001000000110011", -- t[4147] = 0
      "000000" when "0001000000110100", -- t[4148] = 0
      "000000" when "0001000000110101", -- t[4149] = 0
      "000000" when "0001000000110110", -- t[4150] = 0
      "000000" when "0001000000110111", -- t[4151] = 0
      "000000" when "0001000000111000", -- t[4152] = 0
      "000000" when "0001000000111001", -- t[4153] = 0
      "000000" when "0001000000111010", -- t[4154] = 0
      "000000" when "0001000000111011", -- t[4155] = 0
      "000000" when "0001000000111100", -- t[4156] = 0
      "000000" when "0001000000111101", -- t[4157] = 0
      "000000" when "0001000000111110", -- t[4158] = 0
      "000000" when "0001000000111111", -- t[4159] = 0
      "000000" when "0001000001000000", -- t[4160] = 0
      "000000" when "0001000001000001", -- t[4161] = 0
      "000000" when "0001000001000010", -- t[4162] = 0
      "000000" when "0001000001000011", -- t[4163] = 0
      "000000" when "0001000001000100", -- t[4164] = 0
      "000000" when "0001000001000101", -- t[4165] = 0
      "000000" when "0001000001000110", -- t[4166] = 0
      "000000" when "0001000001000111", -- t[4167] = 0
      "000000" when "0001000001001000", -- t[4168] = 0
      "000000" when "0001000001001001", -- t[4169] = 0
      "000000" when "0001000001001010", -- t[4170] = 0
      "000000" when "0001000001001011", -- t[4171] = 0
      "000000" when "0001000001001100", -- t[4172] = 0
      "000000" when "0001000001001101", -- t[4173] = 0
      "000000" when "0001000001001110", -- t[4174] = 0
      "000000" when "0001000001001111", -- t[4175] = 0
      "000000" when "0001000001010000", -- t[4176] = 0
      "000000" when "0001000001010001", -- t[4177] = 0
      "000000" when "0001000001010010", -- t[4178] = 0
      "000000" when "0001000001010011", -- t[4179] = 0
      "000000" when "0001000001010100", -- t[4180] = 0
      "000000" when "0001000001010101", -- t[4181] = 0
      "000000" when "0001000001010110", -- t[4182] = 0
      "000000" when "0001000001010111", -- t[4183] = 0
      "000000" when "0001000001011000", -- t[4184] = 0
      "000000" when "0001000001011001", -- t[4185] = 0
      "000000" when "0001000001011010", -- t[4186] = 0
      "000000" when "0001000001011011", -- t[4187] = 0
      "000000" when "0001000001011100", -- t[4188] = 0
      "000000" when "0001000001011101", -- t[4189] = 0
      "000000" when "0001000001011110", -- t[4190] = 0
      "000000" when "0001000001011111", -- t[4191] = 0
      "000000" when "0001000001100000", -- t[4192] = 0
      "000000" when "0001000001100001", -- t[4193] = 0
      "000000" when "0001000001100010", -- t[4194] = 0
      "000000" when "0001000001100011", -- t[4195] = 0
      "000000" when "0001000001100100", -- t[4196] = 0
      "000000" when "0001000001100101", -- t[4197] = 0
      "000000" when "0001000001100110", -- t[4198] = 0
      "000000" when "0001000001100111", -- t[4199] = 0
      "000000" when "0001000001101000", -- t[4200] = 0
      "000000" when "0001000001101001", -- t[4201] = 0
      "000000" when "0001000001101010", -- t[4202] = 0
      "000000" when "0001000001101011", -- t[4203] = 0
      "000000" when "0001000001101100", -- t[4204] = 0
      "000000" when "0001000001101101", -- t[4205] = 0
      "000000" when "0001000001101110", -- t[4206] = 0
      "000000" when "0001000001101111", -- t[4207] = 0
      "000000" when "0001000001110000", -- t[4208] = 0
      "000000" when "0001000001110001", -- t[4209] = 0
      "000000" when "0001000001110010", -- t[4210] = 0
      "000000" when "0001000001110011", -- t[4211] = 0
      "000000" when "0001000001110100", -- t[4212] = 0
      "000000" when "0001000001110101", -- t[4213] = 0
      "000000" when "0001000001110110", -- t[4214] = 0
      "000000" when "0001000001110111", -- t[4215] = 0
      "000000" when "0001000001111000", -- t[4216] = 0
      "000000" when "0001000001111001", -- t[4217] = 0
      "000000" when "0001000001111010", -- t[4218] = 0
      "000000" when "0001000001111011", -- t[4219] = 0
      "000000" when "0001000001111100", -- t[4220] = 0
      "000000" when "0001000001111101", -- t[4221] = 0
      "000000" when "0001000001111110", -- t[4222] = 0
      "000000" when "0001000001111111", -- t[4223] = 0
      "000000" when "0001000010000000", -- t[4224] = 0
      "000000" when "0001000010000001", -- t[4225] = 0
      "000000" when "0001000010000010", -- t[4226] = 0
      "000000" when "0001000010000011", -- t[4227] = 0
      "000000" when "0001000010000100", -- t[4228] = 0
      "000000" when "0001000010000101", -- t[4229] = 0
      "000000" when "0001000010000110", -- t[4230] = 0
      "000000" when "0001000010000111", -- t[4231] = 0
      "000000" when "0001000010001000", -- t[4232] = 0
      "000000" when "0001000010001001", -- t[4233] = 0
      "000000" when "0001000010001010", -- t[4234] = 0
      "000000" when "0001000010001011", -- t[4235] = 0
      "000000" when "0001000010001100", -- t[4236] = 0
      "000000" when "0001000010001101", -- t[4237] = 0
      "000000" when "0001000010001110", -- t[4238] = 0
      "000000" when "0001000010001111", -- t[4239] = 0
      "000000" when "0001000010010000", -- t[4240] = 0
      "000000" when "0001000010010001", -- t[4241] = 0
      "000000" when "0001000010010010", -- t[4242] = 0
      "000000" when "0001000010010011", -- t[4243] = 0
      "000000" when "0001000010010100", -- t[4244] = 0
      "000000" when "0001000010010101", -- t[4245] = 0
      "000000" when "0001000010010110", -- t[4246] = 0
      "000000" when "0001000010010111", -- t[4247] = 0
      "000000" when "0001000010011000", -- t[4248] = 0
      "000000" when "0001000010011001", -- t[4249] = 0
      "000000" when "0001000010011010", -- t[4250] = 0
      "000000" when "0001000010011011", -- t[4251] = 0
      "000000" when "0001000010011100", -- t[4252] = 0
      "000000" when "0001000010011101", -- t[4253] = 0
      "000000" when "0001000010011110", -- t[4254] = 0
      "000000" when "0001000010011111", -- t[4255] = 0
      "000000" when "0001000010100000", -- t[4256] = 0
      "000000" when "0001000010100001", -- t[4257] = 0
      "000000" when "0001000010100010", -- t[4258] = 0
      "000000" when "0001000010100011", -- t[4259] = 0
      "000000" when "0001000010100100", -- t[4260] = 0
      "000000" when "0001000010100101", -- t[4261] = 0
      "000000" when "0001000010100110", -- t[4262] = 0
      "000000" when "0001000010100111", -- t[4263] = 0
      "000000" when "0001000010101000", -- t[4264] = 0
      "000000" when "0001000010101001", -- t[4265] = 0
      "000000" when "0001000010101010", -- t[4266] = 0
      "000000" when "0001000010101011", -- t[4267] = 0
      "000000" when "0001000010101100", -- t[4268] = 0
      "000000" when "0001000010101101", -- t[4269] = 0
      "000000" when "0001000010101110", -- t[4270] = 0
      "000000" when "0001000010101111", -- t[4271] = 0
      "000000" when "0001000010110000", -- t[4272] = 0
      "000000" when "0001000010110001", -- t[4273] = 0
      "000000" when "0001000010110010", -- t[4274] = 0
      "000000" when "0001000010110011", -- t[4275] = 0
      "000000" when "0001000010110100", -- t[4276] = 0
      "000000" when "0001000010110101", -- t[4277] = 0
      "000000" when "0001000010110110", -- t[4278] = 0
      "000000" when "0001000010110111", -- t[4279] = 0
      "000000" when "0001000010111000", -- t[4280] = 0
      "000000" when "0001000010111001", -- t[4281] = 0
      "000000" when "0001000010111010", -- t[4282] = 0
      "000000" when "0001000010111011", -- t[4283] = 0
      "000000" when "0001000010111100", -- t[4284] = 0
      "000000" when "0001000010111101", -- t[4285] = 0
      "000000" when "0001000010111110", -- t[4286] = 0
      "000000" when "0001000010111111", -- t[4287] = 0
      "000000" when "0001000011000000", -- t[4288] = 0
      "000000" when "0001000011000001", -- t[4289] = 0
      "000000" when "0001000011000010", -- t[4290] = 0
      "000000" when "0001000011000011", -- t[4291] = 0
      "000000" when "0001000011000100", -- t[4292] = 0
      "000000" when "0001000011000101", -- t[4293] = 0
      "000000" when "0001000011000110", -- t[4294] = 0
      "000000" when "0001000011000111", -- t[4295] = 0
      "000000" when "0001000011001000", -- t[4296] = 0
      "000000" when "0001000011001001", -- t[4297] = 0
      "000000" when "0001000011001010", -- t[4298] = 0
      "000000" when "0001000011001011", -- t[4299] = 0
      "000000" when "0001000011001100", -- t[4300] = 0
      "000000" when "0001000011001101", -- t[4301] = 0
      "000000" when "0001000011001110", -- t[4302] = 0
      "000000" when "0001000011001111", -- t[4303] = 0
      "000000" when "0001000011010000", -- t[4304] = 0
      "000000" when "0001000011010001", -- t[4305] = 0
      "000000" when "0001000011010010", -- t[4306] = 0
      "000000" when "0001000011010011", -- t[4307] = 0
      "000000" when "0001000011010100", -- t[4308] = 0
      "000000" when "0001000011010101", -- t[4309] = 0
      "000000" when "0001000011010110", -- t[4310] = 0
      "000000" when "0001000011010111", -- t[4311] = 0
      "000000" when "0001000011011000", -- t[4312] = 0
      "000000" when "0001000011011001", -- t[4313] = 0
      "000000" when "0001000011011010", -- t[4314] = 0
      "000000" when "0001000011011011", -- t[4315] = 0
      "000000" when "0001000011011100", -- t[4316] = 0
      "000000" when "0001000011011101", -- t[4317] = 0
      "000000" when "0001000011011110", -- t[4318] = 0
      "000000" when "0001000011011111", -- t[4319] = 0
      "000000" when "0001000011100000", -- t[4320] = 0
      "000000" when "0001000011100001", -- t[4321] = 0
      "000000" when "0001000011100010", -- t[4322] = 0
      "000000" when "0001000011100011", -- t[4323] = 0
      "000000" when "0001000011100100", -- t[4324] = 0
      "000000" when "0001000011100101", -- t[4325] = 0
      "000000" when "0001000011100110", -- t[4326] = 0
      "000000" when "0001000011100111", -- t[4327] = 0
      "000000" when "0001000011101000", -- t[4328] = 0
      "000000" when "0001000011101001", -- t[4329] = 0
      "000000" when "0001000011101010", -- t[4330] = 0
      "000000" when "0001000011101011", -- t[4331] = 0
      "000000" when "0001000011101100", -- t[4332] = 0
      "000000" when "0001000011101101", -- t[4333] = 0
      "000000" when "0001000011101110", -- t[4334] = 0
      "000000" when "0001000011101111", -- t[4335] = 0
      "000000" when "0001000011110000", -- t[4336] = 0
      "000000" when "0001000011110001", -- t[4337] = 0
      "000000" when "0001000011110010", -- t[4338] = 0
      "000000" when "0001000011110011", -- t[4339] = 0
      "000000" when "0001000011110100", -- t[4340] = 0
      "000000" when "0001000011110101", -- t[4341] = 0
      "000000" when "0001000011110110", -- t[4342] = 0
      "000000" when "0001000011110111", -- t[4343] = 0
      "000000" when "0001000011111000", -- t[4344] = 0
      "000000" when "0001000011111001", -- t[4345] = 0
      "000000" when "0001000011111010", -- t[4346] = 0
      "000000" when "0001000011111011", -- t[4347] = 0
      "000000" when "0001000011111100", -- t[4348] = 0
      "000000" when "0001000011111101", -- t[4349] = 0
      "000000" when "0001000011111110", -- t[4350] = 0
      "000000" when "0001000011111111", -- t[4351] = 0
      "000000" when "0001000100000000", -- t[4352] = 0
      "000000" when "0001000100000001", -- t[4353] = 0
      "000000" when "0001000100000010", -- t[4354] = 0
      "000000" when "0001000100000011", -- t[4355] = 0
      "000000" when "0001000100000100", -- t[4356] = 0
      "000000" when "0001000100000101", -- t[4357] = 0
      "000000" when "0001000100000110", -- t[4358] = 0
      "000000" when "0001000100000111", -- t[4359] = 0
      "000000" when "0001000100001000", -- t[4360] = 0
      "000000" when "0001000100001001", -- t[4361] = 0
      "000000" when "0001000100001010", -- t[4362] = 0
      "000000" when "0001000100001011", -- t[4363] = 0
      "000000" when "0001000100001100", -- t[4364] = 0
      "000000" when "0001000100001101", -- t[4365] = 0
      "000000" when "0001000100001110", -- t[4366] = 0
      "000000" when "0001000100001111", -- t[4367] = 0
      "000000" when "0001000100010000", -- t[4368] = 0
      "000000" when "0001000100010001", -- t[4369] = 0
      "000000" when "0001000100010010", -- t[4370] = 0
      "000000" when "0001000100010011", -- t[4371] = 0
      "000000" when "0001000100010100", -- t[4372] = 0
      "000000" when "0001000100010101", -- t[4373] = 0
      "000000" when "0001000100010110", -- t[4374] = 0
      "000000" when "0001000100010111", -- t[4375] = 0
      "000000" when "0001000100011000", -- t[4376] = 0
      "000000" when "0001000100011001", -- t[4377] = 0
      "000000" when "0001000100011010", -- t[4378] = 0
      "000000" when "0001000100011011", -- t[4379] = 0
      "000000" when "0001000100011100", -- t[4380] = 0
      "000000" when "0001000100011101", -- t[4381] = 0
      "000000" when "0001000100011110", -- t[4382] = 0
      "000000" when "0001000100011111", -- t[4383] = 0
      "000000" when "0001000100100000", -- t[4384] = 0
      "000000" when "0001000100100001", -- t[4385] = 0
      "000000" when "0001000100100010", -- t[4386] = 0
      "000000" when "0001000100100011", -- t[4387] = 0
      "000000" when "0001000100100100", -- t[4388] = 0
      "000000" when "0001000100100101", -- t[4389] = 0
      "000000" when "0001000100100110", -- t[4390] = 0
      "000000" when "0001000100100111", -- t[4391] = 0
      "000000" when "0001000100101000", -- t[4392] = 0
      "000000" when "0001000100101001", -- t[4393] = 0
      "000000" when "0001000100101010", -- t[4394] = 0
      "000000" when "0001000100101011", -- t[4395] = 0
      "000000" when "0001000100101100", -- t[4396] = 0
      "000000" when "0001000100101101", -- t[4397] = 0
      "000000" when "0001000100101110", -- t[4398] = 0
      "000000" when "0001000100101111", -- t[4399] = 0
      "000000" when "0001000100110000", -- t[4400] = 0
      "000000" when "0001000100110001", -- t[4401] = 0
      "000000" when "0001000100110010", -- t[4402] = 0
      "000000" when "0001000100110011", -- t[4403] = 0
      "000000" when "0001000100110100", -- t[4404] = 0
      "000000" when "0001000100110101", -- t[4405] = 0
      "000000" when "0001000100110110", -- t[4406] = 0
      "000000" when "0001000100110111", -- t[4407] = 0
      "000000" when "0001000100111000", -- t[4408] = 0
      "000000" when "0001000100111001", -- t[4409] = 0
      "000000" when "0001000100111010", -- t[4410] = 0
      "000000" when "0001000100111011", -- t[4411] = 0
      "000000" when "0001000100111100", -- t[4412] = 0
      "000000" when "0001000100111101", -- t[4413] = 0
      "000000" when "0001000100111110", -- t[4414] = 0
      "000000" when "0001000100111111", -- t[4415] = 0
      "000000" when "0001000101000000", -- t[4416] = 0
      "000000" when "0001000101000001", -- t[4417] = 0
      "000000" when "0001000101000010", -- t[4418] = 0
      "000000" when "0001000101000011", -- t[4419] = 0
      "000000" when "0001000101000100", -- t[4420] = 0
      "000000" when "0001000101000101", -- t[4421] = 0
      "000000" when "0001000101000110", -- t[4422] = 0
      "000000" when "0001000101000111", -- t[4423] = 0
      "000000" when "0001000101001000", -- t[4424] = 0
      "000000" when "0001000101001001", -- t[4425] = 0
      "000000" when "0001000101001010", -- t[4426] = 0
      "000000" when "0001000101001011", -- t[4427] = 0
      "000000" when "0001000101001100", -- t[4428] = 0
      "000000" when "0001000101001101", -- t[4429] = 0
      "000000" when "0001000101001110", -- t[4430] = 0
      "000000" when "0001000101001111", -- t[4431] = 0
      "000000" when "0001000101010000", -- t[4432] = 0
      "000000" when "0001000101010001", -- t[4433] = 0
      "000000" when "0001000101010010", -- t[4434] = 0
      "000000" when "0001000101010011", -- t[4435] = 0
      "000000" when "0001000101010100", -- t[4436] = 0
      "000000" when "0001000101010101", -- t[4437] = 0
      "000000" when "0001000101010110", -- t[4438] = 0
      "000000" when "0001000101010111", -- t[4439] = 0
      "000000" when "0001000101011000", -- t[4440] = 0
      "000000" when "0001000101011001", -- t[4441] = 0
      "000000" when "0001000101011010", -- t[4442] = 0
      "000000" when "0001000101011011", -- t[4443] = 0
      "000000" when "0001000101011100", -- t[4444] = 0
      "000000" when "0001000101011101", -- t[4445] = 0
      "000000" when "0001000101011110", -- t[4446] = 0
      "000000" when "0001000101011111", -- t[4447] = 0
      "000000" when "0001000101100000", -- t[4448] = 0
      "000000" when "0001000101100001", -- t[4449] = 0
      "000000" when "0001000101100010", -- t[4450] = 0
      "000000" when "0001000101100011", -- t[4451] = 0
      "000000" when "0001000101100100", -- t[4452] = 0
      "000000" when "0001000101100101", -- t[4453] = 0
      "000000" when "0001000101100110", -- t[4454] = 0
      "000000" when "0001000101100111", -- t[4455] = 0
      "000000" when "0001000101101000", -- t[4456] = 0
      "000000" when "0001000101101001", -- t[4457] = 0
      "000000" when "0001000101101010", -- t[4458] = 0
      "000000" when "0001000101101011", -- t[4459] = 0
      "000000" when "0001000101101100", -- t[4460] = 0
      "000000" when "0001000101101101", -- t[4461] = 0
      "000000" when "0001000101101110", -- t[4462] = 0
      "000000" when "0001000101101111", -- t[4463] = 0
      "000000" when "0001000101110000", -- t[4464] = 0
      "000000" when "0001000101110001", -- t[4465] = 0
      "000000" when "0001000101110010", -- t[4466] = 0
      "000000" when "0001000101110011", -- t[4467] = 0
      "000000" when "0001000101110100", -- t[4468] = 0
      "000000" when "0001000101110101", -- t[4469] = 0
      "000000" when "0001000101110110", -- t[4470] = 0
      "000000" when "0001000101110111", -- t[4471] = 0
      "000000" when "0001000101111000", -- t[4472] = 0
      "000000" when "0001000101111001", -- t[4473] = 0
      "000000" when "0001000101111010", -- t[4474] = 0
      "000000" when "0001000101111011", -- t[4475] = 0
      "000000" when "0001000101111100", -- t[4476] = 0
      "000000" when "0001000101111101", -- t[4477] = 0
      "000000" when "0001000101111110", -- t[4478] = 0
      "000000" when "0001000101111111", -- t[4479] = 0
      "000000" when "0001000110000000", -- t[4480] = 0
      "000000" when "0001000110000001", -- t[4481] = 0
      "000000" when "0001000110000010", -- t[4482] = 0
      "000000" when "0001000110000011", -- t[4483] = 0
      "000000" when "0001000110000100", -- t[4484] = 0
      "000000" when "0001000110000101", -- t[4485] = 0
      "000000" when "0001000110000110", -- t[4486] = 0
      "000000" when "0001000110000111", -- t[4487] = 0
      "000000" when "0001000110001000", -- t[4488] = 0
      "000000" when "0001000110001001", -- t[4489] = 0
      "000000" when "0001000110001010", -- t[4490] = 0
      "000000" when "0001000110001011", -- t[4491] = 0
      "000000" when "0001000110001100", -- t[4492] = 0
      "000000" when "0001000110001101", -- t[4493] = 0
      "000000" when "0001000110001110", -- t[4494] = 0
      "000000" when "0001000110001111", -- t[4495] = 0
      "000000" when "0001000110010000", -- t[4496] = 0
      "000000" when "0001000110010001", -- t[4497] = 0
      "000000" when "0001000110010010", -- t[4498] = 0
      "000000" when "0001000110010011", -- t[4499] = 0
      "000000" when "0001000110010100", -- t[4500] = 0
      "000000" when "0001000110010101", -- t[4501] = 0
      "000000" when "0001000110010110", -- t[4502] = 0
      "000000" when "0001000110010111", -- t[4503] = 0
      "000000" when "0001000110011000", -- t[4504] = 0
      "000000" when "0001000110011001", -- t[4505] = 0
      "000000" when "0001000110011010", -- t[4506] = 0
      "000000" when "0001000110011011", -- t[4507] = 0
      "000000" when "0001000110011100", -- t[4508] = 0
      "000000" when "0001000110011101", -- t[4509] = 0
      "000000" when "0001000110011110", -- t[4510] = 0
      "000000" when "0001000110011111", -- t[4511] = 0
      "000000" when "0001000110100000", -- t[4512] = 0
      "000000" when "0001000110100001", -- t[4513] = 0
      "000000" when "0001000110100010", -- t[4514] = 0
      "000000" when "0001000110100011", -- t[4515] = 0
      "000000" when "0001000110100100", -- t[4516] = 0
      "000000" when "0001000110100101", -- t[4517] = 0
      "000000" when "0001000110100110", -- t[4518] = 0
      "000000" when "0001000110100111", -- t[4519] = 0
      "000000" when "0001000110101000", -- t[4520] = 0
      "000000" when "0001000110101001", -- t[4521] = 0
      "000000" when "0001000110101010", -- t[4522] = 0
      "000000" when "0001000110101011", -- t[4523] = 0
      "000000" when "0001000110101100", -- t[4524] = 0
      "000000" when "0001000110101101", -- t[4525] = 0
      "000000" when "0001000110101110", -- t[4526] = 0
      "000000" when "0001000110101111", -- t[4527] = 0
      "000000" when "0001000110110000", -- t[4528] = 0
      "000000" when "0001000110110001", -- t[4529] = 0
      "000000" when "0001000110110010", -- t[4530] = 0
      "000000" when "0001000110110011", -- t[4531] = 0
      "000000" when "0001000110110100", -- t[4532] = 0
      "000000" when "0001000110110101", -- t[4533] = 0
      "000000" when "0001000110110110", -- t[4534] = 0
      "000000" when "0001000110110111", -- t[4535] = 0
      "000000" when "0001000110111000", -- t[4536] = 0
      "000000" when "0001000110111001", -- t[4537] = 0
      "000000" when "0001000110111010", -- t[4538] = 0
      "000000" when "0001000110111011", -- t[4539] = 0
      "000000" when "0001000110111100", -- t[4540] = 0
      "000000" when "0001000110111101", -- t[4541] = 0
      "000000" when "0001000110111110", -- t[4542] = 0
      "000000" when "0001000110111111", -- t[4543] = 0
      "000000" when "0001000111000000", -- t[4544] = 0
      "000000" when "0001000111000001", -- t[4545] = 0
      "000000" when "0001000111000010", -- t[4546] = 0
      "000000" when "0001000111000011", -- t[4547] = 0
      "000000" when "0001000111000100", -- t[4548] = 0
      "000000" when "0001000111000101", -- t[4549] = 0
      "000000" when "0001000111000110", -- t[4550] = 0
      "000000" when "0001000111000111", -- t[4551] = 0
      "000000" when "0001000111001000", -- t[4552] = 0
      "000000" when "0001000111001001", -- t[4553] = 0
      "000000" when "0001000111001010", -- t[4554] = 0
      "000000" when "0001000111001011", -- t[4555] = 0
      "000000" when "0001000111001100", -- t[4556] = 0
      "000000" when "0001000111001101", -- t[4557] = 0
      "000000" when "0001000111001110", -- t[4558] = 0
      "000000" when "0001000111001111", -- t[4559] = 0
      "000000" when "0001000111010000", -- t[4560] = 0
      "000000" when "0001000111010001", -- t[4561] = 0
      "000000" when "0001000111010010", -- t[4562] = 0
      "000000" when "0001000111010011", -- t[4563] = 0
      "000000" when "0001000111010100", -- t[4564] = 0
      "000000" when "0001000111010101", -- t[4565] = 0
      "000000" when "0001000111010110", -- t[4566] = 0
      "000000" when "0001000111010111", -- t[4567] = 0
      "000000" when "0001000111011000", -- t[4568] = 0
      "000000" when "0001000111011001", -- t[4569] = 0
      "000000" when "0001000111011010", -- t[4570] = 0
      "000000" when "0001000111011011", -- t[4571] = 0
      "000000" when "0001000111011100", -- t[4572] = 0
      "000000" when "0001000111011101", -- t[4573] = 0
      "000000" when "0001000111011110", -- t[4574] = 0
      "000000" when "0001000111011111", -- t[4575] = 0
      "000000" when "0001000111100000", -- t[4576] = 0
      "000000" when "0001000111100001", -- t[4577] = 0
      "000000" when "0001000111100010", -- t[4578] = 0
      "000000" when "0001000111100011", -- t[4579] = 0
      "000000" when "0001000111100100", -- t[4580] = 0
      "000000" when "0001000111100101", -- t[4581] = 0
      "000000" when "0001000111100110", -- t[4582] = 0
      "000000" when "0001000111100111", -- t[4583] = 0
      "000000" when "0001000111101000", -- t[4584] = 0
      "000000" when "0001000111101001", -- t[4585] = 0
      "000000" when "0001000111101010", -- t[4586] = 0
      "000000" when "0001000111101011", -- t[4587] = 0
      "000000" when "0001000111101100", -- t[4588] = 0
      "000000" when "0001000111101101", -- t[4589] = 0
      "000000" when "0001000111101110", -- t[4590] = 0
      "000000" when "0001000111101111", -- t[4591] = 0
      "000000" when "0001000111110000", -- t[4592] = 0
      "000000" when "0001000111110001", -- t[4593] = 0
      "000000" when "0001000111110010", -- t[4594] = 0
      "000000" when "0001000111110011", -- t[4595] = 0
      "000000" when "0001000111110100", -- t[4596] = 0
      "000000" when "0001000111110101", -- t[4597] = 0
      "000000" when "0001000111110110", -- t[4598] = 0
      "000000" when "0001000111110111", -- t[4599] = 0
      "000000" when "0001000111111000", -- t[4600] = 0
      "000000" when "0001000111111001", -- t[4601] = 0
      "000000" when "0001000111111010", -- t[4602] = 0
      "000000" when "0001000111111011", -- t[4603] = 0
      "000000" when "0001000111111100", -- t[4604] = 0
      "000000" when "0001000111111101", -- t[4605] = 0
      "000000" when "0001000111111110", -- t[4606] = 0
      "000000" when "0001000111111111", -- t[4607] = 0
      "000000" when "0001001000000000", -- t[4608] = 0
      "000000" when "0001001000000001", -- t[4609] = 0
      "000000" when "0001001000000010", -- t[4610] = 0
      "000000" when "0001001000000011", -- t[4611] = 0
      "000000" when "0001001000000100", -- t[4612] = 0
      "000000" when "0001001000000101", -- t[4613] = 0
      "000000" when "0001001000000110", -- t[4614] = 0
      "000000" when "0001001000000111", -- t[4615] = 0
      "000000" when "0001001000001000", -- t[4616] = 0
      "000000" when "0001001000001001", -- t[4617] = 0
      "000000" when "0001001000001010", -- t[4618] = 0
      "000000" when "0001001000001011", -- t[4619] = 0
      "000000" when "0001001000001100", -- t[4620] = 0
      "000000" when "0001001000001101", -- t[4621] = 0
      "000000" when "0001001000001110", -- t[4622] = 0
      "000000" when "0001001000001111", -- t[4623] = 0
      "000000" when "0001001000010000", -- t[4624] = 0
      "000000" when "0001001000010001", -- t[4625] = 0
      "000000" when "0001001000010010", -- t[4626] = 0
      "000000" when "0001001000010011", -- t[4627] = 0
      "000000" when "0001001000010100", -- t[4628] = 0
      "000000" when "0001001000010101", -- t[4629] = 0
      "000000" when "0001001000010110", -- t[4630] = 0
      "000000" when "0001001000010111", -- t[4631] = 0
      "000000" when "0001001000011000", -- t[4632] = 0
      "000000" when "0001001000011001", -- t[4633] = 0
      "000000" when "0001001000011010", -- t[4634] = 0
      "000000" when "0001001000011011", -- t[4635] = 0
      "000000" when "0001001000011100", -- t[4636] = 0
      "000000" when "0001001000011101", -- t[4637] = 0
      "000000" when "0001001000011110", -- t[4638] = 0
      "000000" when "0001001000011111", -- t[4639] = 0
      "000000" when "0001001000100000", -- t[4640] = 0
      "000000" when "0001001000100001", -- t[4641] = 0
      "000000" when "0001001000100010", -- t[4642] = 0
      "000000" when "0001001000100011", -- t[4643] = 0
      "000000" when "0001001000100100", -- t[4644] = 0
      "000000" when "0001001000100101", -- t[4645] = 0
      "000000" when "0001001000100110", -- t[4646] = 0
      "000000" when "0001001000100111", -- t[4647] = 0
      "000000" when "0001001000101000", -- t[4648] = 0
      "000000" when "0001001000101001", -- t[4649] = 0
      "000000" when "0001001000101010", -- t[4650] = 0
      "000000" when "0001001000101011", -- t[4651] = 0
      "000000" when "0001001000101100", -- t[4652] = 0
      "000000" when "0001001000101101", -- t[4653] = 0
      "000000" when "0001001000101110", -- t[4654] = 0
      "000000" when "0001001000101111", -- t[4655] = 0
      "000000" when "0001001000110000", -- t[4656] = 0
      "000000" when "0001001000110001", -- t[4657] = 0
      "000000" when "0001001000110010", -- t[4658] = 0
      "000000" when "0001001000110011", -- t[4659] = 0
      "000000" when "0001001000110100", -- t[4660] = 0
      "000000" when "0001001000110101", -- t[4661] = 0
      "000000" when "0001001000110110", -- t[4662] = 0
      "000000" when "0001001000110111", -- t[4663] = 0
      "000000" when "0001001000111000", -- t[4664] = 0
      "000000" when "0001001000111001", -- t[4665] = 0
      "000000" when "0001001000111010", -- t[4666] = 0
      "000000" when "0001001000111011", -- t[4667] = 0
      "000000" when "0001001000111100", -- t[4668] = 0
      "000000" when "0001001000111101", -- t[4669] = 0
      "000000" when "0001001000111110", -- t[4670] = 0
      "000000" when "0001001000111111", -- t[4671] = 0
      "000000" when "0001001001000000", -- t[4672] = 0
      "000000" when "0001001001000001", -- t[4673] = 0
      "000000" when "0001001001000010", -- t[4674] = 0
      "000000" when "0001001001000011", -- t[4675] = 0
      "000000" when "0001001001000100", -- t[4676] = 0
      "000000" when "0001001001000101", -- t[4677] = 0
      "000000" when "0001001001000110", -- t[4678] = 0
      "000000" when "0001001001000111", -- t[4679] = 0
      "000000" when "0001001001001000", -- t[4680] = 0
      "000000" when "0001001001001001", -- t[4681] = 0
      "000000" when "0001001001001010", -- t[4682] = 0
      "000000" when "0001001001001011", -- t[4683] = 0
      "000000" when "0001001001001100", -- t[4684] = 0
      "000000" when "0001001001001101", -- t[4685] = 0
      "000000" when "0001001001001110", -- t[4686] = 0
      "000000" when "0001001001001111", -- t[4687] = 0
      "000000" when "0001001001010000", -- t[4688] = 0
      "000000" when "0001001001010001", -- t[4689] = 0
      "000000" when "0001001001010010", -- t[4690] = 0
      "000000" when "0001001001010011", -- t[4691] = 0
      "000000" when "0001001001010100", -- t[4692] = 0
      "000000" when "0001001001010101", -- t[4693] = 0
      "000000" when "0001001001010110", -- t[4694] = 0
      "000000" when "0001001001010111", -- t[4695] = 0
      "000000" when "0001001001011000", -- t[4696] = 0
      "000000" when "0001001001011001", -- t[4697] = 0
      "000000" when "0001001001011010", -- t[4698] = 0
      "000000" when "0001001001011011", -- t[4699] = 0
      "000000" when "0001001001011100", -- t[4700] = 0
      "000000" when "0001001001011101", -- t[4701] = 0
      "000000" when "0001001001011110", -- t[4702] = 0
      "000000" when "0001001001011111", -- t[4703] = 0
      "000000" when "0001001001100000", -- t[4704] = 0
      "000000" when "0001001001100001", -- t[4705] = 0
      "000000" when "0001001001100010", -- t[4706] = 0
      "000000" when "0001001001100011", -- t[4707] = 0
      "000000" when "0001001001100100", -- t[4708] = 0
      "000000" when "0001001001100101", -- t[4709] = 0
      "000000" when "0001001001100110", -- t[4710] = 0
      "000000" when "0001001001100111", -- t[4711] = 0
      "000000" when "0001001001101000", -- t[4712] = 0
      "000000" when "0001001001101001", -- t[4713] = 0
      "000000" when "0001001001101010", -- t[4714] = 0
      "000000" when "0001001001101011", -- t[4715] = 0
      "000000" when "0001001001101100", -- t[4716] = 0
      "000000" when "0001001001101101", -- t[4717] = 0
      "000000" when "0001001001101110", -- t[4718] = 0
      "000000" when "0001001001101111", -- t[4719] = 0
      "000000" when "0001001001110000", -- t[4720] = 0
      "000000" when "0001001001110001", -- t[4721] = 0
      "000000" when "0001001001110010", -- t[4722] = 0
      "000000" when "0001001001110011", -- t[4723] = 0
      "000000" when "0001001001110100", -- t[4724] = 0
      "000000" when "0001001001110101", -- t[4725] = 0
      "000000" when "0001001001110110", -- t[4726] = 0
      "000000" when "0001001001110111", -- t[4727] = 0
      "000000" when "0001001001111000", -- t[4728] = 0
      "000000" when "0001001001111001", -- t[4729] = 0
      "000000" when "0001001001111010", -- t[4730] = 0
      "000000" when "0001001001111011", -- t[4731] = 0
      "000000" when "0001001001111100", -- t[4732] = 0
      "000000" when "0001001001111101", -- t[4733] = 0
      "000000" when "0001001001111110", -- t[4734] = 0
      "000000" when "0001001001111111", -- t[4735] = 0
      "000000" when "0001001010000000", -- t[4736] = 0
      "000000" when "0001001010000001", -- t[4737] = 0
      "000000" when "0001001010000010", -- t[4738] = 0
      "000000" when "0001001010000011", -- t[4739] = 0
      "000000" when "0001001010000100", -- t[4740] = 0
      "000000" when "0001001010000101", -- t[4741] = 0
      "000000" when "0001001010000110", -- t[4742] = 0
      "000000" when "0001001010000111", -- t[4743] = 0
      "000000" when "0001001010001000", -- t[4744] = 0
      "000000" when "0001001010001001", -- t[4745] = 0
      "000000" when "0001001010001010", -- t[4746] = 0
      "000000" when "0001001010001011", -- t[4747] = 0
      "000000" when "0001001010001100", -- t[4748] = 0
      "000000" when "0001001010001101", -- t[4749] = 0
      "000000" when "0001001010001110", -- t[4750] = 0
      "000000" when "0001001010001111", -- t[4751] = 0
      "000000" when "0001001010010000", -- t[4752] = 0
      "000000" when "0001001010010001", -- t[4753] = 0
      "000000" when "0001001010010010", -- t[4754] = 0
      "000000" when "0001001010010011", -- t[4755] = 0
      "000000" when "0001001010010100", -- t[4756] = 0
      "000000" when "0001001010010101", -- t[4757] = 0
      "000000" when "0001001010010110", -- t[4758] = 0
      "000000" when "0001001010010111", -- t[4759] = 0
      "000000" when "0001001010011000", -- t[4760] = 0
      "000000" when "0001001010011001", -- t[4761] = 0
      "000000" when "0001001010011010", -- t[4762] = 0
      "000000" when "0001001010011011", -- t[4763] = 0
      "000000" when "0001001010011100", -- t[4764] = 0
      "000000" when "0001001010011101", -- t[4765] = 0
      "000000" when "0001001010011110", -- t[4766] = 0
      "000000" when "0001001010011111", -- t[4767] = 0
      "000000" when "0001001010100000", -- t[4768] = 0
      "000000" when "0001001010100001", -- t[4769] = 0
      "000000" when "0001001010100010", -- t[4770] = 0
      "000000" when "0001001010100011", -- t[4771] = 0
      "000000" when "0001001010100100", -- t[4772] = 0
      "000000" when "0001001010100101", -- t[4773] = 0
      "000000" when "0001001010100110", -- t[4774] = 0
      "000000" when "0001001010100111", -- t[4775] = 0
      "000000" when "0001001010101000", -- t[4776] = 0
      "000000" when "0001001010101001", -- t[4777] = 0
      "000000" when "0001001010101010", -- t[4778] = 0
      "000000" when "0001001010101011", -- t[4779] = 0
      "000000" when "0001001010101100", -- t[4780] = 0
      "000000" when "0001001010101101", -- t[4781] = 0
      "000000" when "0001001010101110", -- t[4782] = 0
      "000000" when "0001001010101111", -- t[4783] = 0
      "000000" when "0001001010110000", -- t[4784] = 0
      "000000" when "0001001010110001", -- t[4785] = 0
      "000000" when "0001001010110010", -- t[4786] = 0
      "000000" when "0001001010110011", -- t[4787] = 0
      "000000" when "0001001010110100", -- t[4788] = 0
      "000000" when "0001001010110101", -- t[4789] = 0
      "000000" when "0001001010110110", -- t[4790] = 0
      "000000" when "0001001010110111", -- t[4791] = 0
      "000000" when "0001001010111000", -- t[4792] = 0
      "000000" when "0001001010111001", -- t[4793] = 0
      "000000" when "0001001010111010", -- t[4794] = 0
      "000000" when "0001001010111011", -- t[4795] = 0
      "000000" when "0001001010111100", -- t[4796] = 0
      "000000" when "0001001010111101", -- t[4797] = 0
      "000000" when "0001001010111110", -- t[4798] = 0
      "000000" when "0001001010111111", -- t[4799] = 0
      "000000" when "0001001011000000", -- t[4800] = 0
      "000000" when "0001001011000001", -- t[4801] = 0
      "000000" when "0001001011000010", -- t[4802] = 0
      "000000" when "0001001011000011", -- t[4803] = 0
      "000000" when "0001001011000100", -- t[4804] = 0
      "000000" when "0001001011000101", -- t[4805] = 0
      "000000" when "0001001011000110", -- t[4806] = 0
      "000000" when "0001001011000111", -- t[4807] = 0
      "000000" when "0001001011001000", -- t[4808] = 0
      "000000" when "0001001011001001", -- t[4809] = 0
      "000000" when "0001001011001010", -- t[4810] = 0
      "000000" when "0001001011001011", -- t[4811] = 0
      "000000" when "0001001011001100", -- t[4812] = 0
      "000000" when "0001001011001101", -- t[4813] = 0
      "000000" when "0001001011001110", -- t[4814] = 0
      "000000" when "0001001011001111", -- t[4815] = 0
      "000000" when "0001001011010000", -- t[4816] = 0
      "000000" when "0001001011010001", -- t[4817] = 0
      "000000" when "0001001011010010", -- t[4818] = 0
      "000000" when "0001001011010011", -- t[4819] = 0
      "000000" when "0001001011010100", -- t[4820] = 0
      "000000" when "0001001011010101", -- t[4821] = 0
      "000000" when "0001001011010110", -- t[4822] = 0
      "000000" when "0001001011010111", -- t[4823] = 0
      "000000" when "0001001011011000", -- t[4824] = 0
      "000000" when "0001001011011001", -- t[4825] = 0
      "000000" when "0001001011011010", -- t[4826] = 0
      "000000" when "0001001011011011", -- t[4827] = 0
      "000000" when "0001001011011100", -- t[4828] = 0
      "000000" when "0001001011011101", -- t[4829] = 0
      "000000" when "0001001011011110", -- t[4830] = 0
      "000000" when "0001001011011111", -- t[4831] = 0
      "000000" when "0001001011100000", -- t[4832] = 0
      "000000" when "0001001011100001", -- t[4833] = 0
      "000000" when "0001001011100010", -- t[4834] = 0
      "000000" when "0001001011100011", -- t[4835] = 0
      "000000" when "0001001011100100", -- t[4836] = 0
      "000000" when "0001001011100101", -- t[4837] = 0
      "000000" when "0001001011100110", -- t[4838] = 0
      "000000" when "0001001011100111", -- t[4839] = 0
      "000000" when "0001001011101000", -- t[4840] = 0
      "000000" when "0001001011101001", -- t[4841] = 0
      "000000" when "0001001011101010", -- t[4842] = 0
      "000000" when "0001001011101011", -- t[4843] = 0
      "000000" when "0001001011101100", -- t[4844] = 0
      "000000" when "0001001011101101", -- t[4845] = 0
      "000000" when "0001001011101110", -- t[4846] = 0
      "000000" when "0001001011101111", -- t[4847] = 0
      "000000" when "0001001011110000", -- t[4848] = 0
      "000000" when "0001001011110001", -- t[4849] = 0
      "000000" when "0001001011110010", -- t[4850] = 0
      "000000" when "0001001011110011", -- t[4851] = 0
      "000000" when "0001001011110100", -- t[4852] = 0
      "000000" when "0001001011110101", -- t[4853] = 0
      "000000" when "0001001011110110", -- t[4854] = 0
      "000000" when "0001001011110111", -- t[4855] = 0
      "000000" when "0001001011111000", -- t[4856] = 0
      "000000" when "0001001011111001", -- t[4857] = 0
      "000000" when "0001001011111010", -- t[4858] = 0
      "000000" when "0001001011111011", -- t[4859] = 0
      "000000" when "0001001011111100", -- t[4860] = 0
      "000000" when "0001001011111101", -- t[4861] = 0
      "000000" when "0001001011111110", -- t[4862] = 0
      "000000" when "0001001011111111", -- t[4863] = 0
      "000000" when "0001001100000000", -- t[4864] = 0
      "000000" when "0001001100000001", -- t[4865] = 0
      "000000" when "0001001100000010", -- t[4866] = 0
      "000000" when "0001001100000011", -- t[4867] = 0
      "000000" when "0001001100000100", -- t[4868] = 0
      "000000" when "0001001100000101", -- t[4869] = 0
      "000000" when "0001001100000110", -- t[4870] = 0
      "000000" when "0001001100000111", -- t[4871] = 0
      "000000" when "0001001100001000", -- t[4872] = 0
      "000000" when "0001001100001001", -- t[4873] = 0
      "000000" when "0001001100001010", -- t[4874] = 0
      "000000" when "0001001100001011", -- t[4875] = 0
      "000000" when "0001001100001100", -- t[4876] = 0
      "000000" when "0001001100001101", -- t[4877] = 0
      "000000" when "0001001100001110", -- t[4878] = 0
      "000000" when "0001001100001111", -- t[4879] = 0
      "000000" when "0001001100010000", -- t[4880] = 0
      "000000" when "0001001100010001", -- t[4881] = 0
      "000000" when "0001001100010010", -- t[4882] = 0
      "000000" when "0001001100010011", -- t[4883] = 0
      "000000" when "0001001100010100", -- t[4884] = 0
      "000000" when "0001001100010101", -- t[4885] = 0
      "000000" when "0001001100010110", -- t[4886] = 0
      "000000" when "0001001100010111", -- t[4887] = 0
      "000000" when "0001001100011000", -- t[4888] = 0
      "000000" when "0001001100011001", -- t[4889] = 0
      "000000" when "0001001100011010", -- t[4890] = 0
      "000000" when "0001001100011011", -- t[4891] = 0
      "000000" when "0001001100011100", -- t[4892] = 0
      "000000" when "0001001100011101", -- t[4893] = 0
      "000000" when "0001001100011110", -- t[4894] = 0
      "000000" when "0001001100011111", -- t[4895] = 0
      "000000" when "0001001100100000", -- t[4896] = 0
      "000000" when "0001001100100001", -- t[4897] = 0
      "000000" when "0001001100100010", -- t[4898] = 0
      "000000" when "0001001100100011", -- t[4899] = 0
      "000000" when "0001001100100100", -- t[4900] = 0
      "000000" when "0001001100100101", -- t[4901] = 0
      "000000" when "0001001100100110", -- t[4902] = 0
      "000000" when "0001001100100111", -- t[4903] = 0
      "000000" when "0001001100101000", -- t[4904] = 0
      "000000" when "0001001100101001", -- t[4905] = 0
      "000000" when "0001001100101010", -- t[4906] = 0
      "000000" when "0001001100101011", -- t[4907] = 0
      "000000" when "0001001100101100", -- t[4908] = 0
      "000000" when "0001001100101101", -- t[4909] = 0
      "000000" when "0001001100101110", -- t[4910] = 0
      "000000" when "0001001100101111", -- t[4911] = 0
      "000000" when "0001001100110000", -- t[4912] = 0
      "000000" when "0001001100110001", -- t[4913] = 0
      "000000" when "0001001100110010", -- t[4914] = 0
      "000000" when "0001001100110011", -- t[4915] = 0
      "000000" when "0001001100110100", -- t[4916] = 0
      "000000" when "0001001100110101", -- t[4917] = 0
      "000000" when "0001001100110110", -- t[4918] = 0
      "000000" when "0001001100110111", -- t[4919] = 0
      "000000" when "0001001100111000", -- t[4920] = 0
      "000000" when "0001001100111001", -- t[4921] = 0
      "000000" when "0001001100111010", -- t[4922] = 0
      "000000" when "0001001100111011", -- t[4923] = 0
      "000000" when "0001001100111100", -- t[4924] = 0
      "000000" when "0001001100111101", -- t[4925] = 0
      "000000" when "0001001100111110", -- t[4926] = 0
      "000000" when "0001001100111111", -- t[4927] = 0
      "000000" when "0001001101000000", -- t[4928] = 0
      "000000" when "0001001101000001", -- t[4929] = 0
      "000000" when "0001001101000010", -- t[4930] = 0
      "000000" when "0001001101000011", -- t[4931] = 0
      "000000" when "0001001101000100", -- t[4932] = 0
      "000000" when "0001001101000101", -- t[4933] = 0
      "000000" when "0001001101000110", -- t[4934] = 0
      "000000" when "0001001101000111", -- t[4935] = 0
      "000000" when "0001001101001000", -- t[4936] = 0
      "000000" when "0001001101001001", -- t[4937] = 0
      "000000" when "0001001101001010", -- t[4938] = 0
      "000000" when "0001001101001011", -- t[4939] = 0
      "000000" when "0001001101001100", -- t[4940] = 0
      "000000" when "0001001101001101", -- t[4941] = 0
      "000000" when "0001001101001110", -- t[4942] = 0
      "000000" when "0001001101001111", -- t[4943] = 0
      "000000" when "0001001101010000", -- t[4944] = 0
      "000000" when "0001001101010001", -- t[4945] = 0
      "000000" when "0001001101010010", -- t[4946] = 0
      "000000" when "0001001101010011", -- t[4947] = 0
      "000000" when "0001001101010100", -- t[4948] = 0
      "000000" when "0001001101010101", -- t[4949] = 0
      "000000" when "0001001101010110", -- t[4950] = 0
      "000000" when "0001001101010111", -- t[4951] = 0
      "000000" when "0001001101011000", -- t[4952] = 0
      "000000" when "0001001101011001", -- t[4953] = 0
      "000000" when "0001001101011010", -- t[4954] = 0
      "000000" when "0001001101011011", -- t[4955] = 0
      "000000" when "0001001101011100", -- t[4956] = 0
      "000000" when "0001001101011101", -- t[4957] = 0
      "000000" when "0001001101011110", -- t[4958] = 0
      "000000" when "0001001101011111", -- t[4959] = 0
      "000000" when "0001001101100000", -- t[4960] = 0
      "000000" when "0001001101100001", -- t[4961] = 0
      "000000" when "0001001101100010", -- t[4962] = 0
      "000000" when "0001001101100011", -- t[4963] = 0
      "000000" when "0001001101100100", -- t[4964] = 0
      "000000" when "0001001101100101", -- t[4965] = 0
      "000000" when "0001001101100110", -- t[4966] = 0
      "000000" when "0001001101100111", -- t[4967] = 0
      "000000" when "0001001101101000", -- t[4968] = 0
      "000000" when "0001001101101001", -- t[4969] = 0
      "000000" when "0001001101101010", -- t[4970] = 0
      "000000" when "0001001101101011", -- t[4971] = 0
      "000000" when "0001001101101100", -- t[4972] = 0
      "000000" when "0001001101101101", -- t[4973] = 0
      "000000" when "0001001101101110", -- t[4974] = 0
      "000000" when "0001001101101111", -- t[4975] = 0
      "000000" when "0001001101110000", -- t[4976] = 0
      "000000" when "0001001101110001", -- t[4977] = 0
      "000000" when "0001001101110010", -- t[4978] = 0
      "000000" when "0001001101110011", -- t[4979] = 0
      "000000" when "0001001101110100", -- t[4980] = 0
      "000000" when "0001001101110101", -- t[4981] = 0
      "000000" when "0001001101110110", -- t[4982] = 0
      "000000" when "0001001101110111", -- t[4983] = 0
      "000000" when "0001001101111000", -- t[4984] = 0
      "000000" when "0001001101111001", -- t[4985] = 0
      "000000" when "0001001101111010", -- t[4986] = 0
      "000000" when "0001001101111011", -- t[4987] = 0
      "000000" when "0001001101111100", -- t[4988] = 0
      "000000" when "0001001101111101", -- t[4989] = 0
      "000000" when "0001001101111110", -- t[4990] = 0
      "000000" when "0001001101111111", -- t[4991] = 0
      "000000" when "0001001110000000", -- t[4992] = 0
      "000000" when "0001001110000001", -- t[4993] = 0
      "000000" when "0001001110000010", -- t[4994] = 0
      "000000" when "0001001110000011", -- t[4995] = 0
      "000000" when "0001001110000100", -- t[4996] = 0
      "000000" when "0001001110000101", -- t[4997] = 0
      "000000" when "0001001110000110", -- t[4998] = 0
      "000000" when "0001001110000111", -- t[4999] = 0
      "000000" when "0001001110001000", -- t[5000] = 0
      "000000" when "0001001110001001", -- t[5001] = 0
      "000000" when "0001001110001010", -- t[5002] = 0
      "000000" when "0001001110001011", -- t[5003] = 0
      "000000" when "0001001110001100", -- t[5004] = 0
      "000000" when "0001001110001101", -- t[5005] = 0
      "000000" when "0001001110001110", -- t[5006] = 0
      "000000" when "0001001110001111", -- t[5007] = 0
      "000000" when "0001001110010000", -- t[5008] = 0
      "000000" when "0001001110010001", -- t[5009] = 0
      "000000" when "0001001110010010", -- t[5010] = 0
      "000000" when "0001001110010011", -- t[5011] = 0
      "000000" when "0001001110010100", -- t[5012] = 0
      "000000" when "0001001110010101", -- t[5013] = 0
      "000000" when "0001001110010110", -- t[5014] = 0
      "000000" when "0001001110010111", -- t[5015] = 0
      "000000" when "0001001110011000", -- t[5016] = 0
      "000000" when "0001001110011001", -- t[5017] = 0
      "000000" when "0001001110011010", -- t[5018] = 0
      "000000" when "0001001110011011", -- t[5019] = 0
      "000000" when "0001001110011100", -- t[5020] = 0
      "000000" when "0001001110011101", -- t[5021] = 0
      "000000" when "0001001110011110", -- t[5022] = 0
      "000000" when "0001001110011111", -- t[5023] = 0
      "000000" when "0001001110100000", -- t[5024] = 0
      "000000" when "0001001110100001", -- t[5025] = 0
      "000000" when "0001001110100010", -- t[5026] = 0
      "000000" when "0001001110100011", -- t[5027] = 0
      "000000" when "0001001110100100", -- t[5028] = 0
      "000000" when "0001001110100101", -- t[5029] = 0
      "000000" when "0001001110100110", -- t[5030] = 0
      "000000" when "0001001110100111", -- t[5031] = 0
      "000000" when "0001001110101000", -- t[5032] = 0
      "000000" when "0001001110101001", -- t[5033] = 0
      "000000" when "0001001110101010", -- t[5034] = 0
      "000000" when "0001001110101011", -- t[5035] = 0
      "000000" when "0001001110101100", -- t[5036] = 0
      "000000" when "0001001110101101", -- t[5037] = 0
      "000000" when "0001001110101110", -- t[5038] = 0
      "000000" when "0001001110101111", -- t[5039] = 0
      "000000" when "0001001110110000", -- t[5040] = 0
      "000000" when "0001001110110001", -- t[5041] = 0
      "000000" when "0001001110110010", -- t[5042] = 0
      "000000" when "0001001110110011", -- t[5043] = 0
      "000000" when "0001001110110100", -- t[5044] = 0
      "000000" when "0001001110110101", -- t[5045] = 0
      "000000" when "0001001110110110", -- t[5046] = 0
      "000000" when "0001001110110111", -- t[5047] = 0
      "000000" when "0001001110111000", -- t[5048] = 0
      "000000" when "0001001110111001", -- t[5049] = 0
      "000000" when "0001001110111010", -- t[5050] = 0
      "000000" when "0001001110111011", -- t[5051] = 0
      "000000" when "0001001110111100", -- t[5052] = 0
      "000000" when "0001001110111101", -- t[5053] = 0
      "000000" when "0001001110111110", -- t[5054] = 0
      "000000" when "0001001110111111", -- t[5055] = 0
      "000000" when "0001001111000000", -- t[5056] = 0
      "000000" when "0001001111000001", -- t[5057] = 0
      "000000" when "0001001111000010", -- t[5058] = 0
      "000000" when "0001001111000011", -- t[5059] = 0
      "000000" when "0001001111000100", -- t[5060] = 0
      "000000" when "0001001111000101", -- t[5061] = 0
      "000000" when "0001001111000110", -- t[5062] = 0
      "000000" when "0001001111000111", -- t[5063] = 0
      "000000" when "0001001111001000", -- t[5064] = 0
      "000000" when "0001001111001001", -- t[5065] = 0
      "000000" when "0001001111001010", -- t[5066] = 0
      "000000" when "0001001111001011", -- t[5067] = 0
      "000000" when "0001001111001100", -- t[5068] = 0
      "000000" when "0001001111001101", -- t[5069] = 0
      "000000" when "0001001111001110", -- t[5070] = 0
      "000000" when "0001001111001111", -- t[5071] = 0
      "000000" when "0001001111010000", -- t[5072] = 0
      "000000" when "0001001111010001", -- t[5073] = 0
      "000000" when "0001001111010010", -- t[5074] = 0
      "000000" when "0001001111010011", -- t[5075] = 0
      "000000" when "0001001111010100", -- t[5076] = 0
      "000000" when "0001001111010101", -- t[5077] = 0
      "000000" when "0001001111010110", -- t[5078] = 0
      "000000" when "0001001111010111", -- t[5079] = 0
      "000000" when "0001001111011000", -- t[5080] = 0
      "000000" when "0001001111011001", -- t[5081] = 0
      "000000" when "0001001111011010", -- t[5082] = 0
      "000000" when "0001001111011011", -- t[5083] = 0
      "000000" when "0001001111011100", -- t[5084] = 0
      "000000" when "0001001111011101", -- t[5085] = 0
      "000000" when "0001001111011110", -- t[5086] = 0
      "000000" when "0001001111011111", -- t[5087] = 0
      "000000" when "0001001111100000", -- t[5088] = 0
      "000000" when "0001001111100001", -- t[5089] = 0
      "000000" when "0001001111100010", -- t[5090] = 0
      "000000" when "0001001111100011", -- t[5091] = 0
      "000000" when "0001001111100100", -- t[5092] = 0
      "000000" when "0001001111100101", -- t[5093] = 0
      "000000" when "0001001111100110", -- t[5094] = 0
      "000000" when "0001001111100111", -- t[5095] = 0
      "000000" when "0001001111101000", -- t[5096] = 0
      "000000" when "0001001111101001", -- t[5097] = 0
      "000000" when "0001001111101010", -- t[5098] = 0
      "000000" when "0001001111101011", -- t[5099] = 0
      "000000" when "0001001111101100", -- t[5100] = 0
      "000000" when "0001001111101101", -- t[5101] = 0
      "000000" when "0001001111101110", -- t[5102] = 0
      "000000" when "0001001111101111", -- t[5103] = 0
      "000000" when "0001001111110000", -- t[5104] = 0
      "000000" when "0001001111110001", -- t[5105] = 0
      "000000" when "0001001111110010", -- t[5106] = 0
      "000000" when "0001001111110011", -- t[5107] = 0
      "000000" when "0001001111110100", -- t[5108] = 0
      "000000" when "0001001111110101", -- t[5109] = 0
      "000000" when "0001001111110110", -- t[5110] = 0
      "000000" when "0001001111110111", -- t[5111] = 0
      "000000" when "0001001111111000", -- t[5112] = 0
      "000000" when "0001001111111001", -- t[5113] = 0
      "000000" when "0001001111111010", -- t[5114] = 0
      "000000" when "0001001111111011", -- t[5115] = 0
      "000000" when "0001001111111100", -- t[5116] = 0
      "000000" when "0001001111111101", -- t[5117] = 0
      "000000" when "0001001111111110", -- t[5118] = 0
      "000000" when "0001001111111111", -- t[5119] = 0
      "000000" when "0001010000000000", -- t[5120] = 0
      "000000" when "0001010000000001", -- t[5121] = 0
      "000000" when "0001010000000010", -- t[5122] = 0
      "000000" when "0001010000000011", -- t[5123] = 0
      "000000" when "0001010000000100", -- t[5124] = 0
      "000000" when "0001010000000101", -- t[5125] = 0
      "000000" when "0001010000000110", -- t[5126] = 0
      "000000" when "0001010000000111", -- t[5127] = 0
      "000000" when "0001010000001000", -- t[5128] = 0
      "000000" when "0001010000001001", -- t[5129] = 0
      "000000" when "0001010000001010", -- t[5130] = 0
      "000000" when "0001010000001011", -- t[5131] = 0
      "000000" when "0001010000001100", -- t[5132] = 0
      "000000" when "0001010000001101", -- t[5133] = 0
      "000000" when "0001010000001110", -- t[5134] = 0
      "000000" when "0001010000001111", -- t[5135] = 0
      "000000" when "0001010000010000", -- t[5136] = 0
      "000000" when "0001010000010001", -- t[5137] = 0
      "000000" when "0001010000010010", -- t[5138] = 0
      "000000" when "0001010000010011", -- t[5139] = 0
      "000000" when "0001010000010100", -- t[5140] = 0
      "000000" when "0001010000010101", -- t[5141] = 0
      "000000" when "0001010000010110", -- t[5142] = 0
      "000000" when "0001010000010111", -- t[5143] = 0
      "000000" when "0001010000011000", -- t[5144] = 0
      "000000" when "0001010000011001", -- t[5145] = 0
      "000000" when "0001010000011010", -- t[5146] = 0
      "000000" when "0001010000011011", -- t[5147] = 0
      "000000" when "0001010000011100", -- t[5148] = 0
      "000000" when "0001010000011101", -- t[5149] = 0
      "000000" when "0001010000011110", -- t[5150] = 0
      "000000" when "0001010000011111", -- t[5151] = 0
      "000000" when "0001010000100000", -- t[5152] = 0
      "000000" when "0001010000100001", -- t[5153] = 0
      "000000" when "0001010000100010", -- t[5154] = 0
      "000000" when "0001010000100011", -- t[5155] = 0
      "000000" when "0001010000100100", -- t[5156] = 0
      "000000" when "0001010000100101", -- t[5157] = 0
      "000000" when "0001010000100110", -- t[5158] = 0
      "000000" when "0001010000100111", -- t[5159] = 0
      "000000" when "0001010000101000", -- t[5160] = 0
      "000000" when "0001010000101001", -- t[5161] = 0
      "000000" when "0001010000101010", -- t[5162] = 0
      "000000" when "0001010000101011", -- t[5163] = 0
      "000000" when "0001010000101100", -- t[5164] = 0
      "000000" when "0001010000101101", -- t[5165] = 0
      "000000" when "0001010000101110", -- t[5166] = 0
      "000000" when "0001010000101111", -- t[5167] = 0
      "000000" when "0001010000110000", -- t[5168] = 0
      "000000" when "0001010000110001", -- t[5169] = 0
      "000000" when "0001010000110010", -- t[5170] = 0
      "000000" when "0001010000110011", -- t[5171] = 0
      "000000" when "0001010000110100", -- t[5172] = 0
      "000000" when "0001010000110101", -- t[5173] = 0
      "000000" when "0001010000110110", -- t[5174] = 0
      "000000" when "0001010000110111", -- t[5175] = 0
      "000000" when "0001010000111000", -- t[5176] = 0
      "000000" when "0001010000111001", -- t[5177] = 0
      "000000" when "0001010000111010", -- t[5178] = 0
      "000000" when "0001010000111011", -- t[5179] = 0
      "000000" when "0001010000111100", -- t[5180] = 0
      "000000" when "0001010000111101", -- t[5181] = 0
      "000000" when "0001010000111110", -- t[5182] = 0
      "000000" when "0001010000111111", -- t[5183] = 0
      "000000" when "0001010001000000", -- t[5184] = 0
      "000000" when "0001010001000001", -- t[5185] = 0
      "000000" when "0001010001000010", -- t[5186] = 0
      "000000" when "0001010001000011", -- t[5187] = 0
      "000000" when "0001010001000100", -- t[5188] = 0
      "000000" when "0001010001000101", -- t[5189] = 0
      "000000" when "0001010001000110", -- t[5190] = 0
      "000000" when "0001010001000111", -- t[5191] = 0
      "000000" when "0001010001001000", -- t[5192] = 0
      "000000" when "0001010001001001", -- t[5193] = 0
      "000000" when "0001010001001010", -- t[5194] = 0
      "000000" when "0001010001001011", -- t[5195] = 0
      "000000" when "0001010001001100", -- t[5196] = 0
      "000000" when "0001010001001101", -- t[5197] = 0
      "000000" when "0001010001001110", -- t[5198] = 0
      "000000" when "0001010001001111", -- t[5199] = 0
      "000000" when "0001010001010000", -- t[5200] = 0
      "000000" when "0001010001010001", -- t[5201] = 0
      "000000" when "0001010001010010", -- t[5202] = 0
      "000000" when "0001010001010011", -- t[5203] = 0
      "000000" when "0001010001010100", -- t[5204] = 0
      "000000" when "0001010001010101", -- t[5205] = 0
      "000000" when "0001010001010110", -- t[5206] = 0
      "000000" when "0001010001010111", -- t[5207] = 0
      "000000" when "0001010001011000", -- t[5208] = 0
      "000000" when "0001010001011001", -- t[5209] = 0
      "000000" when "0001010001011010", -- t[5210] = 0
      "000000" when "0001010001011011", -- t[5211] = 0
      "000000" when "0001010001011100", -- t[5212] = 0
      "000000" when "0001010001011101", -- t[5213] = 0
      "000000" when "0001010001011110", -- t[5214] = 0
      "000000" when "0001010001011111", -- t[5215] = 0
      "000000" when "0001010001100000", -- t[5216] = 0
      "000000" when "0001010001100001", -- t[5217] = 0
      "000000" when "0001010001100010", -- t[5218] = 0
      "000000" when "0001010001100011", -- t[5219] = 0
      "000000" when "0001010001100100", -- t[5220] = 0
      "000000" when "0001010001100101", -- t[5221] = 0
      "000000" when "0001010001100110", -- t[5222] = 0
      "000000" when "0001010001100111", -- t[5223] = 0
      "000000" when "0001010001101000", -- t[5224] = 0
      "000000" when "0001010001101001", -- t[5225] = 0
      "000000" when "0001010001101010", -- t[5226] = 0
      "000000" when "0001010001101011", -- t[5227] = 0
      "000000" when "0001010001101100", -- t[5228] = 0
      "000000" when "0001010001101101", -- t[5229] = 0
      "000000" when "0001010001101110", -- t[5230] = 0
      "000000" when "0001010001101111", -- t[5231] = 0
      "000000" when "0001010001110000", -- t[5232] = 0
      "000000" when "0001010001110001", -- t[5233] = 0
      "000000" when "0001010001110010", -- t[5234] = 0
      "000000" when "0001010001110011", -- t[5235] = 0
      "000000" when "0001010001110100", -- t[5236] = 0
      "000000" when "0001010001110101", -- t[5237] = 0
      "000000" when "0001010001110110", -- t[5238] = 0
      "000000" when "0001010001110111", -- t[5239] = 0
      "000000" when "0001010001111000", -- t[5240] = 0
      "000000" when "0001010001111001", -- t[5241] = 0
      "000000" when "0001010001111010", -- t[5242] = 0
      "000000" when "0001010001111011", -- t[5243] = 0
      "000000" when "0001010001111100", -- t[5244] = 0
      "000000" when "0001010001111101", -- t[5245] = 0
      "000000" when "0001010001111110", -- t[5246] = 0
      "000000" when "0001010001111111", -- t[5247] = 0
      "000000" when "0001010010000000", -- t[5248] = 0
      "000000" when "0001010010000001", -- t[5249] = 0
      "000000" when "0001010010000010", -- t[5250] = 0
      "000000" when "0001010010000011", -- t[5251] = 0
      "000000" when "0001010010000100", -- t[5252] = 0
      "000000" when "0001010010000101", -- t[5253] = 0
      "000000" when "0001010010000110", -- t[5254] = 0
      "000000" when "0001010010000111", -- t[5255] = 0
      "000000" when "0001010010001000", -- t[5256] = 0
      "000000" when "0001010010001001", -- t[5257] = 0
      "000000" when "0001010010001010", -- t[5258] = 0
      "000000" when "0001010010001011", -- t[5259] = 0
      "000000" when "0001010010001100", -- t[5260] = 0
      "000000" when "0001010010001101", -- t[5261] = 0
      "000000" when "0001010010001110", -- t[5262] = 0
      "000000" when "0001010010001111", -- t[5263] = 0
      "000000" when "0001010010010000", -- t[5264] = 0
      "000000" when "0001010010010001", -- t[5265] = 0
      "000000" when "0001010010010010", -- t[5266] = 0
      "000000" when "0001010010010011", -- t[5267] = 0
      "000000" when "0001010010010100", -- t[5268] = 0
      "000000" when "0001010010010101", -- t[5269] = 0
      "000000" when "0001010010010110", -- t[5270] = 0
      "000000" when "0001010010010111", -- t[5271] = 0
      "000000" when "0001010010011000", -- t[5272] = 0
      "000000" when "0001010010011001", -- t[5273] = 0
      "000000" when "0001010010011010", -- t[5274] = 0
      "000000" when "0001010010011011", -- t[5275] = 0
      "000000" when "0001010010011100", -- t[5276] = 0
      "000000" when "0001010010011101", -- t[5277] = 0
      "000000" when "0001010010011110", -- t[5278] = 0
      "000000" when "0001010010011111", -- t[5279] = 0
      "000000" when "0001010010100000", -- t[5280] = 0
      "000000" when "0001010010100001", -- t[5281] = 0
      "000000" when "0001010010100010", -- t[5282] = 0
      "000000" when "0001010010100011", -- t[5283] = 0
      "000000" when "0001010010100100", -- t[5284] = 0
      "000000" when "0001010010100101", -- t[5285] = 0
      "000000" when "0001010010100110", -- t[5286] = 0
      "000000" when "0001010010100111", -- t[5287] = 0
      "000000" when "0001010010101000", -- t[5288] = 0
      "000000" when "0001010010101001", -- t[5289] = 0
      "000000" when "0001010010101010", -- t[5290] = 0
      "000000" when "0001010010101011", -- t[5291] = 0
      "000000" when "0001010010101100", -- t[5292] = 0
      "000000" when "0001010010101101", -- t[5293] = 0
      "000000" when "0001010010101110", -- t[5294] = 0
      "000000" when "0001010010101111", -- t[5295] = 0
      "000000" when "0001010010110000", -- t[5296] = 0
      "000000" when "0001010010110001", -- t[5297] = 0
      "000000" when "0001010010110010", -- t[5298] = 0
      "000000" when "0001010010110011", -- t[5299] = 0
      "000000" when "0001010010110100", -- t[5300] = 0
      "000000" when "0001010010110101", -- t[5301] = 0
      "000000" when "0001010010110110", -- t[5302] = 0
      "000000" when "0001010010110111", -- t[5303] = 0
      "000000" when "0001010010111000", -- t[5304] = 0
      "000000" when "0001010010111001", -- t[5305] = 0
      "000000" when "0001010010111010", -- t[5306] = 0
      "000000" when "0001010010111011", -- t[5307] = 0
      "000000" when "0001010010111100", -- t[5308] = 0
      "000000" when "0001010010111101", -- t[5309] = 0
      "000000" when "0001010010111110", -- t[5310] = 0
      "000000" when "0001010010111111", -- t[5311] = 0
      "000000" when "0001010011000000", -- t[5312] = 0
      "000000" when "0001010011000001", -- t[5313] = 0
      "000000" when "0001010011000010", -- t[5314] = 0
      "000000" when "0001010011000011", -- t[5315] = 0
      "000000" when "0001010011000100", -- t[5316] = 0
      "000000" when "0001010011000101", -- t[5317] = 0
      "000000" when "0001010011000110", -- t[5318] = 0
      "000000" when "0001010011000111", -- t[5319] = 0
      "000000" when "0001010011001000", -- t[5320] = 0
      "000000" when "0001010011001001", -- t[5321] = 0
      "000000" when "0001010011001010", -- t[5322] = 0
      "000000" when "0001010011001011", -- t[5323] = 0
      "000000" when "0001010011001100", -- t[5324] = 0
      "000000" when "0001010011001101", -- t[5325] = 0
      "000000" when "0001010011001110", -- t[5326] = 0
      "000000" when "0001010011001111", -- t[5327] = 0
      "000000" when "0001010011010000", -- t[5328] = 0
      "000000" when "0001010011010001", -- t[5329] = 0
      "000000" when "0001010011010010", -- t[5330] = 0
      "000000" when "0001010011010011", -- t[5331] = 0
      "000000" when "0001010011010100", -- t[5332] = 0
      "000000" when "0001010011010101", -- t[5333] = 0
      "000000" when "0001010011010110", -- t[5334] = 0
      "000000" when "0001010011010111", -- t[5335] = 0
      "000000" when "0001010011011000", -- t[5336] = 0
      "000000" when "0001010011011001", -- t[5337] = 0
      "000000" when "0001010011011010", -- t[5338] = 0
      "000000" when "0001010011011011", -- t[5339] = 0
      "000000" when "0001010011011100", -- t[5340] = 0
      "000000" when "0001010011011101", -- t[5341] = 0
      "000000" when "0001010011011110", -- t[5342] = 0
      "000000" when "0001010011011111", -- t[5343] = 0
      "000000" when "0001010011100000", -- t[5344] = 0
      "000000" when "0001010011100001", -- t[5345] = 0
      "000000" when "0001010011100010", -- t[5346] = 0
      "000000" when "0001010011100011", -- t[5347] = 0
      "000000" when "0001010011100100", -- t[5348] = 0
      "000000" when "0001010011100101", -- t[5349] = 0
      "000000" when "0001010011100110", -- t[5350] = 0
      "000000" when "0001010011100111", -- t[5351] = 0
      "000000" when "0001010011101000", -- t[5352] = 0
      "000000" when "0001010011101001", -- t[5353] = 0
      "000000" when "0001010011101010", -- t[5354] = 0
      "000000" when "0001010011101011", -- t[5355] = 0
      "000000" when "0001010011101100", -- t[5356] = 0
      "000000" when "0001010011101101", -- t[5357] = 0
      "000000" when "0001010011101110", -- t[5358] = 0
      "000000" when "0001010011101111", -- t[5359] = 0
      "000000" when "0001010011110000", -- t[5360] = 0
      "000000" when "0001010011110001", -- t[5361] = 0
      "000000" when "0001010011110010", -- t[5362] = 0
      "000000" when "0001010011110011", -- t[5363] = 0
      "000000" when "0001010011110100", -- t[5364] = 0
      "000000" when "0001010011110101", -- t[5365] = 0
      "000000" when "0001010011110110", -- t[5366] = 0
      "000000" when "0001010011110111", -- t[5367] = 0
      "000000" when "0001010011111000", -- t[5368] = 0
      "000000" when "0001010011111001", -- t[5369] = 0
      "000000" when "0001010011111010", -- t[5370] = 0
      "000000" when "0001010011111011", -- t[5371] = 0
      "000000" when "0001010011111100", -- t[5372] = 0
      "000000" when "0001010011111101", -- t[5373] = 0
      "000000" when "0001010011111110", -- t[5374] = 0
      "000000" when "0001010011111111", -- t[5375] = 0
      "000000" when "0001010100000000", -- t[5376] = 0
      "000000" when "0001010100000001", -- t[5377] = 0
      "000000" when "0001010100000010", -- t[5378] = 0
      "000000" when "0001010100000011", -- t[5379] = 0
      "000000" when "0001010100000100", -- t[5380] = 0
      "000000" when "0001010100000101", -- t[5381] = 0
      "000000" when "0001010100000110", -- t[5382] = 0
      "000000" when "0001010100000111", -- t[5383] = 0
      "000000" when "0001010100001000", -- t[5384] = 0
      "000000" when "0001010100001001", -- t[5385] = 0
      "000000" when "0001010100001010", -- t[5386] = 0
      "000000" when "0001010100001011", -- t[5387] = 0
      "000000" when "0001010100001100", -- t[5388] = 0
      "000000" when "0001010100001101", -- t[5389] = 0
      "000000" when "0001010100001110", -- t[5390] = 0
      "000000" when "0001010100001111", -- t[5391] = 0
      "000000" when "0001010100010000", -- t[5392] = 0
      "000000" when "0001010100010001", -- t[5393] = 0
      "000000" when "0001010100010010", -- t[5394] = 0
      "000000" when "0001010100010011", -- t[5395] = 0
      "000000" when "0001010100010100", -- t[5396] = 0
      "000000" when "0001010100010101", -- t[5397] = 0
      "000000" when "0001010100010110", -- t[5398] = 0
      "000000" when "0001010100010111", -- t[5399] = 0
      "000000" when "0001010100011000", -- t[5400] = 0
      "000000" when "0001010100011001", -- t[5401] = 0
      "000000" when "0001010100011010", -- t[5402] = 0
      "000000" when "0001010100011011", -- t[5403] = 0
      "000000" when "0001010100011100", -- t[5404] = 0
      "000000" when "0001010100011101", -- t[5405] = 0
      "000000" when "0001010100011110", -- t[5406] = 0
      "000000" when "0001010100011111", -- t[5407] = 0
      "000000" when "0001010100100000", -- t[5408] = 0
      "000000" when "0001010100100001", -- t[5409] = 0
      "000000" when "0001010100100010", -- t[5410] = 0
      "000000" when "0001010100100011", -- t[5411] = 0
      "000000" when "0001010100100100", -- t[5412] = 0
      "000000" when "0001010100100101", -- t[5413] = 0
      "000000" when "0001010100100110", -- t[5414] = 0
      "000000" when "0001010100100111", -- t[5415] = 0
      "000000" when "0001010100101000", -- t[5416] = 0
      "000000" when "0001010100101001", -- t[5417] = 0
      "000000" when "0001010100101010", -- t[5418] = 0
      "000000" when "0001010100101011", -- t[5419] = 0
      "000000" when "0001010100101100", -- t[5420] = 0
      "000000" when "0001010100101101", -- t[5421] = 0
      "000000" when "0001010100101110", -- t[5422] = 0
      "000000" when "0001010100101111", -- t[5423] = 0
      "000000" when "0001010100110000", -- t[5424] = 0
      "000000" when "0001010100110001", -- t[5425] = 0
      "000000" when "0001010100110010", -- t[5426] = 0
      "000000" when "0001010100110011", -- t[5427] = 0
      "000000" when "0001010100110100", -- t[5428] = 0
      "000000" when "0001010100110101", -- t[5429] = 0
      "000000" when "0001010100110110", -- t[5430] = 0
      "000000" when "0001010100110111", -- t[5431] = 0
      "000000" when "0001010100111000", -- t[5432] = 0
      "000000" when "0001010100111001", -- t[5433] = 0
      "000000" when "0001010100111010", -- t[5434] = 0
      "000000" when "0001010100111011", -- t[5435] = 0
      "000000" when "0001010100111100", -- t[5436] = 0
      "000000" when "0001010100111101", -- t[5437] = 0
      "000000" when "0001010100111110", -- t[5438] = 0
      "000000" when "0001010100111111", -- t[5439] = 0
      "000000" when "0001010101000000", -- t[5440] = 0
      "000000" when "0001010101000001", -- t[5441] = 0
      "000000" when "0001010101000010", -- t[5442] = 0
      "000000" when "0001010101000011", -- t[5443] = 0
      "000000" when "0001010101000100", -- t[5444] = 0
      "000000" when "0001010101000101", -- t[5445] = 0
      "000000" when "0001010101000110", -- t[5446] = 0
      "000000" when "0001010101000111", -- t[5447] = 0
      "000000" when "0001010101001000", -- t[5448] = 0
      "000000" when "0001010101001001", -- t[5449] = 0
      "000000" when "0001010101001010", -- t[5450] = 0
      "000000" when "0001010101001011", -- t[5451] = 0
      "000000" when "0001010101001100", -- t[5452] = 0
      "000000" when "0001010101001101", -- t[5453] = 0
      "000000" when "0001010101001110", -- t[5454] = 0
      "000000" when "0001010101001111", -- t[5455] = 0
      "000000" when "0001010101010000", -- t[5456] = 0
      "000000" when "0001010101010001", -- t[5457] = 0
      "000000" when "0001010101010010", -- t[5458] = 0
      "000000" when "0001010101010011", -- t[5459] = 0
      "000000" when "0001010101010100", -- t[5460] = 0
      "000000" when "0001010101010101", -- t[5461] = 0
      "000000" when "0001010101010110", -- t[5462] = 0
      "000000" when "0001010101010111", -- t[5463] = 0
      "000000" when "0001010101011000", -- t[5464] = 0
      "000000" when "0001010101011001", -- t[5465] = 0
      "000000" when "0001010101011010", -- t[5466] = 0
      "000000" when "0001010101011011", -- t[5467] = 0
      "000000" when "0001010101011100", -- t[5468] = 0
      "000000" when "0001010101011101", -- t[5469] = 0
      "000000" when "0001010101011110", -- t[5470] = 0
      "000000" when "0001010101011111", -- t[5471] = 0
      "000000" when "0001010101100000", -- t[5472] = 0
      "000000" when "0001010101100001", -- t[5473] = 0
      "000000" when "0001010101100010", -- t[5474] = 0
      "000000" when "0001010101100011", -- t[5475] = 0
      "000000" when "0001010101100100", -- t[5476] = 0
      "000000" when "0001010101100101", -- t[5477] = 0
      "000000" when "0001010101100110", -- t[5478] = 0
      "000000" when "0001010101100111", -- t[5479] = 0
      "000000" when "0001010101101000", -- t[5480] = 0
      "000000" when "0001010101101001", -- t[5481] = 0
      "000000" when "0001010101101010", -- t[5482] = 0
      "000000" when "0001010101101011", -- t[5483] = 0
      "000000" when "0001010101101100", -- t[5484] = 0
      "000000" when "0001010101101101", -- t[5485] = 0
      "000000" when "0001010101101110", -- t[5486] = 0
      "000000" when "0001010101101111", -- t[5487] = 0
      "000000" when "0001010101110000", -- t[5488] = 0
      "000000" when "0001010101110001", -- t[5489] = 0
      "000000" when "0001010101110010", -- t[5490] = 0
      "000000" when "0001010101110011", -- t[5491] = 0
      "000000" when "0001010101110100", -- t[5492] = 0
      "000000" when "0001010101110101", -- t[5493] = 0
      "000000" when "0001010101110110", -- t[5494] = 0
      "000000" when "0001010101110111", -- t[5495] = 0
      "000000" when "0001010101111000", -- t[5496] = 0
      "000000" when "0001010101111001", -- t[5497] = 0
      "000000" when "0001010101111010", -- t[5498] = 0
      "000000" when "0001010101111011", -- t[5499] = 0
      "000000" when "0001010101111100", -- t[5500] = 0
      "000000" when "0001010101111101", -- t[5501] = 0
      "000000" when "0001010101111110", -- t[5502] = 0
      "000000" when "0001010101111111", -- t[5503] = 0
      "000000" when "0001010110000000", -- t[5504] = 0
      "000000" when "0001010110000001", -- t[5505] = 0
      "000000" when "0001010110000010", -- t[5506] = 0
      "000000" when "0001010110000011", -- t[5507] = 0
      "000000" when "0001010110000100", -- t[5508] = 0
      "000000" when "0001010110000101", -- t[5509] = 0
      "000000" when "0001010110000110", -- t[5510] = 0
      "000000" when "0001010110000111", -- t[5511] = 0
      "000000" when "0001010110001000", -- t[5512] = 0
      "000000" when "0001010110001001", -- t[5513] = 0
      "000000" when "0001010110001010", -- t[5514] = 0
      "000000" when "0001010110001011", -- t[5515] = 0
      "000000" when "0001010110001100", -- t[5516] = 0
      "000000" when "0001010110001101", -- t[5517] = 0
      "000000" when "0001010110001110", -- t[5518] = 0
      "000000" when "0001010110001111", -- t[5519] = 0
      "000000" when "0001010110010000", -- t[5520] = 0
      "000000" when "0001010110010001", -- t[5521] = 0
      "000000" when "0001010110010010", -- t[5522] = 0
      "000000" when "0001010110010011", -- t[5523] = 0
      "000000" when "0001010110010100", -- t[5524] = 0
      "000000" when "0001010110010101", -- t[5525] = 0
      "000000" when "0001010110010110", -- t[5526] = 0
      "000000" when "0001010110010111", -- t[5527] = 0
      "000000" when "0001010110011000", -- t[5528] = 0
      "000000" when "0001010110011001", -- t[5529] = 0
      "000000" when "0001010110011010", -- t[5530] = 0
      "000000" when "0001010110011011", -- t[5531] = 0
      "000000" when "0001010110011100", -- t[5532] = 0
      "000000" when "0001010110011101", -- t[5533] = 0
      "000000" when "0001010110011110", -- t[5534] = 0
      "000000" when "0001010110011111", -- t[5535] = 0
      "000000" when "0001010110100000", -- t[5536] = 0
      "000000" when "0001010110100001", -- t[5537] = 0
      "000000" when "0001010110100010", -- t[5538] = 0
      "000000" when "0001010110100011", -- t[5539] = 0
      "000000" when "0001010110100100", -- t[5540] = 0
      "000000" when "0001010110100101", -- t[5541] = 0
      "000000" when "0001010110100110", -- t[5542] = 0
      "000000" when "0001010110100111", -- t[5543] = 0
      "000000" when "0001010110101000", -- t[5544] = 0
      "000000" when "0001010110101001", -- t[5545] = 0
      "000000" when "0001010110101010", -- t[5546] = 0
      "000000" when "0001010110101011", -- t[5547] = 0
      "000000" when "0001010110101100", -- t[5548] = 0
      "000000" when "0001010110101101", -- t[5549] = 0
      "000000" when "0001010110101110", -- t[5550] = 0
      "000000" when "0001010110101111", -- t[5551] = 0
      "000000" when "0001010110110000", -- t[5552] = 0
      "000000" when "0001010110110001", -- t[5553] = 0
      "000000" when "0001010110110010", -- t[5554] = 0
      "000000" when "0001010110110011", -- t[5555] = 0
      "000000" when "0001010110110100", -- t[5556] = 0
      "000000" when "0001010110110101", -- t[5557] = 0
      "000000" when "0001010110110110", -- t[5558] = 0
      "000000" when "0001010110110111", -- t[5559] = 0
      "000000" when "0001010110111000", -- t[5560] = 0
      "000000" when "0001010110111001", -- t[5561] = 0
      "000000" when "0001010110111010", -- t[5562] = 0
      "000000" when "0001010110111011", -- t[5563] = 0
      "000000" when "0001010110111100", -- t[5564] = 0
      "000000" when "0001010110111101", -- t[5565] = 0
      "000000" when "0001010110111110", -- t[5566] = 0
      "000000" when "0001010110111111", -- t[5567] = 0
      "000000" when "0001010111000000", -- t[5568] = 0
      "000000" when "0001010111000001", -- t[5569] = 0
      "000000" when "0001010111000010", -- t[5570] = 0
      "000000" when "0001010111000011", -- t[5571] = 0
      "000000" when "0001010111000100", -- t[5572] = 0
      "000000" when "0001010111000101", -- t[5573] = 0
      "000000" when "0001010111000110", -- t[5574] = 0
      "000000" when "0001010111000111", -- t[5575] = 0
      "000000" when "0001010111001000", -- t[5576] = 0
      "000000" when "0001010111001001", -- t[5577] = 0
      "000000" when "0001010111001010", -- t[5578] = 0
      "000000" when "0001010111001011", -- t[5579] = 0
      "000000" when "0001010111001100", -- t[5580] = 0
      "000000" when "0001010111001101", -- t[5581] = 0
      "000000" when "0001010111001110", -- t[5582] = 0
      "000000" when "0001010111001111", -- t[5583] = 0
      "000000" when "0001010111010000", -- t[5584] = 0
      "000000" when "0001010111010001", -- t[5585] = 0
      "000000" when "0001010111010010", -- t[5586] = 0
      "000000" when "0001010111010011", -- t[5587] = 0
      "000000" when "0001010111010100", -- t[5588] = 0
      "000000" when "0001010111010101", -- t[5589] = 0
      "000000" when "0001010111010110", -- t[5590] = 0
      "000000" when "0001010111010111", -- t[5591] = 0
      "000000" when "0001010111011000", -- t[5592] = 0
      "000000" when "0001010111011001", -- t[5593] = 0
      "000000" when "0001010111011010", -- t[5594] = 0
      "000000" when "0001010111011011", -- t[5595] = 0
      "000000" when "0001010111011100", -- t[5596] = 0
      "000000" when "0001010111011101", -- t[5597] = 0
      "000000" when "0001010111011110", -- t[5598] = 0
      "000000" when "0001010111011111", -- t[5599] = 0
      "000000" when "0001010111100000", -- t[5600] = 0
      "000000" when "0001010111100001", -- t[5601] = 0
      "000000" when "0001010111100010", -- t[5602] = 0
      "000000" when "0001010111100011", -- t[5603] = 0
      "000000" when "0001010111100100", -- t[5604] = 0
      "000000" when "0001010111100101", -- t[5605] = 0
      "000000" when "0001010111100110", -- t[5606] = 0
      "000000" when "0001010111100111", -- t[5607] = 0
      "000000" when "0001010111101000", -- t[5608] = 0
      "000000" when "0001010111101001", -- t[5609] = 0
      "000000" when "0001010111101010", -- t[5610] = 0
      "000000" when "0001010111101011", -- t[5611] = 0
      "000000" when "0001010111101100", -- t[5612] = 0
      "000000" when "0001010111101101", -- t[5613] = 0
      "000000" when "0001010111101110", -- t[5614] = 0
      "000000" when "0001010111101111", -- t[5615] = 0
      "000000" when "0001010111110000", -- t[5616] = 0
      "000000" when "0001010111110001", -- t[5617] = 0
      "000000" when "0001010111110010", -- t[5618] = 0
      "000000" when "0001010111110011", -- t[5619] = 0
      "000000" when "0001010111110100", -- t[5620] = 0
      "000000" when "0001010111110101", -- t[5621] = 0
      "000000" when "0001010111110110", -- t[5622] = 0
      "000000" when "0001010111110111", -- t[5623] = 0
      "000000" when "0001010111111000", -- t[5624] = 0
      "000000" when "0001010111111001", -- t[5625] = 0
      "000000" when "0001010111111010", -- t[5626] = 0
      "000000" when "0001010111111011", -- t[5627] = 0
      "000000" when "0001010111111100", -- t[5628] = 0
      "000000" when "0001010111111101", -- t[5629] = 0
      "000000" when "0001010111111110", -- t[5630] = 0
      "000000" when "0001010111111111", -- t[5631] = 0
      "000000" when "0001011000000000", -- t[5632] = 0
      "000000" when "0001011000000001", -- t[5633] = 0
      "000000" when "0001011000000010", -- t[5634] = 0
      "000000" when "0001011000000011", -- t[5635] = 0
      "000000" when "0001011000000100", -- t[5636] = 0
      "000000" when "0001011000000101", -- t[5637] = 0
      "000000" when "0001011000000110", -- t[5638] = 0
      "000000" when "0001011000000111", -- t[5639] = 0
      "000000" when "0001011000001000", -- t[5640] = 0
      "000000" when "0001011000001001", -- t[5641] = 0
      "000000" when "0001011000001010", -- t[5642] = 0
      "000000" when "0001011000001011", -- t[5643] = 0
      "000000" when "0001011000001100", -- t[5644] = 0
      "000000" when "0001011000001101", -- t[5645] = 0
      "000000" when "0001011000001110", -- t[5646] = 0
      "000000" when "0001011000001111", -- t[5647] = 0
      "000000" when "0001011000010000", -- t[5648] = 0
      "000000" when "0001011000010001", -- t[5649] = 0
      "000000" when "0001011000010010", -- t[5650] = 0
      "000000" when "0001011000010011", -- t[5651] = 0
      "000000" when "0001011000010100", -- t[5652] = 0
      "000000" when "0001011000010101", -- t[5653] = 0
      "000000" when "0001011000010110", -- t[5654] = 0
      "000000" when "0001011000010111", -- t[5655] = 0
      "000000" when "0001011000011000", -- t[5656] = 0
      "000000" when "0001011000011001", -- t[5657] = 0
      "000000" when "0001011000011010", -- t[5658] = 0
      "000000" when "0001011000011011", -- t[5659] = 0
      "000000" when "0001011000011100", -- t[5660] = 0
      "000000" when "0001011000011101", -- t[5661] = 0
      "000000" when "0001011000011110", -- t[5662] = 0
      "000000" when "0001011000011111", -- t[5663] = 0
      "000000" when "0001011000100000", -- t[5664] = 0
      "000000" when "0001011000100001", -- t[5665] = 0
      "000000" when "0001011000100010", -- t[5666] = 0
      "000000" when "0001011000100011", -- t[5667] = 0
      "000000" when "0001011000100100", -- t[5668] = 0
      "000000" when "0001011000100101", -- t[5669] = 0
      "000000" when "0001011000100110", -- t[5670] = 0
      "000000" when "0001011000100111", -- t[5671] = 0
      "000000" when "0001011000101000", -- t[5672] = 0
      "000000" when "0001011000101001", -- t[5673] = 0
      "000000" when "0001011000101010", -- t[5674] = 0
      "000000" when "0001011000101011", -- t[5675] = 0
      "000000" when "0001011000101100", -- t[5676] = 0
      "000000" when "0001011000101101", -- t[5677] = 0
      "000000" when "0001011000101110", -- t[5678] = 0
      "000000" when "0001011000101111", -- t[5679] = 0
      "000000" when "0001011000110000", -- t[5680] = 0
      "000000" when "0001011000110001", -- t[5681] = 0
      "000000" when "0001011000110010", -- t[5682] = 0
      "000000" when "0001011000110011", -- t[5683] = 0
      "000000" when "0001011000110100", -- t[5684] = 0
      "000000" when "0001011000110101", -- t[5685] = 0
      "000000" when "0001011000110110", -- t[5686] = 0
      "000000" when "0001011000110111", -- t[5687] = 0
      "000000" when "0001011000111000", -- t[5688] = 0
      "000000" when "0001011000111001", -- t[5689] = 0
      "000000" when "0001011000111010", -- t[5690] = 0
      "000000" when "0001011000111011", -- t[5691] = 0
      "000000" when "0001011000111100", -- t[5692] = 0
      "000000" when "0001011000111101", -- t[5693] = 0
      "000000" when "0001011000111110", -- t[5694] = 0
      "000000" when "0001011000111111", -- t[5695] = 0
      "000000" when "0001011001000000", -- t[5696] = 0
      "000000" when "0001011001000001", -- t[5697] = 0
      "000000" when "0001011001000010", -- t[5698] = 0
      "000000" when "0001011001000011", -- t[5699] = 0
      "000000" when "0001011001000100", -- t[5700] = 0
      "000000" when "0001011001000101", -- t[5701] = 0
      "000000" when "0001011001000110", -- t[5702] = 0
      "000000" when "0001011001000111", -- t[5703] = 0
      "000000" when "0001011001001000", -- t[5704] = 0
      "000000" when "0001011001001001", -- t[5705] = 0
      "000000" when "0001011001001010", -- t[5706] = 0
      "000000" when "0001011001001011", -- t[5707] = 0
      "000000" when "0001011001001100", -- t[5708] = 0
      "000000" when "0001011001001101", -- t[5709] = 0
      "000000" when "0001011001001110", -- t[5710] = 0
      "000000" when "0001011001001111", -- t[5711] = 0
      "000000" when "0001011001010000", -- t[5712] = 0
      "000000" when "0001011001010001", -- t[5713] = 0
      "000000" when "0001011001010010", -- t[5714] = 0
      "000000" when "0001011001010011", -- t[5715] = 0
      "000000" when "0001011001010100", -- t[5716] = 0
      "000000" when "0001011001010101", -- t[5717] = 0
      "000000" when "0001011001010110", -- t[5718] = 0
      "000000" when "0001011001010111", -- t[5719] = 0
      "000000" when "0001011001011000", -- t[5720] = 0
      "000000" when "0001011001011001", -- t[5721] = 0
      "000000" when "0001011001011010", -- t[5722] = 0
      "000000" when "0001011001011011", -- t[5723] = 0
      "000000" when "0001011001011100", -- t[5724] = 0
      "000000" when "0001011001011101", -- t[5725] = 0
      "000000" when "0001011001011110", -- t[5726] = 0
      "000000" when "0001011001011111", -- t[5727] = 0
      "000000" when "0001011001100000", -- t[5728] = 0
      "000000" when "0001011001100001", -- t[5729] = 0
      "000000" when "0001011001100010", -- t[5730] = 0
      "000000" when "0001011001100011", -- t[5731] = 0
      "000000" when "0001011001100100", -- t[5732] = 0
      "000000" when "0001011001100101", -- t[5733] = 0
      "000000" when "0001011001100110", -- t[5734] = 0
      "000000" when "0001011001100111", -- t[5735] = 0
      "000000" when "0001011001101000", -- t[5736] = 0
      "000000" when "0001011001101001", -- t[5737] = 0
      "000000" when "0001011001101010", -- t[5738] = 0
      "000000" when "0001011001101011", -- t[5739] = 0
      "000000" when "0001011001101100", -- t[5740] = 0
      "000000" when "0001011001101101", -- t[5741] = 0
      "000000" when "0001011001101110", -- t[5742] = 0
      "000000" when "0001011001101111", -- t[5743] = 0
      "000000" when "0001011001110000", -- t[5744] = 0
      "000000" when "0001011001110001", -- t[5745] = 0
      "000000" when "0001011001110010", -- t[5746] = 0
      "000000" when "0001011001110011", -- t[5747] = 0
      "000000" when "0001011001110100", -- t[5748] = 0
      "000000" when "0001011001110101", -- t[5749] = 0
      "000000" when "0001011001110110", -- t[5750] = 0
      "000000" when "0001011001110111", -- t[5751] = 0
      "000000" when "0001011001111000", -- t[5752] = 0
      "000000" when "0001011001111001", -- t[5753] = 0
      "000000" when "0001011001111010", -- t[5754] = 0
      "000000" when "0001011001111011", -- t[5755] = 0
      "000000" when "0001011001111100", -- t[5756] = 0
      "000000" when "0001011001111101", -- t[5757] = 0
      "000000" when "0001011001111110", -- t[5758] = 0
      "000000" when "0001011001111111", -- t[5759] = 0
      "000000" when "0001011010000000", -- t[5760] = 0
      "000000" when "0001011010000001", -- t[5761] = 0
      "000000" when "0001011010000010", -- t[5762] = 0
      "000000" when "0001011010000011", -- t[5763] = 0
      "000000" when "0001011010000100", -- t[5764] = 0
      "000000" when "0001011010000101", -- t[5765] = 0
      "000000" when "0001011010000110", -- t[5766] = 0
      "000000" when "0001011010000111", -- t[5767] = 0
      "000000" when "0001011010001000", -- t[5768] = 0
      "000000" when "0001011010001001", -- t[5769] = 0
      "000000" when "0001011010001010", -- t[5770] = 0
      "000000" when "0001011010001011", -- t[5771] = 0
      "000000" when "0001011010001100", -- t[5772] = 0
      "000000" when "0001011010001101", -- t[5773] = 0
      "000000" when "0001011010001110", -- t[5774] = 0
      "000000" when "0001011010001111", -- t[5775] = 0
      "000000" when "0001011010010000", -- t[5776] = 0
      "000000" when "0001011010010001", -- t[5777] = 0
      "000000" when "0001011010010010", -- t[5778] = 0
      "000000" when "0001011010010011", -- t[5779] = 0
      "000000" when "0001011010010100", -- t[5780] = 0
      "000000" when "0001011010010101", -- t[5781] = 0
      "000000" when "0001011010010110", -- t[5782] = 0
      "000000" when "0001011010010111", -- t[5783] = 0
      "000000" when "0001011010011000", -- t[5784] = 0
      "000000" when "0001011010011001", -- t[5785] = 0
      "000000" when "0001011010011010", -- t[5786] = 0
      "000000" when "0001011010011011", -- t[5787] = 0
      "000000" when "0001011010011100", -- t[5788] = 0
      "000000" when "0001011010011101", -- t[5789] = 0
      "000000" when "0001011010011110", -- t[5790] = 0
      "000000" when "0001011010011111", -- t[5791] = 0
      "000000" when "0001011010100000", -- t[5792] = 0
      "000000" when "0001011010100001", -- t[5793] = 0
      "000000" when "0001011010100010", -- t[5794] = 0
      "000000" when "0001011010100011", -- t[5795] = 0
      "000000" when "0001011010100100", -- t[5796] = 0
      "000000" when "0001011010100101", -- t[5797] = 0
      "000000" when "0001011010100110", -- t[5798] = 0
      "000000" when "0001011010100111", -- t[5799] = 0
      "000000" when "0001011010101000", -- t[5800] = 0
      "000000" when "0001011010101001", -- t[5801] = 0
      "000000" when "0001011010101010", -- t[5802] = 0
      "000000" when "0001011010101011", -- t[5803] = 0
      "000000" when "0001011010101100", -- t[5804] = 0
      "000000" when "0001011010101101", -- t[5805] = 0
      "000000" when "0001011010101110", -- t[5806] = 0
      "000000" when "0001011010101111", -- t[5807] = 0
      "000000" when "0001011010110000", -- t[5808] = 0
      "000000" when "0001011010110001", -- t[5809] = 0
      "000000" when "0001011010110010", -- t[5810] = 0
      "000000" when "0001011010110011", -- t[5811] = 0
      "000000" when "0001011010110100", -- t[5812] = 0
      "000000" when "0001011010110101", -- t[5813] = 0
      "000000" when "0001011010110110", -- t[5814] = 0
      "000000" when "0001011010110111", -- t[5815] = 0
      "000000" when "0001011010111000", -- t[5816] = 0
      "000000" when "0001011010111001", -- t[5817] = 0
      "000000" when "0001011010111010", -- t[5818] = 0
      "000000" when "0001011010111011", -- t[5819] = 0
      "000000" when "0001011010111100", -- t[5820] = 0
      "000000" when "0001011010111101", -- t[5821] = 0
      "000000" when "0001011010111110", -- t[5822] = 0
      "000000" when "0001011010111111", -- t[5823] = 0
      "000000" when "0001011011000000", -- t[5824] = 0
      "000000" when "0001011011000001", -- t[5825] = 0
      "000000" when "0001011011000010", -- t[5826] = 0
      "000000" when "0001011011000011", -- t[5827] = 0
      "000000" when "0001011011000100", -- t[5828] = 0
      "000000" when "0001011011000101", -- t[5829] = 0
      "000000" when "0001011011000110", -- t[5830] = 0
      "000000" when "0001011011000111", -- t[5831] = 0
      "000000" when "0001011011001000", -- t[5832] = 0
      "000000" when "0001011011001001", -- t[5833] = 0
      "000000" when "0001011011001010", -- t[5834] = 0
      "000000" when "0001011011001011", -- t[5835] = 0
      "000000" when "0001011011001100", -- t[5836] = 0
      "000000" when "0001011011001101", -- t[5837] = 0
      "000000" when "0001011011001110", -- t[5838] = 0
      "000000" when "0001011011001111", -- t[5839] = 0
      "000000" when "0001011011010000", -- t[5840] = 0
      "000000" when "0001011011010001", -- t[5841] = 0
      "000000" when "0001011011010010", -- t[5842] = 0
      "000000" when "0001011011010011", -- t[5843] = 0
      "000000" when "0001011011010100", -- t[5844] = 0
      "000000" when "0001011011010101", -- t[5845] = 0
      "000000" when "0001011011010110", -- t[5846] = 0
      "000000" when "0001011011010111", -- t[5847] = 0
      "000000" when "0001011011011000", -- t[5848] = 0
      "000000" when "0001011011011001", -- t[5849] = 0
      "000000" when "0001011011011010", -- t[5850] = 0
      "000000" when "0001011011011011", -- t[5851] = 0
      "000000" when "0001011011011100", -- t[5852] = 0
      "000000" when "0001011011011101", -- t[5853] = 0
      "000000" when "0001011011011110", -- t[5854] = 0
      "000000" when "0001011011011111", -- t[5855] = 0
      "000000" when "0001011011100000", -- t[5856] = 0
      "000000" when "0001011011100001", -- t[5857] = 0
      "000000" when "0001011011100010", -- t[5858] = 0
      "000000" when "0001011011100011", -- t[5859] = 0
      "000000" when "0001011011100100", -- t[5860] = 0
      "000000" when "0001011011100101", -- t[5861] = 0
      "000000" when "0001011011100110", -- t[5862] = 0
      "000000" when "0001011011100111", -- t[5863] = 0
      "000000" when "0001011011101000", -- t[5864] = 0
      "000000" when "0001011011101001", -- t[5865] = 0
      "000000" when "0001011011101010", -- t[5866] = 0
      "000000" when "0001011011101011", -- t[5867] = 0
      "000000" when "0001011011101100", -- t[5868] = 0
      "000000" when "0001011011101101", -- t[5869] = 0
      "000000" when "0001011011101110", -- t[5870] = 0
      "000000" when "0001011011101111", -- t[5871] = 0
      "000000" when "0001011011110000", -- t[5872] = 0
      "000000" when "0001011011110001", -- t[5873] = 0
      "000000" when "0001011011110010", -- t[5874] = 0
      "000000" when "0001011011110011", -- t[5875] = 0
      "000000" when "0001011011110100", -- t[5876] = 0
      "000000" when "0001011011110101", -- t[5877] = 0
      "000000" when "0001011011110110", -- t[5878] = 0
      "000000" when "0001011011110111", -- t[5879] = 0
      "000000" when "0001011011111000", -- t[5880] = 0
      "000000" when "0001011011111001", -- t[5881] = 0
      "000000" when "0001011011111010", -- t[5882] = 0
      "000000" when "0001011011111011", -- t[5883] = 0
      "000000" when "0001011011111100", -- t[5884] = 0
      "000000" when "0001011011111101", -- t[5885] = 0
      "000000" when "0001011011111110", -- t[5886] = 0
      "000000" when "0001011011111111", -- t[5887] = 0
      "000000" when "0001011100000000", -- t[5888] = 0
      "000000" when "0001011100000001", -- t[5889] = 0
      "000000" when "0001011100000010", -- t[5890] = 0
      "000000" when "0001011100000011", -- t[5891] = 0
      "000000" when "0001011100000100", -- t[5892] = 0
      "000000" when "0001011100000101", -- t[5893] = 0
      "000000" when "0001011100000110", -- t[5894] = 0
      "000000" when "0001011100000111", -- t[5895] = 0
      "000000" when "0001011100001000", -- t[5896] = 0
      "000000" when "0001011100001001", -- t[5897] = 0
      "000000" when "0001011100001010", -- t[5898] = 0
      "000000" when "0001011100001011", -- t[5899] = 0
      "000000" when "0001011100001100", -- t[5900] = 0
      "000000" when "0001011100001101", -- t[5901] = 0
      "000000" when "0001011100001110", -- t[5902] = 0
      "000000" when "0001011100001111", -- t[5903] = 0
      "000000" when "0001011100010000", -- t[5904] = 0
      "000000" when "0001011100010001", -- t[5905] = 0
      "000000" when "0001011100010010", -- t[5906] = 0
      "000000" when "0001011100010011", -- t[5907] = 0
      "000000" when "0001011100010100", -- t[5908] = 0
      "000000" when "0001011100010101", -- t[5909] = 0
      "000000" when "0001011100010110", -- t[5910] = 0
      "000000" when "0001011100010111", -- t[5911] = 0
      "000000" when "0001011100011000", -- t[5912] = 0
      "000000" when "0001011100011001", -- t[5913] = 0
      "000000" when "0001011100011010", -- t[5914] = 0
      "000000" when "0001011100011011", -- t[5915] = 0
      "000000" when "0001011100011100", -- t[5916] = 0
      "000000" when "0001011100011101", -- t[5917] = 0
      "000000" when "0001011100011110", -- t[5918] = 0
      "000000" when "0001011100011111", -- t[5919] = 0
      "000000" when "0001011100100000", -- t[5920] = 0
      "000000" when "0001011100100001", -- t[5921] = 0
      "000000" when "0001011100100010", -- t[5922] = 0
      "000000" when "0001011100100011", -- t[5923] = 0
      "000000" when "0001011100100100", -- t[5924] = 0
      "000000" when "0001011100100101", -- t[5925] = 0
      "000000" when "0001011100100110", -- t[5926] = 0
      "000000" when "0001011100100111", -- t[5927] = 0
      "000000" when "0001011100101000", -- t[5928] = 0
      "000000" when "0001011100101001", -- t[5929] = 0
      "000000" when "0001011100101010", -- t[5930] = 0
      "000000" when "0001011100101011", -- t[5931] = 0
      "000000" when "0001011100101100", -- t[5932] = 0
      "000000" when "0001011100101101", -- t[5933] = 0
      "000000" when "0001011100101110", -- t[5934] = 0
      "000000" when "0001011100101111", -- t[5935] = 0
      "000000" when "0001011100110000", -- t[5936] = 0
      "000000" when "0001011100110001", -- t[5937] = 0
      "000000" when "0001011100110010", -- t[5938] = 0
      "000000" when "0001011100110011", -- t[5939] = 0
      "000000" when "0001011100110100", -- t[5940] = 0
      "000000" when "0001011100110101", -- t[5941] = 0
      "000000" when "0001011100110110", -- t[5942] = 0
      "000000" when "0001011100110111", -- t[5943] = 0
      "000000" when "0001011100111000", -- t[5944] = 0
      "000000" when "0001011100111001", -- t[5945] = 0
      "000000" when "0001011100111010", -- t[5946] = 0
      "000000" when "0001011100111011", -- t[5947] = 0
      "000000" when "0001011100111100", -- t[5948] = 0
      "000000" when "0001011100111101", -- t[5949] = 0
      "000000" when "0001011100111110", -- t[5950] = 0
      "000000" when "0001011100111111", -- t[5951] = 0
      "000000" when "0001011101000000", -- t[5952] = 0
      "000000" when "0001011101000001", -- t[5953] = 0
      "000000" when "0001011101000010", -- t[5954] = 0
      "000000" when "0001011101000011", -- t[5955] = 0
      "000000" when "0001011101000100", -- t[5956] = 0
      "000000" when "0001011101000101", -- t[5957] = 0
      "000000" when "0001011101000110", -- t[5958] = 0
      "000000" when "0001011101000111", -- t[5959] = 0
      "000000" when "0001011101001000", -- t[5960] = 0
      "000000" when "0001011101001001", -- t[5961] = 0
      "000000" when "0001011101001010", -- t[5962] = 0
      "000000" when "0001011101001011", -- t[5963] = 0
      "000000" when "0001011101001100", -- t[5964] = 0
      "000000" when "0001011101001101", -- t[5965] = 0
      "000000" when "0001011101001110", -- t[5966] = 0
      "000000" when "0001011101001111", -- t[5967] = 0
      "000000" when "0001011101010000", -- t[5968] = 0
      "000000" when "0001011101010001", -- t[5969] = 0
      "000000" when "0001011101010010", -- t[5970] = 0
      "000000" when "0001011101010011", -- t[5971] = 0
      "000000" when "0001011101010100", -- t[5972] = 0
      "000000" when "0001011101010101", -- t[5973] = 0
      "000000" when "0001011101010110", -- t[5974] = 0
      "000000" when "0001011101010111", -- t[5975] = 0
      "000000" when "0001011101011000", -- t[5976] = 0
      "000000" when "0001011101011001", -- t[5977] = 0
      "000000" when "0001011101011010", -- t[5978] = 0
      "000000" when "0001011101011011", -- t[5979] = 0
      "000000" when "0001011101011100", -- t[5980] = 0
      "000000" when "0001011101011101", -- t[5981] = 0
      "000000" when "0001011101011110", -- t[5982] = 0
      "000000" when "0001011101011111", -- t[5983] = 0
      "000000" when "0001011101100000", -- t[5984] = 0
      "000000" when "0001011101100001", -- t[5985] = 0
      "000000" when "0001011101100010", -- t[5986] = 0
      "000000" when "0001011101100011", -- t[5987] = 0
      "000000" when "0001011101100100", -- t[5988] = 0
      "000000" when "0001011101100101", -- t[5989] = 0
      "000000" when "0001011101100110", -- t[5990] = 0
      "000000" when "0001011101100111", -- t[5991] = 0
      "000000" when "0001011101101000", -- t[5992] = 0
      "000000" when "0001011101101001", -- t[5993] = 0
      "000000" when "0001011101101010", -- t[5994] = 0
      "000000" when "0001011101101011", -- t[5995] = 0
      "000000" when "0001011101101100", -- t[5996] = 0
      "000000" when "0001011101101101", -- t[5997] = 0
      "000000" when "0001011101101110", -- t[5998] = 0
      "000000" when "0001011101101111", -- t[5999] = 0
      "000000" when "0001011101110000", -- t[6000] = 0
      "000000" when "0001011101110001", -- t[6001] = 0
      "000000" when "0001011101110010", -- t[6002] = 0
      "000000" when "0001011101110011", -- t[6003] = 0
      "000000" when "0001011101110100", -- t[6004] = 0
      "000000" when "0001011101110101", -- t[6005] = 0
      "000000" when "0001011101110110", -- t[6006] = 0
      "000000" when "0001011101110111", -- t[6007] = 0
      "000000" when "0001011101111000", -- t[6008] = 0
      "000000" when "0001011101111001", -- t[6009] = 0
      "000000" when "0001011101111010", -- t[6010] = 0
      "000000" when "0001011101111011", -- t[6011] = 0
      "000000" when "0001011101111100", -- t[6012] = 0
      "000000" when "0001011101111101", -- t[6013] = 0
      "000000" when "0001011101111110", -- t[6014] = 0
      "000000" when "0001011101111111", -- t[6015] = 0
      "000000" when "0001011110000000", -- t[6016] = 0
      "000000" when "0001011110000001", -- t[6017] = 0
      "000000" when "0001011110000010", -- t[6018] = 0
      "000000" when "0001011110000011", -- t[6019] = 0
      "000000" when "0001011110000100", -- t[6020] = 0
      "000000" when "0001011110000101", -- t[6021] = 0
      "000000" when "0001011110000110", -- t[6022] = 0
      "000000" when "0001011110000111", -- t[6023] = 0
      "000000" when "0001011110001000", -- t[6024] = 0
      "000000" when "0001011110001001", -- t[6025] = 0
      "000000" when "0001011110001010", -- t[6026] = 0
      "000000" when "0001011110001011", -- t[6027] = 0
      "000000" when "0001011110001100", -- t[6028] = 0
      "000000" when "0001011110001101", -- t[6029] = 0
      "000000" when "0001011110001110", -- t[6030] = 0
      "000000" when "0001011110001111", -- t[6031] = 0
      "000000" when "0001011110010000", -- t[6032] = 0
      "000000" when "0001011110010001", -- t[6033] = 0
      "000000" when "0001011110010010", -- t[6034] = 0
      "000000" when "0001011110010011", -- t[6035] = 0
      "000000" when "0001011110010100", -- t[6036] = 0
      "000000" when "0001011110010101", -- t[6037] = 0
      "000000" when "0001011110010110", -- t[6038] = 0
      "000000" when "0001011110010111", -- t[6039] = 0
      "000000" when "0001011110011000", -- t[6040] = 0
      "000000" when "0001011110011001", -- t[6041] = 0
      "000000" when "0001011110011010", -- t[6042] = 0
      "000000" when "0001011110011011", -- t[6043] = 0
      "000000" when "0001011110011100", -- t[6044] = 0
      "000000" when "0001011110011101", -- t[6045] = 0
      "000000" when "0001011110011110", -- t[6046] = 0
      "000000" when "0001011110011111", -- t[6047] = 0
      "000000" when "0001011110100000", -- t[6048] = 0
      "000000" when "0001011110100001", -- t[6049] = 0
      "000000" when "0001011110100010", -- t[6050] = 0
      "000000" when "0001011110100011", -- t[6051] = 0
      "000000" when "0001011110100100", -- t[6052] = 0
      "000000" when "0001011110100101", -- t[6053] = 0
      "000000" when "0001011110100110", -- t[6054] = 0
      "000000" when "0001011110100111", -- t[6055] = 0
      "000000" when "0001011110101000", -- t[6056] = 0
      "000000" when "0001011110101001", -- t[6057] = 0
      "000000" when "0001011110101010", -- t[6058] = 0
      "000000" when "0001011110101011", -- t[6059] = 0
      "000000" when "0001011110101100", -- t[6060] = 0
      "000000" when "0001011110101101", -- t[6061] = 0
      "000000" when "0001011110101110", -- t[6062] = 0
      "000000" when "0001011110101111", -- t[6063] = 0
      "000000" when "0001011110110000", -- t[6064] = 0
      "000000" when "0001011110110001", -- t[6065] = 0
      "000000" when "0001011110110010", -- t[6066] = 0
      "000000" when "0001011110110011", -- t[6067] = 0
      "000000" when "0001011110110100", -- t[6068] = 0
      "000000" when "0001011110110101", -- t[6069] = 0
      "000000" when "0001011110110110", -- t[6070] = 0
      "000000" when "0001011110110111", -- t[6071] = 0
      "000000" when "0001011110111000", -- t[6072] = 0
      "000000" when "0001011110111001", -- t[6073] = 0
      "000000" when "0001011110111010", -- t[6074] = 0
      "000000" when "0001011110111011", -- t[6075] = 0
      "000000" when "0001011110111100", -- t[6076] = 0
      "000000" when "0001011110111101", -- t[6077] = 0
      "000000" when "0001011110111110", -- t[6078] = 0
      "000000" when "0001011110111111", -- t[6079] = 0
      "000000" when "0001011111000000", -- t[6080] = 0
      "000000" when "0001011111000001", -- t[6081] = 0
      "000000" when "0001011111000010", -- t[6082] = 0
      "000000" when "0001011111000011", -- t[6083] = 0
      "000000" when "0001011111000100", -- t[6084] = 0
      "000000" when "0001011111000101", -- t[6085] = 0
      "000000" when "0001011111000110", -- t[6086] = 0
      "000000" when "0001011111000111", -- t[6087] = 0
      "000000" when "0001011111001000", -- t[6088] = 0
      "000000" when "0001011111001001", -- t[6089] = 0
      "000000" when "0001011111001010", -- t[6090] = 0
      "000000" when "0001011111001011", -- t[6091] = 0
      "000000" when "0001011111001100", -- t[6092] = 0
      "000000" when "0001011111001101", -- t[6093] = 0
      "000000" when "0001011111001110", -- t[6094] = 0
      "000000" when "0001011111001111", -- t[6095] = 0
      "000000" when "0001011111010000", -- t[6096] = 0
      "000000" when "0001011111010001", -- t[6097] = 0
      "000000" when "0001011111010010", -- t[6098] = 0
      "000000" when "0001011111010011", -- t[6099] = 0
      "000000" when "0001011111010100", -- t[6100] = 0
      "000000" when "0001011111010101", -- t[6101] = 0
      "000000" when "0001011111010110", -- t[6102] = 0
      "000000" when "0001011111010111", -- t[6103] = 0
      "000000" when "0001011111011000", -- t[6104] = 0
      "000000" when "0001011111011001", -- t[6105] = 0
      "000000" when "0001011111011010", -- t[6106] = 0
      "000000" when "0001011111011011", -- t[6107] = 0
      "000000" when "0001011111011100", -- t[6108] = 0
      "000000" when "0001011111011101", -- t[6109] = 0
      "000000" when "0001011111011110", -- t[6110] = 0
      "000000" when "0001011111011111", -- t[6111] = 0
      "000000" when "0001011111100000", -- t[6112] = 0
      "000000" when "0001011111100001", -- t[6113] = 0
      "000000" when "0001011111100010", -- t[6114] = 0
      "000000" when "0001011111100011", -- t[6115] = 0
      "000000" when "0001011111100100", -- t[6116] = 0
      "000000" when "0001011111100101", -- t[6117] = 0
      "000000" when "0001011111100110", -- t[6118] = 0
      "000000" when "0001011111100111", -- t[6119] = 0
      "000000" when "0001011111101000", -- t[6120] = 0
      "000000" when "0001011111101001", -- t[6121] = 0
      "000000" when "0001011111101010", -- t[6122] = 0
      "000000" when "0001011111101011", -- t[6123] = 0
      "000000" when "0001011111101100", -- t[6124] = 0
      "000000" when "0001011111101101", -- t[6125] = 0
      "000000" when "0001011111101110", -- t[6126] = 0
      "000000" when "0001011111101111", -- t[6127] = 0
      "000000" when "0001011111110000", -- t[6128] = 0
      "000000" when "0001011111110001", -- t[6129] = 0
      "000000" when "0001011111110010", -- t[6130] = 0
      "000000" when "0001011111110011", -- t[6131] = 0
      "000000" when "0001011111110100", -- t[6132] = 0
      "000000" when "0001011111110101", -- t[6133] = 0
      "000000" when "0001011111110110", -- t[6134] = 0
      "000000" when "0001011111110111", -- t[6135] = 0
      "000000" when "0001011111111000", -- t[6136] = 0
      "000000" when "0001011111111001", -- t[6137] = 0
      "000000" when "0001011111111010", -- t[6138] = 0
      "000000" when "0001011111111011", -- t[6139] = 0
      "000000" when "0001011111111100", -- t[6140] = 0
      "000000" when "0001011111111101", -- t[6141] = 0
      "000000" when "0001011111111110", -- t[6142] = 0
      "000000" when "0001011111111111", -- t[6143] = 0
      "000000" when "0001100000000000", -- t[6144] = 0
      "000000" when "0001100000000001", -- t[6145] = 0
      "000000" when "0001100000000010", -- t[6146] = 0
      "000000" when "0001100000000011", -- t[6147] = 0
      "000000" when "0001100000000100", -- t[6148] = 0
      "000000" when "0001100000000101", -- t[6149] = 0
      "000000" when "0001100000000110", -- t[6150] = 0
      "000000" when "0001100000000111", -- t[6151] = 0
      "000000" when "0001100000001000", -- t[6152] = 0
      "000000" when "0001100000001001", -- t[6153] = 0
      "000000" when "0001100000001010", -- t[6154] = 0
      "000000" when "0001100000001011", -- t[6155] = 0
      "000000" when "0001100000001100", -- t[6156] = 0
      "000000" when "0001100000001101", -- t[6157] = 0
      "000000" when "0001100000001110", -- t[6158] = 0
      "000000" when "0001100000001111", -- t[6159] = 0
      "000000" when "0001100000010000", -- t[6160] = 0
      "000000" when "0001100000010001", -- t[6161] = 0
      "000000" when "0001100000010010", -- t[6162] = 0
      "000000" when "0001100000010011", -- t[6163] = 0
      "000000" when "0001100000010100", -- t[6164] = 0
      "000000" when "0001100000010101", -- t[6165] = 0
      "000000" when "0001100000010110", -- t[6166] = 0
      "000000" when "0001100000010111", -- t[6167] = 0
      "000000" when "0001100000011000", -- t[6168] = 0
      "000000" when "0001100000011001", -- t[6169] = 0
      "000000" when "0001100000011010", -- t[6170] = 0
      "000000" when "0001100000011011", -- t[6171] = 0
      "000000" when "0001100000011100", -- t[6172] = 0
      "000000" when "0001100000011101", -- t[6173] = 0
      "000000" when "0001100000011110", -- t[6174] = 0
      "000000" when "0001100000011111", -- t[6175] = 0
      "000000" when "0001100000100000", -- t[6176] = 0
      "000000" when "0001100000100001", -- t[6177] = 0
      "000000" when "0001100000100010", -- t[6178] = 0
      "000000" when "0001100000100011", -- t[6179] = 0
      "000000" when "0001100000100100", -- t[6180] = 0
      "000000" when "0001100000100101", -- t[6181] = 0
      "000000" when "0001100000100110", -- t[6182] = 0
      "000000" when "0001100000100111", -- t[6183] = 0
      "000000" when "0001100000101000", -- t[6184] = 0
      "000000" when "0001100000101001", -- t[6185] = 0
      "000000" when "0001100000101010", -- t[6186] = 0
      "000000" when "0001100000101011", -- t[6187] = 0
      "000000" when "0001100000101100", -- t[6188] = 0
      "000000" when "0001100000101101", -- t[6189] = 0
      "000000" when "0001100000101110", -- t[6190] = 0
      "000000" when "0001100000101111", -- t[6191] = 0
      "000000" when "0001100000110000", -- t[6192] = 0
      "000000" when "0001100000110001", -- t[6193] = 0
      "000000" when "0001100000110010", -- t[6194] = 0
      "000000" when "0001100000110011", -- t[6195] = 0
      "000000" when "0001100000110100", -- t[6196] = 0
      "000000" when "0001100000110101", -- t[6197] = 0
      "000000" when "0001100000110110", -- t[6198] = 0
      "000000" when "0001100000110111", -- t[6199] = 0
      "000000" when "0001100000111000", -- t[6200] = 0
      "000000" when "0001100000111001", -- t[6201] = 0
      "000000" when "0001100000111010", -- t[6202] = 0
      "000000" when "0001100000111011", -- t[6203] = 0
      "000000" when "0001100000111100", -- t[6204] = 0
      "000000" when "0001100000111101", -- t[6205] = 0
      "000000" when "0001100000111110", -- t[6206] = 0
      "000000" when "0001100000111111", -- t[6207] = 0
      "000000" when "0001100001000000", -- t[6208] = 0
      "000000" when "0001100001000001", -- t[6209] = 0
      "000000" when "0001100001000010", -- t[6210] = 0
      "000000" when "0001100001000011", -- t[6211] = 0
      "000000" when "0001100001000100", -- t[6212] = 0
      "000000" when "0001100001000101", -- t[6213] = 0
      "000000" when "0001100001000110", -- t[6214] = 0
      "000000" when "0001100001000111", -- t[6215] = 0
      "000000" when "0001100001001000", -- t[6216] = 0
      "000000" when "0001100001001001", -- t[6217] = 0
      "000000" when "0001100001001010", -- t[6218] = 0
      "000000" when "0001100001001011", -- t[6219] = 0
      "000000" when "0001100001001100", -- t[6220] = 0
      "000000" when "0001100001001101", -- t[6221] = 0
      "000000" when "0001100001001110", -- t[6222] = 0
      "000000" when "0001100001001111", -- t[6223] = 0
      "000000" when "0001100001010000", -- t[6224] = 0
      "000000" when "0001100001010001", -- t[6225] = 0
      "000000" when "0001100001010010", -- t[6226] = 0
      "000000" when "0001100001010011", -- t[6227] = 0
      "000000" when "0001100001010100", -- t[6228] = 0
      "000000" when "0001100001010101", -- t[6229] = 0
      "000000" when "0001100001010110", -- t[6230] = 0
      "000000" when "0001100001010111", -- t[6231] = 0
      "000000" when "0001100001011000", -- t[6232] = 0
      "000000" when "0001100001011001", -- t[6233] = 0
      "000000" when "0001100001011010", -- t[6234] = 0
      "000000" when "0001100001011011", -- t[6235] = 0
      "000000" when "0001100001011100", -- t[6236] = 0
      "000000" when "0001100001011101", -- t[6237] = 0
      "000000" when "0001100001011110", -- t[6238] = 0
      "000000" when "0001100001011111", -- t[6239] = 0
      "000000" when "0001100001100000", -- t[6240] = 0
      "000000" when "0001100001100001", -- t[6241] = 0
      "000000" when "0001100001100010", -- t[6242] = 0
      "000000" when "0001100001100011", -- t[6243] = 0
      "000000" when "0001100001100100", -- t[6244] = 0
      "000000" when "0001100001100101", -- t[6245] = 0
      "000000" when "0001100001100110", -- t[6246] = 0
      "000000" when "0001100001100111", -- t[6247] = 0
      "000000" when "0001100001101000", -- t[6248] = 0
      "000000" when "0001100001101001", -- t[6249] = 0
      "000000" when "0001100001101010", -- t[6250] = 0
      "000000" when "0001100001101011", -- t[6251] = 0
      "000000" when "0001100001101100", -- t[6252] = 0
      "000000" when "0001100001101101", -- t[6253] = 0
      "000000" when "0001100001101110", -- t[6254] = 0
      "000000" when "0001100001101111", -- t[6255] = 0
      "000000" when "0001100001110000", -- t[6256] = 0
      "000000" when "0001100001110001", -- t[6257] = 0
      "000000" when "0001100001110010", -- t[6258] = 0
      "000000" when "0001100001110011", -- t[6259] = 0
      "000000" when "0001100001110100", -- t[6260] = 0
      "000000" when "0001100001110101", -- t[6261] = 0
      "000000" when "0001100001110110", -- t[6262] = 0
      "000000" when "0001100001110111", -- t[6263] = 0
      "000000" when "0001100001111000", -- t[6264] = 0
      "000000" when "0001100001111001", -- t[6265] = 0
      "000000" when "0001100001111010", -- t[6266] = 0
      "000000" when "0001100001111011", -- t[6267] = 0
      "000000" when "0001100001111100", -- t[6268] = 0
      "000000" when "0001100001111101", -- t[6269] = 0
      "000000" when "0001100001111110", -- t[6270] = 0
      "000000" when "0001100001111111", -- t[6271] = 0
      "000000" when "0001100010000000", -- t[6272] = 0
      "000000" when "0001100010000001", -- t[6273] = 0
      "000000" when "0001100010000010", -- t[6274] = 0
      "000000" when "0001100010000011", -- t[6275] = 0
      "000000" when "0001100010000100", -- t[6276] = 0
      "000000" when "0001100010000101", -- t[6277] = 0
      "000000" when "0001100010000110", -- t[6278] = 0
      "000000" when "0001100010000111", -- t[6279] = 0
      "000000" when "0001100010001000", -- t[6280] = 0
      "000000" when "0001100010001001", -- t[6281] = 0
      "000000" when "0001100010001010", -- t[6282] = 0
      "000000" when "0001100010001011", -- t[6283] = 0
      "000000" when "0001100010001100", -- t[6284] = 0
      "000000" when "0001100010001101", -- t[6285] = 0
      "000000" when "0001100010001110", -- t[6286] = 0
      "000000" when "0001100010001111", -- t[6287] = 0
      "000000" when "0001100010010000", -- t[6288] = 0
      "000000" when "0001100010010001", -- t[6289] = 0
      "000000" when "0001100010010010", -- t[6290] = 0
      "000000" when "0001100010010011", -- t[6291] = 0
      "000000" when "0001100010010100", -- t[6292] = 0
      "000000" when "0001100010010101", -- t[6293] = 0
      "000000" when "0001100010010110", -- t[6294] = 0
      "000000" when "0001100010010111", -- t[6295] = 0
      "000000" when "0001100010011000", -- t[6296] = 0
      "000000" when "0001100010011001", -- t[6297] = 0
      "000000" when "0001100010011010", -- t[6298] = 0
      "000000" when "0001100010011011", -- t[6299] = 0
      "000000" when "0001100010011100", -- t[6300] = 0
      "000000" when "0001100010011101", -- t[6301] = 0
      "000000" when "0001100010011110", -- t[6302] = 0
      "000000" when "0001100010011111", -- t[6303] = 0
      "000000" when "0001100010100000", -- t[6304] = 0
      "000000" when "0001100010100001", -- t[6305] = 0
      "000000" when "0001100010100010", -- t[6306] = 0
      "000000" when "0001100010100011", -- t[6307] = 0
      "000000" when "0001100010100100", -- t[6308] = 0
      "000000" when "0001100010100101", -- t[6309] = 0
      "000000" when "0001100010100110", -- t[6310] = 0
      "000000" when "0001100010100111", -- t[6311] = 0
      "000000" when "0001100010101000", -- t[6312] = 0
      "000000" when "0001100010101001", -- t[6313] = 0
      "000000" when "0001100010101010", -- t[6314] = 0
      "000000" when "0001100010101011", -- t[6315] = 0
      "000000" when "0001100010101100", -- t[6316] = 0
      "000000" when "0001100010101101", -- t[6317] = 0
      "000000" when "0001100010101110", -- t[6318] = 0
      "000000" when "0001100010101111", -- t[6319] = 0
      "000000" when "0001100010110000", -- t[6320] = 0
      "000000" when "0001100010110001", -- t[6321] = 0
      "000000" when "0001100010110010", -- t[6322] = 0
      "000000" when "0001100010110011", -- t[6323] = 0
      "000000" when "0001100010110100", -- t[6324] = 0
      "000000" when "0001100010110101", -- t[6325] = 0
      "000000" when "0001100010110110", -- t[6326] = 0
      "000000" when "0001100010110111", -- t[6327] = 0
      "000000" when "0001100010111000", -- t[6328] = 0
      "000000" when "0001100010111001", -- t[6329] = 0
      "000000" when "0001100010111010", -- t[6330] = 0
      "000000" when "0001100010111011", -- t[6331] = 0
      "000000" when "0001100010111100", -- t[6332] = 0
      "000000" when "0001100010111101", -- t[6333] = 0
      "000000" when "0001100010111110", -- t[6334] = 0
      "000000" when "0001100010111111", -- t[6335] = 0
      "000000" when "0001100011000000", -- t[6336] = 0
      "000000" when "0001100011000001", -- t[6337] = 0
      "000000" when "0001100011000010", -- t[6338] = 0
      "000000" when "0001100011000011", -- t[6339] = 0
      "000000" when "0001100011000100", -- t[6340] = 0
      "000000" when "0001100011000101", -- t[6341] = 0
      "000000" when "0001100011000110", -- t[6342] = 0
      "000000" when "0001100011000111", -- t[6343] = 0
      "000000" when "0001100011001000", -- t[6344] = 0
      "000000" when "0001100011001001", -- t[6345] = 0
      "000000" when "0001100011001010", -- t[6346] = 0
      "000000" when "0001100011001011", -- t[6347] = 0
      "000000" when "0001100011001100", -- t[6348] = 0
      "000000" when "0001100011001101", -- t[6349] = 0
      "000000" when "0001100011001110", -- t[6350] = 0
      "000000" when "0001100011001111", -- t[6351] = 0
      "000000" when "0001100011010000", -- t[6352] = 0
      "000000" when "0001100011010001", -- t[6353] = 0
      "000000" when "0001100011010010", -- t[6354] = 0
      "000000" when "0001100011010011", -- t[6355] = 0
      "000000" when "0001100011010100", -- t[6356] = 0
      "000000" when "0001100011010101", -- t[6357] = 0
      "000000" when "0001100011010110", -- t[6358] = 0
      "000000" when "0001100011010111", -- t[6359] = 0
      "000000" when "0001100011011000", -- t[6360] = 0
      "000000" when "0001100011011001", -- t[6361] = 0
      "000000" when "0001100011011010", -- t[6362] = 0
      "000000" when "0001100011011011", -- t[6363] = 0
      "000000" when "0001100011011100", -- t[6364] = 0
      "000000" when "0001100011011101", -- t[6365] = 0
      "000000" when "0001100011011110", -- t[6366] = 0
      "000000" when "0001100011011111", -- t[6367] = 0
      "000000" when "0001100011100000", -- t[6368] = 0
      "000000" when "0001100011100001", -- t[6369] = 0
      "000000" when "0001100011100010", -- t[6370] = 0
      "000000" when "0001100011100011", -- t[6371] = 0
      "000000" when "0001100011100100", -- t[6372] = 0
      "000000" when "0001100011100101", -- t[6373] = 0
      "000000" when "0001100011100110", -- t[6374] = 0
      "000000" when "0001100011100111", -- t[6375] = 0
      "000000" when "0001100011101000", -- t[6376] = 0
      "000000" when "0001100011101001", -- t[6377] = 0
      "000000" when "0001100011101010", -- t[6378] = 0
      "000000" when "0001100011101011", -- t[6379] = 0
      "000000" when "0001100011101100", -- t[6380] = 0
      "000000" when "0001100011101101", -- t[6381] = 0
      "000000" when "0001100011101110", -- t[6382] = 0
      "000000" when "0001100011101111", -- t[6383] = 0
      "000000" when "0001100011110000", -- t[6384] = 0
      "000000" when "0001100011110001", -- t[6385] = 0
      "000000" when "0001100011110010", -- t[6386] = 0
      "000000" when "0001100011110011", -- t[6387] = 0
      "000000" when "0001100011110100", -- t[6388] = 0
      "000000" when "0001100011110101", -- t[6389] = 0
      "000000" when "0001100011110110", -- t[6390] = 0
      "000000" when "0001100011110111", -- t[6391] = 0
      "000000" when "0001100011111000", -- t[6392] = 0
      "000000" when "0001100011111001", -- t[6393] = 0
      "000000" when "0001100011111010", -- t[6394] = 0
      "000000" when "0001100011111011", -- t[6395] = 0
      "000000" when "0001100011111100", -- t[6396] = 0
      "000000" when "0001100011111101", -- t[6397] = 0
      "000000" when "0001100011111110", -- t[6398] = 0
      "000000" when "0001100011111111", -- t[6399] = 0
      "000000" when "0001100100000000", -- t[6400] = 0
      "000000" when "0001100100000001", -- t[6401] = 0
      "000000" when "0001100100000010", -- t[6402] = 0
      "000000" when "0001100100000011", -- t[6403] = 0
      "000000" when "0001100100000100", -- t[6404] = 0
      "000000" when "0001100100000101", -- t[6405] = 0
      "000000" when "0001100100000110", -- t[6406] = 0
      "000000" when "0001100100000111", -- t[6407] = 0
      "000000" when "0001100100001000", -- t[6408] = 0
      "000000" when "0001100100001001", -- t[6409] = 0
      "000000" when "0001100100001010", -- t[6410] = 0
      "000000" when "0001100100001011", -- t[6411] = 0
      "000000" when "0001100100001100", -- t[6412] = 0
      "000000" when "0001100100001101", -- t[6413] = 0
      "000000" when "0001100100001110", -- t[6414] = 0
      "000000" when "0001100100001111", -- t[6415] = 0
      "000000" when "0001100100010000", -- t[6416] = 0
      "000000" when "0001100100010001", -- t[6417] = 0
      "000000" when "0001100100010010", -- t[6418] = 0
      "000000" when "0001100100010011", -- t[6419] = 0
      "000000" when "0001100100010100", -- t[6420] = 0
      "000000" when "0001100100010101", -- t[6421] = 0
      "000000" when "0001100100010110", -- t[6422] = 0
      "000000" when "0001100100010111", -- t[6423] = 0
      "000000" when "0001100100011000", -- t[6424] = 0
      "000000" when "0001100100011001", -- t[6425] = 0
      "000000" when "0001100100011010", -- t[6426] = 0
      "000000" when "0001100100011011", -- t[6427] = 0
      "000000" when "0001100100011100", -- t[6428] = 0
      "000000" when "0001100100011101", -- t[6429] = 0
      "000000" when "0001100100011110", -- t[6430] = 0
      "000000" when "0001100100011111", -- t[6431] = 0
      "000000" when "0001100100100000", -- t[6432] = 0
      "000000" when "0001100100100001", -- t[6433] = 0
      "000000" when "0001100100100010", -- t[6434] = 0
      "000000" when "0001100100100011", -- t[6435] = 0
      "000000" when "0001100100100100", -- t[6436] = 0
      "000000" when "0001100100100101", -- t[6437] = 0
      "000000" when "0001100100100110", -- t[6438] = 0
      "000000" when "0001100100100111", -- t[6439] = 0
      "000000" when "0001100100101000", -- t[6440] = 0
      "000000" when "0001100100101001", -- t[6441] = 0
      "000000" when "0001100100101010", -- t[6442] = 0
      "000000" when "0001100100101011", -- t[6443] = 0
      "000000" when "0001100100101100", -- t[6444] = 0
      "000000" when "0001100100101101", -- t[6445] = 0
      "000000" when "0001100100101110", -- t[6446] = 0
      "000000" when "0001100100101111", -- t[6447] = 0
      "000000" when "0001100100110000", -- t[6448] = 0
      "000000" when "0001100100110001", -- t[6449] = 0
      "000000" when "0001100100110010", -- t[6450] = 0
      "000000" when "0001100100110011", -- t[6451] = 0
      "000000" when "0001100100110100", -- t[6452] = 0
      "000000" when "0001100100110101", -- t[6453] = 0
      "000000" when "0001100100110110", -- t[6454] = 0
      "000000" when "0001100100110111", -- t[6455] = 0
      "000000" when "0001100100111000", -- t[6456] = 0
      "000000" when "0001100100111001", -- t[6457] = 0
      "000000" when "0001100100111010", -- t[6458] = 0
      "000000" when "0001100100111011", -- t[6459] = 0
      "000000" when "0001100100111100", -- t[6460] = 0
      "000000" when "0001100100111101", -- t[6461] = 0
      "000000" when "0001100100111110", -- t[6462] = 0
      "000000" when "0001100100111111", -- t[6463] = 0
      "000000" when "0001100101000000", -- t[6464] = 0
      "000000" when "0001100101000001", -- t[6465] = 0
      "000000" when "0001100101000010", -- t[6466] = 0
      "000000" when "0001100101000011", -- t[6467] = 0
      "000000" when "0001100101000100", -- t[6468] = 0
      "000000" when "0001100101000101", -- t[6469] = 0
      "000000" when "0001100101000110", -- t[6470] = 0
      "000000" when "0001100101000111", -- t[6471] = 0
      "000000" when "0001100101001000", -- t[6472] = 0
      "000000" when "0001100101001001", -- t[6473] = 0
      "000000" when "0001100101001010", -- t[6474] = 0
      "000000" when "0001100101001011", -- t[6475] = 0
      "000000" when "0001100101001100", -- t[6476] = 0
      "000000" when "0001100101001101", -- t[6477] = 0
      "000000" when "0001100101001110", -- t[6478] = 0
      "000000" when "0001100101001111", -- t[6479] = 0
      "000000" when "0001100101010000", -- t[6480] = 0
      "000000" when "0001100101010001", -- t[6481] = 0
      "000000" when "0001100101010010", -- t[6482] = 0
      "000000" when "0001100101010011", -- t[6483] = 0
      "000000" when "0001100101010100", -- t[6484] = 0
      "000000" when "0001100101010101", -- t[6485] = 0
      "000000" when "0001100101010110", -- t[6486] = 0
      "000000" when "0001100101010111", -- t[6487] = 0
      "000000" when "0001100101011000", -- t[6488] = 0
      "000000" when "0001100101011001", -- t[6489] = 0
      "000000" when "0001100101011010", -- t[6490] = 0
      "000000" when "0001100101011011", -- t[6491] = 0
      "000000" when "0001100101011100", -- t[6492] = 0
      "000000" when "0001100101011101", -- t[6493] = 0
      "000000" when "0001100101011110", -- t[6494] = 0
      "000000" when "0001100101011111", -- t[6495] = 0
      "000000" when "0001100101100000", -- t[6496] = 0
      "000000" when "0001100101100001", -- t[6497] = 0
      "000000" when "0001100101100010", -- t[6498] = 0
      "000000" when "0001100101100011", -- t[6499] = 0
      "000000" when "0001100101100100", -- t[6500] = 0
      "000000" when "0001100101100101", -- t[6501] = 0
      "000000" when "0001100101100110", -- t[6502] = 0
      "000000" when "0001100101100111", -- t[6503] = 0
      "000000" when "0001100101101000", -- t[6504] = 0
      "000000" when "0001100101101001", -- t[6505] = 0
      "000000" when "0001100101101010", -- t[6506] = 0
      "000000" when "0001100101101011", -- t[6507] = 0
      "000000" when "0001100101101100", -- t[6508] = 0
      "000000" when "0001100101101101", -- t[6509] = 0
      "000000" when "0001100101101110", -- t[6510] = 0
      "000000" when "0001100101101111", -- t[6511] = 0
      "000000" when "0001100101110000", -- t[6512] = 0
      "000000" when "0001100101110001", -- t[6513] = 0
      "000000" when "0001100101110010", -- t[6514] = 0
      "000000" when "0001100101110011", -- t[6515] = 0
      "000000" when "0001100101110100", -- t[6516] = 0
      "000000" when "0001100101110101", -- t[6517] = 0
      "000000" when "0001100101110110", -- t[6518] = 0
      "000000" when "0001100101110111", -- t[6519] = 0
      "000000" when "0001100101111000", -- t[6520] = 0
      "000000" when "0001100101111001", -- t[6521] = 0
      "000000" when "0001100101111010", -- t[6522] = 0
      "000000" when "0001100101111011", -- t[6523] = 0
      "000000" when "0001100101111100", -- t[6524] = 0
      "000000" when "0001100101111101", -- t[6525] = 0
      "000000" when "0001100101111110", -- t[6526] = 0
      "000000" when "0001100101111111", -- t[6527] = 0
      "000000" when "0001100110000000", -- t[6528] = 0
      "000000" when "0001100110000001", -- t[6529] = 0
      "000000" when "0001100110000010", -- t[6530] = 0
      "000000" when "0001100110000011", -- t[6531] = 0
      "000000" when "0001100110000100", -- t[6532] = 0
      "000000" when "0001100110000101", -- t[6533] = 0
      "000000" when "0001100110000110", -- t[6534] = 0
      "000000" when "0001100110000111", -- t[6535] = 0
      "000000" when "0001100110001000", -- t[6536] = 0
      "000000" when "0001100110001001", -- t[6537] = 0
      "000000" when "0001100110001010", -- t[6538] = 0
      "000000" when "0001100110001011", -- t[6539] = 0
      "000000" when "0001100110001100", -- t[6540] = 0
      "000000" when "0001100110001101", -- t[6541] = 0
      "000000" when "0001100110001110", -- t[6542] = 0
      "000000" when "0001100110001111", -- t[6543] = 0
      "000000" when "0001100110010000", -- t[6544] = 0
      "000000" when "0001100110010001", -- t[6545] = 0
      "000000" when "0001100110010010", -- t[6546] = 0
      "000000" when "0001100110010011", -- t[6547] = 0
      "000000" when "0001100110010100", -- t[6548] = 0
      "000000" when "0001100110010101", -- t[6549] = 0
      "000000" when "0001100110010110", -- t[6550] = 0
      "000000" when "0001100110010111", -- t[6551] = 0
      "000000" when "0001100110011000", -- t[6552] = 0
      "000000" when "0001100110011001", -- t[6553] = 0
      "000000" when "0001100110011010", -- t[6554] = 0
      "000000" when "0001100110011011", -- t[6555] = 0
      "000000" when "0001100110011100", -- t[6556] = 0
      "000000" when "0001100110011101", -- t[6557] = 0
      "000000" when "0001100110011110", -- t[6558] = 0
      "000000" when "0001100110011111", -- t[6559] = 0
      "000000" when "0001100110100000", -- t[6560] = 0
      "000000" when "0001100110100001", -- t[6561] = 0
      "000000" when "0001100110100010", -- t[6562] = 0
      "000000" when "0001100110100011", -- t[6563] = 0
      "000000" when "0001100110100100", -- t[6564] = 0
      "000000" when "0001100110100101", -- t[6565] = 0
      "000000" when "0001100110100110", -- t[6566] = 0
      "000000" when "0001100110100111", -- t[6567] = 0
      "000000" when "0001100110101000", -- t[6568] = 0
      "000000" when "0001100110101001", -- t[6569] = 0
      "000000" when "0001100110101010", -- t[6570] = 0
      "000000" when "0001100110101011", -- t[6571] = 0
      "000000" when "0001100110101100", -- t[6572] = 0
      "000000" when "0001100110101101", -- t[6573] = 0
      "000000" when "0001100110101110", -- t[6574] = 0
      "000000" when "0001100110101111", -- t[6575] = 0
      "000000" when "0001100110110000", -- t[6576] = 0
      "000000" when "0001100110110001", -- t[6577] = 0
      "000000" when "0001100110110010", -- t[6578] = 0
      "000000" when "0001100110110011", -- t[6579] = 0
      "000000" when "0001100110110100", -- t[6580] = 0
      "000000" when "0001100110110101", -- t[6581] = 0
      "000000" when "0001100110110110", -- t[6582] = 0
      "000000" when "0001100110110111", -- t[6583] = 0
      "000000" when "0001100110111000", -- t[6584] = 0
      "000000" when "0001100110111001", -- t[6585] = 0
      "000000" when "0001100110111010", -- t[6586] = 0
      "000000" when "0001100110111011", -- t[6587] = 0
      "000000" when "0001100110111100", -- t[6588] = 0
      "000000" when "0001100110111101", -- t[6589] = 0
      "000000" when "0001100110111110", -- t[6590] = 0
      "000000" when "0001100110111111", -- t[6591] = 0
      "000000" when "0001100111000000", -- t[6592] = 0
      "000000" when "0001100111000001", -- t[6593] = 0
      "000000" when "0001100111000010", -- t[6594] = 0
      "000000" when "0001100111000011", -- t[6595] = 0
      "000000" when "0001100111000100", -- t[6596] = 0
      "000000" when "0001100111000101", -- t[6597] = 0
      "000000" when "0001100111000110", -- t[6598] = 0
      "000000" when "0001100111000111", -- t[6599] = 0
      "000000" when "0001100111001000", -- t[6600] = 0
      "000000" when "0001100111001001", -- t[6601] = 0
      "000000" when "0001100111001010", -- t[6602] = 0
      "000000" when "0001100111001011", -- t[6603] = 0
      "000000" when "0001100111001100", -- t[6604] = 0
      "000000" when "0001100111001101", -- t[6605] = 0
      "000000" when "0001100111001110", -- t[6606] = 0
      "000000" when "0001100111001111", -- t[6607] = 0
      "000000" when "0001100111010000", -- t[6608] = 0
      "000000" when "0001100111010001", -- t[6609] = 0
      "000000" when "0001100111010010", -- t[6610] = 0
      "000000" when "0001100111010011", -- t[6611] = 0
      "000000" when "0001100111010100", -- t[6612] = 0
      "000000" when "0001100111010101", -- t[6613] = 0
      "000000" when "0001100111010110", -- t[6614] = 0
      "000000" when "0001100111010111", -- t[6615] = 0
      "000000" when "0001100111011000", -- t[6616] = 0
      "000000" when "0001100111011001", -- t[6617] = 0
      "000000" when "0001100111011010", -- t[6618] = 0
      "000000" when "0001100111011011", -- t[6619] = 0
      "000000" when "0001100111011100", -- t[6620] = 0
      "000000" when "0001100111011101", -- t[6621] = 0
      "000000" when "0001100111011110", -- t[6622] = 0
      "000000" when "0001100111011111", -- t[6623] = 0
      "000000" when "0001100111100000", -- t[6624] = 0
      "000000" when "0001100111100001", -- t[6625] = 0
      "000000" when "0001100111100010", -- t[6626] = 0
      "000000" when "0001100111100011", -- t[6627] = 0
      "000000" when "0001100111100100", -- t[6628] = 0
      "000000" when "0001100111100101", -- t[6629] = 0
      "000000" when "0001100111100110", -- t[6630] = 0
      "000000" when "0001100111100111", -- t[6631] = 0
      "000000" when "0001100111101000", -- t[6632] = 0
      "000000" when "0001100111101001", -- t[6633] = 0
      "000000" when "0001100111101010", -- t[6634] = 0
      "000000" when "0001100111101011", -- t[6635] = 0
      "000000" when "0001100111101100", -- t[6636] = 0
      "000000" when "0001100111101101", -- t[6637] = 0
      "000000" when "0001100111101110", -- t[6638] = 0
      "000000" when "0001100111101111", -- t[6639] = 0
      "000000" when "0001100111110000", -- t[6640] = 0
      "000000" when "0001100111110001", -- t[6641] = 0
      "000000" when "0001100111110010", -- t[6642] = 0
      "000000" when "0001100111110011", -- t[6643] = 0
      "000000" when "0001100111110100", -- t[6644] = 0
      "000000" when "0001100111110101", -- t[6645] = 0
      "000000" when "0001100111110110", -- t[6646] = 0
      "000000" when "0001100111110111", -- t[6647] = 0
      "000000" when "0001100111111000", -- t[6648] = 0
      "000000" when "0001100111111001", -- t[6649] = 0
      "000000" when "0001100111111010", -- t[6650] = 0
      "000000" when "0001100111111011", -- t[6651] = 0
      "000000" when "0001100111111100", -- t[6652] = 0
      "000000" when "0001100111111101", -- t[6653] = 0
      "000000" when "0001100111111110", -- t[6654] = 0
      "000000" when "0001100111111111", -- t[6655] = 0
      "000000" when "0001101000000000", -- t[6656] = 0
      "000000" when "0001101000000001", -- t[6657] = 0
      "000000" when "0001101000000010", -- t[6658] = 0
      "000000" when "0001101000000011", -- t[6659] = 0
      "000000" when "0001101000000100", -- t[6660] = 0
      "000000" when "0001101000000101", -- t[6661] = 0
      "000000" when "0001101000000110", -- t[6662] = 0
      "000000" when "0001101000000111", -- t[6663] = 0
      "000000" when "0001101000001000", -- t[6664] = 0
      "000000" when "0001101000001001", -- t[6665] = 0
      "000000" when "0001101000001010", -- t[6666] = 0
      "000000" when "0001101000001011", -- t[6667] = 0
      "000000" when "0001101000001100", -- t[6668] = 0
      "000000" when "0001101000001101", -- t[6669] = 0
      "000000" when "0001101000001110", -- t[6670] = 0
      "000000" when "0001101000001111", -- t[6671] = 0
      "000000" when "0001101000010000", -- t[6672] = 0
      "000000" when "0001101000010001", -- t[6673] = 0
      "000000" when "0001101000010010", -- t[6674] = 0
      "000000" when "0001101000010011", -- t[6675] = 0
      "000000" when "0001101000010100", -- t[6676] = 0
      "000000" when "0001101000010101", -- t[6677] = 0
      "000000" when "0001101000010110", -- t[6678] = 0
      "000000" when "0001101000010111", -- t[6679] = 0
      "000000" when "0001101000011000", -- t[6680] = 0
      "000000" when "0001101000011001", -- t[6681] = 0
      "000000" when "0001101000011010", -- t[6682] = 0
      "000000" when "0001101000011011", -- t[6683] = 0
      "000000" when "0001101000011100", -- t[6684] = 0
      "000000" when "0001101000011101", -- t[6685] = 0
      "000000" when "0001101000011110", -- t[6686] = 0
      "000000" when "0001101000011111", -- t[6687] = 0
      "000000" when "0001101000100000", -- t[6688] = 0
      "000000" when "0001101000100001", -- t[6689] = 0
      "000000" when "0001101000100010", -- t[6690] = 0
      "000000" when "0001101000100011", -- t[6691] = 0
      "000000" when "0001101000100100", -- t[6692] = 0
      "000000" when "0001101000100101", -- t[6693] = 0
      "000000" when "0001101000100110", -- t[6694] = 0
      "000000" when "0001101000100111", -- t[6695] = 0
      "000000" when "0001101000101000", -- t[6696] = 0
      "000000" when "0001101000101001", -- t[6697] = 0
      "000000" when "0001101000101010", -- t[6698] = 0
      "000000" when "0001101000101011", -- t[6699] = 0
      "000000" when "0001101000101100", -- t[6700] = 0
      "000000" when "0001101000101101", -- t[6701] = 0
      "000000" when "0001101000101110", -- t[6702] = 0
      "000000" when "0001101000101111", -- t[6703] = 0
      "000000" when "0001101000110000", -- t[6704] = 0
      "000000" when "0001101000110001", -- t[6705] = 0
      "000000" when "0001101000110010", -- t[6706] = 0
      "000000" when "0001101000110011", -- t[6707] = 0
      "000000" when "0001101000110100", -- t[6708] = 0
      "000000" when "0001101000110101", -- t[6709] = 0
      "000000" when "0001101000110110", -- t[6710] = 0
      "000000" when "0001101000110111", -- t[6711] = 0
      "000000" when "0001101000111000", -- t[6712] = 0
      "000000" when "0001101000111001", -- t[6713] = 0
      "000000" when "0001101000111010", -- t[6714] = 0
      "000000" when "0001101000111011", -- t[6715] = 0
      "000000" when "0001101000111100", -- t[6716] = 0
      "000000" when "0001101000111101", -- t[6717] = 0
      "000000" when "0001101000111110", -- t[6718] = 0
      "000000" when "0001101000111111", -- t[6719] = 0
      "000000" when "0001101001000000", -- t[6720] = 0
      "000000" when "0001101001000001", -- t[6721] = 0
      "000000" when "0001101001000010", -- t[6722] = 0
      "000000" when "0001101001000011", -- t[6723] = 0
      "000000" when "0001101001000100", -- t[6724] = 0
      "000000" when "0001101001000101", -- t[6725] = 0
      "000000" when "0001101001000110", -- t[6726] = 0
      "000000" when "0001101001000111", -- t[6727] = 0
      "000000" when "0001101001001000", -- t[6728] = 0
      "000000" when "0001101001001001", -- t[6729] = 0
      "000000" when "0001101001001010", -- t[6730] = 0
      "000000" when "0001101001001011", -- t[6731] = 0
      "000000" when "0001101001001100", -- t[6732] = 0
      "000000" when "0001101001001101", -- t[6733] = 0
      "000000" when "0001101001001110", -- t[6734] = 0
      "000000" when "0001101001001111", -- t[6735] = 0
      "000000" when "0001101001010000", -- t[6736] = 0
      "000000" when "0001101001010001", -- t[6737] = 0
      "000000" when "0001101001010010", -- t[6738] = 0
      "000000" when "0001101001010011", -- t[6739] = 0
      "000000" when "0001101001010100", -- t[6740] = 0
      "000000" when "0001101001010101", -- t[6741] = 0
      "000000" when "0001101001010110", -- t[6742] = 0
      "000000" when "0001101001010111", -- t[6743] = 0
      "000000" when "0001101001011000", -- t[6744] = 0
      "000000" when "0001101001011001", -- t[6745] = 0
      "000000" when "0001101001011010", -- t[6746] = 0
      "000000" when "0001101001011011", -- t[6747] = 0
      "000000" when "0001101001011100", -- t[6748] = 0
      "000000" when "0001101001011101", -- t[6749] = 0
      "000000" when "0001101001011110", -- t[6750] = 0
      "000000" when "0001101001011111", -- t[6751] = 0
      "000000" when "0001101001100000", -- t[6752] = 0
      "000000" when "0001101001100001", -- t[6753] = 0
      "000000" when "0001101001100010", -- t[6754] = 0
      "000000" when "0001101001100011", -- t[6755] = 0
      "000000" when "0001101001100100", -- t[6756] = 0
      "000000" when "0001101001100101", -- t[6757] = 0
      "000000" when "0001101001100110", -- t[6758] = 0
      "000000" when "0001101001100111", -- t[6759] = 0
      "000000" when "0001101001101000", -- t[6760] = 0
      "000000" when "0001101001101001", -- t[6761] = 0
      "000000" when "0001101001101010", -- t[6762] = 0
      "000000" when "0001101001101011", -- t[6763] = 0
      "000000" when "0001101001101100", -- t[6764] = 0
      "000000" when "0001101001101101", -- t[6765] = 0
      "000000" when "0001101001101110", -- t[6766] = 0
      "000000" when "0001101001101111", -- t[6767] = 0
      "000000" when "0001101001110000", -- t[6768] = 0
      "000000" when "0001101001110001", -- t[6769] = 0
      "000000" when "0001101001110010", -- t[6770] = 0
      "000000" when "0001101001110011", -- t[6771] = 0
      "000000" when "0001101001110100", -- t[6772] = 0
      "000000" when "0001101001110101", -- t[6773] = 0
      "000000" when "0001101001110110", -- t[6774] = 0
      "000000" when "0001101001110111", -- t[6775] = 0
      "000000" when "0001101001111000", -- t[6776] = 0
      "000000" when "0001101001111001", -- t[6777] = 0
      "000000" when "0001101001111010", -- t[6778] = 0
      "000000" when "0001101001111011", -- t[6779] = 0
      "000000" when "0001101001111100", -- t[6780] = 0
      "000000" when "0001101001111101", -- t[6781] = 0
      "000000" when "0001101001111110", -- t[6782] = 0
      "000000" when "0001101001111111", -- t[6783] = 0
      "000000" when "0001101010000000", -- t[6784] = 0
      "000000" when "0001101010000001", -- t[6785] = 0
      "000000" when "0001101010000010", -- t[6786] = 0
      "000000" when "0001101010000011", -- t[6787] = 0
      "000000" when "0001101010000100", -- t[6788] = 0
      "000000" when "0001101010000101", -- t[6789] = 0
      "000000" when "0001101010000110", -- t[6790] = 0
      "000000" when "0001101010000111", -- t[6791] = 0
      "000000" when "0001101010001000", -- t[6792] = 0
      "000000" when "0001101010001001", -- t[6793] = 0
      "000000" when "0001101010001010", -- t[6794] = 0
      "000000" when "0001101010001011", -- t[6795] = 0
      "000000" when "0001101010001100", -- t[6796] = 0
      "000000" when "0001101010001101", -- t[6797] = 0
      "000000" when "0001101010001110", -- t[6798] = 0
      "000000" when "0001101010001111", -- t[6799] = 0
      "000000" when "0001101010010000", -- t[6800] = 0
      "000000" when "0001101010010001", -- t[6801] = 0
      "000000" when "0001101010010010", -- t[6802] = 0
      "000000" when "0001101010010011", -- t[6803] = 0
      "000000" when "0001101010010100", -- t[6804] = 0
      "000000" when "0001101010010101", -- t[6805] = 0
      "000000" when "0001101010010110", -- t[6806] = 0
      "000000" when "0001101010010111", -- t[6807] = 0
      "000000" when "0001101010011000", -- t[6808] = 0
      "000000" when "0001101010011001", -- t[6809] = 0
      "000000" when "0001101010011010", -- t[6810] = 0
      "000000" when "0001101010011011", -- t[6811] = 0
      "000000" when "0001101010011100", -- t[6812] = 0
      "000000" when "0001101010011101", -- t[6813] = 0
      "000000" when "0001101010011110", -- t[6814] = 0
      "000000" when "0001101010011111", -- t[6815] = 0
      "000000" when "0001101010100000", -- t[6816] = 0
      "000000" when "0001101010100001", -- t[6817] = 0
      "000000" when "0001101010100010", -- t[6818] = 0
      "000000" when "0001101010100011", -- t[6819] = 0
      "000000" when "0001101010100100", -- t[6820] = 0
      "000000" when "0001101010100101", -- t[6821] = 0
      "000000" when "0001101010100110", -- t[6822] = 0
      "000000" when "0001101010100111", -- t[6823] = 0
      "000000" when "0001101010101000", -- t[6824] = 0
      "000000" when "0001101010101001", -- t[6825] = 0
      "000000" when "0001101010101010", -- t[6826] = 0
      "000000" when "0001101010101011", -- t[6827] = 0
      "000000" when "0001101010101100", -- t[6828] = 0
      "000000" when "0001101010101101", -- t[6829] = 0
      "000000" when "0001101010101110", -- t[6830] = 0
      "000000" when "0001101010101111", -- t[6831] = 0
      "000000" when "0001101010110000", -- t[6832] = 0
      "000000" when "0001101010110001", -- t[6833] = 0
      "000000" when "0001101010110010", -- t[6834] = 0
      "000000" when "0001101010110011", -- t[6835] = 0
      "000000" when "0001101010110100", -- t[6836] = 0
      "000000" when "0001101010110101", -- t[6837] = 0
      "000000" when "0001101010110110", -- t[6838] = 0
      "000000" when "0001101010110111", -- t[6839] = 0
      "000000" when "0001101010111000", -- t[6840] = 0
      "000000" when "0001101010111001", -- t[6841] = 0
      "000000" when "0001101010111010", -- t[6842] = 0
      "000000" when "0001101010111011", -- t[6843] = 0
      "000000" when "0001101010111100", -- t[6844] = 0
      "000000" when "0001101010111101", -- t[6845] = 0
      "000000" when "0001101010111110", -- t[6846] = 0
      "000000" when "0001101010111111", -- t[6847] = 0
      "000000" when "0001101011000000", -- t[6848] = 0
      "000000" when "0001101011000001", -- t[6849] = 0
      "000000" when "0001101011000010", -- t[6850] = 0
      "000000" when "0001101011000011", -- t[6851] = 0
      "000000" when "0001101011000100", -- t[6852] = 0
      "000000" when "0001101011000101", -- t[6853] = 0
      "000000" when "0001101011000110", -- t[6854] = 0
      "000000" when "0001101011000111", -- t[6855] = 0
      "000000" when "0001101011001000", -- t[6856] = 0
      "000000" when "0001101011001001", -- t[6857] = 0
      "000000" when "0001101011001010", -- t[6858] = 0
      "000000" when "0001101011001011", -- t[6859] = 0
      "000000" when "0001101011001100", -- t[6860] = 0
      "000000" when "0001101011001101", -- t[6861] = 0
      "000000" when "0001101011001110", -- t[6862] = 0
      "000000" when "0001101011001111", -- t[6863] = 0
      "000000" when "0001101011010000", -- t[6864] = 0
      "000000" when "0001101011010001", -- t[6865] = 0
      "000000" when "0001101011010010", -- t[6866] = 0
      "000000" when "0001101011010011", -- t[6867] = 0
      "000000" when "0001101011010100", -- t[6868] = 0
      "000000" when "0001101011010101", -- t[6869] = 0
      "000000" when "0001101011010110", -- t[6870] = 0
      "000000" when "0001101011010111", -- t[6871] = 0
      "000000" when "0001101011011000", -- t[6872] = 0
      "000000" when "0001101011011001", -- t[6873] = 0
      "000000" when "0001101011011010", -- t[6874] = 0
      "000000" when "0001101011011011", -- t[6875] = 0
      "000000" when "0001101011011100", -- t[6876] = 0
      "000000" when "0001101011011101", -- t[6877] = 0
      "000000" when "0001101011011110", -- t[6878] = 0
      "000000" when "0001101011011111", -- t[6879] = 0
      "000000" when "0001101011100000", -- t[6880] = 0
      "000000" when "0001101011100001", -- t[6881] = 0
      "000000" when "0001101011100010", -- t[6882] = 0
      "000000" when "0001101011100011", -- t[6883] = 0
      "000000" when "0001101011100100", -- t[6884] = 0
      "000000" when "0001101011100101", -- t[6885] = 0
      "000000" when "0001101011100110", -- t[6886] = 0
      "000000" when "0001101011100111", -- t[6887] = 0
      "000000" when "0001101011101000", -- t[6888] = 0
      "000000" when "0001101011101001", -- t[6889] = 0
      "000000" when "0001101011101010", -- t[6890] = 0
      "000000" when "0001101011101011", -- t[6891] = 0
      "000000" when "0001101011101100", -- t[6892] = 0
      "000000" when "0001101011101101", -- t[6893] = 0
      "000000" when "0001101011101110", -- t[6894] = 0
      "000000" when "0001101011101111", -- t[6895] = 0
      "000000" when "0001101011110000", -- t[6896] = 0
      "000000" when "0001101011110001", -- t[6897] = 0
      "000000" when "0001101011110010", -- t[6898] = 0
      "000000" when "0001101011110011", -- t[6899] = 0
      "000000" when "0001101011110100", -- t[6900] = 0
      "000000" when "0001101011110101", -- t[6901] = 0
      "000000" when "0001101011110110", -- t[6902] = 0
      "000000" when "0001101011110111", -- t[6903] = 0
      "000000" when "0001101011111000", -- t[6904] = 0
      "000000" when "0001101011111001", -- t[6905] = 0
      "000000" when "0001101011111010", -- t[6906] = 0
      "000000" when "0001101011111011", -- t[6907] = 0
      "000000" when "0001101011111100", -- t[6908] = 0
      "000000" when "0001101011111101", -- t[6909] = 0
      "000000" when "0001101011111110", -- t[6910] = 0
      "000000" when "0001101011111111", -- t[6911] = 0
      "000000" when "0001101100000000", -- t[6912] = 0
      "000000" when "0001101100000001", -- t[6913] = 0
      "000000" when "0001101100000010", -- t[6914] = 0
      "000000" when "0001101100000011", -- t[6915] = 0
      "000000" when "0001101100000100", -- t[6916] = 0
      "000000" when "0001101100000101", -- t[6917] = 0
      "000000" when "0001101100000110", -- t[6918] = 0
      "000000" when "0001101100000111", -- t[6919] = 0
      "000000" when "0001101100001000", -- t[6920] = 0
      "000000" when "0001101100001001", -- t[6921] = 0
      "000000" when "0001101100001010", -- t[6922] = 0
      "000000" when "0001101100001011", -- t[6923] = 0
      "000000" when "0001101100001100", -- t[6924] = 0
      "000000" when "0001101100001101", -- t[6925] = 0
      "000000" when "0001101100001110", -- t[6926] = 0
      "000000" when "0001101100001111", -- t[6927] = 0
      "000000" when "0001101100010000", -- t[6928] = 0
      "000000" when "0001101100010001", -- t[6929] = 0
      "000000" when "0001101100010010", -- t[6930] = 0
      "000000" when "0001101100010011", -- t[6931] = 0
      "000000" when "0001101100010100", -- t[6932] = 0
      "000000" when "0001101100010101", -- t[6933] = 0
      "000000" when "0001101100010110", -- t[6934] = 0
      "000000" when "0001101100010111", -- t[6935] = 0
      "000000" when "0001101100011000", -- t[6936] = 0
      "000000" when "0001101100011001", -- t[6937] = 0
      "000000" when "0001101100011010", -- t[6938] = 0
      "000000" when "0001101100011011", -- t[6939] = 0
      "000000" when "0001101100011100", -- t[6940] = 0
      "000000" when "0001101100011101", -- t[6941] = 0
      "000000" when "0001101100011110", -- t[6942] = 0
      "000000" when "0001101100011111", -- t[6943] = 0
      "000000" when "0001101100100000", -- t[6944] = 0
      "000000" when "0001101100100001", -- t[6945] = 0
      "000000" when "0001101100100010", -- t[6946] = 0
      "000000" when "0001101100100011", -- t[6947] = 0
      "000000" when "0001101100100100", -- t[6948] = 0
      "000000" when "0001101100100101", -- t[6949] = 0
      "000000" when "0001101100100110", -- t[6950] = 0
      "000000" when "0001101100100111", -- t[6951] = 0
      "000000" when "0001101100101000", -- t[6952] = 0
      "000000" when "0001101100101001", -- t[6953] = 0
      "000000" when "0001101100101010", -- t[6954] = 0
      "000000" when "0001101100101011", -- t[6955] = 0
      "000000" when "0001101100101100", -- t[6956] = 0
      "000000" when "0001101100101101", -- t[6957] = 0
      "000000" when "0001101100101110", -- t[6958] = 0
      "000000" when "0001101100101111", -- t[6959] = 0
      "000000" when "0001101100110000", -- t[6960] = 0
      "000000" when "0001101100110001", -- t[6961] = 0
      "000000" when "0001101100110010", -- t[6962] = 0
      "000000" when "0001101100110011", -- t[6963] = 0
      "000000" when "0001101100110100", -- t[6964] = 0
      "000000" when "0001101100110101", -- t[6965] = 0
      "000000" when "0001101100110110", -- t[6966] = 0
      "000000" when "0001101100110111", -- t[6967] = 0
      "000000" when "0001101100111000", -- t[6968] = 0
      "000000" when "0001101100111001", -- t[6969] = 0
      "000000" when "0001101100111010", -- t[6970] = 0
      "000000" when "0001101100111011", -- t[6971] = 0
      "000000" when "0001101100111100", -- t[6972] = 0
      "000000" when "0001101100111101", -- t[6973] = 0
      "000000" when "0001101100111110", -- t[6974] = 0
      "000000" when "0001101100111111", -- t[6975] = 0
      "000000" when "0001101101000000", -- t[6976] = 0
      "000000" when "0001101101000001", -- t[6977] = 0
      "000000" when "0001101101000010", -- t[6978] = 0
      "000000" when "0001101101000011", -- t[6979] = 0
      "000000" when "0001101101000100", -- t[6980] = 0
      "000000" when "0001101101000101", -- t[6981] = 0
      "000000" when "0001101101000110", -- t[6982] = 0
      "000000" when "0001101101000111", -- t[6983] = 0
      "000000" when "0001101101001000", -- t[6984] = 0
      "000000" when "0001101101001001", -- t[6985] = 0
      "000000" when "0001101101001010", -- t[6986] = 0
      "000000" when "0001101101001011", -- t[6987] = 0
      "000000" when "0001101101001100", -- t[6988] = 0
      "000000" when "0001101101001101", -- t[6989] = 0
      "000000" when "0001101101001110", -- t[6990] = 0
      "000000" when "0001101101001111", -- t[6991] = 0
      "000000" when "0001101101010000", -- t[6992] = 0
      "000000" when "0001101101010001", -- t[6993] = 0
      "000000" when "0001101101010010", -- t[6994] = 0
      "000000" when "0001101101010011", -- t[6995] = 0
      "000000" when "0001101101010100", -- t[6996] = 0
      "000000" when "0001101101010101", -- t[6997] = 0
      "000000" when "0001101101010110", -- t[6998] = 0
      "000000" when "0001101101010111", -- t[6999] = 0
      "000000" when "0001101101011000", -- t[7000] = 0
      "000000" when "0001101101011001", -- t[7001] = 0
      "000000" when "0001101101011010", -- t[7002] = 0
      "000000" when "0001101101011011", -- t[7003] = 0
      "000000" when "0001101101011100", -- t[7004] = 0
      "000000" when "0001101101011101", -- t[7005] = 0
      "000000" when "0001101101011110", -- t[7006] = 0
      "000000" when "0001101101011111", -- t[7007] = 0
      "000000" when "0001101101100000", -- t[7008] = 0
      "000000" when "0001101101100001", -- t[7009] = 0
      "000000" when "0001101101100010", -- t[7010] = 0
      "000000" when "0001101101100011", -- t[7011] = 0
      "000000" when "0001101101100100", -- t[7012] = 0
      "000000" when "0001101101100101", -- t[7013] = 0
      "000000" when "0001101101100110", -- t[7014] = 0
      "000000" when "0001101101100111", -- t[7015] = 0
      "000000" when "0001101101101000", -- t[7016] = 0
      "000000" when "0001101101101001", -- t[7017] = 0
      "000000" when "0001101101101010", -- t[7018] = 0
      "000000" when "0001101101101011", -- t[7019] = 0
      "000000" when "0001101101101100", -- t[7020] = 0
      "000000" when "0001101101101101", -- t[7021] = 0
      "000000" when "0001101101101110", -- t[7022] = 0
      "000000" when "0001101101101111", -- t[7023] = 0
      "000000" when "0001101101110000", -- t[7024] = 0
      "000000" when "0001101101110001", -- t[7025] = 0
      "000000" when "0001101101110010", -- t[7026] = 0
      "000000" when "0001101101110011", -- t[7027] = 0
      "000000" when "0001101101110100", -- t[7028] = 0
      "000000" when "0001101101110101", -- t[7029] = 0
      "000000" when "0001101101110110", -- t[7030] = 0
      "000000" when "0001101101110111", -- t[7031] = 0
      "000000" when "0001101101111000", -- t[7032] = 0
      "000000" when "0001101101111001", -- t[7033] = 0
      "000000" when "0001101101111010", -- t[7034] = 0
      "000000" when "0001101101111011", -- t[7035] = 0
      "000000" when "0001101101111100", -- t[7036] = 0
      "000000" when "0001101101111101", -- t[7037] = 0
      "000000" when "0001101101111110", -- t[7038] = 0
      "000000" when "0001101101111111", -- t[7039] = 0
      "000000" when "0001101110000000", -- t[7040] = 0
      "000000" when "0001101110000001", -- t[7041] = 0
      "000000" when "0001101110000010", -- t[7042] = 0
      "000000" when "0001101110000011", -- t[7043] = 0
      "000000" when "0001101110000100", -- t[7044] = 0
      "000000" when "0001101110000101", -- t[7045] = 0
      "000000" when "0001101110000110", -- t[7046] = 0
      "000000" when "0001101110000111", -- t[7047] = 0
      "000000" when "0001101110001000", -- t[7048] = 0
      "000000" when "0001101110001001", -- t[7049] = 0
      "000000" when "0001101110001010", -- t[7050] = 0
      "000000" when "0001101110001011", -- t[7051] = 0
      "000000" when "0001101110001100", -- t[7052] = 0
      "000000" when "0001101110001101", -- t[7053] = 0
      "000000" when "0001101110001110", -- t[7054] = 0
      "000000" when "0001101110001111", -- t[7055] = 0
      "000000" when "0001101110010000", -- t[7056] = 0
      "000000" when "0001101110010001", -- t[7057] = 0
      "000000" when "0001101110010010", -- t[7058] = 0
      "000000" when "0001101110010011", -- t[7059] = 0
      "000000" when "0001101110010100", -- t[7060] = 0
      "000000" when "0001101110010101", -- t[7061] = 0
      "000000" when "0001101110010110", -- t[7062] = 0
      "000000" when "0001101110010111", -- t[7063] = 0
      "000000" when "0001101110011000", -- t[7064] = 0
      "000000" when "0001101110011001", -- t[7065] = 0
      "000000" when "0001101110011010", -- t[7066] = 0
      "000000" when "0001101110011011", -- t[7067] = 0
      "000000" when "0001101110011100", -- t[7068] = 0
      "000000" when "0001101110011101", -- t[7069] = 0
      "000000" when "0001101110011110", -- t[7070] = 0
      "000000" when "0001101110011111", -- t[7071] = 0
      "000000" when "0001101110100000", -- t[7072] = 0
      "000000" when "0001101110100001", -- t[7073] = 0
      "000000" when "0001101110100010", -- t[7074] = 0
      "000000" when "0001101110100011", -- t[7075] = 0
      "000000" when "0001101110100100", -- t[7076] = 0
      "000000" when "0001101110100101", -- t[7077] = 0
      "000000" when "0001101110100110", -- t[7078] = 0
      "000000" when "0001101110100111", -- t[7079] = 0
      "000000" when "0001101110101000", -- t[7080] = 0
      "000000" when "0001101110101001", -- t[7081] = 0
      "000000" when "0001101110101010", -- t[7082] = 0
      "000000" when "0001101110101011", -- t[7083] = 0
      "000000" when "0001101110101100", -- t[7084] = 0
      "000000" when "0001101110101101", -- t[7085] = 0
      "000000" when "0001101110101110", -- t[7086] = 0
      "000000" when "0001101110101111", -- t[7087] = 0
      "000000" when "0001101110110000", -- t[7088] = 0
      "000000" when "0001101110110001", -- t[7089] = 0
      "000000" when "0001101110110010", -- t[7090] = 0
      "000000" when "0001101110110011", -- t[7091] = 0
      "000000" when "0001101110110100", -- t[7092] = 0
      "000000" when "0001101110110101", -- t[7093] = 0
      "000000" when "0001101110110110", -- t[7094] = 0
      "000000" when "0001101110110111", -- t[7095] = 0
      "000000" when "0001101110111000", -- t[7096] = 0
      "000000" when "0001101110111001", -- t[7097] = 0
      "000000" when "0001101110111010", -- t[7098] = 0
      "000000" when "0001101110111011", -- t[7099] = 0
      "000000" when "0001101110111100", -- t[7100] = 0
      "000000" when "0001101110111101", -- t[7101] = 0
      "000000" when "0001101110111110", -- t[7102] = 0
      "000000" when "0001101110111111", -- t[7103] = 0
      "000000" when "0001101111000000", -- t[7104] = 0
      "000000" when "0001101111000001", -- t[7105] = 0
      "000000" when "0001101111000010", -- t[7106] = 0
      "000000" when "0001101111000011", -- t[7107] = 0
      "000000" when "0001101111000100", -- t[7108] = 0
      "000000" when "0001101111000101", -- t[7109] = 0
      "000000" when "0001101111000110", -- t[7110] = 0
      "000000" when "0001101111000111", -- t[7111] = 0
      "000000" when "0001101111001000", -- t[7112] = 0
      "000000" when "0001101111001001", -- t[7113] = 0
      "000000" when "0001101111001010", -- t[7114] = 0
      "000000" when "0001101111001011", -- t[7115] = 0
      "000000" when "0001101111001100", -- t[7116] = 0
      "000000" when "0001101111001101", -- t[7117] = 0
      "000000" when "0001101111001110", -- t[7118] = 0
      "000000" when "0001101111001111", -- t[7119] = 0
      "000000" when "0001101111010000", -- t[7120] = 0
      "000000" when "0001101111010001", -- t[7121] = 0
      "000000" when "0001101111010010", -- t[7122] = 0
      "000000" when "0001101111010011", -- t[7123] = 0
      "000000" when "0001101111010100", -- t[7124] = 0
      "000000" when "0001101111010101", -- t[7125] = 0
      "000000" when "0001101111010110", -- t[7126] = 0
      "000000" when "0001101111010111", -- t[7127] = 0
      "000000" when "0001101111011000", -- t[7128] = 0
      "000000" when "0001101111011001", -- t[7129] = 0
      "000000" when "0001101111011010", -- t[7130] = 0
      "000000" when "0001101111011011", -- t[7131] = 0
      "000000" when "0001101111011100", -- t[7132] = 0
      "000000" when "0001101111011101", -- t[7133] = 0
      "000000" when "0001101111011110", -- t[7134] = 0
      "000000" when "0001101111011111", -- t[7135] = 0
      "000000" when "0001101111100000", -- t[7136] = 0
      "000000" when "0001101111100001", -- t[7137] = 0
      "000000" when "0001101111100010", -- t[7138] = 0
      "000000" when "0001101111100011", -- t[7139] = 0
      "000000" when "0001101111100100", -- t[7140] = 0
      "000000" when "0001101111100101", -- t[7141] = 0
      "000000" when "0001101111100110", -- t[7142] = 0
      "000000" when "0001101111100111", -- t[7143] = 0
      "000000" when "0001101111101000", -- t[7144] = 0
      "000000" when "0001101111101001", -- t[7145] = 0
      "000000" when "0001101111101010", -- t[7146] = 0
      "000000" when "0001101111101011", -- t[7147] = 0
      "000000" when "0001101111101100", -- t[7148] = 0
      "000000" when "0001101111101101", -- t[7149] = 0
      "000000" when "0001101111101110", -- t[7150] = 0
      "000000" when "0001101111101111", -- t[7151] = 0
      "000000" when "0001101111110000", -- t[7152] = 0
      "000000" when "0001101111110001", -- t[7153] = 0
      "000000" when "0001101111110010", -- t[7154] = 0
      "000000" when "0001101111110011", -- t[7155] = 0
      "000000" when "0001101111110100", -- t[7156] = 0
      "000000" when "0001101111110101", -- t[7157] = 0
      "000000" when "0001101111110110", -- t[7158] = 0
      "000000" when "0001101111110111", -- t[7159] = 0
      "000000" when "0001101111111000", -- t[7160] = 0
      "000000" when "0001101111111001", -- t[7161] = 0
      "000000" when "0001101111111010", -- t[7162] = 0
      "000000" when "0001101111111011", -- t[7163] = 0
      "000000" when "0001101111111100", -- t[7164] = 0
      "000000" when "0001101111111101", -- t[7165] = 0
      "000000" when "0001101111111110", -- t[7166] = 0
      "000000" when "0001101111111111", -- t[7167] = 0
      "000000" when "0001110000000000", -- t[7168] = 0
      "000000" when "0001110000000001", -- t[7169] = 0
      "000000" when "0001110000000010", -- t[7170] = 0
      "000000" when "0001110000000011", -- t[7171] = 0
      "000000" when "0001110000000100", -- t[7172] = 0
      "000000" when "0001110000000101", -- t[7173] = 0
      "000000" when "0001110000000110", -- t[7174] = 0
      "000000" when "0001110000000111", -- t[7175] = 0
      "000000" when "0001110000001000", -- t[7176] = 0
      "000000" when "0001110000001001", -- t[7177] = 0
      "000000" when "0001110000001010", -- t[7178] = 0
      "000000" when "0001110000001011", -- t[7179] = 0
      "000000" when "0001110000001100", -- t[7180] = 0
      "000000" when "0001110000001101", -- t[7181] = 0
      "000000" when "0001110000001110", -- t[7182] = 0
      "000000" when "0001110000001111", -- t[7183] = 0
      "000000" when "0001110000010000", -- t[7184] = 0
      "000000" when "0001110000010001", -- t[7185] = 0
      "000000" when "0001110000010010", -- t[7186] = 0
      "000000" when "0001110000010011", -- t[7187] = 0
      "000000" when "0001110000010100", -- t[7188] = 0
      "000000" when "0001110000010101", -- t[7189] = 0
      "000000" when "0001110000010110", -- t[7190] = 0
      "000000" when "0001110000010111", -- t[7191] = 0
      "000000" when "0001110000011000", -- t[7192] = 0
      "000000" when "0001110000011001", -- t[7193] = 0
      "000000" when "0001110000011010", -- t[7194] = 0
      "000000" when "0001110000011011", -- t[7195] = 0
      "000000" when "0001110000011100", -- t[7196] = 0
      "000000" when "0001110000011101", -- t[7197] = 0
      "000000" when "0001110000011110", -- t[7198] = 0
      "000000" when "0001110000011111", -- t[7199] = 0
      "000000" when "0001110000100000", -- t[7200] = 0
      "000000" when "0001110000100001", -- t[7201] = 0
      "000000" when "0001110000100010", -- t[7202] = 0
      "000000" when "0001110000100011", -- t[7203] = 0
      "000000" when "0001110000100100", -- t[7204] = 0
      "000000" when "0001110000100101", -- t[7205] = 0
      "000000" when "0001110000100110", -- t[7206] = 0
      "000000" when "0001110000100111", -- t[7207] = 0
      "000000" when "0001110000101000", -- t[7208] = 0
      "000000" when "0001110000101001", -- t[7209] = 0
      "000000" when "0001110000101010", -- t[7210] = 0
      "000000" when "0001110000101011", -- t[7211] = 0
      "000000" when "0001110000101100", -- t[7212] = 0
      "000000" when "0001110000101101", -- t[7213] = 0
      "000000" when "0001110000101110", -- t[7214] = 0
      "000000" when "0001110000101111", -- t[7215] = 0
      "000000" when "0001110000110000", -- t[7216] = 0
      "000000" when "0001110000110001", -- t[7217] = 0
      "000000" when "0001110000110010", -- t[7218] = 0
      "000000" when "0001110000110011", -- t[7219] = 0
      "000000" when "0001110000110100", -- t[7220] = 0
      "000000" when "0001110000110101", -- t[7221] = 0
      "000000" when "0001110000110110", -- t[7222] = 0
      "000000" when "0001110000110111", -- t[7223] = 0
      "000000" when "0001110000111000", -- t[7224] = 0
      "000000" when "0001110000111001", -- t[7225] = 0
      "000000" when "0001110000111010", -- t[7226] = 0
      "000000" when "0001110000111011", -- t[7227] = 0
      "000000" when "0001110000111100", -- t[7228] = 0
      "000000" when "0001110000111101", -- t[7229] = 0
      "000000" when "0001110000111110", -- t[7230] = 0
      "000000" when "0001110000111111", -- t[7231] = 0
      "000000" when "0001110001000000", -- t[7232] = 0
      "000000" when "0001110001000001", -- t[7233] = 0
      "000000" when "0001110001000010", -- t[7234] = 0
      "000000" when "0001110001000011", -- t[7235] = 0
      "000000" when "0001110001000100", -- t[7236] = 0
      "000000" when "0001110001000101", -- t[7237] = 0
      "000000" when "0001110001000110", -- t[7238] = 0
      "000000" when "0001110001000111", -- t[7239] = 0
      "000000" when "0001110001001000", -- t[7240] = 0
      "000000" when "0001110001001001", -- t[7241] = 0
      "000000" when "0001110001001010", -- t[7242] = 0
      "000000" when "0001110001001011", -- t[7243] = 0
      "000000" when "0001110001001100", -- t[7244] = 0
      "000000" when "0001110001001101", -- t[7245] = 0
      "000000" when "0001110001001110", -- t[7246] = 0
      "000000" when "0001110001001111", -- t[7247] = 0
      "000000" when "0001110001010000", -- t[7248] = 0
      "000000" when "0001110001010001", -- t[7249] = 0
      "000000" when "0001110001010010", -- t[7250] = 0
      "000000" when "0001110001010011", -- t[7251] = 0
      "000000" when "0001110001010100", -- t[7252] = 0
      "000000" when "0001110001010101", -- t[7253] = 0
      "000000" when "0001110001010110", -- t[7254] = 0
      "000000" when "0001110001010111", -- t[7255] = 0
      "000000" when "0001110001011000", -- t[7256] = 0
      "000000" when "0001110001011001", -- t[7257] = 0
      "000000" when "0001110001011010", -- t[7258] = 0
      "000000" when "0001110001011011", -- t[7259] = 0
      "000000" when "0001110001011100", -- t[7260] = 0
      "000000" when "0001110001011101", -- t[7261] = 0
      "000000" when "0001110001011110", -- t[7262] = 0
      "000000" when "0001110001011111", -- t[7263] = 0
      "000000" when "0001110001100000", -- t[7264] = 0
      "000000" when "0001110001100001", -- t[7265] = 0
      "000000" when "0001110001100010", -- t[7266] = 0
      "000000" when "0001110001100011", -- t[7267] = 0
      "000000" when "0001110001100100", -- t[7268] = 0
      "000000" when "0001110001100101", -- t[7269] = 0
      "000000" when "0001110001100110", -- t[7270] = 0
      "000000" when "0001110001100111", -- t[7271] = 0
      "000000" when "0001110001101000", -- t[7272] = 0
      "000000" when "0001110001101001", -- t[7273] = 0
      "000000" when "0001110001101010", -- t[7274] = 0
      "000000" when "0001110001101011", -- t[7275] = 0
      "000000" when "0001110001101100", -- t[7276] = 0
      "000000" when "0001110001101101", -- t[7277] = 0
      "000000" when "0001110001101110", -- t[7278] = 0
      "000000" when "0001110001101111", -- t[7279] = 0
      "000000" when "0001110001110000", -- t[7280] = 0
      "000000" when "0001110001110001", -- t[7281] = 0
      "000000" when "0001110001110010", -- t[7282] = 0
      "000000" when "0001110001110011", -- t[7283] = 0
      "000000" when "0001110001110100", -- t[7284] = 0
      "000000" when "0001110001110101", -- t[7285] = 0
      "000000" when "0001110001110110", -- t[7286] = 0
      "000000" when "0001110001110111", -- t[7287] = 0
      "000000" when "0001110001111000", -- t[7288] = 0
      "000000" when "0001110001111001", -- t[7289] = 0
      "000000" when "0001110001111010", -- t[7290] = 0
      "000000" when "0001110001111011", -- t[7291] = 0
      "000000" when "0001110001111100", -- t[7292] = 0
      "000000" when "0001110001111101", -- t[7293] = 0
      "000000" when "0001110001111110", -- t[7294] = 0
      "000000" when "0001110001111111", -- t[7295] = 0
      "000000" when "0001110010000000", -- t[7296] = 0
      "000000" when "0001110010000001", -- t[7297] = 0
      "000000" when "0001110010000010", -- t[7298] = 0
      "000000" when "0001110010000011", -- t[7299] = 0
      "000000" when "0001110010000100", -- t[7300] = 0
      "000000" when "0001110010000101", -- t[7301] = 0
      "000000" when "0001110010000110", -- t[7302] = 0
      "000000" when "0001110010000111", -- t[7303] = 0
      "000000" when "0001110010001000", -- t[7304] = 0
      "000000" when "0001110010001001", -- t[7305] = 0
      "000000" when "0001110010001010", -- t[7306] = 0
      "000000" when "0001110010001011", -- t[7307] = 0
      "000000" when "0001110010001100", -- t[7308] = 0
      "000000" when "0001110010001101", -- t[7309] = 0
      "000000" when "0001110010001110", -- t[7310] = 0
      "000000" when "0001110010001111", -- t[7311] = 0
      "000000" when "0001110010010000", -- t[7312] = 0
      "000000" when "0001110010010001", -- t[7313] = 0
      "000000" when "0001110010010010", -- t[7314] = 0
      "000000" when "0001110010010011", -- t[7315] = 0
      "000000" when "0001110010010100", -- t[7316] = 0
      "000000" when "0001110010010101", -- t[7317] = 0
      "000000" when "0001110010010110", -- t[7318] = 0
      "000000" when "0001110010010111", -- t[7319] = 0
      "000000" when "0001110010011000", -- t[7320] = 0
      "000000" when "0001110010011001", -- t[7321] = 0
      "000000" when "0001110010011010", -- t[7322] = 0
      "000000" when "0001110010011011", -- t[7323] = 0
      "000000" when "0001110010011100", -- t[7324] = 0
      "000000" when "0001110010011101", -- t[7325] = 0
      "000000" when "0001110010011110", -- t[7326] = 0
      "000000" when "0001110010011111", -- t[7327] = 0
      "000000" when "0001110010100000", -- t[7328] = 0
      "000000" when "0001110010100001", -- t[7329] = 0
      "000000" when "0001110010100010", -- t[7330] = 0
      "000000" when "0001110010100011", -- t[7331] = 0
      "000000" when "0001110010100100", -- t[7332] = 0
      "000000" when "0001110010100101", -- t[7333] = 0
      "000000" when "0001110010100110", -- t[7334] = 0
      "000000" when "0001110010100111", -- t[7335] = 0
      "000000" when "0001110010101000", -- t[7336] = 0
      "000000" when "0001110010101001", -- t[7337] = 0
      "000000" when "0001110010101010", -- t[7338] = 0
      "000000" when "0001110010101011", -- t[7339] = 0
      "000000" when "0001110010101100", -- t[7340] = 0
      "000000" when "0001110010101101", -- t[7341] = 0
      "000000" when "0001110010101110", -- t[7342] = 0
      "000000" when "0001110010101111", -- t[7343] = 0
      "000000" when "0001110010110000", -- t[7344] = 0
      "000000" when "0001110010110001", -- t[7345] = 0
      "000000" when "0001110010110010", -- t[7346] = 0
      "000000" when "0001110010110011", -- t[7347] = 0
      "000000" when "0001110010110100", -- t[7348] = 0
      "000000" when "0001110010110101", -- t[7349] = 0
      "000000" when "0001110010110110", -- t[7350] = 0
      "000000" when "0001110010110111", -- t[7351] = 0
      "000000" when "0001110010111000", -- t[7352] = 0
      "000000" when "0001110010111001", -- t[7353] = 0
      "000000" when "0001110010111010", -- t[7354] = 0
      "000000" when "0001110010111011", -- t[7355] = 0
      "000000" when "0001110010111100", -- t[7356] = 0
      "000000" when "0001110010111101", -- t[7357] = 0
      "000000" when "0001110010111110", -- t[7358] = 0
      "000000" when "0001110010111111", -- t[7359] = 0
      "000000" when "0001110011000000", -- t[7360] = 0
      "000000" when "0001110011000001", -- t[7361] = 0
      "000000" when "0001110011000010", -- t[7362] = 0
      "000000" when "0001110011000011", -- t[7363] = 0
      "000000" when "0001110011000100", -- t[7364] = 0
      "000000" when "0001110011000101", -- t[7365] = 0
      "000000" when "0001110011000110", -- t[7366] = 0
      "000000" when "0001110011000111", -- t[7367] = 0
      "000000" when "0001110011001000", -- t[7368] = 0
      "000000" when "0001110011001001", -- t[7369] = 0
      "000000" when "0001110011001010", -- t[7370] = 0
      "000000" when "0001110011001011", -- t[7371] = 0
      "000000" when "0001110011001100", -- t[7372] = 0
      "000000" when "0001110011001101", -- t[7373] = 0
      "000000" when "0001110011001110", -- t[7374] = 0
      "000000" when "0001110011001111", -- t[7375] = 0
      "000000" when "0001110011010000", -- t[7376] = 0
      "000000" when "0001110011010001", -- t[7377] = 0
      "000000" when "0001110011010010", -- t[7378] = 0
      "000000" when "0001110011010011", -- t[7379] = 0
      "000000" when "0001110011010100", -- t[7380] = 0
      "000000" when "0001110011010101", -- t[7381] = 0
      "000000" when "0001110011010110", -- t[7382] = 0
      "000000" when "0001110011010111", -- t[7383] = 0
      "000000" when "0001110011011000", -- t[7384] = 0
      "000000" when "0001110011011001", -- t[7385] = 0
      "000000" when "0001110011011010", -- t[7386] = 0
      "000000" when "0001110011011011", -- t[7387] = 0
      "000000" when "0001110011011100", -- t[7388] = 0
      "000000" when "0001110011011101", -- t[7389] = 0
      "000000" when "0001110011011110", -- t[7390] = 0
      "000000" when "0001110011011111", -- t[7391] = 0
      "000000" when "0001110011100000", -- t[7392] = 0
      "000000" when "0001110011100001", -- t[7393] = 0
      "000000" when "0001110011100010", -- t[7394] = 0
      "000000" when "0001110011100011", -- t[7395] = 0
      "000000" when "0001110011100100", -- t[7396] = 0
      "000000" when "0001110011100101", -- t[7397] = 0
      "000000" when "0001110011100110", -- t[7398] = 0
      "000000" when "0001110011100111", -- t[7399] = 0
      "000000" when "0001110011101000", -- t[7400] = 0
      "000000" when "0001110011101001", -- t[7401] = 0
      "000000" when "0001110011101010", -- t[7402] = 0
      "000000" when "0001110011101011", -- t[7403] = 0
      "000000" when "0001110011101100", -- t[7404] = 0
      "000000" when "0001110011101101", -- t[7405] = 0
      "000000" when "0001110011101110", -- t[7406] = 0
      "000000" when "0001110011101111", -- t[7407] = 0
      "000000" when "0001110011110000", -- t[7408] = 0
      "000000" when "0001110011110001", -- t[7409] = 0
      "000000" when "0001110011110010", -- t[7410] = 0
      "000000" when "0001110011110011", -- t[7411] = 0
      "000000" when "0001110011110100", -- t[7412] = 0
      "000000" when "0001110011110101", -- t[7413] = 0
      "000000" when "0001110011110110", -- t[7414] = 0
      "000000" when "0001110011110111", -- t[7415] = 0
      "000000" when "0001110011111000", -- t[7416] = 0
      "000000" when "0001110011111001", -- t[7417] = 0
      "000000" when "0001110011111010", -- t[7418] = 0
      "000000" when "0001110011111011", -- t[7419] = 0
      "000000" when "0001110011111100", -- t[7420] = 0
      "000000" when "0001110011111101", -- t[7421] = 0
      "000000" when "0001110011111110", -- t[7422] = 0
      "000000" when "0001110011111111", -- t[7423] = 0
      "000000" when "0001110100000000", -- t[7424] = 0
      "000000" when "0001110100000001", -- t[7425] = 0
      "000000" when "0001110100000010", -- t[7426] = 0
      "000000" when "0001110100000011", -- t[7427] = 0
      "000000" when "0001110100000100", -- t[7428] = 0
      "000000" when "0001110100000101", -- t[7429] = 0
      "000000" when "0001110100000110", -- t[7430] = 0
      "000000" when "0001110100000111", -- t[7431] = 0
      "000000" when "0001110100001000", -- t[7432] = 0
      "000000" when "0001110100001001", -- t[7433] = 0
      "000000" when "0001110100001010", -- t[7434] = 0
      "000000" when "0001110100001011", -- t[7435] = 0
      "000000" when "0001110100001100", -- t[7436] = 0
      "000000" when "0001110100001101", -- t[7437] = 0
      "000000" when "0001110100001110", -- t[7438] = 0
      "000000" when "0001110100001111", -- t[7439] = 0
      "000000" when "0001110100010000", -- t[7440] = 0
      "000000" when "0001110100010001", -- t[7441] = 0
      "000000" when "0001110100010010", -- t[7442] = 0
      "000000" when "0001110100010011", -- t[7443] = 0
      "000000" when "0001110100010100", -- t[7444] = 0
      "000000" when "0001110100010101", -- t[7445] = 0
      "000000" when "0001110100010110", -- t[7446] = 0
      "000000" when "0001110100010111", -- t[7447] = 0
      "000000" when "0001110100011000", -- t[7448] = 0
      "000000" when "0001110100011001", -- t[7449] = 0
      "000000" when "0001110100011010", -- t[7450] = 0
      "000000" when "0001110100011011", -- t[7451] = 0
      "000000" when "0001110100011100", -- t[7452] = 0
      "000000" when "0001110100011101", -- t[7453] = 0
      "000000" when "0001110100011110", -- t[7454] = 0
      "000000" when "0001110100011111", -- t[7455] = 0
      "000000" when "0001110100100000", -- t[7456] = 0
      "000000" when "0001110100100001", -- t[7457] = 0
      "000000" when "0001110100100010", -- t[7458] = 0
      "000000" when "0001110100100011", -- t[7459] = 0
      "000000" when "0001110100100100", -- t[7460] = 0
      "000000" when "0001110100100101", -- t[7461] = 0
      "000000" when "0001110100100110", -- t[7462] = 0
      "000000" when "0001110100100111", -- t[7463] = 0
      "000000" when "0001110100101000", -- t[7464] = 0
      "000000" when "0001110100101001", -- t[7465] = 0
      "000000" when "0001110100101010", -- t[7466] = 0
      "000000" when "0001110100101011", -- t[7467] = 0
      "000000" when "0001110100101100", -- t[7468] = 0
      "000000" when "0001110100101101", -- t[7469] = 0
      "000000" when "0001110100101110", -- t[7470] = 0
      "000000" when "0001110100101111", -- t[7471] = 0
      "000000" when "0001110100110000", -- t[7472] = 0
      "000000" when "0001110100110001", -- t[7473] = 0
      "000000" when "0001110100110010", -- t[7474] = 0
      "000000" when "0001110100110011", -- t[7475] = 0
      "000000" when "0001110100110100", -- t[7476] = 0
      "000000" when "0001110100110101", -- t[7477] = 0
      "000000" when "0001110100110110", -- t[7478] = 0
      "000000" when "0001110100110111", -- t[7479] = 0
      "000000" when "0001110100111000", -- t[7480] = 0
      "000000" when "0001110100111001", -- t[7481] = 0
      "000000" when "0001110100111010", -- t[7482] = 0
      "000000" when "0001110100111011", -- t[7483] = 0
      "000000" when "0001110100111100", -- t[7484] = 0
      "000000" when "0001110100111101", -- t[7485] = 0
      "000000" when "0001110100111110", -- t[7486] = 0
      "000000" when "0001110100111111", -- t[7487] = 0
      "000000" when "0001110101000000", -- t[7488] = 0
      "000000" when "0001110101000001", -- t[7489] = 0
      "000000" when "0001110101000010", -- t[7490] = 0
      "000000" when "0001110101000011", -- t[7491] = 0
      "000000" when "0001110101000100", -- t[7492] = 0
      "000000" when "0001110101000101", -- t[7493] = 0
      "000000" when "0001110101000110", -- t[7494] = 0
      "000000" when "0001110101000111", -- t[7495] = 0
      "000000" when "0001110101001000", -- t[7496] = 0
      "000000" when "0001110101001001", -- t[7497] = 0
      "000000" when "0001110101001010", -- t[7498] = 0
      "000000" when "0001110101001011", -- t[7499] = 0
      "000000" when "0001110101001100", -- t[7500] = 0
      "000000" when "0001110101001101", -- t[7501] = 0
      "000000" when "0001110101001110", -- t[7502] = 0
      "000000" when "0001110101001111", -- t[7503] = 0
      "000000" when "0001110101010000", -- t[7504] = 0
      "000000" when "0001110101010001", -- t[7505] = 0
      "000000" when "0001110101010010", -- t[7506] = 0
      "000000" when "0001110101010011", -- t[7507] = 0
      "000000" when "0001110101010100", -- t[7508] = 0
      "000000" when "0001110101010101", -- t[7509] = 0
      "000000" when "0001110101010110", -- t[7510] = 0
      "000000" when "0001110101010111", -- t[7511] = 0
      "000000" when "0001110101011000", -- t[7512] = 0
      "000000" when "0001110101011001", -- t[7513] = 0
      "000000" when "0001110101011010", -- t[7514] = 0
      "000000" when "0001110101011011", -- t[7515] = 0
      "000000" when "0001110101011100", -- t[7516] = 0
      "000000" when "0001110101011101", -- t[7517] = 0
      "000000" when "0001110101011110", -- t[7518] = 0
      "000000" when "0001110101011111", -- t[7519] = 0
      "000000" when "0001110101100000", -- t[7520] = 0
      "000000" when "0001110101100001", -- t[7521] = 0
      "000000" when "0001110101100010", -- t[7522] = 0
      "000000" when "0001110101100011", -- t[7523] = 0
      "000000" when "0001110101100100", -- t[7524] = 0
      "000000" when "0001110101100101", -- t[7525] = 0
      "000000" when "0001110101100110", -- t[7526] = 0
      "000000" when "0001110101100111", -- t[7527] = 0
      "000000" when "0001110101101000", -- t[7528] = 0
      "000000" when "0001110101101001", -- t[7529] = 0
      "000000" when "0001110101101010", -- t[7530] = 0
      "000000" when "0001110101101011", -- t[7531] = 0
      "000000" when "0001110101101100", -- t[7532] = 0
      "000000" when "0001110101101101", -- t[7533] = 0
      "000000" when "0001110101101110", -- t[7534] = 0
      "000000" when "0001110101101111", -- t[7535] = 0
      "000000" when "0001110101110000", -- t[7536] = 0
      "000000" when "0001110101110001", -- t[7537] = 0
      "000000" when "0001110101110010", -- t[7538] = 0
      "000000" when "0001110101110011", -- t[7539] = 0
      "000000" when "0001110101110100", -- t[7540] = 0
      "000000" when "0001110101110101", -- t[7541] = 0
      "000000" when "0001110101110110", -- t[7542] = 0
      "000000" when "0001110101110111", -- t[7543] = 0
      "000000" when "0001110101111000", -- t[7544] = 0
      "000000" when "0001110101111001", -- t[7545] = 0
      "000000" when "0001110101111010", -- t[7546] = 0
      "000000" when "0001110101111011", -- t[7547] = 0
      "000000" when "0001110101111100", -- t[7548] = 0
      "000000" when "0001110101111101", -- t[7549] = 0
      "000000" when "0001110101111110", -- t[7550] = 0
      "000000" when "0001110101111111", -- t[7551] = 0
      "000000" when "0001110110000000", -- t[7552] = 0
      "000000" when "0001110110000001", -- t[7553] = 0
      "000000" when "0001110110000010", -- t[7554] = 0
      "000000" when "0001110110000011", -- t[7555] = 0
      "000000" when "0001110110000100", -- t[7556] = 0
      "000000" when "0001110110000101", -- t[7557] = 0
      "000000" when "0001110110000110", -- t[7558] = 0
      "000000" when "0001110110000111", -- t[7559] = 0
      "000000" when "0001110110001000", -- t[7560] = 0
      "000000" when "0001110110001001", -- t[7561] = 0
      "000000" when "0001110110001010", -- t[7562] = 0
      "000000" when "0001110110001011", -- t[7563] = 0
      "000000" when "0001110110001100", -- t[7564] = 0
      "000000" when "0001110110001101", -- t[7565] = 0
      "000000" when "0001110110001110", -- t[7566] = 0
      "000000" when "0001110110001111", -- t[7567] = 0
      "000000" when "0001110110010000", -- t[7568] = 0
      "000000" when "0001110110010001", -- t[7569] = 0
      "000000" when "0001110110010010", -- t[7570] = 0
      "000000" when "0001110110010011", -- t[7571] = 0
      "000000" when "0001110110010100", -- t[7572] = 0
      "000000" when "0001110110010101", -- t[7573] = 0
      "000000" when "0001110110010110", -- t[7574] = 0
      "000000" when "0001110110010111", -- t[7575] = 0
      "000000" when "0001110110011000", -- t[7576] = 0
      "000000" when "0001110110011001", -- t[7577] = 0
      "000000" when "0001110110011010", -- t[7578] = 0
      "000000" when "0001110110011011", -- t[7579] = 0
      "000000" when "0001110110011100", -- t[7580] = 0
      "000000" when "0001110110011101", -- t[7581] = 0
      "000000" when "0001110110011110", -- t[7582] = 0
      "000000" when "0001110110011111", -- t[7583] = 0
      "000000" when "0001110110100000", -- t[7584] = 0
      "000000" when "0001110110100001", -- t[7585] = 0
      "000000" when "0001110110100010", -- t[7586] = 0
      "000000" when "0001110110100011", -- t[7587] = 0
      "000000" when "0001110110100100", -- t[7588] = 0
      "000000" when "0001110110100101", -- t[7589] = 0
      "000000" when "0001110110100110", -- t[7590] = 0
      "000000" when "0001110110100111", -- t[7591] = 0
      "000000" when "0001110110101000", -- t[7592] = 0
      "000000" when "0001110110101001", -- t[7593] = 0
      "000000" when "0001110110101010", -- t[7594] = 0
      "000000" when "0001110110101011", -- t[7595] = 0
      "000000" when "0001110110101100", -- t[7596] = 0
      "000000" when "0001110110101101", -- t[7597] = 0
      "000000" when "0001110110101110", -- t[7598] = 0
      "000000" when "0001110110101111", -- t[7599] = 0
      "000000" when "0001110110110000", -- t[7600] = 0
      "000000" when "0001110110110001", -- t[7601] = 0
      "000000" when "0001110110110010", -- t[7602] = 0
      "000000" when "0001110110110011", -- t[7603] = 0
      "000000" when "0001110110110100", -- t[7604] = 0
      "000000" when "0001110110110101", -- t[7605] = 0
      "000000" when "0001110110110110", -- t[7606] = 0
      "000000" when "0001110110110111", -- t[7607] = 0
      "000000" when "0001110110111000", -- t[7608] = 0
      "000000" when "0001110110111001", -- t[7609] = 0
      "000000" when "0001110110111010", -- t[7610] = 0
      "000000" when "0001110110111011", -- t[7611] = 0
      "000000" when "0001110110111100", -- t[7612] = 0
      "000000" when "0001110110111101", -- t[7613] = 0
      "000000" when "0001110110111110", -- t[7614] = 0
      "000000" when "0001110110111111", -- t[7615] = 0
      "000000" when "0001110111000000", -- t[7616] = 0
      "000000" when "0001110111000001", -- t[7617] = 0
      "000000" when "0001110111000010", -- t[7618] = 0
      "000000" when "0001110111000011", -- t[7619] = 0
      "000000" when "0001110111000100", -- t[7620] = 0
      "000000" when "0001110111000101", -- t[7621] = 0
      "000000" when "0001110111000110", -- t[7622] = 0
      "000000" when "0001110111000111", -- t[7623] = 0
      "000000" when "0001110111001000", -- t[7624] = 0
      "000000" when "0001110111001001", -- t[7625] = 0
      "000000" when "0001110111001010", -- t[7626] = 0
      "000000" when "0001110111001011", -- t[7627] = 0
      "000000" when "0001110111001100", -- t[7628] = 0
      "000000" when "0001110111001101", -- t[7629] = 0
      "000000" when "0001110111001110", -- t[7630] = 0
      "000000" when "0001110111001111", -- t[7631] = 0
      "000000" when "0001110111010000", -- t[7632] = 0
      "000000" when "0001110111010001", -- t[7633] = 0
      "000000" when "0001110111010010", -- t[7634] = 0
      "000000" when "0001110111010011", -- t[7635] = 0
      "000000" when "0001110111010100", -- t[7636] = 0
      "000000" when "0001110111010101", -- t[7637] = 0
      "000000" when "0001110111010110", -- t[7638] = 0
      "000000" when "0001110111010111", -- t[7639] = 0
      "000000" when "0001110111011000", -- t[7640] = 0
      "000000" when "0001110111011001", -- t[7641] = 0
      "000000" when "0001110111011010", -- t[7642] = 0
      "000000" when "0001110111011011", -- t[7643] = 0
      "000000" when "0001110111011100", -- t[7644] = 0
      "000000" when "0001110111011101", -- t[7645] = 0
      "000000" when "0001110111011110", -- t[7646] = 0
      "000000" when "0001110111011111", -- t[7647] = 0
      "000000" when "0001110111100000", -- t[7648] = 0
      "000000" when "0001110111100001", -- t[7649] = 0
      "000000" when "0001110111100010", -- t[7650] = 0
      "000000" when "0001110111100011", -- t[7651] = 0
      "000000" when "0001110111100100", -- t[7652] = 0
      "000000" when "0001110111100101", -- t[7653] = 0
      "000000" when "0001110111100110", -- t[7654] = 0
      "000000" when "0001110111100111", -- t[7655] = 0
      "000000" when "0001110111101000", -- t[7656] = 0
      "000000" when "0001110111101001", -- t[7657] = 0
      "000000" when "0001110111101010", -- t[7658] = 0
      "000000" when "0001110111101011", -- t[7659] = 0
      "000000" when "0001110111101100", -- t[7660] = 0
      "000000" when "0001110111101101", -- t[7661] = 0
      "000000" when "0001110111101110", -- t[7662] = 0
      "000000" when "0001110111101111", -- t[7663] = 0
      "000000" when "0001110111110000", -- t[7664] = 0
      "000000" when "0001110111110001", -- t[7665] = 0
      "000000" when "0001110111110010", -- t[7666] = 0
      "000000" when "0001110111110011", -- t[7667] = 0
      "000000" when "0001110111110100", -- t[7668] = 0
      "000000" when "0001110111110101", -- t[7669] = 0
      "000000" when "0001110111110110", -- t[7670] = 0
      "000000" when "0001110111110111", -- t[7671] = 0
      "000000" when "0001110111111000", -- t[7672] = 0
      "000000" when "0001110111111001", -- t[7673] = 0
      "000000" when "0001110111111010", -- t[7674] = 0
      "000000" when "0001110111111011", -- t[7675] = 0
      "000000" when "0001110111111100", -- t[7676] = 0
      "000000" when "0001110111111101", -- t[7677] = 0
      "000000" when "0001110111111110", -- t[7678] = 0
      "000000" when "0001110111111111", -- t[7679] = 0
      "000000" when "0001111000000000", -- t[7680] = 0
      "000000" when "0001111000000001", -- t[7681] = 0
      "000000" when "0001111000000010", -- t[7682] = 0
      "000000" when "0001111000000011", -- t[7683] = 0
      "000000" when "0001111000000100", -- t[7684] = 0
      "000000" when "0001111000000101", -- t[7685] = 0
      "000000" when "0001111000000110", -- t[7686] = 0
      "000000" when "0001111000000111", -- t[7687] = 0
      "000000" when "0001111000001000", -- t[7688] = 0
      "000000" when "0001111000001001", -- t[7689] = 0
      "000000" when "0001111000001010", -- t[7690] = 0
      "000000" when "0001111000001011", -- t[7691] = 0
      "000000" when "0001111000001100", -- t[7692] = 0
      "000000" when "0001111000001101", -- t[7693] = 0
      "000000" when "0001111000001110", -- t[7694] = 0
      "000000" when "0001111000001111", -- t[7695] = 0
      "000000" when "0001111000010000", -- t[7696] = 0
      "000000" when "0001111000010001", -- t[7697] = 0
      "000000" when "0001111000010010", -- t[7698] = 0
      "000000" when "0001111000010011", -- t[7699] = 0
      "000000" when "0001111000010100", -- t[7700] = 0
      "000000" when "0001111000010101", -- t[7701] = 0
      "000000" when "0001111000010110", -- t[7702] = 0
      "000000" when "0001111000010111", -- t[7703] = 0
      "000000" when "0001111000011000", -- t[7704] = 0
      "000000" when "0001111000011001", -- t[7705] = 0
      "000000" when "0001111000011010", -- t[7706] = 0
      "000000" when "0001111000011011", -- t[7707] = 0
      "000000" when "0001111000011100", -- t[7708] = 0
      "000000" when "0001111000011101", -- t[7709] = 0
      "000000" when "0001111000011110", -- t[7710] = 0
      "000000" when "0001111000011111", -- t[7711] = 0
      "000000" when "0001111000100000", -- t[7712] = 0
      "000000" when "0001111000100001", -- t[7713] = 0
      "000000" when "0001111000100010", -- t[7714] = 0
      "000000" when "0001111000100011", -- t[7715] = 0
      "000000" when "0001111000100100", -- t[7716] = 0
      "000000" when "0001111000100101", -- t[7717] = 0
      "000000" when "0001111000100110", -- t[7718] = 0
      "000000" when "0001111000100111", -- t[7719] = 0
      "000000" when "0001111000101000", -- t[7720] = 0
      "000000" when "0001111000101001", -- t[7721] = 0
      "000000" when "0001111000101010", -- t[7722] = 0
      "000000" when "0001111000101011", -- t[7723] = 0
      "000000" when "0001111000101100", -- t[7724] = 0
      "000000" when "0001111000101101", -- t[7725] = 0
      "000000" when "0001111000101110", -- t[7726] = 0
      "000000" when "0001111000101111", -- t[7727] = 0
      "000000" when "0001111000110000", -- t[7728] = 0
      "000000" when "0001111000110001", -- t[7729] = 0
      "000000" when "0001111000110010", -- t[7730] = 0
      "000000" when "0001111000110011", -- t[7731] = 0
      "000000" when "0001111000110100", -- t[7732] = 0
      "000000" when "0001111000110101", -- t[7733] = 0
      "000000" when "0001111000110110", -- t[7734] = 0
      "000000" when "0001111000110111", -- t[7735] = 0
      "000000" when "0001111000111000", -- t[7736] = 0
      "000000" when "0001111000111001", -- t[7737] = 0
      "000000" when "0001111000111010", -- t[7738] = 0
      "000000" when "0001111000111011", -- t[7739] = 0
      "000000" when "0001111000111100", -- t[7740] = 0
      "000000" when "0001111000111101", -- t[7741] = 0
      "000000" when "0001111000111110", -- t[7742] = 0
      "000000" when "0001111000111111", -- t[7743] = 0
      "000000" when "0001111001000000", -- t[7744] = 0
      "000000" when "0001111001000001", -- t[7745] = 0
      "000000" when "0001111001000010", -- t[7746] = 0
      "000000" when "0001111001000011", -- t[7747] = 0
      "000000" when "0001111001000100", -- t[7748] = 0
      "000000" when "0001111001000101", -- t[7749] = 0
      "000000" when "0001111001000110", -- t[7750] = 0
      "000000" when "0001111001000111", -- t[7751] = 0
      "000000" when "0001111001001000", -- t[7752] = 0
      "000000" when "0001111001001001", -- t[7753] = 0
      "000000" when "0001111001001010", -- t[7754] = 0
      "000000" when "0001111001001011", -- t[7755] = 0
      "000000" when "0001111001001100", -- t[7756] = 0
      "000000" when "0001111001001101", -- t[7757] = 0
      "000000" when "0001111001001110", -- t[7758] = 0
      "000000" when "0001111001001111", -- t[7759] = 0
      "000000" when "0001111001010000", -- t[7760] = 0
      "000000" when "0001111001010001", -- t[7761] = 0
      "000000" when "0001111001010010", -- t[7762] = 0
      "000000" when "0001111001010011", -- t[7763] = 0
      "000000" when "0001111001010100", -- t[7764] = 0
      "000000" when "0001111001010101", -- t[7765] = 0
      "000000" when "0001111001010110", -- t[7766] = 0
      "000000" when "0001111001010111", -- t[7767] = 0
      "000000" when "0001111001011000", -- t[7768] = 0
      "000000" when "0001111001011001", -- t[7769] = 0
      "000000" when "0001111001011010", -- t[7770] = 0
      "000000" when "0001111001011011", -- t[7771] = 0
      "000000" when "0001111001011100", -- t[7772] = 0
      "000000" when "0001111001011101", -- t[7773] = 0
      "000000" when "0001111001011110", -- t[7774] = 0
      "000000" when "0001111001011111", -- t[7775] = 0
      "000000" when "0001111001100000", -- t[7776] = 0
      "000000" when "0001111001100001", -- t[7777] = 0
      "000000" when "0001111001100010", -- t[7778] = 0
      "000000" when "0001111001100011", -- t[7779] = 0
      "000000" when "0001111001100100", -- t[7780] = 0
      "000000" when "0001111001100101", -- t[7781] = 0
      "000000" when "0001111001100110", -- t[7782] = 0
      "000000" when "0001111001100111", -- t[7783] = 0
      "000000" when "0001111001101000", -- t[7784] = 0
      "000000" when "0001111001101001", -- t[7785] = 0
      "000000" when "0001111001101010", -- t[7786] = 0
      "000000" when "0001111001101011", -- t[7787] = 0
      "000000" when "0001111001101100", -- t[7788] = 0
      "000000" when "0001111001101101", -- t[7789] = 0
      "000000" when "0001111001101110", -- t[7790] = 0
      "000000" when "0001111001101111", -- t[7791] = 0
      "000000" when "0001111001110000", -- t[7792] = 0
      "000000" when "0001111001110001", -- t[7793] = 0
      "000000" when "0001111001110010", -- t[7794] = 0
      "000000" when "0001111001110011", -- t[7795] = 0
      "000000" when "0001111001110100", -- t[7796] = 0
      "000000" when "0001111001110101", -- t[7797] = 0
      "000000" when "0001111001110110", -- t[7798] = 0
      "000000" when "0001111001110111", -- t[7799] = 0
      "000000" when "0001111001111000", -- t[7800] = 0
      "000000" when "0001111001111001", -- t[7801] = 0
      "000000" when "0001111001111010", -- t[7802] = 0
      "000000" when "0001111001111011", -- t[7803] = 0
      "000000" when "0001111001111100", -- t[7804] = 0
      "000000" when "0001111001111101", -- t[7805] = 0
      "000000" when "0001111001111110", -- t[7806] = 0
      "000000" when "0001111001111111", -- t[7807] = 0
      "000000" when "0001111010000000", -- t[7808] = 0
      "000000" when "0001111010000001", -- t[7809] = 0
      "000000" when "0001111010000010", -- t[7810] = 0
      "000000" when "0001111010000011", -- t[7811] = 0
      "000000" when "0001111010000100", -- t[7812] = 0
      "000000" when "0001111010000101", -- t[7813] = 0
      "000000" when "0001111010000110", -- t[7814] = 0
      "000000" when "0001111010000111", -- t[7815] = 0
      "000000" when "0001111010001000", -- t[7816] = 0
      "000000" when "0001111010001001", -- t[7817] = 0
      "000000" when "0001111010001010", -- t[7818] = 0
      "000000" when "0001111010001011", -- t[7819] = 0
      "000000" when "0001111010001100", -- t[7820] = 0
      "000000" when "0001111010001101", -- t[7821] = 0
      "000000" when "0001111010001110", -- t[7822] = 0
      "000000" when "0001111010001111", -- t[7823] = 0
      "000000" when "0001111010010000", -- t[7824] = 0
      "000000" when "0001111010010001", -- t[7825] = 0
      "000000" when "0001111010010010", -- t[7826] = 0
      "000000" when "0001111010010011", -- t[7827] = 0
      "000000" when "0001111010010100", -- t[7828] = 0
      "000000" when "0001111010010101", -- t[7829] = 0
      "000000" when "0001111010010110", -- t[7830] = 0
      "000000" when "0001111010010111", -- t[7831] = 0
      "000000" when "0001111010011000", -- t[7832] = 0
      "000000" when "0001111010011001", -- t[7833] = 0
      "000000" when "0001111010011010", -- t[7834] = 0
      "000000" when "0001111010011011", -- t[7835] = 0
      "000000" when "0001111010011100", -- t[7836] = 0
      "000000" when "0001111010011101", -- t[7837] = 0
      "000000" when "0001111010011110", -- t[7838] = 0
      "000000" when "0001111010011111", -- t[7839] = 0
      "000000" when "0001111010100000", -- t[7840] = 0
      "000000" when "0001111010100001", -- t[7841] = 0
      "000000" when "0001111010100010", -- t[7842] = 0
      "000000" when "0001111010100011", -- t[7843] = 0
      "000000" when "0001111010100100", -- t[7844] = 0
      "000000" when "0001111010100101", -- t[7845] = 0
      "000000" when "0001111010100110", -- t[7846] = 0
      "000000" when "0001111010100111", -- t[7847] = 0
      "000000" when "0001111010101000", -- t[7848] = 0
      "000000" when "0001111010101001", -- t[7849] = 0
      "000000" when "0001111010101010", -- t[7850] = 0
      "000000" when "0001111010101011", -- t[7851] = 0
      "000000" when "0001111010101100", -- t[7852] = 0
      "000000" when "0001111010101101", -- t[7853] = 0
      "000000" when "0001111010101110", -- t[7854] = 0
      "000000" when "0001111010101111", -- t[7855] = 0
      "000000" when "0001111010110000", -- t[7856] = 0
      "000000" when "0001111010110001", -- t[7857] = 0
      "000000" when "0001111010110010", -- t[7858] = 0
      "000000" when "0001111010110011", -- t[7859] = 0
      "000000" when "0001111010110100", -- t[7860] = 0
      "000000" when "0001111010110101", -- t[7861] = 0
      "000000" when "0001111010110110", -- t[7862] = 0
      "000000" when "0001111010110111", -- t[7863] = 0
      "000000" when "0001111010111000", -- t[7864] = 0
      "000000" when "0001111010111001", -- t[7865] = 0
      "000000" when "0001111010111010", -- t[7866] = 0
      "000000" when "0001111010111011", -- t[7867] = 0
      "000000" when "0001111010111100", -- t[7868] = 0
      "000000" when "0001111010111101", -- t[7869] = 0
      "000000" when "0001111010111110", -- t[7870] = 0
      "000000" when "0001111010111111", -- t[7871] = 0
      "000000" when "0001111011000000", -- t[7872] = 0
      "000000" when "0001111011000001", -- t[7873] = 0
      "000000" when "0001111011000010", -- t[7874] = 0
      "000000" when "0001111011000011", -- t[7875] = 0
      "000000" when "0001111011000100", -- t[7876] = 0
      "000000" when "0001111011000101", -- t[7877] = 0
      "000000" when "0001111011000110", -- t[7878] = 0
      "000000" when "0001111011000111", -- t[7879] = 0
      "000000" when "0001111011001000", -- t[7880] = 0
      "000000" when "0001111011001001", -- t[7881] = 0
      "000000" when "0001111011001010", -- t[7882] = 0
      "000000" when "0001111011001011", -- t[7883] = 0
      "000000" when "0001111011001100", -- t[7884] = 0
      "000000" when "0001111011001101", -- t[7885] = 0
      "000000" when "0001111011001110", -- t[7886] = 0
      "000000" when "0001111011001111", -- t[7887] = 0
      "000000" when "0001111011010000", -- t[7888] = 0
      "000000" when "0001111011010001", -- t[7889] = 0
      "000000" when "0001111011010010", -- t[7890] = 0
      "000000" when "0001111011010011", -- t[7891] = 0
      "000000" when "0001111011010100", -- t[7892] = 0
      "000000" when "0001111011010101", -- t[7893] = 0
      "000000" when "0001111011010110", -- t[7894] = 0
      "000000" when "0001111011010111", -- t[7895] = 0
      "000000" when "0001111011011000", -- t[7896] = 0
      "000000" when "0001111011011001", -- t[7897] = 0
      "000000" when "0001111011011010", -- t[7898] = 0
      "000000" when "0001111011011011", -- t[7899] = 0
      "000000" when "0001111011011100", -- t[7900] = 0
      "000000" when "0001111011011101", -- t[7901] = 0
      "000000" when "0001111011011110", -- t[7902] = 0
      "000000" when "0001111011011111", -- t[7903] = 0
      "000000" when "0001111011100000", -- t[7904] = 0
      "000000" when "0001111011100001", -- t[7905] = 0
      "000000" when "0001111011100010", -- t[7906] = 0
      "000000" when "0001111011100011", -- t[7907] = 0
      "000000" when "0001111011100100", -- t[7908] = 0
      "000000" when "0001111011100101", -- t[7909] = 0
      "000000" when "0001111011100110", -- t[7910] = 0
      "000000" when "0001111011100111", -- t[7911] = 0
      "000000" when "0001111011101000", -- t[7912] = 0
      "000000" when "0001111011101001", -- t[7913] = 0
      "000000" when "0001111011101010", -- t[7914] = 0
      "000000" when "0001111011101011", -- t[7915] = 0
      "000000" when "0001111011101100", -- t[7916] = 0
      "000000" when "0001111011101101", -- t[7917] = 0
      "000000" when "0001111011101110", -- t[7918] = 0
      "000000" when "0001111011101111", -- t[7919] = 0
      "000000" when "0001111011110000", -- t[7920] = 0
      "000000" when "0001111011110001", -- t[7921] = 0
      "000000" when "0001111011110010", -- t[7922] = 0
      "000000" when "0001111011110011", -- t[7923] = 0
      "000000" when "0001111011110100", -- t[7924] = 0
      "000000" when "0001111011110101", -- t[7925] = 0
      "000000" when "0001111011110110", -- t[7926] = 0
      "000000" when "0001111011110111", -- t[7927] = 0
      "000000" when "0001111011111000", -- t[7928] = 0
      "000000" when "0001111011111001", -- t[7929] = 0
      "000000" when "0001111011111010", -- t[7930] = 0
      "000000" when "0001111011111011", -- t[7931] = 0
      "000000" when "0001111011111100", -- t[7932] = 0
      "000000" when "0001111011111101", -- t[7933] = 0
      "000000" when "0001111011111110", -- t[7934] = 0
      "000000" when "0001111011111111", -- t[7935] = 0
      "000000" when "0001111100000000", -- t[7936] = 0
      "000000" when "0001111100000001", -- t[7937] = 0
      "000000" when "0001111100000010", -- t[7938] = 0
      "000000" when "0001111100000011", -- t[7939] = 0
      "000000" when "0001111100000100", -- t[7940] = 0
      "000000" when "0001111100000101", -- t[7941] = 0
      "000000" when "0001111100000110", -- t[7942] = 0
      "000000" when "0001111100000111", -- t[7943] = 0
      "000000" when "0001111100001000", -- t[7944] = 0
      "000000" when "0001111100001001", -- t[7945] = 0
      "000000" when "0001111100001010", -- t[7946] = 0
      "000000" when "0001111100001011", -- t[7947] = 0
      "000000" when "0001111100001100", -- t[7948] = 0
      "000000" when "0001111100001101", -- t[7949] = 0
      "000000" when "0001111100001110", -- t[7950] = 0
      "000000" when "0001111100001111", -- t[7951] = 0
      "000000" when "0001111100010000", -- t[7952] = 0
      "000000" when "0001111100010001", -- t[7953] = 0
      "000000" when "0001111100010010", -- t[7954] = 0
      "000000" when "0001111100010011", -- t[7955] = 0
      "000000" when "0001111100010100", -- t[7956] = 0
      "000000" when "0001111100010101", -- t[7957] = 0
      "000000" when "0001111100010110", -- t[7958] = 0
      "000000" when "0001111100010111", -- t[7959] = 0
      "000000" when "0001111100011000", -- t[7960] = 0
      "000000" when "0001111100011001", -- t[7961] = 0
      "000000" when "0001111100011010", -- t[7962] = 0
      "000000" when "0001111100011011", -- t[7963] = 0
      "000000" when "0001111100011100", -- t[7964] = 0
      "000000" when "0001111100011101", -- t[7965] = 0
      "000000" when "0001111100011110", -- t[7966] = 0
      "000000" when "0001111100011111", -- t[7967] = 0
      "000000" when "0001111100100000", -- t[7968] = 0
      "000000" when "0001111100100001", -- t[7969] = 0
      "000000" when "0001111100100010", -- t[7970] = 0
      "000000" when "0001111100100011", -- t[7971] = 0
      "000000" when "0001111100100100", -- t[7972] = 0
      "000000" when "0001111100100101", -- t[7973] = 0
      "000000" when "0001111100100110", -- t[7974] = 0
      "000000" when "0001111100100111", -- t[7975] = 0
      "000000" when "0001111100101000", -- t[7976] = 0
      "000000" when "0001111100101001", -- t[7977] = 0
      "000000" when "0001111100101010", -- t[7978] = 0
      "000000" when "0001111100101011", -- t[7979] = 0
      "000000" when "0001111100101100", -- t[7980] = 0
      "000000" when "0001111100101101", -- t[7981] = 0
      "000000" when "0001111100101110", -- t[7982] = 0
      "000000" when "0001111100101111", -- t[7983] = 0
      "000000" when "0001111100110000", -- t[7984] = 0
      "000000" when "0001111100110001", -- t[7985] = 0
      "000000" when "0001111100110010", -- t[7986] = 0
      "000000" when "0001111100110011", -- t[7987] = 0
      "000000" when "0001111100110100", -- t[7988] = 0
      "000000" when "0001111100110101", -- t[7989] = 0
      "000000" when "0001111100110110", -- t[7990] = 0
      "000000" when "0001111100110111", -- t[7991] = 0
      "000000" when "0001111100111000", -- t[7992] = 0
      "000000" when "0001111100111001", -- t[7993] = 0
      "000000" when "0001111100111010", -- t[7994] = 0
      "000000" when "0001111100111011", -- t[7995] = 0
      "000000" when "0001111100111100", -- t[7996] = 0
      "000000" when "0001111100111101", -- t[7997] = 0
      "000000" when "0001111100111110", -- t[7998] = 0
      "000000" when "0001111100111111", -- t[7999] = 0
      "000000" when "0001111101000000", -- t[8000] = 0
      "000000" when "0001111101000001", -- t[8001] = 0
      "000000" when "0001111101000010", -- t[8002] = 0
      "000000" when "0001111101000011", -- t[8003] = 0
      "000000" when "0001111101000100", -- t[8004] = 0
      "000000" when "0001111101000101", -- t[8005] = 0
      "000000" when "0001111101000110", -- t[8006] = 0
      "000000" when "0001111101000111", -- t[8007] = 0
      "000000" when "0001111101001000", -- t[8008] = 0
      "000000" when "0001111101001001", -- t[8009] = 0
      "000000" when "0001111101001010", -- t[8010] = 0
      "000000" when "0001111101001011", -- t[8011] = 0
      "000000" when "0001111101001100", -- t[8012] = 0
      "000000" when "0001111101001101", -- t[8013] = 0
      "000000" when "0001111101001110", -- t[8014] = 0
      "000000" when "0001111101001111", -- t[8015] = 0
      "000000" when "0001111101010000", -- t[8016] = 0
      "000000" when "0001111101010001", -- t[8017] = 0
      "000000" when "0001111101010010", -- t[8018] = 0
      "000000" when "0001111101010011", -- t[8019] = 0
      "000000" when "0001111101010100", -- t[8020] = 0
      "000000" when "0001111101010101", -- t[8021] = 0
      "000000" when "0001111101010110", -- t[8022] = 0
      "000000" when "0001111101010111", -- t[8023] = 0
      "000000" when "0001111101011000", -- t[8024] = 0
      "000000" when "0001111101011001", -- t[8025] = 0
      "000000" when "0001111101011010", -- t[8026] = 0
      "000000" when "0001111101011011", -- t[8027] = 0
      "000000" when "0001111101011100", -- t[8028] = 0
      "000000" when "0001111101011101", -- t[8029] = 0
      "000000" when "0001111101011110", -- t[8030] = 0
      "000000" when "0001111101011111", -- t[8031] = 0
      "000000" when "0001111101100000", -- t[8032] = 0
      "000000" when "0001111101100001", -- t[8033] = 0
      "000000" when "0001111101100010", -- t[8034] = 0
      "000000" when "0001111101100011", -- t[8035] = 0
      "000000" when "0001111101100100", -- t[8036] = 0
      "000000" when "0001111101100101", -- t[8037] = 0
      "000000" when "0001111101100110", -- t[8038] = 0
      "000000" when "0001111101100111", -- t[8039] = 0
      "000000" when "0001111101101000", -- t[8040] = 0
      "000000" when "0001111101101001", -- t[8041] = 0
      "000000" when "0001111101101010", -- t[8042] = 0
      "000000" when "0001111101101011", -- t[8043] = 0
      "000000" when "0001111101101100", -- t[8044] = 0
      "000000" when "0001111101101101", -- t[8045] = 0
      "000000" when "0001111101101110", -- t[8046] = 0
      "000000" when "0001111101101111", -- t[8047] = 0
      "000000" when "0001111101110000", -- t[8048] = 0
      "000000" when "0001111101110001", -- t[8049] = 0
      "000000" when "0001111101110010", -- t[8050] = 0
      "000000" when "0001111101110011", -- t[8051] = 0
      "000000" when "0001111101110100", -- t[8052] = 0
      "000000" when "0001111101110101", -- t[8053] = 0
      "000000" when "0001111101110110", -- t[8054] = 0
      "000000" when "0001111101110111", -- t[8055] = 0
      "000000" when "0001111101111000", -- t[8056] = 0
      "000000" when "0001111101111001", -- t[8057] = 0
      "000000" when "0001111101111010", -- t[8058] = 0
      "000000" when "0001111101111011", -- t[8059] = 0
      "000000" when "0001111101111100", -- t[8060] = 0
      "000000" when "0001111101111101", -- t[8061] = 0
      "000000" when "0001111101111110", -- t[8062] = 0
      "000000" when "0001111101111111", -- t[8063] = 0
      "000000" when "0001111110000000", -- t[8064] = 0
      "000000" when "0001111110000001", -- t[8065] = 0
      "000000" when "0001111110000010", -- t[8066] = 0
      "000000" when "0001111110000011", -- t[8067] = 0
      "000000" when "0001111110000100", -- t[8068] = 0
      "000000" when "0001111110000101", -- t[8069] = 0
      "000000" when "0001111110000110", -- t[8070] = 0
      "000000" when "0001111110000111", -- t[8071] = 0
      "000000" when "0001111110001000", -- t[8072] = 0
      "000000" when "0001111110001001", -- t[8073] = 0
      "000000" when "0001111110001010", -- t[8074] = 0
      "000000" when "0001111110001011", -- t[8075] = 0
      "000000" when "0001111110001100", -- t[8076] = 0
      "000000" when "0001111110001101", -- t[8077] = 0
      "000000" when "0001111110001110", -- t[8078] = 0
      "000000" when "0001111110001111", -- t[8079] = 0
      "000000" when "0001111110010000", -- t[8080] = 0
      "000000" when "0001111110010001", -- t[8081] = 0
      "000000" when "0001111110010010", -- t[8082] = 0
      "000000" when "0001111110010011", -- t[8083] = 0
      "000000" when "0001111110010100", -- t[8084] = 0
      "000000" when "0001111110010101", -- t[8085] = 0
      "000000" when "0001111110010110", -- t[8086] = 0
      "000000" when "0001111110010111", -- t[8087] = 0
      "000000" when "0001111110011000", -- t[8088] = 0
      "000000" when "0001111110011001", -- t[8089] = 0
      "000000" when "0001111110011010", -- t[8090] = 0
      "000000" when "0001111110011011", -- t[8091] = 0
      "000000" when "0001111110011100", -- t[8092] = 0
      "000000" when "0001111110011101", -- t[8093] = 0
      "000000" when "0001111110011110", -- t[8094] = 0
      "000000" when "0001111110011111", -- t[8095] = 0
      "000000" when "0001111110100000", -- t[8096] = 0
      "000000" when "0001111110100001", -- t[8097] = 0
      "000000" when "0001111110100010", -- t[8098] = 0
      "000000" when "0001111110100011", -- t[8099] = 0
      "000000" when "0001111110100100", -- t[8100] = 0
      "000000" when "0001111110100101", -- t[8101] = 0
      "000000" when "0001111110100110", -- t[8102] = 0
      "000000" when "0001111110100111", -- t[8103] = 0
      "000000" when "0001111110101000", -- t[8104] = 0
      "000000" when "0001111110101001", -- t[8105] = 0
      "000000" when "0001111110101010", -- t[8106] = 0
      "000000" when "0001111110101011", -- t[8107] = 0
      "000000" when "0001111110101100", -- t[8108] = 0
      "000000" when "0001111110101101", -- t[8109] = 0
      "000000" when "0001111110101110", -- t[8110] = 0
      "000000" when "0001111110101111", -- t[8111] = 0
      "000000" when "0001111110110000", -- t[8112] = 0
      "000000" when "0001111110110001", -- t[8113] = 0
      "000000" when "0001111110110010", -- t[8114] = 0
      "000000" when "0001111110110011", -- t[8115] = 0
      "000000" when "0001111110110100", -- t[8116] = 0
      "000000" when "0001111110110101", -- t[8117] = 0
      "000000" when "0001111110110110", -- t[8118] = 0
      "000000" when "0001111110110111", -- t[8119] = 0
      "000000" when "0001111110111000", -- t[8120] = 0
      "000000" when "0001111110111001", -- t[8121] = 0
      "000000" when "0001111110111010", -- t[8122] = 0
      "000000" when "0001111110111011", -- t[8123] = 0
      "000000" when "0001111110111100", -- t[8124] = 0
      "000000" when "0001111110111101", -- t[8125] = 0
      "000000" when "0001111110111110", -- t[8126] = 0
      "000000" when "0001111110111111", -- t[8127] = 0
      "000000" when "0001111111000000", -- t[8128] = 0
      "000000" when "0001111111000001", -- t[8129] = 0
      "000000" when "0001111111000010", -- t[8130] = 0
      "000000" when "0001111111000011", -- t[8131] = 0
      "000000" when "0001111111000100", -- t[8132] = 0
      "000000" when "0001111111000101", -- t[8133] = 0
      "000000" when "0001111111000110", -- t[8134] = 0
      "000000" when "0001111111000111", -- t[8135] = 0
      "000000" when "0001111111001000", -- t[8136] = 0
      "000000" when "0001111111001001", -- t[8137] = 0
      "000000" when "0001111111001010", -- t[8138] = 0
      "000000" when "0001111111001011", -- t[8139] = 0
      "000000" when "0001111111001100", -- t[8140] = 0
      "000000" when "0001111111001101", -- t[8141] = 0
      "000000" when "0001111111001110", -- t[8142] = 0
      "000000" when "0001111111001111", -- t[8143] = 0
      "000000" when "0001111111010000", -- t[8144] = 0
      "000000" when "0001111111010001", -- t[8145] = 0
      "000000" when "0001111111010010", -- t[8146] = 0
      "000000" when "0001111111010011", -- t[8147] = 0
      "000000" when "0001111111010100", -- t[8148] = 0
      "000000" when "0001111111010101", -- t[8149] = 0
      "000000" when "0001111111010110", -- t[8150] = 0
      "000000" when "0001111111010111", -- t[8151] = 0
      "000000" when "0001111111011000", -- t[8152] = 0
      "000000" when "0001111111011001", -- t[8153] = 0
      "000000" when "0001111111011010", -- t[8154] = 0
      "000000" when "0001111111011011", -- t[8155] = 0
      "000000" when "0001111111011100", -- t[8156] = 0
      "000000" when "0001111111011101", -- t[8157] = 0
      "000000" when "0001111111011110", -- t[8158] = 0
      "000000" when "0001111111011111", -- t[8159] = 0
      "000000" when "0001111111100000", -- t[8160] = 0
      "000000" when "0001111111100001", -- t[8161] = 0
      "000000" when "0001111111100010", -- t[8162] = 0
      "000000" when "0001111111100011", -- t[8163] = 0
      "000000" when "0001111111100100", -- t[8164] = 0
      "000000" when "0001111111100101", -- t[8165] = 0
      "000000" when "0001111111100110", -- t[8166] = 0
      "000000" when "0001111111100111", -- t[8167] = 0
      "000000" when "0001111111101000", -- t[8168] = 0
      "000000" when "0001111111101001", -- t[8169] = 0
      "000000" when "0001111111101010", -- t[8170] = 0
      "000000" when "0001111111101011", -- t[8171] = 0
      "000000" when "0001111111101100", -- t[8172] = 0
      "000000" when "0001111111101101", -- t[8173] = 0
      "000000" when "0001111111101110", -- t[8174] = 0
      "000000" when "0001111111101111", -- t[8175] = 0
      "000000" when "0001111111110000", -- t[8176] = 0
      "000000" when "0001111111110001", -- t[8177] = 0
      "000000" when "0001111111110010", -- t[8178] = 0
      "000000" when "0001111111110011", -- t[8179] = 0
      "000000" when "0001111111110100", -- t[8180] = 0
      "000000" when "0001111111110101", -- t[8181] = 0
      "000000" when "0001111111110110", -- t[8182] = 0
      "000000" when "0001111111110111", -- t[8183] = 0
      "000000" when "0001111111111000", -- t[8184] = 0
      "000000" when "0001111111111001", -- t[8185] = 0
      "000000" when "0001111111111010", -- t[8186] = 0
      "000000" when "0001111111111011", -- t[8187] = 0
      "000000" when "0001111111111100", -- t[8188] = 0
      "000000" when "0001111111111101", -- t[8189] = 0
      "000000" when "0001111111111110", -- t[8190] = 0
      "000000" when "0001111111111111", -- t[8191] = 0
      "000000" when "0010000000000000", -- t[8192] = 0
      "000000" when "0010000000000001", -- t[8193] = 0
      "000000" when "0010000000000010", -- t[8194] = 0
      "000000" when "0010000000000011", -- t[8195] = 0
      "000000" when "0010000000000100", -- t[8196] = 0
      "000000" when "0010000000000101", -- t[8197] = 0
      "000000" when "0010000000000110", -- t[8198] = 0
      "000000" when "0010000000000111", -- t[8199] = 0
      "000000" when "0010000000001000", -- t[8200] = 0
      "000000" when "0010000000001001", -- t[8201] = 0
      "000000" when "0010000000001010", -- t[8202] = 0
      "000000" when "0010000000001011", -- t[8203] = 0
      "000000" when "0010000000001100", -- t[8204] = 0
      "000000" when "0010000000001101", -- t[8205] = 0
      "000000" when "0010000000001110", -- t[8206] = 0
      "000000" when "0010000000001111", -- t[8207] = 0
      "000000" when "0010000000010000", -- t[8208] = 0
      "000000" when "0010000000010001", -- t[8209] = 0
      "000000" when "0010000000010010", -- t[8210] = 0
      "000000" when "0010000000010011", -- t[8211] = 0
      "000000" when "0010000000010100", -- t[8212] = 0
      "000000" when "0010000000010101", -- t[8213] = 0
      "000000" when "0010000000010110", -- t[8214] = 0
      "000000" when "0010000000010111", -- t[8215] = 0
      "000000" when "0010000000011000", -- t[8216] = 0
      "000000" when "0010000000011001", -- t[8217] = 0
      "000000" when "0010000000011010", -- t[8218] = 0
      "000000" when "0010000000011011", -- t[8219] = 0
      "000000" when "0010000000011100", -- t[8220] = 0
      "000000" when "0010000000011101", -- t[8221] = 0
      "000000" when "0010000000011110", -- t[8222] = 0
      "000000" when "0010000000011111", -- t[8223] = 0
      "000000" when "0010000000100000", -- t[8224] = 0
      "000000" when "0010000000100001", -- t[8225] = 0
      "000000" when "0010000000100010", -- t[8226] = 0
      "000000" when "0010000000100011", -- t[8227] = 0
      "000000" when "0010000000100100", -- t[8228] = 0
      "000000" when "0010000000100101", -- t[8229] = 0
      "000000" when "0010000000100110", -- t[8230] = 0
      "000000" when "0010000000100111", -- t[8231] = 0
      "000000" when "0010000000101000", -- t[8232] = 0
      "000000" when "0010000000101001", -- t[8233] = 0
      "000000" when "0010000000101010", -- t[8234] = 0
      "000000" when "0010000000101011", -- t[8235] = 0
      "000000" when "0010000000101100", -- t[8236] = 0
      "000000" when "0010000000101101", -- t[8237] = 0
      "000000" when "0010000000101110", -- t[8238] = 0
      "000000" when "0010000000101111", -- t[8239] = 0
      "000000" when "0010000000110000", -- t[8240] = 0
      "000000" when "0010000000110001", -- t[8241] = 0
      "000000" when "0010000000110010", -- t[8242] = 0
      "000000" when "0010000000110011", -- t[8243] = 0
      "000000" when "0010000000110100", -- t[8244] = 0
      "000000" when "0010000000110101", -- t[8245] = 0
      "000000" when "0010000000110110", -- t[8246] = 0
      "000000" when "0010000000110111", -- t[8247] = 0
      "000000" when "0010000000111000", -- t[8248] = 0
      "000000" when "0010000000111001", -- t[8249] = 0
      "000000" when "0010000000111010", -- t[8250] = 0
      "000000" when "0010000000111011", -- t[8251] = 0
      "000000" when "0010000000111100", -- t[8252] = 0
      "000000" when "0010000000111101", -- t[8253] = 0
      "000000" when "0010000000111110", -- t[8254] = 0
      "000000" when "0010000000111111", -- t[8255] = 0
      "000000" when "0010000001000000", -- t[8256] = 0
      "000000" when "0010000001000001", -- t[8257] = 0
      "000000" when "0010000001000010", -- t[8258] = 0
      "000000" when "0010000001000011", -- t[8259] = 0
      "000000" when "0010000001000100", -- t[8260] = 0
      "000000" when "0010000001000101", -- t[8261] = 0
      "000000" when "0010000001000110", -- t[8262] = 0
      "000000" when "0010000001000111", -- t[8263] = 0
      "000000" when "0010000001001000", -- t[8264] = 0
      "000000" when "0010000001001001", -- t[8265] = 0
      "000000" when "0010000001001010", -- t[8266] = 0
      "000000" when "0010000001001011", -- t[8267] = 0
      "000000" when "0010000001001100", -- t[8268] = 0
      "000000" when "0010000001001101", -- t[8269] = 0
      "000000" when "0010000001001110", -- t[8270] = 0
      "000000" when "0010000001001111", -- t[8271] = 0
      "000000" when "0010000001010000", -- t[8272] = 0
      "000000" when "0010000001010001", -- t[8273] = 0
      "000000" when "0010000001010010", -- t[8274] = 0
      "000000" when "0010000001010011", -- t[8275] = 0
      "000000" when "0010000001010100", -- t[8276] = 0
      "000000" when "0010000001010101", -- t[8277] = 0
      "000000" when "0010000001010110", -- t[8278] = 0
      "000000" when "0010000001010111", -- t[8279] = 0
      "000000" when "0010000001011000", -- t[8280] = 0
      "000000" when "0010000001011001", -- t[8281] = 0
      "000000" when "0010000001011010", -- t[8282] = 0
      "000000" when "0010000001011011", -- t[8283] = 0
      "000000" when "0010000001011100", -- t[8284] = 0
      "000000" when "0010000001011101", -- t[8285] = 0
      "000000" when "0010000001011110", -- t[8286] = 0
      "000000" when "0010000001011111", -- t[8287] = 0
      "000000" when "0010000001100000", -- t[8288] = 0
      "000000" when "0010000001100001", -- t[8289] = 0
      "000000" when "0010000001100010", -- t[8290] = 0
      "000000" when "0010000001100011", -- t[8291] = 0
      "000000" when "0010000001100100", -- t[8292] = 0
      "000000" when "0010000001100101", -- t[8293] = 0
      "000000" when "0010000001100110", -- t[8294] = 0
      "000000" when "0010000001100111", -- t[8295] = 0
      "000000" when "0010000001101000", -- t[8296] = 0
      "000000" when "0010000001101001", -- t[8297] = 0
      "000000" when "0010000001101010", -- t[8298] = 0
      "000000" when "0010000001101011", -- t[8299] = 0
      "000000" when "0010000001101100", -- t[8300] = 0
      "000000" when "0010000001101101", -- t[8301] = 0
      "000000" when "0010000001101110", -- t[8302] = 0
      "000000" when "0010000001101111", -- t[8303] = 0
      "000000" when "0010000001110000", -- t[8304] = 0
      "000000" when "0010000001110001", -- t[8305] = 0
      "000000" when "0010000001110010", -- t[8306] = 0
      "000000" when "0010000001110011", -- t[8307] = 0
      "000000" when "0010000001110100", -- t[8308] = 0
      "000000" when "0010000001110101", -- t[8309] = 0
      "000000" when "0010000001110110", -- t[8310] = 0
      "000000" when "0010000001110111", -- t[8311] = 0
      "000000" when "0010000001111000", -- t[8312] = 0
      "000000" when "0010000001111001", -- t[8313] = 0
      "000000" when "0010000001111010", -- t[8314] = 0
      "000000" when "0010000001111011", -- t[8315] = 0
      "000000" when "0010000001111100", -- t[8316] = 0
      "000000" when "0010000001111101", -- t[8317] = 0
      "000000" when "0010000001111110", -- t[8318] = 0
      "000000" when "0010000001111111", -- t[8319] = 0
      "000000" when "0010000010000000", -- t[8320] = 0
      "000000" when "0010000010000001", -- t[8321] = 0
      "000000" when "0010000010000010", -- t[8322] = 0
      "000000" when "0010000010000011", -- t[8323] = 0
      "000000" when "0010000010000100", -- t[8324] = 0
      "000000" when "0010000010000101", -- t[8325] = 0
      "000000" when "0010000010000110", -- t[8326] = 0
      "000000" when "0010000010000111", -- t[8327] = 0
      "000000" when "0010000010001000", -- t[8328] = 0
      "000000" when "0010000010001001", -- t[8329] = 0
      "000000" when "0010000010001010", -- t[8330] = 0
      "000000" when "0010000010001011", -- t[8331] = 0
      "000000" when "0010000010001100", -- t[8332] = 0
      "000000" when "0010000010001101", -- t[8333] = 0
      "000000" when "0010000010001110", -- t[8334] = 0
      "000000" when "0010000010001111", -- t[8335] = 0
      "000000" when "0010000010010000", -- t[8336] = 0
      "000000" when "0010000010010001", -- t[8337] = 0
      "000000" when "0010000010010010", -- t[8338] = 0
      "000000" when "0010000010010011", -- t[8339] = 0
      "000000" when "0010000010010100", -- t[8340] = 0
      "000000" when "0010000010010101", -- t[8341] = 0
      "000000" when "0010000010010110", -- t[8342] = 0
      "000000" when "0010000010010111", -- t[8343] = 0
      "000000" when "0010000010011000", -- t[8344] = 0
      "000000" when "0010000010011001", -- t[8345] = 0
      "000000" when "0010000010011010", -- t[8346] = 0
      "000000" when "0010000010011011", -- t[8347] = 0
      "000000" when "0010000010011100", -- t[8348] = 0
      "000000" when "0010000010011101", -- t[8349] = 0
      "000000" when "0010000010011110", -- t[8350] = 0
      "000000" when "0010000010011111", -- t[8351] = 0
      "000000" when "0010000010100000", -- t[8352] = 0
      "000000" when "0010000010100001", -- t[8353] = 0
      "000000" when "0010000010100010", -- t[8354] = 0
      "000000" when "0010000010100011", -- t[8355] = 0
      "000000" when "0010000010100100", -- t[8356] = 0
      "000000" when "0010000010100101", -- t[8357] = 0
      "000000" when "0010000010100110", -- t[8358] = 0
      "000000" when "0010000010100111", -- t[8359] = 0
      "000000" when "0010000010101000", -- t[8360] = 0
      "000000" when "0010000010101001", -- t[8361] = 0
      "000000" when "0010000010101010", -- t[8362] = 0
      "000000" when "0010000010101011", -- t[8363] = 0
      "000000" when "0010000010101100", -- t[8364] = 0
      "000000" when "0010000010101101", -- t[8365] = 0
      "000000" when "0010000010101110", -- t[8366] = 0
      "000000" when "0010000010101111", -- t[8367] = 0
      "000000" when "0010000010110000", -- t[8368] = 0
      "000000" when "0010000010110001", -- t[8369] = 0
      "000000" when "0010000010110010", -- t[8370] = 0
      "000000" when "0010000010110011", -- t[8371] = 0
      "000000" when "0010000010110100", -- t[8372] = 0
      "000000" when "0010000010110101", -- t[8373] = 0
      "000000" when "0010000010110110", -- t[8374] = 0
      "000000" when "0010000010110111", -- t[8375] = 0
      "000000" when "0010000010111000", -- t[8376] = 0
      "000000" when "0010000010111001", -- t[8377] = 0
      "000000" when "0010000010111010", -- t[8378] = 0
      "000000" when "0010000010111011", -- t[8379] = 0
      "000000" when "0010000010111100", -- t[8380] = 0
      "000000" when "0010000010111101", -- t[8381] = 0
      "000000" when "0010000010111110", -- t[8382] = 0
      "000000" when "0010000010111111", -- t[8383] = 0
      "000000" when "0010000011000000", -- t[8384] = 0
      "000000" when "0010000011000001", -- t[8385] = 0
      "000000" when "0010000011000010", -- t[8386] = 0
      "000000" when "0010000011000011", -- t[8387] = 0
      "000000" when "0010000011000100", -- t[8388] = 0
      "000000" when "0010000011000101", -- t[8389] = 0
      "000000" when "0010000011000110", -- t[8390] = 0
      "000000" when "0010000011000111", -- t[8391] = 0
      "000000" when "0010000011001000", -- t[8392] = 0
      "000000" when "0010000011001001", -- t[8393] = 0
      "000000" when "0010000011001010", -- t[8394] = 0
      "000000" when "0010000011001011", -- t[8395] = 0
      "000000" when "0010000011001100", -- t[8396] = 0
      "000000" when "0010000011001101", -- t[8397] = 0
      "000000" when "0010000011001110", -- t[8398] = 0
      "000000" when "0010000011001111", -- t[8399] = 0
      "000000" when "0010000011010000", -- t[8400] = 0
      "000000" when "0010000011010001", -- t[8401] = 0
      "000000" when "0010000011010010", -- t[8402] = 0
      "000000" when "0010000011010011", -- t[8403] = 0
      "000000" when "0010000011010100", -- t[8404] = 0
      "000000" when "0010000011010101", -- t[8405] = 0
      "000000" when "0010000011010110", -- t[8406] = 0
      "000000" when "0010000011010111", -- t[8407] = 0
      "000000" when "0010000011011000", -- t[8408] = 0
      "000000" when "0010000011011001", -- t[8409] = 0
      "000000" when "0010000011011010", -- t[8410] = 0
      "000000" when "0010000011011011", -- t[8411] = 0
      "000000" when "0010000011011100", -- t[8412] = 0
      "000000" when "0010000011011101", -- t[8413] = 0
      "000000" when "0010000011011110", -- t[8414] = 0
      "000000" when "0010000011011111", -- t[8415] = 0
      "000000" when "0010000011100000", -- t[8416] = 0
      "000000" when "0010000011100001", -- t[8417] = 0
      "000000" when "0010000011100010", -- t[8418] = 0
      "000000" when "0010000011100011", -- t[8419] = 0
      "000000" when "0010000011100100", -- t[8420] = 0
      "000000" when "0010000011100101", -- t[8421] = 0
      "000000" when "0010000011100110", -- t[8422] = 0
      "000000" when "0010000011100111", -- t[8423] = 0
      "000000" when "0010000011101000", -- t[8424] = 0
      "000000" when "0010000011101001", -- t[8425] = 0
      "000000" when "0010000011101010", -- t[8426] = 0
      "000000" when "0010000011101011", -- t[8427] = 0
      "000000" when "0010000011101100", -- t[8428] = 0
      "000000" when "0010000011101101", -- t[8429] = 0
      "000000" when "0010000011101110", -- t[8430] = 0
      "000000" when "0010000011101111", -- t[8431] = 0
      "000000" when "0010000011110000", -- t[8432] = 0
      "000000" when "0010000011110001", -- t[8433] = 0
      "000000" when "0010000011110010", -- t[8434] = 0
      "000000" when "0010000011110011", -- t[8435] = 0
      "000000" when "0010000011110100", -- t[8436] = 0
      "000000" when "0010000011110101", -- t[8437] = 0
      "000000" when "0010000011110110", -- t[8438] = 0
      "000000" when "0010000011110111", -- t[8439] = 0
      "000000" when "0010000011111000", -- t[8440] = 0
      "000000" when "0010000011111001", -- t[8441] = 0
      "000000" when "0010000011111010", -- t[8442] = 0
      "000000" when "0010000011111011", -- t[8443] = 0
      "000000" when "0010000011111100", -- t[8444] = 0
      "000000" when "0010000011111101", -- t[8445] = 0
      "000000" when "0010000011111110", -- t[8446] = 0
      "000000" when "0010000011111111", -- t[8447] = 0
      "000000" when "0010000100000000", -- t[8448] = 0
      "000000" when "0010000100000001", -- t[8449] = 0
      "000000" when "0010000100000010", -- t[8450] = 0
      "000000" when "0010000100000011", -- t[8451] = 0
      "000000" when "0010000100000100", -- t[8452] = 0
      "000000" when "0010000100000101", -- t[8453] = 0
      "000000" when "0010000100000110", -- t[8454] = 0
      "000000" when "0010000100000111", -- t[8455] = 0
      "000000" when "0010000100001000", -- t[8456] = 0
      "000000" when "0010000100001001", -- t[8457] = 0
      "000000" when "0010000100001010", -- t[8458] = 0
      "000000" when "0010000100001011", -- t[8459] = 0
      "000000" when "0010000100001100", -- t[8460] = 0
      "000000" when "0010000100001101", -- t[8461] = 0
      "000000" when "0010000100001110", -- t[8462] = 0
      "000000" when "0010000100001111", -- t[8463] = 0
      "000000" when "0010000100010000", -- t[8464] = 0
      "000000" when "0010000100010001", -- t[8465] = 0
      "000000" when "0010000100010010", -- t[8466] = 0
      "000000" when "0010000100010011", -- t[8467] = 0
      "000000" when "0010000100010100", -- t[8468] = 0
      "000000" when "0010000100010101", -- t[8469] = 0
      "000000" when "0010000100010110", -- t[8470] = 0
      "000000" when "0010000100010111", -- t[8471] = 0
      "000000" when "0010000100011000", -- t[8472] = 0
      "000000" when "0010000100011001", -- t[8473] = 0
      "000000" when "0010000100011010", -- t[8474] = 0
      "000000" when "0010000100011011", -- t[8475] = 0
      "000000" when "0010000100011100", -- t[8476] = 0
      "000000" when "0010000100011101", -- t[8477] = 0
      "000000" when "0010000100011110", -- t[8478] = 0
      "000000" when "0010000100011111", -- t[8479] = 0
      "000000" when "0010000100100000", -- t[8480] = 0
      "000000" when "0010000100100001", -- t[8481] = 0
      "000000" when "0010000100100010", -- t[8482] = 0
      "000000" when "0010000100100011", -- t[8483] = 0
      "000000" when "0010000100100100", -- t[8484] = 0
      "000000" when "0010000100100101", -- t[8485] = 0
      "000000" when "0010000100100110", -- t[8486] = 0
      "000000" when "0010000100100111", -- t[8487] = 0
      "000000" when "0010000100101000", -- t[8488] = 0
      "000000" when "0010000100101001", -- t[8489] = 0
      "000000" when "0010000100101010", -- t[8490] = 0
      "000000" when "0010000100101011", -- t[8491] = 0
      "000000" when "0010000100101100", -- t[8492] = 0
      "000000" when "0010000100101101", -- t[8493] = 0
      "000000" when "0010000100101110", -- t[8494] = 0
      "000000" when "0010000100101111", -- t[8495] = 0
      "000000" when "0010000100110000", -- t[8496] = 0
      "000000" when "0010000100110001", -- t[8497] = 0
      "000000" when "0010000100110010", -- t[8498] = 0
      "000000" when "0010000100110011", -- t[8499] = 0
      "000000" when "0010000100110100", -- t[8500] = 0
      "000000" when "0010000100110101", -- t[8501] = 0
      "000000" when "0010000100110110", -- t[8502] = 0
      "000000" when "0010000100110111", -- t[8503] = 0
      "000000" when "0010000100111000", -- t[8504] = 0
      "000000" when "0010000100111001", -- t[8505] = 0
      "000000" when "0010000100111010", -- t[8506] = 0
      "000000" when "0010000100111011", -- t[8507] = 0
      "000000" when "0010000100111100", -- t[8508] = 0
      "000000" when "0010000100111101", -- t[8509] = 0
      "000000" when "0010000100111110", -- t[8510] = 0
      "000000" when "0010000100111111", -- t[8511] = 0
      "000000" when "0010000101000000", -- t[8512] = 0
      "000000" when "0010000101000001", -- t[8513] = 0
      "000000" when "0010000101000010", -- t[8514] = 0
      "000000" when "0010000101000011", -- t[8515] = 0
      "000000" when "0010000101000100", -- t[8516] = 0
      "000000" when "0010000101000101", -- t[8517] = 0
      "000000" when "0010000101000110", -- t[8518] = 0
      "000000" when "0010000101000111", -- t[8519] = 0
      "000000" when "0010000101001000", -- t[8520] = 0
      "000000" when "0010000101001001", -- t[8521] = 0
      "000000" when "0010000101001010", -- t[8522] = 0
      "000000" when "0010000101001011", -- t[8523] = 0
      "000000" when "0010000101001100", -- t[8524] = 0
      "000000" when "0010000101001101", -- t[8525] = 0
      "000000" when "0010000101001110", -- t[8526] = 0
      "000000" when "0010000101001111", -- t[8527] = 0
      "000000" when "0010000101010000", -- t[8528] = 0
      "000000" when "0010000101010001", -- t[8529] = 0
      "000000" when "0010000101010010", -- t[8530] = 0
      "000000" when "0010000101010011", -- t[8531] = 0
      "000000" when "0010000101010100", -- t[8532] = 0
      "000000" when "0010000101010101", -- t[8533] = 0
      "000000" when "0010000101010110", -- t[8534] = 0
      "000000" when "0010000101010111", -- t[8535] = 0
      "000000" when "0010000101011000", -- t[8536] = 0
      "000000" when "0010000101011001", -- t[8537] = 0
      "000000" when "0010000101011010", -- t[8538] = 0
      "000000" when "0010000101011011", -- t[8539] = 0
      "000000" when "0010000101011100", -- t[8540] = 0
      "000000" when "0010000101011101", -- t[8541] = 0
      "000000" when "0010000101011110", -- t[8542] = 0
      "000000" when "0010000101011111", -- t[8543] = 0
      "000000" when "0010000101100000", -- t[8544] = 0
      "000000" when "0010000101100001", -- t[8545] = 0
      "000000" when "0010000101100010", -- t[8546] = 0
      "000000" when "0010000101100011", -- t[8547] = 0
      "000000" when "0010000101100100", -- t[8548] = 0
      "000000" when "0010000101100101", -- t[8549] = 0
      "000000" when "0010000101100110", -- t[8550] = 0
      "000000" when "0010000101100111", -- t[8551] = 0
      "000000" when "0010000101101000", -- t[8552] = 0
      "000000" when "0010000101101001", -- t[8553] = 0
      "000000" when "0010000101101010", -- t[8554] = 0
      "000000" when "0010000101101011", -- t[8555] = 0
      "000000" when "0010000101101100", -- t[8556] = 0
      "000000" when "0010000101101101", -- t[8557] = 0
      "000000" when "0010000101101110", -- t[8558] = 0
      "000000" when "0010000101101111", -- t[8559] = 0
      "000000" when "0010000101110000", -- t[8560] = 0
      "000000" when "0010000101110001", -- t[8561] = 0
      "000000" when "0010000101110010", -- t[8562] = 0
      "000000" when "0010000101110011", -- t[8563] = 0
      "000000" when "0010000101110100", -- t[8564] = 0
      "000000" when "0010000101110101", -- t[8565] = 0
      "000000" when "0010000101110110", -- t[8566] = 0
      "000000" when "0010000101110111", -- t[8567] = 0
      "000000" when "0010000101111000", -- t[8568] = 0
      "000000" when "0010000101111001", -- t[8569] = 0
      "000000" when "0010000101111010", -- t[8570] = 0
      "000000" when "0010000101111011", -- t[8571] = 0
      "000000" when "0010000101111100", -- t[8572] = 0
      "000000" when "0010000101111101", -- t[8573] = 0
      "000000" when "0010000101111110", -- t[8574] = 0
      "000000" when "0010000101111111", -- t[8575] = 0
      "000000" when "0010000110000000", -- t[8576] = 0
      "000000" when "0010000110000001", -- t[8577] = 0
      "000000" when "0010000110000010", -- t[8578] = 0
      "000000" when "0010000110000011", -- t[8579] = 0
      "000000" when "0010000110000100", -- t[8580] = 0
      "000000" when "0010000110000101", -- t[8581] = 0
      "000000" when "0010000110000110", -- t[8582] = 0
      "000000" when "0010000110000111", -- t[8583] = 0
      "000000" when "0010000110001000", -- t[8584] = 0
      "000000" when "0010000110001001", -- t[8585] = 0
      "000000" when "0010000110001010", -- t[8586] = 0
      "000000" when "0010000110001011", -- t[8587] = 0
      "000000" when "0010000110001100", -- t[8588] = 0
      "000000" when "0010000110001101", -- t[8589] = 0
      "000000" when "0010000110001110", -- t[8590] = 0
      "000000" when "0010000110001111", -- t[8591] = 0
      "000000" when "0010000110010000", -- t[8592] = 0
      "000000" when "0010000110010001", -- t[8593] = 0
      "000000" when "0010000110010010", -- t[8594] = 0
      "000000" when "0010000110010011", -- t[8595] = 0
      "000000" when "0010000110010100", -- t[8596] = 0
      "000000" when "0010000110010101", -- t[8597] = 0
      "000000" when "0010000110010110", -- t[8598] = 0
      "000000" when "0010000110010111", -- t[8599] = 0
      "000000" when "0010000110011000", -- t[8600] = 0
      "000000" when "0010000110011001", -- t[8601] = 0
      "000000" when "0010000110011010", -- t[8602] = 0
      "000000" when "0010000110011011", -- t[8603] = 0
      "000000" when "0010000110011100", -- t[8604] = 0
      "000000" when "0010000110011101", -- t[8605] = 0
      "000000" when "0010000110011110", -- t[8606] = 0
      "000000" when "0010000110011111", -- t[8607] = 0
      "000000" when "0010000110100000", -- t[8608] = 0
      "000000" when "0010000110100001", -- t[8609] = 0
      "000000" when "0010000110100010", -- t[8610] = 0
      "000000" when "0010000110100011", -- t[8611] = 0
      "000000" when "0010000110100100", -- t[8612] = 0
      "000000" when "0010000110100101", -- t[8613] = 0
      "000000" when "0010000110100110", -- t[8614] = 0
      "000000" when "0010000110100111", -- t[8615] = 0
      "000000" when "0010000110101000", -- t[8616] = 0
      "000000" when "0010000110101001", -- t[8617] = 0
      "000000" when "0010000110101010", -- t[8618] = 0
      "000000" when "0010000110101011", -- t[8619] = 0
      "000000" when "0010000110101100", -- t[8620] = 0
      "000000" when "0010000110101101", -- t[8621] = 0
      "000000" when "0010000110101110", -- t[8622] = 0
      "000000" when "0010000110101111", -- t[8623] = 0
      "000000" when "0010000110110000", -- t[8624] = 0
      "000000" when "0010000110110001", -- t[8625] = 0
      "000000" when "0010000110110010", -- t[8626] = 0
      "000000" when "0010000110110011", -- t[8627] = 0
      "000000" when "0010000110110100", -- t[8628] = 0
      "000000" when "0010000110110101", -- t[8629] = 0
      "000000" when "0010000110110110", -- t[8630] = 0
      "000000" when "0010000110110111", -- t[8631] = 0
      "000000" when "0010000110111000", -- t[8632] = 0
      "000000" when "0010000110111001", -- t[8633] = 0
      "000000" when "0010000110111010", -- t[8634] = 0
      "000000" when "0010000110111011", -- t[8635] = 0
      "000000" when "0010000110111100", -- t[8636] = 0
      "000000" when "0010000110111101", -- t[8637] = 0
      "000000" when "0010000110111110", -- t[8638] = 0
      "000000" when "0010000110111111", -- t[8639] = 0
      "000000" when "0010000111000000", -- t[8640] = 0
      "000000" when "0010000111000001", -- t[8641] = 0
      "000000" when "0010000111000010", -- t[8642] = 0
      "000000" when "0010000111000011", -- t[8643] = 0
      "000000" when "0010000111000100", -- t[8644] = 0
      "000000" when "0010000111000101", -- t[8645] = 0
      "000000" when "0010000111000110", -- t[8646] = 0
      "000000" when "0010000111000111", -- t[8647] = 0
      "000000" when "0010000111001000", -- t[8648] = 0
      "000000" when "0010000111001001", -- t[8649] = 0
      "000000" when "0010000111001010", -- t[8650] = 0
      "000000" when "0010000111001011", -- t[8651] = 0
      "000000" when "0010000111001100", -- t[8652] = 0
      "000000" when "0010000111001101", -- t[8653] = 0
      "000000" when "0010000111001110", -- t[8654] = 0
      "000000" when "0010000111001111", -- t[8655] = 0
      "000000" when "0010000111010000", -- t[8656] = 0
      "000000" when "0010000111010001", -- t[8657] = 0
      "000000" when "0010000111010010", -- t[8658] = 0
      "000000" when "0010000111010011", -- t[8659] = 0
      "000000" when "0010000111010100", -- t[8660] = 0
      "000000" when "0010000111010101", -- t[8661] = 0
      "000000" when "0010000111010110", -- t[8662] = 0
      "000000" when "0010000111010111", -- t[8663] = 0
      "000000" when "0010000111011000", -- t[8664] = 0
      "000000" when "0010000111011001", -- t[8665] = 0
      "000000" when "0010000111011010", -- t[8666] = 0
      "000000" when "0010000111011011", -- t[8667] = 0
      "000000" when "0010000111011100", -- t[8668] = 0
      "000000" when "0010000111011101", -- t[8669] = 0
      "000000" when "0010000111011110", -- t[8670] = 0
      "000000" when "0010000111011111", -- t[8671] = 0
      "000000" when "0010000111100000", -- t[8672] = 0
      "000000" when "0010000111100001", -- t[8673] = 0
      "000000" when "0010000111100010", -- t[8674] = 0
      "000000" when "0010000111100011", -- t[8675] = 0
      "000000" when "0010000111100100", -- t[8676] = 0
      "000000" when "0010000111100101", -- t[8677] = 0
      "000000" when "0010000111100110", -- t[8678] = 0
      "000000" when "0010000111100111", -- t[8679] = 0
      "000000" when "0010000111101000", -- t[8680] = 0
      "000000" when "0010000111101001", -- t[8681] = 0
      "000000" when "0010000111101010", -- t[8682] = 0
      "000000" when "0010000111101011", -- t[8683] = 0
      "000000" when "0010000111101100", -- t[8684] = 0
      "000000" when "0010000111101101", -- t[8685] = 0
      "000000" when "0010000111101110", -- t[8686] = 0
      "000000" when "0010000111101111", -- t[8687] = 0
      "000000" when "0010000111110000", -- t[8688] = 0
      "000000" when "0010000111110001", -- t[8689] = 0
      "000000" when "0010000111110010", -- t[8690] = 0
      "000000" when "0010000111110011", -- t[8691] = 0
      "000000" when "0010000111110100", -- t[8692] = 0
      "000000" when "0010000111110101", -- t[8693] = 0
      "000000" when "0010000111110110", -- t[8694] = 0
      "000000" when "0010000111110111", -- t[8695] = 0
      "000000" when "0010000111111000", -- t[8696] = 0
      "000000" when "0010000111111001", -- t[8697] = 0
      "000000" when "0010000111111010", -- t[8698] = 0
      "000000" when "0010000111111011", -- t[8699] = 0
      "000000" when "0010000111111100", -- t[8700] = 0
      "000000" when "0010000111111101", -- t[8701] = 0
      "000000" when "0010000111111110", -- t[8702] = 0
      "000000" when "0010000111111111", -- t[8703] = 0
      "000000" when "0010001000000000", -- t[8704] = 0
      "000000" when "0010001000000001", -- t[8705] = 0
      "000000" when "0010001000000010", -- t[8706] = 0
      "000000" when "0010001000000011", -- t[8707] = 0
      "000000" when "0010001000000100", -- t[8708] = 0
      "000000" when "0010001000000101", -- t[8709] = 0
      "000000" when "0010001000000110", -- t[8710] = 0
      "000000" when "0010001000000111", -- t[8711] = 0
      "000000" when "0010001000001000", -- t[8712] = 0
      "000000" when "0010001000001001", -- t[8713] = 0
      "000000" when "0010001000001010", -- t[8714] = 0
      "000000" when "0010001000001011", -- t[8715] = 0
      "000000" when "0010001000001100", -- t[8716] = 0
      "000000" when "0010001000001101", -- t[8717] = 0
      "000000" when "0010001000001110", -- t[8718] = 0
      "000000" when "0010001000001111", -- t[8719] = 0
      "000000" when "0010001000010000", -- t[8720] = 0
      "000000" when "0010001000010001", -- t[8721] = 0
      "000000" when "0010001000010010", -- t[8722] = 0
      "000000" when "0010001000010011", -- t[8723] = 0
      "000000" when "0010001000010100", -- t[8724] = 0
      "000000" when "0010001000010101", -- t[8725] = 0
      "000000" when "0010001000010110", -- t[8726] = 0
      "000000" when "0010001000010111", -- t[8727] = 0
      "000000" when "0010001000011000", -- t[8728] = 0
      "000000" when "0010001000011001", -- t[8729] = 0
      "000000" when "0010001000011010", -- t[8730] = 0
      "000000" when "0010001000011011", -- t[8731] = 0
      "000000" when "0010001000011100", -- t[8732] = 0
      "000000" when "0010001000011101", -- t[8733] = 0
      "000000" when "0010001000011110", -- t[8734] = 0
      "000000" when "0010001000011111", -- t[8735] = 0
      "000000" when "0010001000100000", -- t[8736] = 0
      "000000" when "0010001000100001", -- t[8737] = 0
      "000000" when "0010001000100010", -- t[8738] = 0
      "000000" when "0010001000100011", -- t[8739] = 0
      "000000" when "0010001000100100", -- t[8740] = 0
      "000000" when "0010001000100101", -- t[8741] = 0
      "000000" when "0010001000100110", -- t[8742] = 0
      "000000" when "0010001000100111", -- t[8743] = 0
      "000000" when "0010001000101000", -- t[8744] = 0
      "000000" when "0010001000101001", -- t[8745] = 0
      "000000" when "0010001000101010", -- t[8746] = 0
      "000000" when "0010001000101011", -- t[8747] = 0
      "000000" when "0010001000101100", -- t[8748] = 0
      "000000" when "0010001000101101", -- t[8749] = 0
      "000000" when "0010001000101110", -- t[8750] = 0
      "000000" when "0010001000101111", -- t[8751] = 0
      "000000" when "0010001000110000", -- t[8752] = 0
      "000000" when "0010001000110001", -- t[8753] = 0
      "000000" when "0010001000110010", -- t[8754] = 0
      "000000" when "0010001000110011", -- t[8755] = 0
      "000000" when "0010001000110100", -- t[8756] = 0
      "000000" when "0010001000110101", -- t[8757] = 0
      "000000" when "0010001000110110", -- t[8758] = 0
      "000000" when "0010001000110111", -- t[8759] = 0
      "000000" when "0010001000111000", -- t[8760] = 0
      "000000" when "0010001000111001", -- t[8761] = 0
      "000000" when "0010001000111010", -- t[8762] = 0
      "000000" when "0010001000111011", -- t[8763] = 0
      "000000" when "0010001000111100", -- t[8764] = 0
      "000000" when "0010001000111101", -- t[8765] = 0
      "000000" when "0010001000111110", -- t[8766] = 0
      "000000" when "0010001000111111", -- t[8767] = 0
      "000000" when "0010001001000000", -- t[8768] = 0
      "000000" when "0010001001000001", -- t[8769] = 0
      "000000" when "0010001001000010", -- t[8770] = 0
      "000000" when "0010001001000011", -- t[8771] = 0
      "000000" when "0010001001000100", -- t[8772] = 0
      "000000" when "0010001001000101", -- t[8773] = 0
      "000000" when "0010001001000110", -- t[8774] = 0
      "000000" when "0010001001000111", -- t[8775] = 0
      "000000" when "0010001001001000", -- t[8776] = 0
      "000000" when "0010001001001001", -- t[8777] = 0
      "000000" when "0010001001001010", -- t[8778] = 0
      "000000" when "0010001001001011", -- t[8779] = 0
      "000000" when "0010001001001100", -- t[8780] = 0
      "000000" when "0010001001001101", -- t[8781] = 0
      "000000" when "0010001001001110", -- t[8782] = 0
      "000000" when "0010001001001111", -- t[8783] = 0
      "000000" when "0010001001010000", -- t[8784] = 0
      "000000" when "0010001001010001", -- t[8785] = 0
      "000000" when "0010001001010010", -- t[8786] = 0
      "000000" when "0010001001010011", -- t[8787] = 0
      "000000" when "0010001001010100", -- t[8788] = 0
      "000000" when "0010001001010101", -- t[8789] = 0
      "000000" when "0010001001010110", -- t[8790] = 0
      "000000" when "0010001001010111", -- t[8791] = 0
      "000000" when "0010001001011000", -- t[8792] = 0
      "000000" when "0010001001011001", -- t[8793] = 0
      "000000" when "0010001001011010", -- t[8794] = 0
      "000000" when "0010001001011011", -- t[8795] = 0
      "000000" when "0010001001011100", -- t[8796] = 0
      "000000" when "0010001001011101", -- t[8797] = 0
      "000000" when "0010001001011110", -- t[8798] = 0
      "000000" when "0010001001011111", -- t[8799] = 0
      "000000" when "0010001001100000", -- t[8800] = 0
      "000000" when "0010001001100001", -- t[8801] = 0
      "000000" when "0010001001100010", -- t[8802] = 0
      "000000" when "0010001001100011", -- t[8803] = 0
      "000000" when "0010001001100100", -- t[8804] = 0
      "000000" when "0010001001100101", -- t[8805] = 0
      "000000" when "0010001001100110", -- t[8806] = 0
      "000000" when "0010001001100111", -- t[8807] = 0
      "000000" when "0010001001101000", -- t[8808] = 0
      "000000" when "0010001001101001", -- t[8809] = 0
      "000000" when "0010001001101010", -- t[8810] = 0
      "000000" when "0010001001101011", -- t[8811] = 0
      "000000" when "0010001001101100", -- t[8812] = 0
      "000000" when "0010001001101101", -- t[8813] = 0
      "000000" when "0010001001101110", -- t[8814] = 0
      "000000" when "0010001001101111", -- t[8815] = 0
      "000000" when "0010001001110000", -- t[8816] = 0
      "000000" when "0010001001110001", -- t[8817] = 0
      "000000" when "0010001001110010", -- t[8818] = 0
      "000000" when "0010001001110011", -- t[8819] = 0
      "000000" when "0010001001110100", -- t[8820] = 0
      "000000" when "0010001001110101", -- t[8821] = 0
      "000000" when "0010001001110110", -- t[8822] = 0
      "000000" when "0010001001110111", -- t[8823] = 0
      "000000" when "0010001001111000", -- t[8824] = 0
      "000000" when "0010001001111001", -- t[8825] = 0
      "000000" when "0010001001111010", -- t[8826] = 0
      "000000" when "0010001001111011", -- t[8827] = 0
      "000000" when "0010001001111100", -- t[8828] = 0
      "000000" when "0010001001111101", -- t[8829] = 0
      "000000" when "0010001001111110", -- t[8830] = 0
      "000000" when "0010001001111111", -- t[8831] = 0
      "000000" when "0010001010000000", -- t[8832] = 0
      "000000" when "0010001010000001", -- t[8833] = 0
      "000000" when "0010001010000010", -- t[8834] = 0
      "000000" when "0010001010000011", -- t[8835] = 0
      "000000" when "0010001010000100", -- t[8836] = 0
      "000000" when "0010001010000101", -- t[8837] = 0
      "000000" when "0010001010000110", -- t[8838] = 0
      "000000" when "0010001010000111", -- t[8839] = 0
      "000000" when "0010001010001000", -- t[8840] = 0
      "000000" when "0010001010001001", -- t[8841] = 0
      "000000" when "0010001010001010", -- t[8842] = 0
      "000000" when "0010001010001011", -- t[8843] = 0
      "000000" when "0010001010001100", -- t[8844] = 0
      "000000" when "0010001010001101", -- t[8845] = 0
      "000000" when "0010001010001110", -- t[8846] = 0
      "000000" when "0010001010001111", -- t[8847] = 0
      "000000" when "0010001010010000", -- t[8848] = 0
      "000000" when "0010001010010001", -- t[8849] = 0
      "000000" when "0010001010010010", -- t[8850] = 0
      "000000" when "0010001010010011", -- t[8851] = 0
      "000000" when "0010001010010100", -- t[8852] = 0
      "000000" when "0010001010010101", -- t[8853] = 0
      "000000" when "0010001010010110", -- t[8854] = 0
      "000000" when "0010001010010111", -- t[8855] = 0
      "000000" when "0010001010011000", -- t[8856] = 0
      "000000" when "0010001010011001", -- t[8857] = 0
      "000000" when "0010001010011010", -- t[8858] = 0
      "000000" when "0010001010011011", -- t[8859] = 0
      "000000" when "0010001010011100", -- t[8860] = 0
      "000000" when "0010001010011101", -- t[8861] = 0
      "000000" when "0010001010011110", -- t[8862] = 0
      "000000" when "0010001010011111", -- t[8863] = 0
      "000000" when "0010001010100000", -- t[8864] = 0
      "000000" when "0010001010100001", -- t[8865] = 0
      "000000" when "0010001010100010", -- t[8866] = 0
      "000000" when "0010001010100011", -- t[8867] = 0
      "000000" when "0010001010100100", -- t[8868] = 0
      "000000" when "0010001010100101", -- t[8869] = 0
      "000000" when "0010001010100110", -- t[8870] = 0
      "000000" when "0010001010100111", -- t[8871] = 0
      "000000" when "0010001010101000", -- t[8872] = 0
      "000000" when "0010001010101001", -- t[8873] = 0
      "000000" when "0010001010101010", -- t[8874] = 0
      "000000" when "0010001010101011", -- t[8875] = 0
      "000000" when "0010001010101100", -- t[8876] = 0
      "000000" when "0010001010101101", -- t[8877] = 0
      "000000" when "0010001010101110", -- t[8878] = 0
      "000000" when "0010001010101111", -- t[8879] = 0
      "000000" when "0010001010110000", -- t[8880] = 0
      "000000" when "0010001010110001", -- t[8881] = 0
      "000000" when "0010001010110010", -- t[8882] = 0
      "000000" when "0010001010110011", -- t[8883] = 0
      "000000" when "0010001010110100", -- t[8884] = 0
      "000000" when "0010001010110101", -- t[8885] = 0
      "000000" when "0010001010110110", -- t[8886] = 0
      "000000" when "0010001010110111", -- t[8887] = 0
      "000000" when "0010001010111000", -- t[8888] = 0
      "000000" when "0010001010111001", -- t[8889] = 0
      "000000" when "0010001010111010", -- t[8890] = 0
      "000000" when "0010001010111011", -- t[8891] = 0
      "000000" when "0010001010111100", -- t[8892] = 0
      "000000" when "0010001010111101", -- t[8893] = 0
      "000000" when "0010001010111110", -- t[8894] = 0
      "000000" when "0010001010111111", -- t[8895] = 0
      "000000" when "0010001011000000", -- t[8896] = 0
      "000000" when "0010001011000001", -- t[8897] = 0
      "000000" when "0010001011000010", -- t[8898] = 0
      "000000" when "0010001011000011", -- t[8899] = 0
      "000000" when "0010001011000100", -- t[8900] = 0
      "000000" when "0010001011000101", -- t[8901] = 0
      "000000" when "0010001011000110", -- t[8902] = 0
      "000000" when "0010001011000111", -- t[8903] = 0
      "000000" when "0010001011001000", -- t[8904] = 0
      "000000" when "0010001011001001", -- t[8905] = 0
      "000000" when "0010001011001010", -- t[8906] = 0
      "000000" when "0010001011001011", -- t[8907] = 0
      "000000" when "0010001011001100", -- t[8908] = 0
      "000000" when "0010001011001101", -- t[8909] = 0
      "000000" when "0010001011001110", -- t[8910] = 0
      "000000" when "0010001011001111", -- t[8911] = 0
      "000000" when "0010001011010000", -- t[8912] = 0
      "000000" when "0010001011010001", -- t[8913] = 0
      "000000" when "0010001011010010", -- t[8914] = 0
      "000000" when "0010001011010011", -- t[8915] = 0
      "000000" when "0010001011010100", -- t[8916] = 0
      "000000" when "0010001011010101", -- t[8917] = 0
      "000000" when "0010001011010110", -- t[8918] = 0
      "000000" when "0010001011010111", -- t[8919] = 0
      "000000" when "0010001011011000", -- t[8920] = 0
      "000000" when "0010001011011001", -- t[8921] = 0
      "000000" when "0010001011011010", -- t[8922] = 0
      "000000" when "0010001011011011", -- t[8923] = 0
      "000000" when "0010001011011100", -- t[8924] = 0
      "000000" when "0010001011011101", -- t[8925] = 0
      "000000" when "0010001011011110", -- t[8926] = 0
      "000000" when "0010001011011111", -- t[8927] = 0
      "000000" when "0010001011100000", -- t[8928] = 0
      "000000" when "0010001011100001", -- t[8929] = 0
      "000000" when "0010001011100010", -- t[8930] = 0
      "000000" when "0010001011100011", -- t[8931] = 0
      "000000" when "0010001011100100", -- t[8932] = 0
      "000000" when "0010001011100101", -- t[8933] = 0
      "000000" when "0010001011100110", -- t[8934] = 0
      "000000" when "0010001011100111", -- t[8935] = 0
      "000000" when "0010001011101000", -- t[8936] = 0
      "000000" when "0010001011101001", -- t[8937] = 0
      "000000" when "0010001011101010", -- t[8938] = 0
      "000000" when "0010001011101011", -- t[8939] = 0
      "000000" when "0010001011101100", -- t[8940] = 0
      "000000" when "0010001011101101", -- t[8941] = 0
      "000000" when "0010001011101110", -- t[8942] = 0
      "000000" when "0010001011101111", -- t[8943] = 0
      "000000" when "0010001011110000", -- t[8944] = 0
      "000000" when "0010001011110001", -- t[8945] = 0
      "000000" when "0010001011110010", -- t[8946] = 0
      "000000" when "0010001011110011", -- t[8947] = 0
      "000000" when "0010001011110100", -- t[8948] = 0
      "000000" when "0010001011110101", -- t[8949] = 0
      "000000" when "0010001011110110", -- t[8950] = 0
      "000000" when "0010001011110111", -- t[8951] = 0
      "000000" when "0010001011111000", -- t[8952] = 0
      "000000" when "0010001011111001", -- t[8953] = 0
      "000000" when "0010001011111010", -- t[8954] = 0
      "000000" when "0010001011111011", -- t[8955] = 0
      "000000" when "0010001011111100", -- t[8956] = 0
      "000000" when "0010001011111101", -- t[8957] = 0
      "000000" when "0010001011111110", -- t[8958] = 0
      "000000" when "0010001011111111", -- t[8959] = 0
      "000000" when "0010001100000000", -- t[8960] = 0
      "000000" when "0010001100000001", -- t[8961] = 0
      "000000" when "0010001100000010", -- t[8962] = 0
      "000000" when "0010001100000011", -- t[8963] = 0
      "000000" when "0010001100000100", -- t[8964] = 0
      "000000" when "0010001100000101", -- t[8965] = 0
      "000000" when "0010001100000110", -- t[8966] = 0
      "000000" when "0010001100000111", -- t[8967] = 0
      "000000" when "0010001100001000", -- t[8968] = 0
      "000000" when "0010001100001001", -- t[8969] = 0
      "000000" when "0010001100001010", -- t[8970] = 0
      "000000" when "0010001100001011", -- t[8971] = 0
      "000000" when "0010001100001100", -- t[8972] = 0
      "000000" when "0010001100001101", -- t[8973] = 0
      "000000" when "0010001100001110", -- t[8974] = 0
      "000000" when "0010001100001111", -- t[8975] = 0
      "000000" when "0010001100010000", -- t[8976] = 0
      "000000" when "0010001100010001", -- t[8977] = 0
      "000000" when "0010001100010010", -- t[8978] = 0
      "000000" when "0010001100010011", -- t[8979] = 0
      "000000" when "0010001100010100", -- t[8980] = 0
      "000000" when "0010001100010101", -- t[8981] = 0
      "000000" when "0010001100010110", -- t[8982] = 0
      "000000" when "0010001100010111", -- t[8983] = 0
      "000000" when "0010001100011000", -- t[8984] = 0
      "000000" when "0010001100011001", -- t[8985] = 0
      "000000" when "0010001100011010", -- t[8986] = 0
      "000000" when "0010001100011011", -- t[8987] = 0
      "000000" when "0010001100011100", -- t[8988] = 0
      "000000" when "0010001100011101", -- t[8989] = 0
      "000000" when "0010001100011110", -- t[8990] = 0
      "000000" when "0010001100011111", -- t[8991] = 0
      "000000" when "0010001100100000", -- t[8992] = 0
      "000000" when "0010001100100001", -- t[8993] = 0
      "000000" when "0010001100100010", -- t[8994] = 0
      "000000" when "0010001100100011", -- t[8995] = 0
      "000000" when "0010001100100100", -- t[8996] = 0
      "000000" when "0010001100100101", -- t[8997] = 0
      "000000" when "0010001100100110", -- t[8998] = 0
      "000000" when "0010001100100111", -- t[8999] = 0
      "000000" when "0010001100101000", -- t[9000] = 0
      "000000" when "0010001100101001", -- t[9001] = 0
      "000000" when "0010001100101010", -- t[9002] = 0
      "000000" when "0010001100101011", -- t[9003] = 0
      "000000" when "0010001100101100", -- t[9004] = 0
      "000000" when "0010001100101101", -- t[9005] = 0
      "000000" when "0010001100101110", -- t[9006] = 0
      "000000" when "0010001100101111", -- t[9007] = 0
      "000000" when "0010001100110000", -- t[9008] = 0
      "000000" when "0010001100110001", -- t[9009] = 0
      "000000" when "0010001100110010", -- t[9010] = 0
      "000000" when "0010001100110011", -- t[9011] = 0
      "000000" when "0010001100110100", -- t[9012] = 0
      "000000" when "0010001100110101", -- t[9013] = 0
      "000000" when "0010001100110110", -- t[9014] = 0
      "000000" when "0010001100110111", -- t[9015] = 0
      "000000" when "0010001100111000", -- t[9016] = 0
      "000000" when "0010001100111001", -- t[9017] = 0
      "000000" when "0010001100111010", -- t[9018] = 0
      "000000" when "0010001100111011", -- t[9019] = 0
      "000000" when "0010001100111100", -- t[9020] = 0
      "000000" when "0010001100111101", -- t[9021] = 0
      "000000" when "0010001100111110", -- t[9022] = 0
      "000000" when "0010001100111111", -- t[9023] = 0
      "000000" when "0010001101000000", -- t[9024] = 0
      "000000" when "0010001101000001", -- t[9025] = 0
      "000000" when "0010001101000010", -- t[9026] = 0
      "000000" when "0010001101000011", -- t[9027] = 0
      "000000" when "0010001101000100", -- t[9028] = 0
      "000000" when "0010001101000101", -- t[9029] = 0
      "000000" when "0010001101000110", -- t[9030] = 0
      "000000" when "0010001101000111", -- t[9031] = 0
      "000000" when "0010001101001000", -- t[9032] = 0
      "000000" when "0010001101001001", -- t[9033] = 0
      "000000" when "0010001101001010", -- t[9034] = 0
      "000000" when "0010001101001011", -- t[9035] = 0
      "000000" when "0010001101001100", -- t[9036] = 0
      "000000" when "0010001101001101", -- t[9037] = 0
      "000000" when "0010001101001110", -- t[9038] = 0
      "000000" when "0010001101001111", -- t[9039] = 0
      "000000" when "0010001101010000", -- t[9040] = 0
      "000000" when "0010001101010001", -- t[9041] = 0
      "000000" when "0010001101010010", -- t[9042] = 0
      "000000" when "0010001101010011", -- t[9043] = 0
      "000000" when "0010001101010100", -- t[9044] = 0
      "000000" when "0010001101010101", -- t[9045] = 0
      "000000" when "0010001101010110", -- t[9046] = 0
      "000000" when "0010001101010111", -- t[9047] = 0
      "000000" when "0010001101011000", -- t[9048] = 0
      "000000" when "0010001101011001", -- t[9049] = 0
      "000000" when "0010001101011010", -- t[9050] = 0
      "000000" when "0010001101011011", -- t[9051] = 0
      "000000" when "0010001101011100", -- t[9052] = 0
      "000000" when "0010001101011101", -- t[9053] = 0
      "000000" when "0010001101011110", -- t[9054] = 0
      "000000" when "0010001101011111", -- t[9055] = 0
      "000000" when "0010001101100000", -- t[9056] = 0
      "000000" when "0010001101100001", -- t[9057] = 0
      "000000" when "0010001101100010", -- t[9058] = 0
      "000000" when "0010001101100011", -- t[9059] = 0
      "000000" when "0010001101100100", -- t[9060] = 0
      "000000" when "0010001101100101", -- t[9061] = 0
      "000000" when "0010001101100110", -- t[9062] = 0
      "000000" when "0010001101100111", -- t[9063] = 0
      "000000" when "0010001101101000", -- t[9064] = 0
      "000000" when "0010001101101001", -- t[9065] = 0
      "000000" when "0010001101101010", -- t[9066] = 0
      "000000" when "0010001101101011", -- t[9067] = 0
      "000000" when "0010001101101100", -- t[9068] = 0
      "000000" when "0010001101101101", -- t[9069] = 0
      "000000" when "0010001101101110", -- t[9070] = 0
      "000000" when "0010001101101111", -- t[9071] = 0
      "000000" when "0010001101110000", -- t[9072] = 0
      "000000" when "0010001101110001", -- t[9073] = 0
      "000000" when "0010001101110010", -- t[9074] = 0
      "000000" when "0010001101110011", -- t[9075] = 0
      "000000" when "0010001101110100", -- t[9076] = 0
      "000000" when "0010001101110101", -- t[9077] = 0
      "000000" when "0010001101110110", -- t[9078] = 0
      "000000" when "0010001101110111", -- t[9079] = 0
      "000000" when "0010001101111000", -- t[9080] = 0
      "000000" when "0010001101111001", -- t[9081] = 0
      "000000" when "0010001101111010", -- t[9082] = 0
      "000000" when "0010001101111011", -- t[9083] = 0
      "000000" when "0010001101111100", -- t[9084] = 0
      "000000" when "0010001101111101", -- t[9085] = 0
      "000000" when "0010001101111110", -- t[9086] = 0
      "000000" when "0010001101111111", -- t[9087] = 0
      "000000" when "0010001110000000", -- t[9088] = 0
      "000000" when "0010001110000001", -- t[9089] = 0
      "000000" when "0010001110000010", -- t[9090] = 0
      "000000" when "0010001110000011", -- t[9091] = 0
      "000000" when "0010001110000100", -- t[9092] = 0
      "000000" when "0010001110000101", -- t[9093] = 0
      "000000" when "0010001110000110", -- t[9094] = 0
      "000000" when "0010001110000111", -- t[9095] = 0
      "000000" when "0010001110001000", -- t[9096] = 0
      "000000" when "0010001110001001", -- t[9097] = 0
      "000000" when "0010001110001010", -- t[9098] = 0
      "000000" when "0010001110001011", -- t[9099] = 0
      "000000" when "0010001110001100", -- t[9100] = 0
      "000000" when "0010001110001101", -- t[9101] = 0
      "000000" when "0010001110001110", -- t[9102] = 0
      "000000" when "0010001110001111", -- t[9103] = 0
      "000000" when "0010001110010000", -- t[9104] = 0
      "000000" when "0010001110010001", -- t[9105] = 0
      "000000" when "0010001110010010", -- t[9106] = 0
      "000000" when "0010001110010011", -- t[9107] = 0
      "000000" when "0010001110010100", -- t[9108] = 0
      "000000" when "0010001110010101", -- t[9109] = 0
      "000000" when "0010001110010110", -- t[9110] = 0
      "000000" when "0010001110010111", -- t[9111] = 0
      "000000" when "0010001110011000", -- t[9112] = 0
      "000000" when "0010001110011001", -- t[9113] = 0
      "000000" when "0010001110011010", -- t[9114] = 0
      "000000" when "0010001110011011", -- t[9115] = 0
      "000000" when "0010001110011100", -- t[9116] = 0
      "000000" when "0010001110011101", -- t[9117] = 0
      "000000" when "0010001110011110", -- t[9118] = 0
      "000000" when "0010001110011111", -- t[9119] = 0
      "000000" when "0010001110100000", -- t[9120] = 0
      "000000" when "0010001110100001", -- t[9121] = 0
      "000000" when "0010001110100010", -- t[9122] = 0
      "000000" when "0010001110100011", -- t[9123] = 0
      "000000" when "0010001110100100", -- t[9124] = 0
      "000000" when "0010001110100101", -- t[9125] = 0
      "000000" when "0010001110100110", -- t[9126] = 0
      "000000" when "0010001110100111", -- t[9127] = 0
      "000000" when "0010001110101000", -- t[9128] = 0
      "000000" when "0010001110101001", -- t[9129] = 0
      "000000" when "0010001110101010", -- t[9130] = 0
      "000000" when "0010001110101011", -- t[9131] = 0
      "000000" when "0010001110101100", -- t[9132] = 0
      "000000" when "0010001110101101", -- t[9133] = 0
      "000000" when "0010001110101110", -- t[9134] = 0
      "000000" when "0010001110101111", -- t[9135] = 0
      "000000" when "0010001110110000", -- t[9136] = 0
      "000000" when "0010001110110001", -- t[9137] = 0
      "000000" when "0010001110110010", -- t[9138] = 0
      "000000" when "0010001110110011", -- t[9139] = 0
      "000000" when "0010001110110100", -- t[9140] = 0
      "000000" when "0010001110110101", -- t[9141] = 0
      "000000" when "0010001110110110", -- t[9142] = 0
      "000000" when "0010001110110111", -- t[9143] = 0
      "000000" when "0010001110111000", -- t[9144] = 0
      "000000" when "0010001110111001", -- t[9145] = 0
      "000000" when "0010001110111010", -- t[9146] = 0
      "000000" when "0010001110111011", -- t[9147] = 0
      "000000" when "0010001110111100", -- t[9148] = 0
      "000000" when "0010001110111101", -- t[9149] = 0
      "000000" when "0010001110111110", -- t[9150] = 0
      "000000" when "0010001110111111", -- t[9151] = 0
      "000000" when "0010001111000000", -- t[9152] = 0
      "000000" when "0010001111000001", -- t[9153] = 0
      "000000" when "0010001111000010", -- t[9154] = 0
      "000000" when "0010001111000011", -- t[9155] = 0
      "000000" when "0010001111000100", -- t[9156] = 0
      "000000" when "0010001111000101", -- t[9157] = 0
      "000000" when "0010001111000110", -- t[9158] = 0
      "000000" when "0010001111000111", -- t[9159] = 0
      "000000" when "0010001111001000", -- t[9160] = 0
      "000000" when "0010001111001001", -- t[9161] = 0
      "000000" when "0010001111001010", -- t[9162] = 0
      "000000" when "0010001111001011", -- t[9163] = 0
      "000000" when "0010001111001100", -- t[9164] = 0
      "000000" when "0010001111001101", -- t[9165] = 0
      "000000" when "0010001111001110", -- t[9166] = 0
      "000000" when "0010001111001111", -- t[9167] = 0
      "000000" when "0010001111010000", -- t[9168] = 0
      "000000" when "0010001111010001", -- t[9169] = 0
      "000000" when "0010001111010010", -- t[9170] = 0
      "000000" when "0010001111010011", -- t[9171] = 0
      "000000" when "0010001111010100", -- t[9172] = 0
      "000000" when "0010001111010101", -- t[9173] = 0
      "000000" when "0010001111010110", -- t[9174] = 0
      "000000" when "0010001111010111", -- t[9175] = 0
      "000000" when "0010001111011000", -- t[9176] = 0
      "000000" when "0010001111011001", -- t[9177] = 0
      "000000" when "0010001111011010", -- t[9178] = 0
      "000000" when "0010001111011011", -- t[9179] = 0
      "000000" when "0010001111011100", -- t[9180] = 0
      "000000" when "0010001111011101", -- t[9181] = 0
      "000000" when "0010001111011110", -- t[9182] = 0
      "000000" when "0010001111011111", -- t[9183] = 0
      "000000" when "0010001111100000", -- t[9184] = 0
      "000000" when "0010001111100001", -- t[9185] = 0
      "000000" when "0010001111100010", -- t[9186] = 0
      "000000" when "0010001111100011", -- t[9187] = 0
      "000000" when "0010001111100100", -- t[9188] = 0
      "000000" when "0010001111100101", -- t[9189] = 0
      "000000" when "0010001111100110", -- t[9190] = 0
      "000000" when "0010001111100111", -- t[9191] = 0
      "000000" when "0010001111101000", -- t[9192] = 0
      "000000" when "0010001111101001", -- t[9193] = 0
      "000000" when "0010001111101010", -- t[9194] = 0
      "000000" when "0010001111101011", -- t[9195] = 0
      "000000" when "0010001111101100", -- t[9196] = 0
      "000000" when "0010001111101101", -- t[9197] = 0
      "000000" when "0010001111101110", -- t[9198] = 0
      "000000" when "0010001111101111", -- t[9199] = 0
      "000000" when "0010001111110000", -- t[9200] = 0
      "000000" when "0010001111110001", -- t[9201] = 0
      "000000" when "0010001111110010", -- t[9202] = 0
      "000000" when "0010001111110011", -- t[9203] = 0
      "000000" when "0010001111110100", -- t[9204] = 0
      "000000" when "0010001111110101", -- t[9205] = 0
      "000000" when "0010001111110110", -- t[9206] = 0
      "000000" when "0010001111110111", -- t[9207] = 0
      "000000" when "0010001111111000", -- t[9208] = 0
      "000000" when "0010001111111001", -- t[9209] = 0
      "000000" when "0010001111111010", -- t[9210] = 0
      "000000" when "0010001111111011", -- t[9211] = 0
      "000000" when "0010001111111100", -- t[9212] = 0
      "000000" when "0010001111111101", -- t[9213] = 0
      "000000" when "0010001111111110", -- t[9214] = 0
      "000000" when "0010001111111111", -- t[9215] = 0
      "000000" when "0010010000000000", -- t[9216] = 0
      "000000" when "0010010000000001", -- t[9217] = 0
      "000000" when "0010010000000010", -- t[9218] = 0
      "000000" when "0010010000000011", -- t[9219] = 0
      "000000" when "0010010000000100", -- t[9220] = 0
      "000000" when "0010010000000101", -- t[9221] = 0
      "000000" when "0010010000000110", -- t[9222] = 0
      "000000" when "0010010000000111", -- t[9223] = 0
      "000000" when "0010010000001000", -- t[9224] = 0
      "000000" when "0010010000001001", -- t[9225] = 0
      "000000" when "0010010000001010", -- t[9226] = 0
      "000000" when "0010010000001011", -- t[9227] = 0
      "000000" when "0010010000001100", -- t[9228] = 0
      "000000" when "0010010000001101", -- t[9229] = 0
      "000000" when "0010010000001110", -- t[9230] = 0
      "000000" when "0010010000001111", -- t[9231] = 0
      "000000" when "0010010000010000", -- t[9232] = 0
      "000000" when "0010010000010001", -- t[9233] = 0
      "000000" when "0010010000010010", -- t[9234] = 0
      "000000" when "0010010000010011", -- t[9235] = 0
      "000000" when "0010010000010100", -- t[9236] = 0
      "000000" when "0010010000010101", -- t[9237] = 0
      "000000" when "0010010000010110", -- t[9238] = 0
      "000000" when "0010010000010111", -- t[9239] = 0
      "000000" when "0010010000011000", -- t[9240] = 0
      "000000" when "0010010000011001", -- t[9241] = 0
      "000000" when "0010010000011010", -- t[9242] = 0
      "000000" when "0010010000011011", -- t[9243] = 0
      "000000" when "0010010000011100", -- t[9244] = 0
      "000000" when "0010010000011101", -- t[9245] = 0
      "000000" when "0010010000011110", -- t[9246] = 0
      "000000" when "0010010000011111", -- t[9247] = 0
      "000000" when "0010010000100000", -- t[9248] = 0
      "000000" when "0010010000100001", -- t[9249] = 0
      "000000" when "0010010000100010", -- t[9250] = 0
      "000000" when "0010010000100011", -- t[9251] = 0
      "000000" when "0010010000100100", -- t[9252] = 0
      "000000" when "0010010000100101", -- t[9253] = 0
      "000000" when "0010010000100110", -- t[9254] = 0
      "000000" when "0010010000100111", -- t[9255] = 0
      "000000" when "0010010000101000", -- t[9256] = 0
      "000000" when "0010010000101001", -- t[9257] = 0
      "000000" when "0010010000101010", -- t[9258] = 0
      "000000" when "0010010000101011", -- t[9259] = 0
      "000000" when "0010010000101100", -- t[9260] = 0
      "000000" when "0010010000101101", -- t[9261] = 0
      "000000" when "0010010000101110", -- t[9262] = 0
      "000000" when "0010010000101111", -- t[9263] = 0
      "000000" when "0010010000110000", -- t[9264] = 0
      "000000" when "0010010000110001", -- t[9265] = 0
      "000000" when "0010010000110010", -- t[9266] = 0
      "000000" when "0010010000110011", -- t[9267] = 0
      "000000" when "0010010000110100", -- t[9268] = 0
      "000000" when "0010010000110101", -- t[9269] = 0
      "000000" when "0010010000110110", -- t[9270] = 0
      "000000" when "0010010000110111", -- t[9271] = 0
      "000000" when "0010010000111000", -- t[9272] = 0
      "000000" when "0010010000111001", -- t[9273] = 0
      "000000" when "0010010000111010", -- t[9274] = 0
      "000000" when "0010010000111011", -- t[9275] = 0
      "000000" when "0010010000111100", -- t[9276] = 0
      "000000" when "0010010000111101", -- t[9277] = 0
      "000000" when "0010010000111110", -- t[9278] = 0
      "000000" when "0010010000111111", -- t[9279] = 0
      "000000" when "0010010001000000", -- t[9280] = 0
      "000000" when "0010010001000001", -- t[9281] = 0
      "000000" when "0010010001000010", -- t[9282] = 0
      "000000" when "0010010001000011", -- t[9283] = 0
      "000000" when "0010010001000100", -- t[9284] = 0
      "000000" when "0010010001000101", -- t[9285] = 0
      "000000" when "0010010001000110", -- t[9286] = 0
      "000000" when "0010010001000111", -- t[9287] = 0
      "000000" when "0010010001001000", -- t[9288] = 0
      "000000" when "0010010001001001", -- t[9289] = 0
      "000000" when "0010010001001010", -- t[9290] = 0
      "000000" when "0010010001001011", -- t[9291] = 0
      "000000" when "0010010001001100", -- t[9292] = 0
      "000000" when "0010010001001101", -- t[9293] = 0
      "000000" when "0010010001001110", -- t[9294] = 0
      "000000" when "0010010001001111", -- t[9295] = 0
      "000000" when "0010010001010000", -- t[9296] = 0
      "000000" when "0010010001010001", -- t[9297] = 0
      "000000" when "0010010001010010", -- t[9298] = 0
      "000000" when "0010010001010011", -- t[9299] = 0
      "000000" when "0010010001010100", -- t[9300] = 0
      "000000" when "0010010001010101", -- t[9301] = 0
      "000000" when "0010010001010110", -- t[9302] = 0
      "000000" when "0010010001010111", -- t[9303] = 0
      "000000" when "0010010001011000", -- t[9304] = 0
      "000000" when "0010010001011001", -- t[9305] = 0
      "000000" when "0010010001011010", -- t[9306] = 0
      "000000" when "0010010001011011", -- t[9307] = 0
      "000000" when "0010010001011100", -- t[9308] = 0
      "000000" when "0010010001011101", -- t[9309] = 0
      "000000" when "0010010001011110", -- t[9310] = 0
      "000000" when "0010010001011111", -- t[9311] = 0
      "000000" when "0010010001100000", -- t[9312] = 0
      "000000" when "0010010001100001", -- t[9313] = 0
      "000000" when "0010010001100010", -- t[9314] = 0
      "000000" when "0010010001100011", -- t[9315] = 0
      "000000" when "0010010001100100", -- t[9316] = 0
      "000000" when "0010010001100101", -- t[9317] = 0
      "000000" when "0010010001100110", -- t[9318] = 0
      "000000" when "0010010001100111", -- t[9319] = 0
      "000000" when "0010010001101000", -- t[9320] = 0
      "000000" when "0010010001101001", -- t[9321] = 0
      "000000" when "0010010001101010", -- t[9322] = 0
      "000000" when "0010010001101011", -- t[9323] = 0
      "000000" when "0010010001101100", -- t[9324] = 0
      "000000" when "0010010001101101", -- t[9325] = 0
      "000000" when "0010010001101110", -- t[9326] = 0
      "000000" when "0010010001101111", -- t[9327] = 0
      "000000" when "0010010001110000", -- t[9328] = 0
      "000000" when "0010010001110001", -- t[9329] = 0
      "000000" when "0010010001110010", -- t[9330] = 0
      "000000" when "0010010001110011", -- t[9331] = 0
      "000000" when "0010010001110100", -- t[9332] = 0
      "000000" when "0010010001110101", -- t[9333] = 0
      "000000" when "0010010001110110", -- t[9334] = 0
      "000000" when "0010010001110111", -- t[9335] = 0
      "000000" when "0010010001111000", -- t[9336] = 0
      "000000" when "0010010001111001", -- t[9337] = 0
      "000000" when "0010010001111010", -- t[9338] = 0
      "000000" when "0010010001111011", -- t[9339] = 0
      "000000" when "0010010001111100", -- t[9340] = 0
      "000000" when "0010010001111101", -- t[9341] = 0
      "000000" when "0010010001111110", -- t[9342] = 0
      "000000" when "0010010001111111", -- t[9343] = 0
      "000000" when "0010010010000000", -- t[9344] = 0
      "000000" when "0010010010000001", -- t[9345] = 0
      "000000" when "0010010010000010", -- t[9346] = 0
      "000000" when "0010010010000011", -- t[9347] = 0
      "000000" when "0010010010000100", -- t[9348] = 0
      "000000" when "0010010010000101", -- t[9349] = 0
      "000000" when "0010010010000110", -- t[9350] = 0
      "000000" when "0010010010000111", -- t[9351] = 0
      "000000" when "0010010010001000", -- t[9352] = 0
      "000000" when "0010010010001001", -- t[9353] = 0
      "000000" when "0010010010001010", -- t[9354] = 0
      "000000" when "0010010010001011", -- t[9355] = 0
      "000000" when "0010010010001100", -- t[9356] = 0
      "000000" when "0010010010001101", -- t[9357] = 0
      "000000" when "0010010010001110", -- t[9358] = 0
      "000000" when "0010010010001111", -- t[9359] = 0
      "000000" when "0010010010010000", -- t[9360] = 0
      "000000" when "0010010010010001", -- t[9361] = 0
      "000000" when "0010010010010010", -- t[9362] = 0
      "000000" when "0010010010010011", -- t[9363] = 0
      "000000" when "0010010010010100", -- t[9364] = 0
      "000000" when "0010010010010101", -- t[9365] = 0
      "000000" when "0010010010010110", -- t[9366] = 0
      "000000" when "0010010010010111", -- t[9367] = 0
      "000000" when "0010010010011000", -- t[9368] = 0
      "000000" when "0010010010011001", -- t[9369] = 0
      "000000" when "0010010010011010", -- t[9370] = 0
      "000000" when "0010010010011011", -- t[9371] = 0
      "000000" when "0010010010011100", -- t[9372] = 0
      "000000" when "0010010010011101", -- t[9373] = 0
      "000000" when "0010010010011110", -- t[9374] = 0
      "000000" when "0010010010011111", -- t[9375] = 0
      "000000" when "0010010010100000", -- t[9376] = 0
      "000000" when "0010010010100001", -- t[9377] = 0
      "000000" when "0010010010100010", -- t[9378] = 0
      "000000" when "0010010010100011", -- t[9379] = 0
      "000000" when "0010010010100100", -- t[9380] = 0
      "000000" when "0010010010100101", -- t[9381] = 0
      "000000" when "0010010010100110", -- t[9382] = 0
      "000000" when "0010010010100111", -- t[9383] = 0
      "000000" when "0010010010101000", -- t[9384] = 0
      "000000" when "0010010010101001", -- t[9385] = 0
      "000000" when "0010010010101010", -- t[9386] = 0
      "000000" when "0010010010101011", -- t[9387] = 0
      "000000" when "0010010010101100", -- t[9388] = 0
      "000000" when "0010010010101101", -- t[9389] = 0
      "000000" when "0010010010101110", -- t[9390] = 0
      "000000" when "0010010010101111", -- t[9391] = 0
      "000000" when "0010010010110000", -- t[9392] = 0
      "000000" when "0010010010110001", -- t[9393] = 0
      "000000" when "0010010010110010", -- t[9394] = 0
      "000000" when "0010010010110011", -- t[9395] = 0
      "000000" when "0010010010110100", -- t[9396] = 0
      "000000" when "0010010010110101", -- t[9397] = 0
      "000000" when "0010010010110110", -- t[9398] = 0
      "000000" when "0010010010110111", -- t[9399] = 0
      "000000" when "0010010010111000", -- t[9400] = 0
      "000000" when "0010010010111001", -- t[9401] = 0
      "000000" when "0010010010111010", -- t[9402] = 0
      "000000" when "0010010010111011", -- t[9403] = 0
      "000000" when "0010010010111100", -- t[9404] = 0
      "000000" when "0010010010111101", -- t[9405] = 0
      "000000" when "0010010010111110", -- t[9406] = 0
      "000000" when "0010010010111111", -- t[9407] = 0
      "000000" when "0010010011000000", -- t[9408] = 0
      "000000" when "0010010011000001", -- t[9409] = 0
      "000000" when "0010010011000010", -- t[9410] = 0
      "000000" when "0010010011000011", -- t[9411] = 0
      "000000" when "0010010011000100", -- t[9412] = 0
      "000000" when "0010010011000101", -- t[9413] = 0
      "000000" when "0010010011000110", -- t[9414] = 0
      "000000" when "0010010011000111", -- t[9415] = 0
      "000000" when "0010010011001000", -- t[9416] = 0
      "000000" when "0010010011001001", -- t[9417] = 0
      "000000" when "0010010011001010", -- t[9418] = 0
      "000000" when "0010010011001011", -- t[9419] = 0
      "000000" when "0010010011001100", -- t[9420] = 0
      "000000" when "0010010011001101", -- t[9421] = 0
      "000000" when "0010010011001110", -- t[9422] = 0
      "000000" when "0010010011001111", -- t[9423] = 0
      "000000" when "0010010011010000", -- t[9424] = 0
      "000000" when "0010010011010001", -- t[9425] = 0
      "000000" when "0010010011010010", -- t[9426] = 0
      "000000" when "0010010011010011", -- t[9427] = 0
      "000000" when "0010010011010100", -- t[9428] = 0
      "000000" when "0010010011010101", -- t[9429] = 0
      "000000" when "0010010011010110", -- t[9430] = 0
      "000000" when "0010010011010111", -- t[9431] = 0
      "000000" when "0010010011011000", -- t[9432] = 0
      "000000" when "0010010011011001", -- t[9433] = 0
      "000000" when "0010010011011010", -- t[9434] = 0
      "000000" when "0010010011011011", -- t[9435] = 0
      "000000" when "0010010011011100", -- t[9436] = 0
      "000000" when "0010010011011101", -- t[9437] = 0
      "000000" when "0010010011011110", -- t[9438] = 0
      "000000" when "0010010011011111", -- t[9439] = 0
      "000000" when "0010010011100000", -- t[9440] = 0
      "000000" when "0010010011100001", -- t[9441] = 0
      "000000" when "0010010011100010", -- t[9442] = 0
      "000000" when "0010010011100011", -- t[9443] = 0
      "000000" when "0010010011100100", -- t[9444] = 0
      "000000" when "0010010011100101", -- t[9445] = 0
      "000000" when "0010010011100110", -- t[9446] = 0
      "000000" when "0010010011100111", -- t[9447] = 0
      "000000" when "0010010011101000", -- t[9448] = 0
      "000000" when "0010010011101001", -- t[9449] = 0
      "000000" when "0010010011101010", -- t[9450] = 0
      "000000" when "0010010011101011", -- t[9451] = 0
      "000000" when "0010010011101100", -- t[9452] = 0
      "000000" when "0010010011101101", -- t[9453] = 0
      "000000" when "0010010011101110", -- t[9454] = 0
      "000000" when "0010010011101111", -- t[9455] = 0
      "000000" when "0010010011110000", -- t[9456] = 0
      "000000" when "0010010011110001", -- t[9457] = 0
      "000000" when "0010010011110010", -- t[9458] = 0
      "000000" when "0010010011110011", -- t[9459] = 0
      "000000" when "0010010011110100", -- t[9460] = 0
      "000000" when "0010010011110101", -- t[9461] = 0
      "000000" when "0010010011110110", -- t[9462] = 0
      "000000" when "0010010011110111", -- t[9463] = 0
      "000000" when "0010010011111000", -- t[9464] = 0
      "000000" when "0010010011111001", -- t[9465] = 0
      "000000" when "0010010011111010", -- t[9466] = 0
      "000000" when "0010010011111011", -- t[9467] = 0
      "000000" when "0010010011111100", -- t[9468] = 0
      "000000" when "0010010011111101", -- t[9469] = 0
      "000000" when "0010010011111110", -- t[9470] = 0
      "000000" when "0010010011111111", -- t[9471] = 0
      "000000" when "0010010100000000", -- t[9472] = 0
      "000000" when "0010010100000001", -- t[9473] = 0
      "000000" when "0010010100000010", -- t[9474] = 0
      "000000" when "0010010100000011", -- t[9475] = 0
      "000000" when "0010010100000100", -- t[9476] = 0
      "000000" when "0010010100000101", -- t[9477] = 0
      "000000" when "0010010100000110", -- t[9478] = 0
      "000000" when "0010010100000111", -- t[9479] = 0
      "000000" when "0010010100001000", -- t[9480] = 0
      "000000" when "0010010100001001", -- t[9481] = 0
      "000000" when "0010010100001010", -- t[9482] = 0
      "000000" when "0010010100001011", -- t[9483] = 0
      "000000" when "0010010100001100", -- t[9484] = 0
      "000000" when "0010010100001101", -- t[9485] = 0
      "000000" when "0010010100001110", -- t[9486] = 0
      "000000" when "0010010100001111", -- t[9487] = 0
      "000000" when "0010010100010000", -- t[9488] = 0
      "000000" when "0010010100010001", -- t[9489] = 0
      "000000" when "0010010100010010", -- t[9490] = 0
      "000000" when "0010010100010011", -- t[9491] = 0
      "000000" when "0010010100010100", -- t[9492] = 0
      "000000" when "0010010100010101", -- t[9493] = 0
      "000000" when "0010010100010110", -- t[9494] = 0
      "000000" when "0010010100010111", -- t[9495] = 0
      "000000" when "0010010100011000", -- t[9496] = 0
      "000000" when "0010010100011001", -- t[9497] = 0
      "000000" when "0010010100011010", -- t[9498] = 0
      "000000" when "0010010100011011", -- t[9499] = 0
      "000000" when "0010010100011100", -- t[9500] = 0
      "000000" when "0010010100011101", -- t[9501] = 0
      "000000" when "0010010100011110", -- t[9502] = 0
      "000000" when "0010010100011111", -- t[9503] = 0
      "000000" when "0010010100100000", -- t[9504] = 0
      "000000" when "0010010100100001", -- t[9505] = 0
      "000000" when "0010010100100010", -- t[9506] = 0
      "000000" when "0010010100100011", -- t[9507] = 0
      "000000" when "0010010100100100", -- t[9508] = 0
      "000000" when "0010010100100101", -- t[9509] = 0
      "000000" when "0010010100100110", -- t[9510] = 0
      "000000" when "0010010100100111", -- t[9511] = 0
      "000000" when "0010010100101000", -- t[9512] = 0
      "000000" when "0010010100101001", -- t[9513] = 0
      "000000" when "0010010100101010", -- t[9514] = 0
      "000000" when "0010010100101011", -- t[9515] = 0
      "000000" when "0010010100101100", -- t[9516] = 0
      "000000" when "0010010100101101", -- t[9517] = 0
      "000000" when "0010010100101110", -- t[9518] = 0
      "000000" when "0010010100101111", -- t[9519] = 0
      "000000" when "0010010100110000", -- t[9520] = 0
      "000000" when "0010010100110001", -- t[9521] = 0
      "000000" when "0010010100110010", -- t[9522] = 0
      "000000" when "0010010100110011", -- t[9523] = 0
      "000000" when "0010010100110100", -- t[9524] = 0
      "000000" when "0010010100110101", -- t[9525] = 0
      "000000" when "0010010100110110", -- t[9526] = 0
      "000000" when "0010010100110111", -- t[9527] = 0
      "000000" when "0010010100111000", -- t[9528] = 0
      "000000" when "0010010100111001", -- t[9529] = 0
      "000000" when "0010010100111010", -- t[9530] = 0
      "000000" when "0010010100111011", -- t[9531] = 0
      "000000" when "0010010100111100", -- t[9532] = 0
      "000000" when "0010010100111101", -- t[9533] = 0
      "000000" when "0010010100111110", -- t[9534] = 0
      "000000" when "0010010100111111", -- t[9535] = 0
      "000000" when "0010010101000000", -- t[9536] = 0
      "000000" when "0010010101000001", -- t[9537] = 0
      "000000" when "0010010101000010", -- t[9538] = 0
      "000000" when "0010010101000011", -- t[9539] = 0
      "000000" when "0010010101000100", -- t[9540] = 0
      "000000" when "0010010101000101", -- t[9541] = 0
      "000000" when "0010010101000110", -- t[9542] = 0
      "000000" when "0010010101000111", -- t[9543] = 0
      "000000" when "0010010101001000", -- t[9544] = 0
      "000000" when "0010010101001001", -- t[9545] = 0
      "000000" when "0010010101001010", -- t[9546] = 0
      "000000" when "0010010101001011", -- t[9547] = 0
      "000000" when "0010010101001100", -- t[9548] = 0
      "000000" when "0010010101001101", -- t[9549] = 0
      "000000" when "0010010101001110", -- t[9550] = 0
      "000000" when "0010010101001111", -- t[9551] = 0
      "000000" when "0010010101010000", -- t[9552] = 0
      "000000" when "0010010101010001", -- t[9553] = 0
      "000000" when "0010010101010010", -- t[9554] = 0
      "000000" when "0010010101010011", -- t[9555] = 0
      "000000" when "0010010101010100", -- t[9556] = 0
      "000000" when "0010010101010101", -- t[9557] = 0
      "000000" when "0010010101010110", -- t[9558] = 0
      "000000" when "0010010101010111", -- t[9559] = 0
      "000000" when "0010010101011000", -- t[9560] = 0
      "000000" when "0010010101011001", -- t[9561] = 0
      "000000" when "0010010101011010", -- t[9562] = 0
      "000000" when "0010010101011011", -- t[9563] = 0
      "000000" when "0010010101011100", -- t[9564] = 0
      "000000" when "0010010101011101", -- t[9565] = 0
      "000000" when "0010010101011110", -- t[9566] = 0
      "000000" when "0010010101011111", -- t[9567] = 0
      "000000" when "0010010101100000", -- t[9568] = 0
      "000000" when "0010010101100001", -- t[9569] = 0
      "000000" when "0010010101100010", -- t[9570] = 0
      "000000" when "0010010101100011", -- t[9571] = 0
      "000000" when "0010010101100100", -- t[9572] = 0
      "000000" when "0010010101100101", -- t[9573] = 0
      "000000" when "0010010101100110", -- t[9574] = 0
      "000000" when "0010010101100111", -- t[9575] = 0
      "000000" when "0010010101101000", -- t[9576] = 0
      "000000" when "0010010101101001", -- t[9577] = 0
      "000000" when "0010010101101010", -- t[9578] = 0
      "000000" when "0010010101101011", -- t[9579] = 0
      "000000" when "0010010101101100", -- t[9580] = 0
      "000000" when "0010010101101101", -- t[9581] = 0
      "000000" when "0010010101101110", -- t[9582] = 0
      "000000" when "0010010101101111", -- t[9583] = 0
      "000000" when "0010010101110000", -- t[9584] = 0
      "000000" when "0010010101110001", -- t[9585] = 0
      "000000" when "0010010101110010", -- t[9586] = 0
      "000000" when "0010010101110011", -- t[9587] = 0
      "000000" when "0010010101110100", -- t[9588] = 0
      "000000" when "0010010101110101", -- t[9589] = 0
      "000000" when "0010010101110110", -- t[9590] = 0
      "000000" when "0010010101110111", -- t[9591] = 0
      "000000" when "0010010101111000", -- t[9592] = 0
      "000000" when "0010010101111001", -- t[9593] = 0
      "000000" when "0010010101111010", -- t[9594] = 0
      "000000" when "0010010101111011", -- t[9595] = 0
      "000000" when "0010010101111100", -- t[9596] = 0
      "000000" when "0010010101111101", -- t[9597] = 0
      "000000" when "0010010101111110", -- t[9598] = 0
      "000000" when "0010010101111111", -- t[9599] = 0
      "000000" when "0010010110000000", -- t[9600] = 0
      "000000" when "0010010110000001", -- t[9601] = 0
      "000000" when "0010010110000010", -- t[9602] = 0
      "000000" when "0010010110000011", -- t[9603] = 0
      "000000" when "0010010110000100", -- t[9604] = 0
      "000000" when "0010010110000101", -- t[9605] = 0
      "000000" when "0010010110000110", -- t[9606] = 0
      "000000" when "0010010110000111", -- t[9607] = 0
      "000000" when "0010010110001000", -- t[9608] = 0
      "000000" when "0010010110001001", -- t[9609] = 0
      "000000" when "0010010110001010", -- t[9610] = 0
      "000000" when "0010010110001011", -- t[9611] = 0
      "000000" when "0010010110001100", -- t[9612] = 0
      "000000" when "0010010110001101", -- t[9613] = 0
      "000000" when "0010010110001110", -- t[9614] = 0
      "000000" when "0010010110001111", -- t[9615] = 0
      "000000" when "0010010110010000", -- t[9616] = 0
      "000000" when "0010010110010001", -- t[9617] = 0
      "000000" when "0010010110010010", -- t[9618] = 0
      "000000" when "0010010110010011", -- t[9619] = 0
      "000000" when "0010010110010100", -- t[9620] = 0
      "000000" when "0010010110010101", -- t[9621] = 0
      "000000" when "0010010110010110", -- t[9622] = 0
      "000000" when "0010010110010111", -- t[9623] = 0
      "000000" when "0010010110011000", -- t[9624] = 0
      "000000" when "0010010110011001", -- t[9625] = 0
      "000000" when "0010010110011010", -- t[9626] = 0
      "000000" when "0010010110011011", -- t[9627] = 0
      "000000" when "0010010110011100", -- t[9628] = 0
      "000000" when "0010010110011101", -- t[9629] = 0
      "000000" when "0010010110011110", -- t[9630] = 0
      "000000" when "0010010110011111", -- t[9631] = 0
      "000000" when "0010010110100000", -- t[9632] = 0
      "000000" when "0010010110100001", -- t[9633] = 0
      "000000" when "0010010110100010", -- t[9634] = 0
      "000000" when "0010010110100011", -- t[9635] = 0
      "000000" when "0010010110100100", -- t[9636] = 0
      "000000" when "0010010110100101", -- t[9637] = 0
      "000000" when "0010010110100110", -- t[9638] = 0
      "000000" when "0010010110100111", -- t[9639] = 0
      "000000" when "0010010110101000", -- t[9640] = 0
      "000000" when "0010010110101001", -- t[9641] = 0
      "000000" when "0010010110101010", -- t[9642] = 0
      "000000" when "0010010110101011", -- t[9643] = 0
      "000000" when "0010010110101100", -- t[9644] = 0
      "000000" when "0010010110101101", -- t[9645] = 0
      "000000" when "0010010110101110", -- t[9646] = 0
      "000000" when "0010010110101111", -- t[9647] = 0
      "000000" when "0010010110110000", -- t[9648] = 0
      "000000" when "0010010110110001", -- t[9649] = 0
      "000000" when "0010010110110010", -- t[9650] = 0
      "000000" when "0010010110110011", -- t[9651] = 0
      "000000" when "0010010110110100", -- t[9652] = 0
      "000000" when "0010010110110101", -- t[9653] = 0
      "000000" when "0010010110110110", -- t[9654] = 0
      "000000" when "0010010110110111", -- t[9655] = 0
      "000000" when "0010010110111000", -- t[9656] = 0
      "000000" when "0010010110111001", -- t[9657] = 0
      "000000" when "0010010110111010", -- t[9658] = 0
      "000000" when "0010010110111011", -- t[9659] = 0
      "000000" when "0010010110111100", -- t[9660] = 0
      "000000" when "0010010110111101", -- t[9661] = 0
      "000000" when "0010010110111110", -- t[9662] = 0
      "000000" when "0010010110111111", -- t[9663] = 0
      "000000" when "0010010111000000", -- t[9664] = 0
      "000000" when "0010010111000001", -- t[9665] = 0
      "000000" when "0010010111000010", -- t[9666] = 0
      "000000" when "0010010111000011", -- t[9667] = 0
      "000000" when "0010010111000100", -- t[9668] = 0
      "000000" when "0010010111000101", -- t[9669] = 0
      "000000" when "0010010111000110", -- t[9670] = 0
      "000000" when "0010010111000111", -- t[9671] = 0
      "000000" when "0010010111001000", -- t[9672] = 0
      "000000" when "0010010111001001", -- t[9673] = 0
      "000000" when "0010010111001010", -- t[9674] = 0
      "000000" when "0010010111001011", -- t[9675] = 0
      "000000" when "0010010111001100", -- t[9676] = 0
      "000000" when "0010010111001101", -- t[9677] = 0
      "000000" when "0010010111001110", -- t[9678] = 0
      "000000" when "0010010111001111", -- t[9679] = 0
      "000000" when "0010010111010000", -- t[9680] = 0
      "000000" when "0010010111010001", -- t[9681] = 0
      "000000" when "0010010111010010", -- t[9682] = 0
      "000000" when "0010010111010011", -- t[9683] = 0
      "000000" when "0010010111010100", -- t[9684] = 0
      "000000" when "0010010111010101", -- t[9685] = 0
      "000000" when "0010010111010110", -- t[9686] = 0
      "000000" when "0010010111010111", -- t[9687] = 0
      "000000" when "0010010111011000", -- t[9688] = 0
      "000000" when "0010010111011001", -- t[9689] = 0
      "000000" when "0010010111011010", -- t[9690] = 0
      "000000" when "0010010111011011", -- t[9691] = 0
      "000000" when "0010010111011100", -- t[9692] = 0
      "000000" when "0010010111011101", -- t[9693] = 0
      "000000" when "0010010111011110", -- t[9694] = 0
      "000000" when "0010010111011111", -- t[9695] = 0
      "000000" when "0010010111100000", -- t[9696] = 0
      "000000" when "0010010111100001", -- t[9697] = 0
      "000000" when "0010010111100010", -- t[9698] = 0
      "000000" when "0010010111100011", -- t[9699] = 0
      "000000" when "0010010111100100", -- t[9700] = 0
      "000000" when "0010010111100101", -- t[9701] = 0
      "000000" when "0010010111100110", -- t[9702] = 0
      "000000" when "0010010111100111", -- t[9703] = 0
      "000000" when "0010010111101000", -- t[9704] = 0
      "000000" when "0010010111101001", -- t[9705] = 0
      "000000" when "0010010111101010", -- t[9706] = 0
      "000000" when "0010010111101011", -- t[9707] = 0
      "000000" when "0010010111101100", -- t[9708] = 0
      "000000" when "0010010111101101", -- t[9709] = 0
      "000000" when "0010010111101110", -- t[9710] = 0
      "000000" when "0010010111101111", -- t[9711] = 0
      "000000" when "0010010111110000", -- t[9712] = 0
      "000000" when "0010010111110001", -- t[9713] = 0
      "000000" when "0010010111110010", -- t[9714] = 0
      "000000" when "0010010111110011", -- t[9715] = 0
      "000000" when "0010010111110100", -- t[9716] = 0
      "000000" when "0010010111110101", -- t[9717] = 0
      "000000" when "0010010111110110", -- t[9718] = 0
      "000000" when "0010010111110111", -- t[9719] = 0
      "000000" when "0010010111111000", -- t[9720] = 0
      "000000" when "0010010111111001", -- t[9721] = 0
      "000000" when "0010010111111010", -- t[9722] = 0
      "000000" when "0010010111111011", -- t[9723] = 0
      "000000" when "0010010111111100", -- t[9724] = 0
      "000000" when "0010010111111101", -- t[9725] = 0
      "000000" when "0010010111111110", -- t[9726] = 0
      "000000" when "0010010111111111", -- t[9727] = 0
      "000000" when "0010011000000000", -- t[9728] = 0
      "000000" when "0010011000000001", -- t[9729] = 0
      "000000" when "0010011000000010", -- t[9730] = 0
      "000000" when "0010011000000011", -- t[9731] = 0
      "000000" when "0010011000000100", -- t[9732] = 0
      "000000" when "0010011000000101", -- t[9733] = 0
      "000000" when "0010011000000110", -- t[9734] = 0
      "000000" when "0010011000000111", -- t[9735] = 0
      "000000" when "0010011000001000", -- t[9736] = 0
      "000000" when "0010011000001001", -- t[9737] = 0
      "000000" when "0010011000001010", -- t[9738] = 0
      "000000" when "0010011000001011", -- t[9739] = 0
      "000000" when "0010011000001100", -- t[9740] = 0
      "000000" when "0010011000001101", -- t[9741] = 0
      "000000" when "0010011000001110", -- t[9742] = 0
      "000000" when "0010011000001111", -- t[9743] = 0
      "000000" when "0010011000010000", -- t[9744] = 0
      "000000" when "0010011000010001", -- t[9745] = 0
      "000000" when "0010011000010010", -- t[9746] = 0
      "000000" when "0010011000010011", -- t[9747] = 0
      "000000" when "0010011000010100", -- t[9748] = 0
      "000000" when "0010011000010101", -- t[9749] = 0
      "000000" when "0010011000010110", -- t[9750] = 0
      "000000" when "0010011000010111", -- t[9751] = 0
      "000000" when "0010011000011000", -- t[9752] = 0
      "000000" when "0010011000011001", -- t[9753] = 0
      "000000" when "0010011000011010", -- t[9754] = 0
      "000000" when "0010011000011011", -- t[9755] = 0
      "000000" when "0010011000011100", -- t[9756] = 0
      "000000" when "0010011000011101", -- t[9757] = 0
      "000000" when "0010011000011110", -- t[9758] = 0
      "000000" when "0010011000011111", -- t[9759] = 0
      "000000" when "0010011000100000", -- t[9760] = 0
      "000000" when "0010011000100001", -- t[9761] = 0
      "000000" when "0010011000100010", -- t[9762] = 0
      "000000" when "0010011000100011", -- t[9763] = 0
      "000000" when "0010011000100100", -- t[9764] = 0
      "000000" when "0010011000100101", -- t[9765] = 0
      "000000" when "0010011000100110", -- t[9766] = 0
      "000000" when "0010011000100111", -- t[9767] = 0
      "000000" when "0010011000101000", -- t[9768] = 0
      "000000" when "0010011000101001", -- t[9769] = 0
      "000000" when "0010011000101010", -- t[9770] = 0
      "000000" when "0010011000101011", -- t[9771] = 0
      "000000" when "0010011000101100", -- t[9772] = 0
      "000000" when "0010011000101101", -- t[9773] = 0
      "000000" when "0010011000101110", -- t[9774] = 0
      "000000" when "0010011000101111", -- t[9775] = 0
      "000000" when "0010011000110000", -- t[9776] = 0
      "000000" when "0010011000110001", -- t[9777] = 0
      "000000" when "0010011000110010", -- t[9778] = 0
      "000000" when "0010011000110011", -- t[9779] = 0
      "000000" when "0010011000110100", -- t[9780] = 0
      "000000" when "0010011000110101", -- t[9781] = 0
      "000000" when "0010011000110110", -- t[9782] = 0
      "000000" when "0010011000110111", -- t[9783] = 0
      "000000" when "0010011000111000", -- t[9784] = 0
      "000000" when "0010011000111001", -- t[9785] = 0
      "000000" when "0010011000111010", -- t[9786] = 0
      "000000" when "0010011000111011", -- t[9787] = 0
      "000000" when "0010011000111100", -- t[9788] = 0
      "000000" when "0010011000111101", -- t[9789] = 0
      "000000" when "0010011000111110", -- t[9790] = 0
      "000000" when "0010011000111111", -- t[9791] = 0
      "000000" when "0010011001000000", -- t[9792] = 0
      "000000" when "0010011001000001", -- t[9793] = 0
      "000000" when "0010011001000010", -- t[9794] = 0
      "000000" when "0010011001000011", -- t[9795] = 0
      "000000" when "0010011001000100", -- t[9796] = 0
      "000000" when "0010011001000101", -- t[9797] = 0
      "000000" when "0010011001000110", -- t[9798] = 0
      "000000" when "0010011001000111", -- t[9799] = 0
      "000000" when "0010011001001000", -- t[9800] = 0
      "000000" when "0010011001001001", -- t[9801] = 0
      "000000" when "0010011001001010", -- t[9802] = 0
      "000000" when "0010011001001011", -- t[9803] = 0
      "000000" when "0010011001001100", -- t[9804] = 0
      "000000" when "0010011001001101", -- t[9805] = 0
      "000000" when "0010011001001110", -- t[9806] = 0
      "000000" when "0010011001001111", -- t[9807] = 0
      "000000" when "0010011001010000", -- t[9808] = 0
      "000000" when "0010011001010001", -- t[9809] = 0
      "000000" when "0010011001010010", -- t[9810] = 0
      "000000" when "0010011001010011", -- t[9811] = 0
      "000000" when "0010011001010100", -- t[9812] = 0
      "000000" when "0010011001010101", -- t[9813] = 0
      "000000" when "0010011001010110", -- t[9814] = 0
      "000000" when "0010011001010111", -- t[9815] = 0
      "000000" when "0010011001011000", -- t[9816] = 0
      "000000" when "0010011001011001", -- t[9817] = 0
      "000000" when "0010011001011010", -- t[9818] = 0
      "000000" when "0010011001011011", -- t[9819] = 0
      "000000" when "0010011001011100", -- t[9820] = 0
      "000000" when "0010011001011101", -- t[9821] = 0
      "000000" when "0010011001011110", -- t[9822] = 0
      "000000" when "0010011001011111", -- t[9823] = 0
      "000000" when "0010011001100000", -- t[9824] = 0
      "000000" when "0010011001100001", -- t[9825] = 0
      "000000" when "0010011001100010", -- t[9826] = 0
      "000000" when "0010011001100011", -- t[9827] = 0
      "000000" when "0010011001100100", -- t[9828] = 0
      "000000" when "0010011001100101", -- t[9829] = 0
      "000000" when "0010011001100110", -- t[9830] = 0
      "000000" when "0010011001100111", -- t[9831] = 0
      "000000" when "0010011001101000", -- t[9832] = 0
      "000000" when "0010011001101001", -- t[9833] = 0
      "000000" when "0010011001101010", -- t[9834] = 0
      "000000" when "0010011001101011", -- t[9835] = 0
      "000000" when "0010011001101100", -- t[9836] = 0
      "000000" when "0010011001101101", -- t[9837] = 0
      "000000" when "0010011001101110", -- t[9838] = 0
      "000000" when "0010011001101111", -- t[9839] = 0
      "000000" when "0010011001110000", -- t[9840] = 0
      "000000" when "0010011001110001", -- t[9841] = 0
      "000000" when "0010011001110010", -- t[9842] = 0
      "000000" when "0010011001110011", -- t[9843] = 0
      "000000" when "0010011001110100", -- t[9844] = 0
      "000000" when "0010011001110101", -- t[9845] = 0
      "000000" when "0010011001110110", -- t[9846] = 0
      "000000" when "0010011001110111", -- t[9847] = 0
      "000000" when "0010011001111000", -- t[9848] = 0
      "000000" when "0010011001111001", -- t[9849] = 0
      "000000" when "0010011001111010", -- t[9850] = 0
      "000000" when "0010011001111011", -- t[9851] = 0
      "000000" when "0010011001111100", -- t[9852] = 0
      "000000" when "0010011001111101", -- t[9853] = 0
      "000000" when "0010011001111110", -- t[9854] = 0
      "000000" when "0010011001111111", -- t[9855] = 0
      "000000" when "0010011010000000", -- t[9856] = 0
      "000000" when "0010011010000001", -- t[9857] = 0
      "000000" when "0010011010000010", -- t[9858] = 0
      "000000" when "0010011010000011", -- t[9859] = 0
      "000000" when "0010011010000100", -- t[9860] = 0
      "000000" when "0010011010000101", -- t[9861] = 0
      "000000" when "0010011010000110", -- t[9862] = 0
      "000000" when "0010011010000111", -- t[9863] = 0
      "000000" when "0010011010001000", -- t[9864] = 0
      "000000" when "0010011010001001", -- t[9865] = 0
      "000000" when "0010011010001010", -- t[9866] = 0
      "000000" when "0010011010001011", -- t[9867] = 0
      "000000" when "0010011010001100", -- t[9868] = 0
      "000000" when "0010011010001101", -- t[9869] = 0
      "000000" when "0010011010001110", -- t[9870] = 0
      "000000" when "0010011010001111", -- t[9871] = 0
      "000000" when "0010011010010000", -- t[9872] = 0
      "000000" when "0010011010010001", -- t[9873] = 0
      "000000" when "0010011010010010", -- t[9874] = 0
      "000000" when "0010011010010011", -- t[9875] = 0
      "000000" when "0010011010010100", -- t[9876] = 0
      "000000" when "0010011010010101", -- t[9877] = 0
      "000000" when "0010011010010110", -- t[9878] = 0
      "000000" when "0010011010010111", -- t[9879] = 0
      "000000" when "0010011010011000", -- t[9880] = 0
      "000000" when "0010011010011001", -- t[9881] = 0
      "000000" when "0010011010011010", -- t[9882] = 0
      "000000" when "0010011010011011", -- t[9883] = 0
      "000000" when "0010011010011100", -- t[9884] = 0
      "000000" when "0010011010011101", -- t[9885] = 0
      "000000" when "0010011010011110", -- t[9886] = 0
      "000000" when "0010011010011111", -- t[9887] = 0
      "000000" when "0010011010100000", -- t[9888] = 0
      "000000" when "0010011010100001", -- t[9889] = 0
      "000000" when "0010011010100010", -- t[9890] = 0
      "000000" when "0010011010100011", -- t[9891] = 0
      "000000" when "0010011010100100", -- t[9892] = 0
      "000000" when "0010011010100101", -- t[9893] = 0
      "000000" when "0010011010100110", -- t[9894] = 0
      "000000" when "0010011010100111", -- t[9895] = 0
      "000000" when "0010011010101000", -- t[9896] = 0
      "000000" when "0010011010101001", -- t[9897] = 0
      "000000" when "0010011010101010", -- t[9898] = 0
      "000000" when "0010011010101011", -- t[9899] = 0
      "000000" when "0010011010101100", -- t[9900] = 0
      "000000" when "0010011010101101", -- t[9901] = 0
      "000000" when "0010011010101110", -- t[9902] = 0
      "000000" when "0010011010101111", -- t[9903] = 0
      "000000" when "0010011010110000", -- t[9904] = 0
      "000000" when "0010011010110001", -- t[9905] = 0
      "000000" when "0010011010110010", -- t[9906] = 0
      "000000" when "0010011010110011", -- t[9907] = 0
      "000000" when "0010011010110100", -- t[9908] = 0
      "000000" when "0010011010110101", -- t[9909] = 0
      "000000" when "0010011010110110", -- t[9910] = 0
      "000000" when "0010011010110111", -- t[9911] = 0
      "000000" when "0010011010111000", -- t[9912] = 0
      "000000" when "0010011010111001", -- t[9913] = 0
      "000000" when "0010011010111010", -- t[9914] = 0
      "000000" when "0010011010111011", -- t[9915] = 0
      "000000" when "0010011010111100", -- t[9916] = 0
      "000000" when "0010011010111101", -- t[9917] = 0
      "000000" when "0010011010111110", -- t[9918] = 0
      "000000" when "0010011010111111", -- t[9919] = 0
      "000000" when "0010011011000000", -- t[9920] = 0
      "000000" when "0010011011000001", -- t[9921] = 0
      "000000" when "0010011011000010", -- t[9922] = 0
      "000000" when "0010011011000011", -- t[9923] = 0
      "000000" when "0010011011000100", -- t[9924] = 0
      "000000" when "0010011011000101", -- t[9925] = 0
      "000000" when "0010011011000110", -- t[9926] = 0
      "000000" when "0010011011000111", -- t[9927] = 0
      "000000" when "0010011011001000", -- t[9928] = 0
      "000000" when "0010011011001001", -- t[9929] = 0
      "000000" when "0010011011001010", -- t[9930] = 0
      "000000" when "0010011011001011", -- t[9931] = 0
      "000000" when "0010011011001100", -- t[9932] = 0
      "000000" when "0010011011001101", -- t[9933] = 0
      "000000" when "0010011011001110", -- t[9934] = 0
      "000000" when "0010011011001111", -- t[9935] = 0
      "000000" when "0010011011010000", -- t[9936] = 0
      "000000" when "0010011011010001", -- t[9937] = 0
      "000000" when "0010011011010010", -- t[9938] = 0
      "000000" when "0010011011010011", -- t[9939] = 0
      "000000" when "0010011011010100", -- t[9940] = 0
      "000000" when "0010011011010101", -- t[9941] = 0
      "000000" when "0010011011010110", -- t[9942] = 0
      "000000" when "0010011011010111", -- t[9943] = 0
      "000000" when "0010011011011000", -- t[9944] = 0
      "000000" when "0010011011011001", -- t[9945] = 0
      "000000" when "0010011011011010", -- t[9946] = 0
      "000000" when "0010011011011011", -- t[9947] = 0
      "000000" when "0010011011011100", -- t[9948] = 0
      "000000" when "0010011011011101", -- t[9949] = 0
      "000000" when "0010011011011110", -- t[9950] = 0
      "000000" when "0010011011011111", -- t[9951] = 0
      "000000" when "0010011011100000", -- t[9952] = 0
      "000000" when "0010011011100001", -- t[9953] = 0
      "000000" when "0010011011100010", -- t[9954] = 0
      "000000" when "0010011011100011", -- t[9955] = 0
      "000000" when "0010011011100100", -- t[9956] = 0
      "000000" when "0010011011100101", -- t[9957] = 0
      "000000" when "0010011011100110", -- t[9958] = 0
      "000000" when "0010011011100111", -- t[9959] = 0
      "000000" when "0010011011101000", -- t[9960] = 0
      "000000" when "0010011011101001", -- t[9961] = 0
      "000000" when "0010011011101010", -- t[9962] = 0
      "000000" when "0010011011101011", -- t[9963] = 0
      "000000" when "0010011011101100", -- t[9964] = 0
      "000000" when "0010011011101101", -- t[9965] = 0
      "000000" when "0010011011101110", -- t[9966] = 0
      "000000" when "0010011011101111", -- t[9967] = 0
      "000000" when "0010011011110000", -- t[9968] = 0
      "000000" when "0010011011110001", -- t[9969] = 0
      "000000" when "0010011011110010", -- t[9970] = 0
      "000000" when "0010011011110011", -- t[9971] = 0
      "000000" when "0010011011110100", -- t[9972] = 0
      "000000" when "0010011011110101", -- t[9973] = 0
      "000000" when "0010011011110110", -- t[9974] = 0
      "000000" when "0010011011110111", -- t[9975] = 0
      "000000" when "0010011011111000", -- t[9976] = 0
      "000000" when "0010011011111001", -- t[9977] = 0
      "000000" when "0010011011111010", -- t[9978] = 0
      "000000" when "0010011011111011", -- t[9979] = 0
      "000000" when "0010011011111100", -- t[9980] = 0
      "000000" when "0010011011111101", -- t[9981] = 0
      "000000" when "0010011011111110", -- t[9982] = 0
      "000000" when "0010011011111111", -- t[9983] = 0
      "000000" when "0010011100000000", -- t[9984] = 0
      "000000" when "0010011100000001", -- t[9985] = 0
      "000000" when "0010011100000010", -- t[9986] = 0
      "000000" when "0010011100000011", -- t[9987] = 0
      "000000" when "0010011100000100", -- t[9988] = 0
      "000000" when "0010011100000101", -- t[9989] = 0
      "000000" when "0010011100000110", -- t[9990] = 0
      "000000" when "0010011100000111", -- t[9991] = 0
      "000000" when "0010011100001000", -- t[9992] = 0
      "000000" when "0010011100001001", -- t[9993] = 0
      "000000" when "0010011100001010", -- t[9994] = 0
      "000000" when "0010011100001011", -- t[9995] = 0
      "000000" when "0010011100001100", -- t[9996] = 0
      "000000" when "0010011100001101", -- t[9997] = 0
      "000000" when "0010011100001110", -- t[9998] = 0
      "000000" when "0010011100001111", -- t[9999] = 0
      "000000" when "0010011100010000", -- t[10000] = 0
      "000000" when "0010011100010001", -- t[10001] = 0
      "000000" when "0010011100010010", -- t[10002] = 0
      "000000" when "0010011100010011", -- t[10003] = 0
      "000000" when "0010011100010100", -- t[10004] = 0
      "000000" when "0010011100010101", -- t[10005] = 0
      "000000" when "0010011100010110", -- t[10006] = 0
      "000000" when "0010011100010111", -- t[10007] = 0
      "000000" when "0010011100011000", -- t[10008] = 0
      "000000" when "0010011100011001", -- t[10009] = 0
      "000000" when "0010011100011010", -- t[10010] = 0
      "000000" when "0010011100011011", -- t[10011] = 0
      "000000" when "0010011100011100", -- t[10012] = 0
      "000000" when "0010011100011101", -- t[10013] = 0
      "000000" when "0010011100011110", -- t[10014] = 0
      "000000" when "0010011100011111", -- t[10015] = 0
      "000000" when "0010011100100000", -- t[10016] = 0
      "000000" when "0010011100100001", -- t[10017] = 0
      "000000" when "0010011100100010", -- t[10018] = 0
      "000000" when "0010011100100011", -- t[10019] = 0
      "000000" when "0010011100100100", -- t[10020] = 0
      "000000" when "0010011100100101", -- t[10021] = 0
      "000000" when "0010011100100110", -- t[10022] = 0
      "000000" when "0010011100100111", -- t[10023] = 0
      "000000" when "0010011100101000", -- t[10024] = 0
      "000000" when "0010011100101001", -- t[10025] = 0
      "000000" when "0010011100101010", -- t[10026] = 0
      "000000" when "0010011100101011", -- t[10027] = 0
      "000000" when "0010011100101100", -- t[10028] = 0
      "000000" when "0010011100101101", -- t[10029] = 0
      "000000" when "0010011100101110", -- t[10030] = 0
      "000000" when "0010011100101111", -- t[10031] = 0
      "000000" when "0010011100110000", -- t[10032] = 0
      "000000" when "0010011100110001", -- t[10033] = 0
      "000000" when "0010011100110010", -- t[10034] = 0
      "000000" when "0010011100110011", -- t[10035] = 0
      "000000" when "0010011100110100", -- t[10036] = 0
      "000000" when "0010011100110101", -- t[10037] = 0
      "000000" when "0010011100110110", -- t[10038] = 0
      "000000" when "0010011100110111", -- t[10039] = 0
      "000000" when "0010011100111000", -- t[10040] = 0
      "000000" when "0010011100111001", -- t[10041] = 0
      "000000" when "0010011100111010", -- t[10042] = 0
      "000000" when "0010011100111011", -- t[10043] = 0
      "000000" when "0010011100111100", -- t[10044] = 0
      "000000" when "0010011100111101", -- t[10045] = 0
      "000000" when "0010011100111110", -- t[10046] = 0
      "000000" when "0010011100111111", -- t[10047] = 0
      "000000" when "0010011101000000", -- t[10048] = 0
      "000000" when "0010011101000001", -- t[10049] = 0
      "000000" when "0010011101000010", -- t[10050] = 0
      "000000" when "0010011101000011", -- t[10051] = 0
      "000000" when "0010011101000100", -- t[10052] = 0
      "000000" when "0010011101000101", -- t[10053] = 0
      "000000" when "0010011101000110", -- t[10054] = 0
      "000000" when "0010011101000111", -- t[10055] = 0
      "000000" when "0010011101001000", -- t[10056] = 0
      "000000" when "0010011101001001", -- t[10057] = 0
      "000000" when "0010011101001010", -- t[10058] = 0
      "000000" when "0010011101001011", -- t[10059] = 0
      "000000" when "0010011101001100", -- t[10060] = 0
      "000000" when "0010011101001101", -- t[10061] = 0
      "000000" when "0010011101001110", -- t[10062] = 0
      "000000" when "0010011101001111", -- t[10063] = 0
      "000000" when "0010011101010000", -- t[10064] = 0
      "000000" when "0010011101010001", -- t[10065] = 0
      "000000" when "0010011101010010", -- t[10066] = 0
      "000000" when "0010011101010011", -- t[10067] = 0
      "000000" when "0010011101010100", -- t[10068] = 0
      "000000" when "0010011101010101", -- t[10069] = 0
      "000000" when "0010011101010110", -- t[10070] = 0
      "000000" when "0010011101010111", -- t[10071] = 0
      "000000" when "0010011101011000", -- t[10072] = 0
      "000000" when "0010011101011001", -- t[10073] = 0
      "000000" when "0010011101011010", -- t[10074] = 0
      "000000" when "0010011101011011", -- t[10075] = 0
      "000000" when "0010011101011100", -- t[10076] = 0
      "000000" when "0010011101011101", -- t[10077] = 0
      "000000" when "0010011101011110", -- t[10078] = 0
      "000000" when "0010011101011111", -- t[10079] = 0
      "000000" when "0010011101100000", -- t[10080] = 0
      "000000" when "0010011101100001", -- t[10081] = 0
      "000000" when "0010011101100010", -- t[10082] = 0
      "000000" when "0010011101100011", -- t[10083] = 0
      "000000" when "0010011101100100", -- t[10084] = 0
      "000000" when "0010011101100101", -- t[10085] = 0
      "000000" when "0010011101100110", -- t[10086] = 0
      "000000" when "0010011101100111", -- t[10087] = 0
      "000000" when "0010011101101000", -- t[10088] = 0
      "000000" when "0010011101101001", -- t[10089] = 0
      "000000" when "0010011101101010", -- t[10090] = 0
      "000000" when "0010011101101011", -- t[10091] = 0
      "000000" when "0010011101101100", -- t[10092] = 0
      "000000" when "0010011101101101", -- t[10093] = 0
      "000000" when "0010011101101110", -- t[10094] = 0
      "000000" when "0010011101101111", -- t[10095] = 0
      "000000" when "0010011101110000", -- t[10096] = 0
      "000000" when "0010011101110001", -- t[10097] = 0
      "000000" when "0010011101110010", -- t[10098] = 0
      "000000" when "0010011101110011", -- t[10099] = 0
      "000000" when "0010011101110100", -- t[10100] = 0
      "000000" when "0010011101110101", -- t[10101] = 0
      "000000" when "0010011101110110", -- t[10102] = 0
      "000000" when "0010011101110111", -- t[10103] = 0
      "000000" when "0010011101111000", -- t[10104] = 0
      "000000" when "0010011101111001", -- t[10105] = 0
      "000000" when "0010011101111010", -- t[10106] = 0
      "000000" when "0010011101111011", -- t[10107] = 0
      "000000" when "0010011101111100", -- t[10108] = 0
      "000000" when "0010011101111101", -- t[10109] = 0
      "000000" when "0010011101111110", -- t[10110] = 0
      "000000" when "0010011101111111", -- t[10111] = 0
      "000000" when "0010011110000000", -- t[10112] = 0
      "000000" when "0010011110000001", -- t[10113] = 0
      "000000" when "0010011110000010", -- t[10114] = 0
      "000000" when "0010011110000011", -- t[10115] = 0
      "000000" when "0010011110000100", -- t[10116] = 0
      "000000" when "0010011110000101", -- t[10117] = 0
      "000000" when "0010011110000110", -- t[10118] = 0
      "000000" when "0010011110000111", -- t[10119] = 0
      "000000" when "0010011110001000", -- t[10120] = 0
      "000000" when "0010011110001001", -- t[10121] = 0
      "000001" when "0010011110001010", -- t[10122] = 1
      "000001" when "0010011110001011", -- t[10123] = 1
      "000001" when "0010011110001100", -- t[10124] = 1
      "000001" when "0010011110001101", -- t[10125] = 1
      "000001" when "0010011110001110", -- t[10126] = 1
      "000001" when "0010011110001111", -- t[10127] = 1
      "000001" when "0010011110010000", -- t[10128] = 1
      "000001" when "0010011110010001", -- t[10129] = 1
      "000001" when "0010011110010010", -- t[10130] = 1
      "000001" when "0010011110010011", -- t[10131] = 1
      "000001" when "0010011110010100", -- t[10132] = 1
      "000001" when "0010011110010101", -- t[10133] = 1
      "000001" when "0010011110010110", -- t[10134] = 1
      "000001" when "0010011110010111", -- t[10135] = 1
      "000001" when "0010011110011000", -- t[10136] = 1
      "000001" when "0010011110011001", -- t[10137] = 1
      "000001" when "0010011110011010", -- t[10138] = 1
      "000001" when "0010011110011011", -- t[10139] = 1
      "000001" when "0010011110011100", -- t[10140] = 1
      "000001" when "0010011110011101", -- t[10141] = 1
      "000001" when "0010011110011110", -- t[10142] = 1
      "000001" when "0010011110011111", -- t[10143] = 1
      "000001" when "0010011110100000", -- t[10144] = 1
      "000001" when "0010011110100001", -- t[10145] = 1
      "000001" when "0010011110100010", -- t[10146] = 1
      "000001" when "0010011110100011", -- t[10147] = 1
      "000001" when "0010011110100100", -- t[10148] = 1
      "000001" when "0010011110100101", -- t[10149] = 1
      "000001" when "0010011110100110", -- t[10150] = 1
      "000001" when "0010011110100111", -- t[10151] = 1
      "000001" when "0010011110101000", -- t[10152] = 1
      "000001" when "0010011110101001", -- t[10153] = 1
      "000001" when "0010011110101010", -- t[10154] = 1
      "000001" when "0010011110101011", -- t[10155] = 1
      "000001" when "0010011110101100", -- t[10156] = 1
      "000001" when "0010011110101101", -- t[10157] = 1
      "000001" when "0010011110101110", -- t[10158] = 1
      "000001" when "0010011110101111", -- t[10159] = 1
      "000001" when "0010011110110000", -- t[10160] = 1
      "000001" when "0010011110110001", -- t[10161] = 1
      "000001" when "0010011110110010", -- t[10162] = 1
      "000001" when "0010011110110011", -- t[10163] = 1
      "000001" when "0010011110110100", -- t[10164] = 1
      "000001" when "0010011110110101", -- t[10165] = 1
      "000001" when "0010011110110110", -- t[10166] = 1
      "000001" when "0010011110110111", -- t[10167] = 1
      "000001" when "0010011110111000", -- t[10168] = 1
      "000001" when "0010011110111001", -- t[10169] = 1
      "000001" when "0010011110111010", -- t[10170] = 1
      "000001" when "0010011110111011", -- t[10171] = 1
      "000001" when "0010011110111100", -- t[10172] = 1
      "000001" when "0010011110111101", -- t[10173] = 1
      "000001" when "0010011110111110", -- t[10174] = 1
      "000001" when "0010011110111111", -- t[10175] = 1
      "000001" when "0010011111000000", -- t[10176] = 1
      "000001" when "0010011111000001", -- t[10177] = 1
      "000001" when "0010011111000010", -- t[10178] = 1
      "000001" when "0010011111000011", -- t[10179] = 1
      "000001" when "0010011111000100", -- t[10180] = 1
      "000001" when "0010011111000101", -- t[10181] = 1
      "000001" when "0010011111000110", -- t[10182] = 1
      "000001" when "0010011111000111", -- t[10183] = 1
      "000001" when "0010011111001000", -- t[10184] = 1
      "000001" when "0010011111001001", -- t[10185] = 1
      "000001" when "0010011111001010", -- t[10186] = 1
      "000001" when "0010011111001011", -- t[10187] = 1
      "000001" when "0010011111001100", -- t[10188] = 1
      "000001" when "0010011111001101", -- t[10189] = 1
      "000001" when "0010011111001110", -- t[10190] = 1
      "000001" when "0010011111001111", -- t[10191] = 1
      "000001" when "0010011111010000", -- t[10192] = 1
      "000001" when "0010011111010001", -- t[10193] = 1
      "000001" when "0010011111010010", -- t[10194] = 1
      "000001" when "0010011111010011", -- t[10195] = 1
      "000001" when "0010011111010100", -- t[10196] = 1
      "000001" when "0010011111010101", -- t[10197] = 1
      "000001" when "0010011111010110", -- t[10198] = 1
      "000001" when "0010011111010111", -- t[10199] = 1
      "000001" when "0010011111011000", -- t[10200] = 1
      "000001" when "0010011111011001", -- t[10201] = 1
      "000001" when "0010011111011010", -- t[10202] = 1
      "000001" when "0010011111011011", -- t[10203] = 1
      "000001" when "0010011111011100", -- t[10204] = 1
      "000001" when "0010011111011101", -- t[10205] = 1
      "000001" when "0010011111011110", -- t[10206] = 1
      "000001" when "0010011111011111", -- t[10207] = 1
      "000001" when "0010011111100000", -- t[10208] = 1
      "000001" when "0010011111100001", -- t[10209] = 1
      "000001" when "0010011111100010", -- t[10210] = 1
      "000001" when "0010011111100011", -- t[10211] = 1
      "000001" when "0010011111100100", -- t[10212] = 1
      "000001" when "0010011111100101", -- t[10213] = 1
      "000001" when "0010011111100110", -- t[10214] = 1
      "000001" when "0010011111100111", -- t[10215] = 1
      "000001" when "0010011111101000", -- t[10216] = 1
      "000001" when "0010011111101001", -- t[10217] = 1
      "000001" when "0010011111101010", -- t[10218] = 1
      "000001" when "0010011111101011", -- t[10219] = 1
      "000001" when "0010011111101100", -- t[10220] = 1
      "000001" when "0010011111101101", -- t[10221] = 1
      "000001" when "0010011111101110", -- t[10222] = 1
      "000001" when "0010011111101111", -- t[10223] = 1
      "000001" when "0010011111110000", -- t[10224] = 1
      "000001" when "0010011111110001", -- t[10225] = 1
      "000001" when "0010011111110010", -- t[10226] = 1
      "000001" when "0010011111110011", -- t[10227] = 1
      "000001" when "0010011111110100", -- t[10228] = 1
      "000001" when "0010011111110101", -- t[10229] = 1
      "000001" when "0010011111110110", -- t[10230] = 1
      "000001" when "0010011111110111", -- t[10231] = 1
      "000001" when "0010011111111000", -- t[10232] = 1
      "000001" when "0010011111111001", -- t[10233] = 1
      "000001" when "0010011111111010", -- t[10234] = 1
      "000001" when "0010011111111011", -- t[10235] = 1
      "000001" when "0010011111111100", -- t[10236] = 1
      "000001" when "0010011111111101", -- t[10237] = 1
      "000001" when "0010011111111110", -- t[10238] = 1
      "000001" when "0010011111111111", -- t[10239] = 1
      "000001" when "0010100000000000", -- t[10240] = 1
      "000001" when "0010100000000001", -- t[10241] = 1
      "000001" when "0010100000000010", -- t[10242] = 1
      "000001" when "0010100000000011", -- t[10243] = 1
      "000001" when "0010100000000100", -- t[10244] = 1
      "000001" when "0010100000000101", -- t[10245] = 1
      "000001" when "0010100000000110", -- t[10246] = 1
      "000001" when "0010100000000111", -- t[10247] = 1
      "000001" when "0010100000001000", -- t[10248] = 1
      "000001" when "0010100000001001", -- t[10249] = 1
      "000001" when "0010100000001010", -- t[10250] = 1
      "000001" when "0010100000001011", -- t[10251] = 1
      "000001" when "0010100000001100", -- t[10252] = 1
      "000001" when "0010100000001101", -- t[10253] = 1
      "000001" when "0010100000001110", -- t[10254] = 1
      "000001" when "0010100000001111", -- t[10255] = 1
      "000001" when "0010100000010000", -- t[10256] = 1
      "000001" when "0010100000010001", -- t[10257] = 1
      "000001" when "0010100000010010", -- t[10258] = 1
      "000001" when "0010100000010011", -- t[10259] = 1
      "000001" when "0010100000010100", -- t[10260] = 1
      "000001" when "0010100000010101", -- t[10261] = 1
      "000001" when "0010100000010110", -- t[10262] = 1
      "000001" when "0010100000010111", -- t[10263] = 1
      "000001" when "0010100000011000", -- t[10264] = 1
      "000001" when "0010100000011001", -- t[10265] = 1
      "000001" when "0010100000011010", -- t[10266] = 1
      "000001" when "0010100000011011", -- t[10267] = 1
      "000001" when "0010100000011100", -- t[10268] = 1
      "000001" when "0010100000011101", -- t[10269] = 1
      "000001" when "0010100000011110", -- t[10270] = 1
      "000001" when "0010100000011111", -- t[10271] = 1
      "000001" when "0010100000100000", -- t[10272] = 1
      "000001" when "0010100000100001", -- t[10273] = 1
      "000001" when "0010100000100010", -- t[10274] = 1
      "000001" when "0010100000100011", -- t[10275] = 1
      "000001" when "0010100000100100", -- t[10276] = 1
      "000001" when "0010100000100101", -- t[10277] = 1
      "000001" when "0010100000100110", -- t[10278] = 1
      "000001" when "0010100000100111", -- t[10279] = 1
      "000001" when "0010100000101000", -- t[10280] = 1
      "000001" when "0010100000101001", -- t[10281] = 1
      "000001" when "0010100000101010", -- t[10282] = 1
      "000001" when "0010100000101011", -- t[10283] = 1
      "000001" when "0010100000101100", -- t[10284] = 1
      "000001" when "0010100000101101", -- t[10285] = 1
      "000001" when "0010100000101110", -- t[10286] = 1
      "000001" when "0010100000101111", -- t[10287] = 1
      "000001" when "0010100000110000", -- t[10288] = 1
      "000001" when "0010100000110001", -- t[10289] = 1
      "000001" when "0010100000110010", -- t[10290] = 1
      "000001" when "0010100000110011", -- t[10291] = 1
      "000001" when "0010100000110100", -- t[10292] = 1
      "000001" when "0010100000110101", -- t[10293] = 1
      "000001" when "0010100000110110", -- t[10294] = 1
      "000001" when "0010100000110111", -- t[10295] = 1
      "000001" when "0010100000111000", -- t[10296] = 1
      "000001" when "0010100000111001", -- t[10297] = 1
      "000001" when "0010100000111010", -- t[10298] = 1
      "000001" when "0010100000111011", -- t[10299] = 1
      "000001" when "0010100000111100", -- t[10300] = 1
      "000001" when "0010100000111101", -- t[10301] = 1
      "000001" when "0010100000111110", -- t[10302] = 1
      "000001" when "0010100000111111", -- t[10303] = 1
      "000001" when "0010100001000000", -- t[10304] = 1
      "000001" when "0010100001000001", -- t[10305] = 1
      "000001" when "0010100001000010", -- t[10306] = 1
      "000001" when "0010100001000011", -- t[10307] = 1
      "000001" when "0010100001000100", -- t[10308] = 1
      "000001" when "0010100001000101", -- t[10309] = 1
      "000001" when "0010100001000110", -- t[10310] = 1
      "000001" when "0010100001000111", -- t[10311] = 1
      "000001" when "0010100001001000", -- t[10312] = 1
      "000001" when "0010100001001001", -- t[10313] = 1
      "000001" when "0010100001001010", -- t[10314] = 1
      "000001" when "0010100001001011", -- t[10315] = 1
      "000001" when "0010100001001100", -- t[10316] = 1
      "000001" when "0010100001001101", -- t[10317] = 1
      "000001" when "0010100001001110", -- t[10318] = 1
      "000001" when "0010100001001111", -- t[10319] = 1
      "000001" when "0010100001010000", -- t[10320] = 1
      "000001" when "0010100001010001", -- t[10321] = 1
      "000001" when "0010100001010010", -- t[10322] = 1
      "000001" when "0010100001010011", -- t[10323] = 1
      "000001" when "0010100001010100", -- t[10324] = 1
      "000001" when "0010100001010101", -- t[10325] = 1
      "000001" when "0010100001010110", -- t[10326] = 1
      "000001" when "0010100001010111", -- t[10327] = 1
      "000001" when "0010100001011000", -- t[10328] = 1
      "000001" when "0010100001011001", -- t[10329] = 1
      "000001" when "0010100001011010", -- t[10330] = 1
      "000001" when "0010100001011011", -- t[10331] = 1
      "000001" when "0010100001011100", -- t[10332] = 1
      "000001" when "0010100001011101", -- t[10333] = 1
      "000001" when "0010100001011110", -- t[10334] = 1
      "000001" when "0010100001011111", -- t[10335] = 1
      "000001" when "0010100001100000", -- t[10336] = 1
      "000001" when "0010100001100001", -- t[10337] = 1
      "000001" when "0010100001100010", -- t[10338] = 1
      "000001" when "0010100001100011", -- t[10339] = 1
      "000001" when "0010100001100100", -- t[10340] = 1
      "000001" when "0010100001100101", -- t[10341] = 1
      "000001" when "0010100001100110", -- t[10342] = 1
      "000001" when "0010100001100111", -- t[10343] = 1
      "000001" when "0010100001101000", -- t[10344] = 1
      "000001" when "0010100001101001", -- t[10345] = 1
      "000001" when "0010100001101010", -- t[10346] = 1
      "000001" when "0010100001101011", -- t[10347] = 1
      "000001" when "0010100001101100", -- t[10348] = 1
      "000001" when "0010100001101101", -- t[10349] = 1
      "000001" when "0010100001101110", -- t[10350] = 1
      "000001" when "0010100001101111", -- t[10351] = 1
      "000001" when "0010100001110000", -- t[10352] = 1
      "000001" when "0010100001110001", -- t[10353] = 1
      "000001" when "0010100001110010", -- t[10354] = 1
      "000001" when "0010100001110011", -- t[10355] = 1
      "000001" when "0010100001110100", -- t[10356] = 1
      "000001" when "0010100001110101", -- t[10357] = 1
      "000001" when "0010100001110110", -- t[10358] = 1
      "000001" when "0010100001110111", -- t[10359] = 1
      "000001" when "0010100001111000", -- t[10360] = 1
      "000001" when "0010100001111001", -- t[10361] = 1
      "000001" when "0010100001111010", -- t[10362] = 1
      "000001" when "0010100001111011", -- t[10363] = 1
      "000001" when "0010100001111100", -- t[10364] = 1
      "000001" when "0010100001111101", -- t[10365] = 1
      "000001" when "0010100001111110", -- t[10366] = 1
      "000001" when "0010100001111111", -- t[10367] = 1
      "000001" when "0010100010000000", -- t[10368] = 1
      "000001" when "0010100010000001", -- t[10369] = 1
      "000001" when "0010100010000010", -- t[10370] = 1
      "000001" when "0010100010000011", -- t[10371] = 1
      "000001" when "0010100010000100", -- t[10372] = 1
      "000001" when "0010100010000101", -- t[10373] = 1
      "000001" when "0010100010000110", -- t[10374] = 1
      "000001" when "0010100010000111", -- t[10375] = 1
      "000001" when "0010100010001000", -- t[10376] = 1
      "000001" when "0010100010001001", -- t[10377] = 1
      "000001" when "0010100010001010", -- t[10378] = 1
      "000001" when "0010100010001011", -- t[10379] = 1
      "000001" when "0010100010001100", -- t[10380] = 1
      "000001" when "0010100010001101", -- t[10381] = 1
      "000001" when "0010100010001110", -- t[10382] = 1
      "000001" when "0010100010001111", -- t[10383] = 1
      "000001" when "0010100010010000", -- t[10384] = 1
      "000001" when "0010100010010001", -- t[10385] = 1
      "000001" when "0010100010010010", -- t[10386] = 1
      "000001" when "0010100010010011", -- t[10387] = 1
      "000001" when "0010100010010100", -- t[10388] = 1
      "000001" when "0010100010010101", -- t[10389] = 1
      "000001" when "0010100010010110", -- t[10390] = 1
      "000001" when "0010100010010111", -- t[10391] = 1
      "000001" when "0010100010011000", -- t[10392] = 1
      "000001" when "0010100010011001", -- t[10393] = 1
      "000001" when "0010100010011010", -- t[10394] = 1
      "000001" when "0010100010011011", -- t[10395] = 1
      "000001" when "0010100010011100", -- t[10396] = 1
      "000001" when "0010100010011101", -- t[10397] = 1
      "000001" when "0010100010011110", -- t[10398] = 1
      "000001" when "0010100010011111", -- t[10399] = 1
      "000001" when "0010100010100000", -- t[10400] = 1
      "000001" when "0010100010100001", -- t[10401] = 1
      "000001" when "0010100010100010", -- t[10402] = 1
      "000001" when "0010100010100011", -- t[10403] = 1
      "000001" when "0010100010100100", -- t[10404] = 1
      "000001" when "0010100010100101", -- t[10405] = 1
      "000001" when "0010100010100110", -- t[10406] = 1
      "000001" when "0010100010100111", -- t[10407] = 1
      "000001" when "0010100010101000", -- t[10408] = 1
      "000001" when "0010100010101001", -- t[10409] = 1
      "000001" when "0010100010101010", -- t[10410] = 1
      "000001" when "0010100010101011", -- t[10411] = 1
      "000001" when "0010100010101100", -- t[10412] = 1
      "000001" when "0010100010101101", -- t[10413] = 1
      "000001" when "0010100010101110", -- t[10414] = 1
      "000001" when "0010100010101111", -- t[10415] = 1
      "000001" when "0010100010110000", -- t[10416] = 1
      "000001" when "0010100010110001", -- t[10417] = 1
      "000001" when "0010100010110010", -- t[10418] = 1
      "000001" when "0010100010110011", -- t[10419] = 1
      "000001" when "0010100010110100", -- t[10420] = 1
      "000001" when "0010100010110101", -- t[10421] = 1
      "000001" when "0010100010110110", -- t[10422] = 1
      "000001" when "0010100010110111", -- t[10423] = 1
      "000001" when "0010100010111000", -- t[10424] = 1
      "000001" when "0010100010111001", -- t[10425] = 1
      "000001" when "0010100010111010", -- t[10426] = 1
      "000001" when "0010100010111011", -- t[10427] = 1
      "000001" when "0010100010111100", -- t[10428] = 1
      "000001" when "0010100010111101", -- t[10429] = 1
      "000001" when "0010100010111110", -- t[10430] = 1
      "000001" when "0010100010111111", -- t[10431] = 1
      "000001" when "0010100011000000", -- t[10432] = 1
      "000001" when "0010100011000001", -- t[10433] = 1
      "000001" when "0010100011000010", -- t[10434] = 1
      "000001" when "0010100011000011", -- t[10435] = 1
      "000001" when "0010100011000100", -- t[10436] = 1
      "000001" when "0010100011000101", -- t[10437] = 1
      "000001" when "0010100011000110", -- t[10438] = 1
      "000001" when "0010100011000111", -- t[10439] = 1
      "000001" when "0010100011001000", -- t[10440] = 1
      "000001" when "0010100011001001", -- t[10441] = 1
      "000001" when "0010100011001010", -- t[10442] = 1
      "000001" when "0010100011001011", -- t[10443] = 1
      "000001" when "0010100011001100", -- t[10444] = 1
      "000001" when "0010100011001101", -- t[10445] = 1
      "000001" when "0010100011001110", -- t[10446] = 1
      "000001" when "0010100011001111", -- t[10447] = 1
      "000001" when "0010100011010000", -- t[10448] = 1
      "000001" when "0010100011010001", -- t[10449] = 1
      "000001" when "0010100011010010", -- t[10450] = 1
      "000001" when "0010100011010011", -- t[10451] = 1
      "000001" when "0010100011010100", -- t[10452] = 1
      "000001" when "0010100011010101", -- t[10453] = 1
      "000001" when "0010100011010110", -- t[10454] = 1
      "000001" when "0010100011010111", -- t[10455] = 1
      "000001" when "0010100011011000", -- t[10456] = 1
      "000001" when "0010100011011001", -- t[10457] = 1
      "000001" when "0010100011011010", -- t[10458] = 1
      "000001" when "0010100011011011", -- t[10459] = 1
      "000001" when "0010100011011100", -- t[10460] = 1
      "000001" when "0010100011011101", -- t[10461] = 1
      "000001" when "0010100011011110", -- t[10462] = 1
      "000001" when "0010100011011111", -- t[10463] = 1
      "000001" when "0010100011100000", -- t[10464] = 1
      "000001" when "0010100011100001", -- t[10465] = 1
      "000001" when "0010100011100010", -- t[10466] = 1
      "000001" when "0010100011100011", -- t[10467] = 1
      "000001" when "0010100011100100", -- t[10468] = 1
      "000001" when "0010100011100101", -- t[10469] = 1
      "000001" when "0010100011100110", -- t[10470] = 1
      "000001" when "0010100011100111", -- t[10471] = 1
      "000001" when "0010100011101000", -- t[10472] = 1
      "000001" when "0010100011101001", -- t[10473] = 1
      "000001" when "0010100011101010", -- t[10474] = 1
      "000001" when "0010100011101011", -- t[10475] = 1
      "000001" when "0010100011101100", -- t[10476] = 1
      "000001" when "0010100011101101", -- t[10477] = 1
      "000001" when "0010100011101110", -- t[10478] = 1
      "000001" when "0010100011101111", -- t[10479] = 1
      "000001" when "0010100011110000", -- t[10480] = 1
      "000001" when "0010100011110001", -- t[10481] = 1
      "000001" when "0010100011110010", -- t[10482] = 1
      "000001" when "0010100011110011", -- t[10483] = 1
      "000001" when "0010100011110100", -- t[10484] = 1
      "000001" when "0010100011110101", -- t[10485] = 1
      "000001" when "0010100011110110", -- t[10486] = 1
      "000001" when "0010100011110111", -- t[10487] = 1
      "000001" when "0010100011111000", -- t[10488] = 1
      "000001" when "0010100011111001", -- t[10489] = 1
      "000001" when "0010100011111010", -- t[10490] = 1
      "000001" when "0010100011111011", -- t[10491] = 1
      "000001" when "0010100011111100", -- t[10492] = 1
      "000001" when "0010100011111101", -- t[10493] = 1
      "000001" when "0010100011111110", -- t[10494] = 1
      "000001" when "0010100011111111", -- t[10495] = 1
      "000001" when "0010100100000000", -- t[10496] = 1
      "000001" when "0010100100000001", -- t[10497] = 1
      "000001" when "0010100100000010", -- t[10498] = 1
      "000001" when "0010100100000011", -- t[10499] = 1
      "000001" when "0010100100000100", -- t[10500] = 1
      "000001" when "0010100100000101", -- t[10501] = 1
      "000001" when "0010100100000110", -- t[10502] = 1
      "000001" when "0010100100000111", -- t[10503] = 1
      "000001" when "0010100100001000", -- t[10504] = 1
      "000001" when "0010100100001001", -- t[10505] = 1
      "000001" when "0010100100001010", -- t[10506] = 1
      "000001" when "0010100100001011", -- t[10507] = 1
      "000001" when "0010100100001100", -- t[10508] = 1
      "000001" when "0010100100001101", -- t[10509] = 1
      "000001" when "0010100100001110", -- t[10510] = 1
      "000001" when "0010100100001111", -- t[10511] = 1
      "000001" when "0010100100010000", -- t[10512] = 1
      "000001" when "0010100100010001", -- t[10513] = 1
      "000001" when "0010100100010010", -- t[10514] = 1
      "000001" when "0010100100010011", -- t[10515] = 1
      "000001" when "0010100100010100", -- t[10516] = 1
      "000001" when "0010100100010101", -- t[10517] = 1
      "000001" when "0010100100010110", -- t[10518] = 1
      "000001" when "0010100100010111", -- t[10519] = 1
      "000001" when "0010100100011000", -- t[10520] = 1
      "000001" when "0010100100011001", -- t[10521] = 1
      "000001" when "0010100100011010", -- t[10522] = 1
      "000001" when "0010100100011011", -- t[10523] = 1
      "000001" when "0010100100011100", -- t[10524] = 1
      "000001" when "0010100100011101", -- t[10525] = 1
      "000001" when "0010100100011110", -- t[10526] = 1
      "000001" when "0010100100011111", -- t[10527] = 1
      "000001" when "0010100100100000", -- t[10528] = 1
      "000001" when "0010100100100001", -- t[10529] = 1
      "000001" when "0010100100100010", -- t[10530] = 1
      "000001" when "0010100100100011", -- t[10531] = 1
      "000001" when "0010100100100100", -- t[10532] = 1
      "000001" when "0010100100100101", -- t[10533] = 1
      "000001" when "0010100100100110", -- t[10534] = 1
      "000001" when "0010100100100111", -- t[10535] = 1
      "000001" when "0010100100101000", -- t[10536] = 1
      "000001" when "0010100100101001", -- t[10537] = 1
      "000001" when "0010100100101010", -- t[10538] = 1
      "000001" when "0010100100101011", -- t[10539] = 1
      "000001" when "0010100100101100", -- t[10540] = 1
      "000001" when "0010100100101101", -- t[10541] = 1
      "000001" when "0010100100101110", -- t[10542] = 1
      "000001" when "0010100100101111", -- t[10543] = 1
      "000001" when "0010100100110000", -- t[10544] = 1
      "000001" when "0010100100110001", -- t[10545] = 1
      "000001" when "0010100100110010", -- t[10546] = 1
      "000001" when "0010100100110011", -- t[10547] = 1
      "000001" when "0010100100110100", -- t[10548] = 1
      "000001" when "0010100100110101", -- t[10549] = 1
      "000001" when "0010100100110110", -- t[10550] = 1
      "000001" when "0010100100110111", -- t[10551] = 1
      "000001" when "0010100100111000", -- t[10552] = 1
      "000001" when "0010100100111001", -- t[10553] = 1
      "000001" when "0010100100111010", -- t[10554] = 1
      "000001" when "0010100100111011", -- t[10555] = 1
      "000001" when "0010100100111100", -- t[10556] = 1
      "000001" when "0010100100111101", -- t[10557] = 1
      "000001" when "0010100100111110", -- t[10558] = 1
      "000001" when "0010100100111111", -- t[10559] = 1
      "000001" when "0010100101000000", -- t[10560] = 1
      "000001" when "0010100101000001", -- t[10561] = 1
      "000001" when "0010100101000010", -- t[10562] = 1
      "000001" when "0010100101000011", -- t[10563] = 1
      "000001" when "0010100101000100", -- t[10564] = 1
      "000001" when "0010100101000101", -- t[10565] = 1
      "000001" when "0010100101000110", -- t[10566] = 1
      "000001" when "0010100101000111", -- t[10567] = 1
      "000001" when "0010100101001000", -- t[10568] = 1
      "000001" when "0010100101001001", -- t[10569] = 1
      "000001" when "0010100101001010", -- t[10570] = 1
      "000001" when "0010100101001011", -- t[10571] = 1
      "000001" when "0010100101001100", -- t[10572] = 1
      "000001" when "0010100101001101", -- t[10573] = 1
      "000001" when "0010100101001110", -- t[10574] = 1
      "000001" when "0010100101001111", -- t[10575] = 1
      "000001" when "0010100101010000", -- t[10576] = 1
      "000001" when "0010100101010001", -- t[10577] = 1
      "000001" when "0010100101010010", -- t[10578] = 1
      "000001" when "0010100101010011", -- t[10579] = 1
      "000001" when "0010100101010100", -- t[10580] = 1
      "000001" when "0010100101010101", -- t[10581] = 1
      "000001" when "0010100101010110", -- t[10582] = 1
      "000001" when "0010100101010111", -- t[10583] = 1
      "000001" when "0010100101011000", -- t[10584] = 1
      "000001" when "0010100101011001", -- t[10585] = 1
      "000001" when "0010100101011010", -- t[10586] = 1
      "000001" when "0010100101011011", -- t[10587] = 1
      "000001" when "0010100101011100", -- t[10588] = 1
      "000001" when "0010100101011101", -- t[10589] = 1
      "000001" when "0010100101011110", -- t[10590] = 1
      "000001" when "0010100101011111", -- t[10591] = 1
      "000001" when "0010100101100000", -- t[10592] = 1
      "000001" when "0010100101100001", -- t[10593] = 1
      "000001" when "0010100101100010", -- t[10594] = 1
      "000001" when "0010100101100011", -- t[10595] = 1
      "000001" when "0010100101100100", -- t[10596] = 1
      "000001" when "0010100101100101", -- t[10597] = 1
      "000001" when "0010100101100110", -- t[10598] = 1
      "000001" when "0010100101100111", -- t[10599] = 1
      "000001" when "0010100101101000", -- t[10600] = 1
      "000001" when "0010100101101001", -- t[10601] = 1
      "000001" when "0010100101101010", -- t[10602] = 1
      "000001" when "0010100101101011", -- t[10603] = 1
      "000001" when "0010100101101100", -- t[10604] = 1
      "000001" when "0010100101101101", -- t[10605] = 1
      "000001" when "0010100101101110", -- t[10606] = 1
      "000001" when "0010100101101111", -- t[10607] = 1
      "000001" when "0010100101110000", -- t[10608] = 1
      "000001" when "0010100101110001", -- t[10609] = 1
      "000001" when "0010100101110010", -- t[10610] = 1
      "000001" when "0010100101110011", -- t[10611] = 1
      "000001" when "0010100101110100", -- t[10612] = 1
      "000001" when "0010100101110101", -- t[10613] = 1
      "000001" when "0010100101110110", -- t[10614] = 1
      "000001" when "0010100101110111", -- t[10615] = 1
      "000001" when "0010100101111000", -- t[10616] = 1
      "000001" when "0010100101111001", -- t[10617] = 1
      "000001" when "0010100101111010", -- t[10618] = 1
      "000001" when "0010100101111011", -- t[10619] = 1
      "000001" when "0010100101111100", -- t[10620] = 1
      "000001" when "0010100101111101", -- t[10621] = 1
      "000001" when "0010100101111110", -- t[10622] = 1
      "000001" when "0010100101111111", -- t[10623] = 1
      "000001" when "0010100110000000", -- t[10624] = 1
      "000001" when "0010100110000001", -- t[10625] = 1
      "000001" when "0010100110000010", -- t[10626] = 1
      "000001" when "0010100110000011", -- t[10627] = 1
      "000001" when "0010100110000100", -- t[10628] = 1
      "000001" when "0010100110000101", -- t[10629] = 1
      "000001" when "0010100110000110", -- t[10630] = 1
      "000001" when "0010100110000111", -- t[10631] = 1
      "000001" when "0010100110001000", -- t[10632] = 1
      "000001" when "0010100110001001", -- t[10633] = 1
      "000001" when "0010100110001010", -- t[10634] = 1
      "000001" when "0010100110001011", -- t[10635] = 1
      "000001" when "0010100110001100", -- t[10636] = 1
      "000001" when "0010100110001101", -- t[10637] = 1
      "000001" when "0010100110001110", -- t[10638] = 1
      "000001" when "0010100110001111", -- t[10639] = 1
      "000001" when "0010100110010000", -- t[10640] = 1
      "000001" when "0010100110010001", -- t[10641] = 1
      "000001" when "0010100110010010", -- t[10642] = 1
      "000001" when "0010100110010011", -- t[10643] = 1
      "000001" when "0010100110010100", -- t[10644] = 1
      "000001" when "0010100110010101", -- t[10645] = 1
      "000001" when "0010100110010110", -- t[10646] = 1
      "000001" when "0010100110010111", -- t[10647] = 1
      "000001" when "0010100110011000", -- t[10648] = 1
      "000001" when "0010100110011001", -- t[10649] = 1
      "000001" when "0010100110011010", -- t[10650] = 1
      "000001" when "0010100110011011", -- t[10651] = 1
      "000001" when "0010100110011100", -- t[10652] = 1
      "000001" when "0010100110011101", -- t[10653] = 1
      "000001" when "0010100110011110", -- t[10654] = 1
      "000001" when "0010100110011111", -- t[10655] = 1
      "000001" when "0010100110100000", -- t[10656] = 1
      "000001" when "0010100110100001", -- t[10657] = 1
      "000001" when "0010100110100010", -- t[10658] = 1
      "000001" when "0010100110100011", -- t[10659] = 1
      "000001" when "0010100110100100", -- t[10660] = 1
      "000001" when "0010100110100101", -- t[10661] = 1
      "000001" when "0010100110100110", -- t[10662] = 1
      "000001" when "0010100110100111", -- t[10663] = 1
      "000001" when "0010100110101000", -- t[10664] = 1
      "000001" when "0010100110101001", -- t[10665] = 1
      "000001" when "0010100110101010", -- t[10666] = 1
      "000001" when "0010100110101011", -- t[10667] = 1
      "000001" when "0010100110101100", -- t[10668] = 1
      "000001" when "0010100110101101", -- t[10669] = 1
      "000001" when "0010100110101110", -- t[10670] = 1
      "000001" when "0010100110101111", -- t[10671] = 1
      "000001" when "0010100110110000", -- t[10672] = 1
      "000001" when "0010100110110001", -- t[10673] = 1
      "000001" when "0010100110110010", -- t[10674] = 1
      "000001" when "0010100110110011", -- t[10675] = 1
      "000001" when "0010100110110100", -- t[10676] = 1
      "000001" when "0010100110110101", -- t[10677] = 1
      "000001" when "0010100110110110", -- t[10678] = 1
      "000001" when "0010100110110111", -- t[10679] = 1
      "000001" when "0010100110111000", -- t[10680] = 1
      "000001" when "0010100110111001", -- t[10681] = 1
      "000001" when "0010100110111010", -- t[10682] = 1
      "000001" when "0010100110111011", -- t[10683] = 1
      "000001" when "0010100110111100", -- t[10684] = 1
      "000001" when "0010100110111101", -- t[10685] = 1
      "000001" when "0010100110111110", -- t[10686] = 1
      "000001" when "0010100110111111", -- t[10687] = 1
      "000001" when "0010100111000000", -- t[10688] = 1
      "000001" when "0010100111000001", -- t[10689] = 1
      "000001" when "0010100111000010", -- t[10690] = 1
      "000001" when "0010100111000011", -- t[10691] = 1
      "000001" when "0010100111000100", -- t[10692] = 1
      "000001" when "0010100111000101", -- t[10693] = 1
      "000001" when "0010100111000110", -- t[10694] = 1
      "000001" when "0010100111000111", -- t[10695] = 1
      "000001" when "0010100111001000", -- t[10696] = 1
      "000001" when "0010100111001001", -- t[10697] = 1
      "000001" when "0010100111001010", -- t[10698] = 1
      "000001" when "0010100111001011", -- t[10699] = 1
      "000001" when "0010100111001100", -- t[10700] = 1
      "000001" when "0010100111001101", -- t[10701] = 1
      "000001" when "0010100111001110", -- t[10702] = 1
      "000001" when "0010100111001111", -- t[10703] = 1
      "000001" when "0010100111010000", -- t[10704] = 1
      "000001" when "0010100111010001", -- t[10705] = 1
      "000001" when "0010100111010010", -- t[10706] = 1
      "000001" when "0010100111010011", -- t[10707] = 1
      "000001" when "0010100111010100", -- t[10708] = 1
      "000001" when "0010100111010101", -- t[10709] = 1
      "000001" when "0010100111010110", -- t[10710] = 1
      "000001" when "0010100111010111", -- t[10711] = 1
      "000001" when "0010100111011000", -- t[10712] = 1
      "000001" when "0010100111011001", -- t[10713] = 1
      "000001" when "0010100111011010", -- t[10714] = 1
      "000001" when "0010100111011011", -- t[10715] = 1
      "000001" when "0010100111011100", -- t[10716] = 1
      "000001" when "0010100111011101", -- t[10717] = 1
      "000001" when "0010100111011110", -- t[10718] = 1
      "000001" when "0010100111011111", -- t[10719] = 1
      "000001" when "0010100111100000", -- t[10720] = 1
      "000001" when "0010100111100001", -- t[10721] = 1
      "000001" when "0010100111100010", -- t[10722] = 1
      "000001" when "0010100111100011", -- t[10723] = 1
      "000001" when "0010100111100100", -- t[10724] = 1
      "000001" when "0010100111100101", -- t[10725] = 1
      "000001" when "0010100111100110", -- t[10726] = 1
      "000001" when "0010100111100111", -- t[10727] = 1
      "000001" when "0010100111101000", -- t[10728] = 1
      "000001" when "0010100111101001", -- t[10729] = 1
      "000001" when "0010100111101010", -- t[10730] = 1
      "000001" when "0010100111101011", -- t[10731] = 1
      "000001" when "0010100111101100", -- t[10732] = 1
      "000001" when "0010100111101101", -- t[10733] = 1
      "000001" when "0010100111101110", -- t[10734] = 1
      "000001" when "0010100111101111", -- t[10735] = 1
      "000001" when "0010100111110000", -- t[10736] = 1
      "000001" when "0010100111110001", -- t[10737] = 1
      "000001" when "0010100111110010", -- t[10738] = 1
      "000001" when "0010100111110011", -- t[10739] = 1
      "000001" when "0010100111110100", -- t[10740] = 1
      "000001" when "0010100111110101", -- t[10741] = 1
      "000001" when "0010100111110110", -- t[10742] = 1
      "000001" when "0010100111110111", -- t[10743] = 1
      "000001" when "0010100111111000", -- t[10744] = 1
      "000001" when "0010100111111001", -- t[10745] = 1
      "000001" when "0010100111111010", -- t[10746] = 1
      "000001" when "0010100111111011", -- t[10747] = 1
      "000001" when "0010100111111100", -- t[10748] = 1
      "000001" when "0010100111111101", -- t[10749] = 1
      "000001" when "0010100111111110", -- t[10750] = 1
      "000001" when "0010100111111111", -- t[10751] = 1
      "000001" when "0010101000000000", -- t[10752] = 1
      "000001" when "0010101000000001", -- t[10753] = 1
      "000001" when "0010101000000010", -- t[10754] = 1
      "000001" when "0010101000000011", -- t[10755] = 1
      "000001" when "0010101000000100", -- t[10756] = 1
      "000001" when "0010101000000101", -- t[10757] = 1
      "000001" when "0010101000000110", -- t[10758] = 1
      "000001" when "0010101000000111", -- t[10759] = 1
      "000001" when "0010101000001000", -- t[10760] = 1
      "000001" when "0010101000001001", -- t[10761] = 1
      "000001" when "0010101000001010", -- t[10762] = 1
      "000001" when "0010101000001011", -- t[10763] = 1
      "000001" when "0010101000001100", -- t[10764] = 1
      "000001" when "0010101000001101", -- t[10765] = 1
      "000001" when "0010101000001110", -- t[10766] = 1
      "000001" when "0010101000001111", -- t[10767] = 1
      "000001" when "0010101000010000", -- t[10768] = 1
      "000001" when "0010101000010001", -- t[10769] = 1
      "000001" when "0010101000010010", -- t[10770] = 1
      "000001" when "0010101000010011", -- t[10771] = 1
      "000001" when "0010101000010100", -- t[10772] = 1
      "000001" when "0010101000010101", -- t[10773] = 1
      "000001" when "0010101000010110", -- t[10774] = 1
      "000001" when "0010101000010111", -- t[10775] = 1
      "000001" when "0010101000011000", -- t[10776] = 1
      "000001" when "0010101000011001", -- t[10777] = 1
      "000001" when "0010101000011010", -- t[10778] = 1
      "000001" when "0010101000011011", -- t[10779] = 1
      "000001" when "0010101000011100", -- t[10780] = 1
      "000001" when "0010101000011101", -- t[10781] = 1
      "000001" when "0010101000011110", -- t[10782] = 1
      "000001" when "0010101000011111", -- t[10783] = 1
      "000001" when "0010101000100000", -- t[10784] = 1
      "000001" when "0010101000100001", -- t[10785] = 1
      "000001" when "0010101000100010", -- t[10786] = 1
      "000001" when "0010101000100011", -- t[10787] = 1
      "000001" when "0010101000100100", -- t[10788] = 1
      "000001" when "0010101000100101", -- t[10789] = 1
      "000001" when "0010101000100110", -- t[10790] = 1
      "000001" when "0010101000100111", -- t[10791] = 1
      "000001" when "0010101000101000", -- t[10792] = 1
      "000001" when "0010101000101001", -- t[10793] = 1
      "000001" when "0010101000101010", -- t[10794] = 1
      "000001" when "0010101000101011", -- t[10795] = 1
      "000001" when "0010101000101100", -- t[10796] = 1
      "000001" when "0010101000101101", -- t[10797] = 1
      "000001" when "0010101000101110", -- t[10798] = 1
      "000001" when "0010101000101111", -- t[10799] = 1
      "000001" when "0010101000110000", -- t[10800] = 1
      "000001" when "0010101000110001", -- t[10801] = 1
      "000001" when "0010101000110010", -- t[10802] = 1
      "000001" when "0010101000110011", -- t[10803] = 1
      "000001" when "0010101000110100", -- t[10804] = 1
      "000001" when "0010101000110101", -- t[10805] = 1
      "000001" when "0010101000110110", -- t[10806] = 1
      "000001" when "0010101000110111", -- t[10807] = 1
      "000001" when "0010101000111000", -- t[10808] = 1
      "000001" when "0010101000111001", -- t[10809] = 1
      "000001" when "0010101000111010", -- t[10810] = 1
      "000001" when "0010101000111011", -- t[10811] = 1
      "000001" when "0010101000111100", -- t[10812] = 1
      "000001" when "0010101000111101", -- t[10813] = 1
      "000001" when "0010101000111110", -- t[10814] = 1
      "000001" when "0010101000111111", -- t[10815] = 1
      "000001" when "0010101001000000", -- t[10816] = 1
      "000001" when "0010101001000001", -- t[10817] = 1
      "000001" when "0010101001000010", -- t[10818] = 1
      "000001" when "0010101001000011", -- t[10819] = 1
      "000001" when "0010101001000100", -- t[10820] = 1
      "000001" when "0010101001000101", -- t[10821] = 1
      "000001" when "0010101001000110", -- t[10822] = 1
      "000001" when "0010101001000111", -- t[10823] = 1
      "000001" when "0010101001001000", -- t[10824] = 1
      "000001" when "0010101001001001", -- t[10825] = 1
      "000001" when "0010101001001010", -- t[10826] = 1
      "000001" when "0010101001001011", -- t[10827] = 1
      "000001" when "0010101001001100", -- t[10828] = 1
      "000001" when "0010101001001101", -- t[10829] = 1
      "000001" when "0010101001001110", -- t[10830] = 1
      "000001" when "0010101001001111", -- t[10831] = 1
      "000001" when "0010101001010000", -- t[10832] = 1
      "000001" when "0010101001010001", -- t[10833] = 1
      "000001" when "0010101001010010", -- t[10834] = 1
      "000001" when "0010101001010011", -- t[10835] = 1
      "000001" when "0010101001010100", -- t[10836] = 1
      "000001" when "0010101001010101", -- t[10837] = 1
      "000001" when "0010101001010110", -- t[10838] = 1
      "000001" when "0010101001010111", -- t[10839] = 1
      "000001" when "0010101001011000", -- t[10840] = 1
      "000001" when "0010101001011001", -- t[10841] = 1
      "000001" when "0010101001011010", -- t[10842] = 1
      "000001" when "0010101001011011", -- t[10843] = 1
      "000001" when "0010101001011100", -- t[10844] = 1
      "000001" when "0010101001011101", -- t[10845] = 1
      "000001" when "0010101001011110", -- t[10846] = 1
      "000001" when "0010101001011111", -- t[10847] = 1
      "000001" when "0010101001100000", -- t[10848] = 1
      "000001" when "0010101001100001", -- t[10849] = 1
      "000001" when "0010101001100010", -- t[10850] = 1
      "000001" when "0010101001100011", -- t[10851] = 1
      "000001" when "0010101001100100", -- t[10852] = 1
      "000001" when "0010101001100101", -- t[10853] = 1
      "000001" when "0010101001100110", -- t[10854] = 1
      "000001" when "0010101001100111", -- t[10855] = 1
      "000001" when "0010101001101000", -- t[10856] = 1
      "000001" when "0010101001101001", -- t[10857] = 1
      "000001" when "0010101001101010", -- t[10858] = 1
      "000001" when "0010101001101011", -- t[10859] = 1
      "000001" when "0010101001101100", -- t[10860] = 1
      "000001" when "0010101001101101", -- t[10861] = 1
      "000001" when "0010101001101110", -- t[10862] = 1
      "000001" when "0010101001101111", -- t[10863] = 1
      "000001" when "0010101001110000", -- t[10864] = 1
      "000001" when "0010101001110001", -- t[10865] = 1
      "000001" when "0010101001110010", -- t[10866] = 1
      "000001" when "0010101001110011", -- t[10867] = 1
      "000001" when "0010101001110100", -- t[10868] = 1
      "000001" when "0010101001110101", -- t[10869] = 1
      "000001" when "0010101001110110", -- t[10870] = 1
      "000001" when "0010101001110111", -- t[10871] = 1
      "000001" when "0010101001111000", -- t[10872] = 1
      "000001" when "0010101001111001", -- t[10873] = 1
      "000001" when "0010101001111010", -- t[10874] = 1
      "000001" when "0010101001111011", -- t[10875] = 1
      "000001" when "0010101001111100", -- t[10876] = 1
      "000001" when "0010101001111101", -- t[10877] = 1
      "000001" when "0010101001111110", -- t[10878] = 1
      "000001" when "0010101001111111", -- t[10879] = 1
      "000001" when "0010101010000000", -- t[10880] = 1
      "000001" when "0010101010000001", -- t[10881] = 1
      "000001" when "0010101010000010", -- t[10882] = 1
      "000001" when "0010101010000011", -- t[10883] = 1
      "000001" when "0010101010000100", -- t[10884] = 1
      "000001" when "0010101010000101", -- t[10885] = 1
      "000001" when "0010101010000110", -- t[10886] = 1
      "000001" when "0010101010000111", -- t[10887] = 1
      "000001" when "0010101010001000", -- t[10888] = 1
      "000001" when "0010101010001001", -- t[10889] = 1
      "000001" when "0010101010001010", -- t[10890] = 1
      "000001" when "0010101010001011", -- t[10891] = 1
      "000001" when "0010101010001100", -- t[10892] = 1
      "000001" when "0010101010001101", -- t[10893] = 1
      "000001" when "0010101010001110", -- t[10894] = 1
      "000001" when "0010101010001111", -- t[10895] = 1
      "000001" when "0010101010010000", -- t[10896] = 1
      "000001" when "0010101010010001", -- t[10897] = 1
      "000001" when "0010101010010010", -- t[10898] = 1
      "000001" when "0010101010010011", -- t[10899] = 1
      "000001" when "0010101010010100", -- t[10900] = 1
      "000001" when "0010101010010101", -- t[10901] = 1
      "000001" when "0010101010010110", -- t[10902] = 1
      "000001" when "0010101010010111", -- t[10903] = 1
      "000001" when "0010101010011000", -- t[10904] = 1
      "000001" when "0010101010011001", -- t[10905] = 1
      "000001" when "0010101010011010", -- t[10906] = 1
      "000001" when "0010101010011011", -- t[10907] = 1
      "000001" when "0010101010011100", -- t[10908] = 1
      "000001" when "0010101010011101", -- t[10909] = 1
      "000001" when "0010101010011110", -- t[10910] = 1
      "000001" when "0010101010011111", -- t[10911] = 1
      "000001" when "0010101010100000", -- t[10912] = 1
      "000001" when "0010101010100001", -- t[10913] = 1
      "000001" when "0010101010100010", -- t[10914] = 1
      "000001" when "0010101010100011", -- t[10915] = 1
      "000001" when "0010101010100100", -- t[10916] = 1
      "000001" when "0010101010100101", -- t[10917] = 1
      "000001" when "0010101010100110", -- t[10918] = 1
      "000001" when "0010101010100111", -- t[10919] = 1
      "000001" when "0010101010101000", -- t[10920] = 1
      "000001" when "0010101010101001", -- t[10921] = 1
      "000001" when "0010101010101010", -- t[10922] = 1
      "000001" when "0010101010101011", -- t[10923] = 1
      "000001" when "0010101010101100", -- t[10924] = 1
      "000001" when "0010101010101101", -- t[10925] = 1
      "000001" when "0010101010101110", -- t[10926] = 1
      "000001" when "0010101010101111", -- t[10927] = 1
      "000001" when "0010101010110000", -- t[10928] = 1
      "000001" when "0010101010110001", -- t[10929] = 1
      "000001" when "0010101010110010", -- t[10930] = 1
      "000001" when "0010101010110011", -- t[10931] = 1
      "000001" when "0010101010110100", -- t[10932] = 1
      "000001" when "0010101010110101", -- t[10933] = 1
      "000001" when "0010101010110110", -- t[10934] = 1
      "000001" when "0010101010110111", -- t[10935] = 1
      "000001" when "0010101010111000", -- t[10936] = 1
      "000001" when "0010101010111001", -- t[10937] = 1
      "000001" when "0010101010111010", -- t[10938] = 1
      "000001" when "0010101010111011", -- t[10939] = 1
      "000001" when "0010101010111100", -- t[10940] = 1
      "000001" when "0010101010111101", -- t[10941] = 1
      "000001" when "0010101010111110", -- t[10942] = 1
      "000001" when "0010101010111111", -- t[10943] = 1
      "000001" when "0010101011000000", -- t[10944] = 1
      "000001" when "0010101011000001", -- t[10945] = 1
      "000001" when "0010101011000010", -- t[10946] = 1
      "000001" when "0010101011000011", -- t[10947] = 1
      "000001" when "0010101011000100", -- t[10948] = 1
      "000001" when "0010101011000101", -- t[10949] = 1
      "000001" when "0010101011000110", -- t[10950] = 1
      "000001" when "0010101011000111", -- t[10951] = 1
      "000001" when "0010101011001000", -- t[10952] = 1
      "000001" when "0010101011001001", -- t[10953] = 1
      "000001" when "0010101011001010", -- t[10954] = 1
      "000001" when "0010101011001011", -- t[10955] = 1
      "000001" when "0010101011001100", -- t[10956] = 1
      "000001" when "0010101011001101", -- t[10957] = 1
      "000001" when "0010101011001110", -- t[10958] = 1
      "000001" when "0010101011001111", -- t[10959] = 1
      "000001" when "0010101011010000", -- t[10960] = 1
      "000001" when "0010101011010001", -- t[10961] = 1
      "000001" when "0010101011010010", -- t[10962] = 1
      "000001" when "0010101011010011", -- t[10963] = 1
      "000001" when "0010101011010100", -- t[10964] = 1
      "000001" when "0010101011010101", -- t[10965] = 1
      "000001" when "0010101011010110", -- t[10966] = 1
      "000001" when "0010101011010111", -- t[10967] = 1
      "000001" when "0010101011011000", -- t[10968] = 1
      "000001" when "0010101011011001", -- t[10969] = 1
      "000001" when "0010101011011010", -- t[10970] = 1
      "000001" when "0010101011011011", -- t[10971] = 1
      "000001" when "0010101011011100", -- t[10972] = 1
      "000001" when "0010101011011101", -- t[10973] = 1
      "000001" when "0010101011011110", -- t[10974] = 1
      "000001" when "0010101011011111", -- t[10975] = 1
      "000001" when "0010101011100000", -- t[10976] = 1
      "000001" when "0010101011100001", -- t[10977] = 1
      "000001" when "0010101011100010", -- t[10978] = 1
      "000001" when "0010101011100011", -- t[10979] = 1
      "000001" when "0010101011100100", -- t[10980] = 1
      "000001" when "0010101011100101", -- t[10981] = 1
      "000001" when "0010101011100110", -- t[10982] = 1
      "000001" when "0010101011100111", -- t[10983] = 1
      "000001" when "0010101011101000", -- t[10984] = 1
      "000001" when "0010101011101001", -- t[10985] = 1
      "000001" when "0010101011101010", -- t[10986] = 1
      "000001" when "0010101011101011", -- t[10987] = 1
      "000001" when "0010101011101100", -- t[10988] = 1
      "000001" when "0010101011101101", -- t[10989] = 1
      "000001" when "0010101011101110", -- t[10990] = 1
      "000001" when "0010101011101111", -- t[10991] = 1
      "000001" when "0010101011110000", -- t[10992] = 1
      "000001" when "0010101011110001", -- t[10993] = 1
      "000001" when "0010101011110010", -- t[10994] = 1
      "000001" when "0010101011110011", -- t[10995] = 1
      "000001" when "0010101011110100", -- t[10996] = 1
      "000001" when "0010101011110101", -- t[10997] = 1
      "000001" when "0010101011110110", -- t[10998] = 1
      "000001" when "0010101011110111", -- t[10999] = 1
      "000001" when "0010101011111000", -- t[11000] = 1
      "000001" when "0010101011111001", -- t[11001] = 1
      "000001" when "0010101011111010", -- t[11002] = 1
      "000001" when "0010101011111011", -- t[11003] = 1
      "000001" when "0010101011111100", -- t[11004] = 1
      "000001" when "0010101011111101", -- t[11005] = 1
      "000001" when "0010101011111110", -- t[11006] = 1
      "000001" when "0010101011111111", -- t[11007] = 1
      "000001" when "0010101100000000", -- t[11008] = 1
      "000001" when "0010101100000001", -- t[11009] = 1
      "000001" when "0010101100000010", -- t[11010] = 1
      "000001" when "0010101100000011", -- t[11011] = 1
      "000001" when "0010101100000100", -- t[11012] = 1
      "000001" when "0010101100000101", -- t[11013] = 1
      "000001" when "0010101100000110", -- t[11014] = 1
      "000001" when "0010101100000111", -- t[11015] = 1
      "000001" when "0010101100001000", -- t[11016] = 1
      "000001" when "0010101100001001", -- t[11017] = 1
      "000001" when "0010101100001010", -- t[11018] = 1
      "000001" when "0010101100001011", -- t[11019] = 1
      "000001" when "0010101100001100", -- t[11020] = 1
      "000001" when "0010101100001101", -- t[11021] = 1
      "000001" when "0010101100001110", -- t[11022] = 1
      "000001" when "0010101100001111", -- t[11023] = 1
      "000001" when "0010101100010000", -- t[11024] = 1
      "000001" when "0010101100010001", -- t[11025] = 1
      "000001" when "0010101100010010", -- t[11026] = 1
      "000001" when "0010101100010011", -- t[11027] = 1
      "000001" when "0010101100010100", -- t[11028] = 1
      "000001" when "0010101100010101", -- t[11029] = 1
      "000001" when "0010101100010110", -- t[11030] = 1
      "000001" when "0010101100010111", -- t[11031] = 1
      "000001" when "0010101100011000", -- t[11032] = 1
      "000001" when "0010101100011001", -- t[11033] = 1
      "000001" when "0010101100011010", -- t[11034] = 1
      "000001" when "0010101100011011", -- t[11035] = 1
      "000001" when "0010101100011100", -- t[11036] = 1
      "000001" when "0010101100011101", -- t[11037] = 1
      "000001" when "0010101100011110", -- t[11038] = 1
      "000001" when "0010101100011111", -- t[11039] = 1
      "000001" when "0010101100100000", -- t[11040] = 1
      "000001" when "0010101100100001", -- t[11041] = 1
      "000001" when "0010101100100010", -- t[11042] = 1
      "000001" when "0010101100100011", -- t[11043] = 1
      "000001" when "0010101100100100", -- t[11044] = 1
      "000001" when "0010101100100101", -- t[11045] = 1
      "000001" when "0010101100100110", -- t[11046] = 1
      "000001" when "0010101100100111", -- t[11047] = 1
      "000001" when "0010101100101000", -- t[11048] = 1
      "000001" when "0010101100101001", -- t[11049] = 1
      "000001" when "0010101100101010", -- t[11050] = 1
      "000001" when "0010101100101011", -- t[11051] = 1
      "000001" when "0010101100101100", -- t[11052] = 1
      "000001" when "0010101100101101", -- t[11053] = 1
      "000001" when "0010101100101110", -- t[11054] = 1
      "000001" when "0010101100101111", -- t[11055] = 1
      "000001" when "0010101100110000", -- t[11056] = 1
      "000001" when "0010101100110001", -- t[11057] = 1
      "000001" when "0010101100110010", -- t[11058] = 1
      "000001" when "0010101100110011", -- t[11059] = 1
      "000001" when "0010101100110100", -- t[11060] = 1
      "000001" when "0010101100110101", -- t[11061] = 1
      "000001" when "0010101100110110", -- t[11062] = 1
      "000001" when "0010101100110111", -- t[11063] = 1
      "000001" when "0010101100111000", -- t[11064] = 1
      "000001" when "0010101100111001", -- t[11065] = 1
      "000001" when "0010101100111010", -- t[11066] = 1
      "000001" when "0010101100111011", -- t[11067] = 1
      "000001" when "0010101100111100", -- t[11068] = 1
      "000001" when "0010101100111101", -- t[11069] = 1
      "000001" when "0010101100111110", -- t[11070] = 1
      "000001" when "0010101100111111", -- t[11071] = 1
      "000001" when "0010101101000000", -- t[11072] = 1
      "000001" when "0010101101000001", -- t[11073] = 1
      "000001" when "0010101101000010", -- t[11074] = 1
      "000001" when "0010101101000011", -- t[11075] = 1
      "000001" when "0010101101000100", -- t[11076] = 1
      "000001" when "0010101101000101", -- t[11077] = 1
      "000001" when "0010101101000110", -- t[11078] = 1
      "000001" when "0010101101000111", -- t[11079] = 1
      "000001" when "0010101101001000", -- t[11080] = 1
      "000001" when "0010101101001001", -- t[11081] = 1
      "000001" when "0010101101001010", -- t[11082] = 1
      "000001" when "0010101101001011", -- t[11083] = 1
      "000001" when "0010101101001100", -- t[11084] = 1
      "000001" when "0010101101001101", -- t[11085] = 1
      "000001" when "0010101101001110", -- t[11086] = 1
      "000001" when "0010101101001111", -- t[11087] = 1
      "000001" when "0010101101010000", -- t[11088] = 1
      "000001" when "0010101101010001", -- t[11089] = 1
      "000001" when "0010101101010010", -- t[11090] = 1
      "000001" when "0010101101010011", -- t[11091] = 1
      "000001" when "0010101101010100", -- t[11092] = 1
      "000001" when "0010101101010101", -- t[11093] = 1
      "000001" when "0010101101010110", -- t[11094] = 1
      "000001" when "0010101101010111", -- t[11095] = 1
      "000001" when "0010101101011000", -- t[11096] = 1
      "000001" when "0010101101011001", -- t[11097] = 1
      "000001" when "0010101101011010", -- t[11098] = 1
      "000001" when "0010101101011011", -- t[11099] = 1
      "000001" when "0010101101011100", -- t[11100] = 1
      "000001" when "0010101101011101", -- t[11101] = 1
      "000001" when "0010101101011110", -- t[11102] = 1
      "000001" when "0010101101011111", -- t[11103] = 1
      "000001" when "0010101101100000", -- t[11104] = 1
      "000001" when "0010101101100001", -- t[11105] = 1
      "000001" when "0010101101100010", -- t[11106] = 1
      "000001" when "0010101101100011", -- t[11107] = 1
      "000001" when "0010101101100100", -- t[11108] = 1
      "000001" when "0010101101100101", -- t[11109] = 1
      "000001" when "0010101101100110", -- t[11110] = 1
      "000001" when "0010101101100111", -- t[11111] = 1
      "000001" when "0010101101101000", -- t[11112] = 1
      "000001" when "0010101101101001", -- t[11113] = 1
      "000001" when "0010101101101010", -- t[11114] = 1
      "000001" when "0010101101101011", -- t[11115] = 1
      "000001" when "0010101101101100", -- t[11116] = 1
      "000001" when "0010101101101101", -- t[11117] = 1
      "000001" when "0010101101101110", -- t[11118] = 1
      "000001" when "0010101101101111", -- t[11119] = 1
      "000001" when "0010101101110000", -- t[11120] = 1
      "000001" when "0010101101110001", -- t[11121] = 1
      "000001" when "0010101101110010", -- t[11122] = 1
      "000001" when "0010101101110011", -- t[11123] = 1
      "000001" when "0010101101110100", -- t[11124] = 1
      "000001" when "0010101101110101", -- t[11125] = 1
      "000001" when "0010101101110110", -- t[11126] = 1
      "000001" when "0010101101110111", -- t[11127] = 1
      "000001" when "0010101101111000", -- t[11128] = 1
      "000001" when "0010101101111001", -- t[11129] = 1
      "000001" when "0010101101111010", -- t[11130] = 1
      "000001" when "0010101101111011", -- t[11131] = 1
      "000001" when "0010101101111100", -- t[11132] = 1
      "000001" when "0010101101111101", -- t[11133] = 1
      "000001" when "0010101101111110", -- t[11134] = 1
      "000001" when "0010101101111111", -- t[11135] = 1
      "000001" when "0010101110000000", -- t[11136] = 1
      "000001" when "0010101110000001", -- t[11137] = 1
      "000001" when "0010101110000010", -- t[11138] = 1
      "000001" when "0010101110000011", -- t[11139] = 1
      "000001" when "0010101110000100", -- t[11140] = 1
      "000001" when "0010101110000101", -- t[11141] = 1
      "000001" when "0010101110000110", -- t[11142] = 1
      "000001" when "0010101110000111", -- t[11143] = 1
      "000001" when "0010101110001000", -- t[11144] = 1
      "000001" when "0010101110001001", -- t[11145] = 1
      "000001" when "0010101110001010", -- t[11146] = 1
      "000001" when "0010101110001011", -- t[11147] = 1
      "000001" when "0010101110001100", -- t[11148] = 1
      "000001" when "0010101110001101", -- t[11149] = 1
      "000001" when "0010101110001110", -- t[11150] = 1
      "000001" when "0010101110001111", -- t[11151] = 1
      "000001" when "0010101110010000", -- t[11152] = 1
      "000001" when "0010101110010001", -- t[11153] = 1
      "000001" when "0010101110010010", -- t[11154] = 1
      "000001" when "0010101110010011", -- t[11155] = 1
      "000001" when "0010101110010100", -- t[11156] = 1
      "000001" when "0010101110010101", -- t[11157] = 1
      "000001" when "0010101110010110", -- t[11158] = 1
      "000001" when "0010101110010111", -- t[11159] = 1
      "000001" when "0010101110011000", -- t[11160] = 1
      "000001" when "0010101110011001", -- t[11161] = 1
      "000001" when "0010101110011010", -- t[11162] = 1
      "000001" when "0010101110011011", -- t[11163] = 1
      "000001" when "0010101110011100", -- t[11164] = 1
      "000001" when "0010101110011101", -- t[11165] = 1
      "000001" when "0010101110011110", -- t[11166] = 1
      "000001" when "0010101110011111", -- t[11167] = 1
      "000001" when "0010101110100000", -- t[11168] = 1
      "000001" when "0010101110100001", -- t[11169] = 1
      "000001" when "0010101110100010", -- t[11170] = 1
      "000001" when "0010101110100011", -- t[11171] = 1
      "000001" when "0010101110100100", -- t[11172] = 1
      "000001" when "0010101110100101", -- t[11173] = 1
      "000001" when "0010101110100110", -- t[11174] = 1
      "000001" when "0010101110100111", -- t[11175] = 1
      "000001" when "0010101110101000", -- t[11176] = 1
      "000001" when "0010101110101001", -- t[11177] = 1
      "000001" when "0010101110101010", -- t[11178] = 1
      "000001" when "0010101110101011", -- t[11179] = 1
      "000001" when "0010101110101100", -- t[11180] = 1
      "000001" when "0010101110101101", -- t[11181] = 1
      "000001" when "0010101110101110", -- t[11182] = 1
      "000001" when "0010101110101111", -- t[11183] = 1
      "000001" when "0010101110110000", -- t[11184] = 1
      "000001" when "0010101110110001", -- t[11185] = 1
      "000001" when "0010101110110010", -- t[11186] = 1
      "000001" when "0010101110110011", -- t[11187] = 1
      "000001" when "0010101110110100", -- t[11188] = 1
      "000001" when "0010101110110101", -- t[11189] = 1
      "000001" when "0010101110110110", -- t[11190] = 1
      "000001" when "0010101110110111", -- t[11191] = 1
      "000001" when "0010101110111000", -- t[11192] = 1
      "000001" when "0010101110111001", -- t[11193] = 1
      "000001" when "0010101110111010", -- t[11194] = 1
      "000001" when "0010101110111011", -- t[11195] = 1
      "000001" when "0010101110111100", -- t[11196] = 1
      "000001" when "0010101110111101", -- t[11197] = 1
      "000001" when "0010101110111110", -- t[11198] = 1
      "000001" when "0010101110111111", -- t[11199] = 1
      "000001" when "0010101111000000", -- t[11200] = 1
      "000001" when "0010101111000001", -- t[11201] = 1
      "000001" when "0010101111000010", -- t[11202] = 1
      "000001" when "0010101111000011", -- t[11203] = 1
      "000001" when "0010101111000100", -- t[11204] = 1
      "000001" when "0010101111000101", -- t[11205] = 1
      "000001" when "0010101111000110", -- t[11206] = 1
      "000001" when "0010101111000111", -- t[11207] = 1
      "000001" when "0010101111001000", -- t[11208] = 1
      "000001" when "0010101111001001", -- t[11209] = 1
      "000001" when "0010101111001010", -- t[11210] = 1
      "000001" when "0010101111001011", -- t[11211] = 1
      "000001" when "0010101111001100", -- t[11212] = 1
      "000001" when "0010101111001101", -- t[11213] = 1
      "000001" when "0010101111001110", -- t[11214] = 1
      "000001" when "0010101111001111", -- t[11215] = 1
      "000001" when "0010101111010000", -- t[11216] = 1
      "000001" when "0010101111010001", -- t[11217] = 1
      "000001" when "0010101111010010", -- t[11218] = 1
      "000001" when "0010101111010011", -- t[11219] = 1
      "000001" when "0010101111010100", -- t[11220] = 1
      "000001" when "0010101111010101", -- t[11221] = 1
      "000001" when "0010101111010110", -- t[11222] = 1
      "000001" when "0010101111010111", -- t[11223] = 1
      "000001" when "0010101111011000", -- t[11224] = 1
      "000001" when "0010101111011001", -- t[11225] = 1
      "000001" when "0010101111011010", -- t[11226] = 1
      "000001" when "0010101111011011", -- t[11227] = 1
      "000001" when "0010101111011100", -- t[11228] = 1
      "000001" when "0010101111011101", -- t[11229] = 1
      "000001" when "0010101111011110", -- t[11230] = 1
      "000001" when "0010101111011111", -- t[11231] = 1
      "000001" when "0010101111100000", -- t[11232] = 1
      "000001" when "0010101111100001", -- t[11233] = 1
      "000001" when "0010101111100010", -- t[11234] = 1
      "000001" when "0010101111100011", -- t[11235] = 1
      "000001" when "0010101111100100", -- t[11236] = 1
      "000001" when "0010101111100101", -- t[11237] = 1
      "000001" when "0010101111100110", -- t[11238] = 1
      "000001" when "0010101111100111", -- t[11239] = 1
      "000001" when "0010101111101000", -- t[11240] = 1
      "000001" when "0010101111101001", -- t[11241] = 1
      "000001" when "0010101111101010", -- t[11242] = 1
      "000001" when "0010101111101011", -- t[11243] = 1
      "000001" when "0010101111101100", -- t[11244] = 1
      "000001" when "0010101111101101", -- t[11245] = 1
      "000001" when "0010101111101110", -- t[11246] = 1
      "000001" when "0010101111101111", -- t[11247] = 1
      "000001" when "0010101111110000", -- t[11248] = 1
      "000001" when "0010101111110001", -- t[11249] = 1
      "000001" when "0010101111110010", -- t[11250] = 1
      "000001" when "0010101111110011", -- t[11251] = 1
      "000001" when "0010101111110100", -- t[11252] = 1
      "000001" when "0010101111110101", -- t[11253] = 1
      "000001" when "0010101111110110", -- t[11254] = 1
      "000001" when "0010101111110111", -- t[11255] = 1
      "000001" when "0010101111111000", -- t[11256] = 1
      "000001" when "0010101111111001", -- t[11257] = 1
      "000001" when "0010101111111010", -- t[11258] = 1
      "000001" when "0010101111111011", -- t[11259] = 1
      "000001" when "0010101111111100", -- t[11260] = 1
      "000001" when "0010101111111101", -- t[11261] = 1
      "000001" when "0010101111111110", -- t[11262] = 1
      "000001" when "0010101111111111", -- t[11263] = 1
      "000001" when "0010110000000000", -- t[11264] = 1
      "000001" when "0010110000000001", -- t[11265] = 1
      "000001" when "0010110000000010", -- t[11266] = 1
      "000001" when "0010110000000011", -- t[11267] = 1
      "000001" when "0010110000000100", -- t[11268] = 1
      "000001" when "0010110000000101", -- t[11269] = 1
      "000001" when "0010110000000110", -- t[11270] = 1
      "000001" when "0010110000000111", -- t[11271] = 1
      "000001" when "0010110000001000", -- t[11272] = 1
      "000001" when "0010110000001001", -- t[11273] = 1
      "000001" when "0010110000001010", -- t[11274] = 1
      "000001" when "0010110000001011", -- t[11275] = 1
      "000001" when "0010110000001100", -- t[11276] = 1
      "000001" when "0010110000001101", -- t[11277] = 1
      "000001" when "0010110000001110", -- t[11278] = 1
      "000001" when "0010110000001111", -- t[11279] = 1
      "000001" when "0010110000010000", -- t[11280] = 1
      "000001" when "0010110000010001", -- t[11281] = 1
      "000001" when "0010110000010010", -- t[11282] = 1
      "000001" when "0010110000010011", -- t[11283] = 1
      "000001" when "0010110000010100", -- t[11284] = 1
      "000001" when "0010110000010101", -- t[11285] = 1
      "000001" when "0010110000010110", -- t[11286] = 1
      "000001" when "0010110000010111", -- t[11287] = 1
      "000001" when "0010110000011000", -- t[11288] = 1
      "000001" when "0010110000011001", -- t[11289] = 1
      "000001" when "0010110000011010", -- t[11290] = 1
      "000001" when "0010110000011011", -- t[11291] = 1
      "000001" when "0010110000011100", -- t[11292] = 1
      "000001" when "0010110000011101", -- t[11293] = 1
      "000001" when "0010110000011110", -- t[11294] = 1
      "000001" when "0010110000011111", -- t[11295] = 1
      "000001" when "0010110000100000", -- t[11296] = 1
      "000001" when "0010110000100001", -- t[11297] = 1
      "000001" when "0010110000100010", -- t[11298] = 1
      "000001" when "0010110000100011", -- t[11299] = 1
      "000001" when "0010110000100100", -- t[11300] = 1
      "000001" when "0010110000100101", -- t[11301] = 1
      "000001" when "0010110000100110", -- t[11302] = 1
      "000001" when "0010110000100111", -- t[11303] = 1
      "000001" when "0010110000101000", -- t[11304] = 1
      "000001" when "0010110000101001", -- t[11305] = 1
      "000001" when "0010110000101010", -- t[11306] = 1
      "000001" when "0010110000101011", -- t[11307] = 1
      "000001" when "0010110000101100", -- t[11308] = 1
      "000001" when "0010110000101101", -- t[11309] = 1
      "000001" when "0010110000101110", -- t[11310] = 1
      "000001" when "0010110000101111", -- t[11311] = 1
      "000001" when "0010110000110000", -- t[11312] = 1
      "000001" when "0010110000110001", -- t[11313] = 1
      "000001" when "0010110000110010", -- t[11314] = 1
      "000001" when "0010110000110011", -- t[11315] = 1
      "000001" when "0010110000110100", -- t[11316] = 1
      "000001" when "0010110000110101", -- t[11317] = 1
      "000001" when "0010110000110110", -- t[11318] = 1
      "000001" when "0010110000110111", -- t[11319] = 1
      "000001" when "0010110000111000", -- t[11320] = 1
      "000001" when "0010110000111001", -- t[11321] = 1
      "000001" when "0010110000111010", -- t[11322] = 1
      "000001" when "0010110000111011", -- t[11323] = 1
      "000001" when "0010110000111100", -- t[11324] = 1
      "000001" when "0010110000111101", -- t[11325] = 1
      "000001" when "0010110000111110", -- t[11326] = 1
      "000001" when "0010110000111111", -- t[11327] = 1
      "000001" when "0010110001000000", -- t[11328] = 1
      "000001" when "0010110001000001", -- t[11329] = 1
      "000001" when "0010110001000010", -- t[11330] = 1
      "000001" when "0010110001000011", -- t[11331] = 1
      "000001" when "0010110001000100", -- t[11332] = 1
      "000001" when "0010110001000101", -- t[11333] = 1
      "000001" when "0010110001000110", -- t[11334] = 1
      "000001" when "0010110001000111", -- t[11335] = 1
      "000001" when "0010110001001000", -- t[11336] = 1
      "000001" when "0010110001001001", -- t[11337] = 1
      "000001" when "0010110001001010", -- t[11338] = 1
      "000001" when "0010110001001011", -- t[11339] = 1
      "000001" when "0010110001001100", -- t[11340] = 1
      "000001" when "0010110001001101", -- t[11341] = 1
      "000001" when "0010110001001110", -- t[11342] = 1
      "000001" when "0010110001001111", -- t[11343] = 1
      "000001" when "0010110001010000", -- t[11344] = 1
      "000001" when "0010110001010001", -- t[11345] = 1
      "000001" when "0010110001010010", -- t[11346] = 1
      "000001" when "0010110001010011", -- t[11347] = 1
      "000001" when "0010110001010100", -- t[11348] = 1
      "000001" when "0010110001010101", -- t[11349] = 1
      "000001" when "0010110001010110", -- t[11350] = 1
      "000001" when "0010110001010111", -- t[11351] = 1
      "000001" when "0010110001011000", -- t[11352] = 1
      "000001" when "0010110001011001", -- t[11353] = 1
      "000001" when "0010110001011010", -- t[11354] = 1
      "000001" when "0010110001011011", -- t[11355] = 1
      "000001" when "0010110001011100", -- t[11356] = 1
      "000001" when "0010110001011101", -- t[11357] = 1
      "000001" when "0010110001011110", -- t[11358] = 1
      "000001" when "0010110001011111", -- t[11359] = 1
      "000001" when "0010110001100000", -- t[11360] = 1
      "000001" when "0010110001100001", -- t[11361] = 1
      "000001" when "0010110001100010", -- t[11362] = 1
      "000001" when "0010110001100011", -- t[11363] = 1
      "000001" when "0010110001100100", -- t[11364] = 1
      "000001" when "0010110001100101", -- t[11365] = 1
      "000001" when "0010110001100110", -- t[11366] = 1
      "000001" when "0010110001100111", -- t[11367] = 1
      "000001" when "0010110001101000", -- t[11368] = 1
      "000001" when "0010110001101001", -- t[11369] = 1
      "000001" when "0010110001101010", -- t[11370] = 1
      "000001" when "0010110001101011", -- t[11371] = 1
      "000001" when "0010110001101100", -- t[11372] = 1
      "000001" when "0010110001101101", -- t[11373] = 1
      "000001" when "0010110001101110", -- t[11374] = 1
      "000001" when "0010110001101111", -- t[11375] = 1
      "000001" when "0010110001110000", -- t[11376] = 1
      "000001" when "0010110001110001", -- t[11377] = 1
      "000001" when "0010110001110010", -- t[11378] = 1
      "000001" when "0010110001110011", -- t[11379] = 1
      "000001" when "0010110001110100", -- t[11380] = 1
      "000001" when "0010110001110101", -- t[11381] = 1
      "000001" when "0010110001110110", -- t[11382] = 1
      "000001" when "0010110001110111", -- t[11383] = 1
      "000001" when "0010110001111000", -- t[11384] = 1
      "000001" when "0010110001111001", -- t[11385] = 1
      "000001" when "0010110001111010", -- t[11386] = 1
      "000001" when "0010110001111011", -- t[11387] = 1
      "000001" when "0010110001111100", -- t[11388] = 1
      "000001" when "0010110001111101", -- t[11389] = 1
      "000001" when "0010110001111110", -- t[11390] = 1
      "000001" when "0010110001111111", -- t[11391] = 1
      "000001" when "0010110010000000", -- t[11392] = 1
      "000001" when "0010110010000001", -- t[11393] = 1
      "000001" when "0010110010000010", -- t[11394] = 1
      "000001" when "0010110010000011", -- t[11395] = 1
      "000001" when "0010110010000100", -- t[11396] = 1
      "000001" when "0010110010000101", -- t[11397] = 1
      "000001" when "0010110010000110", -- t[11398] = 1
      "000001" when "0010110010000111", -- t[11399] = 1
      "000001" when "0010110010001000", -- t[11400] = 1
      "000001" when "0010110010001001", -- t[11401] = 1
      "000001" when "0010110010001010", -- t[11402] = 1
      "000001" when "0010110010001011", -- t[11403] = 1
      "000001" when "0010110010001100", -- t[11404] = 1
      "000001" when "0010110010001101", -- t[11405] = 1
      "000001" when "0010110010001110", -- t[11406] = 1
      "000001" when "0010110010001111", -- t[11407] = 1
      "000001" when "0010110010010000", -- t[11408] = 1
      "000001" when "0010110010010001", -- t[11409] = 1
      "000001" when "0010110010010010", -- t[11410] = 1
      "000001" when "0010110010010011", -- t[11411] = 1
      "000001" when "0010110010010100", -- t[11412] = 1
      "000001" when "0010110010010101", -- t[11413] = 1
      "000001" when "0010110010010110", -- t[11414] = 1
      "000001" when "0010110010010111", -- t[11415] = 1
      "000001" when "0010110010011000", -- t[11416] = 1
      "000001" when "0010110010011001", -- t[11417] = 1
      "000001" when "0010110010011010", -- t[11418] = 1
      "000001" when "0010110010011011", -- t[11419] = 1
      "000001" when "0010110010011100", -- t[11420] = 1
      "000001" when "0010110010011101", -- t[11421] = 1
      "000001" when "0010110010011110", -- t[11422] = 1
      "000001" when "0010110010011111", -- t[11423] = 1
      "000001" when "0010110010100000", -- t[11424] = 1
      "000001" when "0010110010100001", -- t[11425] = 1
      "000001" when "0010110010100010", -- t[11426] = 1
      "000001" when "0010110010100011", -- t[11427] = 1
      "000001" when "0010110010100100", -- t[11428] = 1
      "000001" when "0010110010100101", -- t[11429] = 1
      "000001" when "0010110010100110", -- t[11430] = 1
      "000001" when "0010110010100111", -- t[11431] = 1
      "000001" when "0010110010101000", -- t[11432] = 1
      "000001" when "0010110010101001", -- t[11433] = 1
      "000001" when "0010110010101010", -- t[11434] = 1
      "000001" when "0010110010101011", -- t[11435] = 1
      "000001" when "0010110010101100", -- t[11436] = 1
      "000001" when "0010110010101101", -- t[11437] = 1
      "000001" when "0010110010101110", -- t[11438] = 1
      "000001" when "0010110010101111", -- t[11439] = 1
      "000001" when "0010110010110000", -- t[11440] = 1
      "000001" when "0010110010110001", -- t[11441] = 1
      "000001" when "0010110010110010", -- t[11442] = 1
      "000001" when "0010110010110011", -- t[11443] = 1
      "000001" when "0010110010110100", -- t[11444] = 1
      "000001" when "0010110010110101", -- t[11445] = 1
      "000001" when "0010110010110110", -- t[11446] = 1
      "000001" when "0010110010110111", -- t[11447] = 1
      "000001" when "0010110010111000", -- t[11448] = 1
      "000001" when "0010110010111001", -- t[11449] = 1
      "000001" when "0010110010111010", -- t[11450] = 1
      "000001" when "0010110010111011", -- t[11451] = 1
      "000001" when "0010110010111100", -- t[11452] = 1
      "000001" when "0010110010111101", -- t[11453] = 1
      "000001" when "0010110010111110", -- t[11454] = 1
      "000001" when "0010110010111111", -- t[11455] = 1
      "000001" when "0010110011000000", -- t[11456] = 1
      "000001" when "0010110011000001", -- t[11457] = 1
      "000001" when "0010110011000010", -- t[11458] = 1
      "000001" when "0010110011000011", -- t[11459] = 1
      "000001" when "0010110011000100", -- t[11460] = 1
      "000001" when "0010110011000101", -- t[11461] = 1
      "000001" when "0010110011000110", -- t[11462] = 1
      "000001" when "0010110011000111", -- t[11463] = 1
      "000001" when "0010110011001000", -- t[11464] = 1
      "000001" when "0010110011001001", -- t[11465] = 1
      "000001" when "0010110011001010", -- t[11466] = 1
      "000001" when "0010110011001011", -- t[11467] = 1
      "000001" when "0010110011001100", -- t[11468] = 1
      "000001" when "0010110011001101", -- t[11469] = 1
      "000001" when "0010110011001110", -- t[11470] = 1
      "000001" when "0010110011001111", -- t[11471] = 1
      "000001" when "0010110011010000", -- t[11472] = 1
      "000001" when "0010110011010001", -- t[11473] = 1
      "000001" when "0010110011010010", -- t[11474] = 1
      "000001" when "0010110011010011", -- t[11475] = 1
      "000001" when "0010110011010100", -- t[11476] = 1
      "000001" when "0010110011010101", -- t[11477] = 1
      "000001" when "0010110011010110", -- t[11478] = 1
      "000001" when "0010110011010111", -- t[11479] = 1
      "000001" when "0010110011011000", -- t[11480] = 1
      "000001" when "0010110011011001", -- t[11481] = 1
      "000001" when "0010110011011010", -- t[11482] = 1
      "000001" when "0010110011011011", -- t[11483] = 1
      "000001" when "0010110011011100", -- t[11484] = 1
      "000001" when "0010110011011101", -- t[11485] = 1
      "000001" when "0010110011011110", -- t[11486] = 1
      "000001" when "0010110011011111", -- t[11487] = 1
      "000001" when "0010110011100000", -- t[11488] = 1
      "000001" when "0010110011100001", -- t[11489] = 1
      "000001" when "0010110011100010", -- t[11490] = 1
      "000001" when "0010110011100011", -- t[11491] = 1
      "000001" when "0010110011100100", -- t[11492] = 1
      "000001" when "0010110011100101", -- t[11493] = 1
      "000001" when "0010110011100110", -- t[11494] = 1
      "000001" when "0010110011100111", -- t[11495] = 1
      "000001" when "0010110011101000", -- t[11496] = 1
      "000001" when "0010110011101001", -- t[11497] = 1
      "000001" when "0010110011101010", -- t[11498] = 1
      "000001" when "0010110011101011", -- t[11499] = 1
      "000001" when "0010110011101100", -- t[11500] = 1
      "000001" when "0010110011101101", -- t[11501] = 1
      "000001" when "0010110011101110", -- t[11502] = 1
      "000001" when "0010110011101111", -- t[11503] = 1
      "000001" when "0010110011110000", -- t[11504] = 1
      "000001" when "0010110011110001", -- t[11505] = 1
      "000001" when "0010110011110010", -- t[11506] = 1
      "000001" when "0010110011110011", -- t[11507] = 1
      "000001" when "0010110011110100", -- t[11508] = 1
      "000001" when "0010110011110101", -- t[11509] = 1
      "000001" when "0010110011110110", -- t[11510] = 1
      "000001" when "0010110011110111", -- t[11511] = 1
      "000001" when "0010110011111000", -- t[11512] = 1
      "000001" when "0010110011111001", -- t[11513] = 1
      "000001" when "0010110011111010", -- t[11514] = 1
      "000001" when "0010110011111011", -- t[11515] = 1
      "000001" when "0010110011111100", -- t[11516] = 1
      "000001" when "0010110011111101", -- t[11517] = 1
      "000001" when "0010110011111110", -- t[11518] = 1
      "000001" when "0010110011111111", -- t[11519] = 1
      "000001" when "0010110100000000", -- t[11520] = 1
      "000001" when "0010110100000001", -- t[11521] = 1
      "000001" when "0010110100000010", -- t[11522] = 1
      "000001" when "0010110100000011", -- t[11523] = 1
      "000001" when "0010110100000100", -- t[11524] = 1
      "000001" when "0010110100000101", -- t[11525] = 1
      "000001" when "0010110100000110", -- t[11526] = 1
      "000001" when "0010110100000111", -- t[11527] = 1
      "000001" when "0010110100001000", -- t[11528] = 1
      "000001" when "0010110100001001", -- t[11529] = 1
      "000001" when "0010110100001010", -- t[11530] = 1
      "000001" when "0010110100001011", -- t[11531] = 1
      "000001" when "0010110100001100", -- t[11532] = 1
      "000001" when "0010110100001101", -- t[11533] = 1
      "000001" when "0010110100001110", -- t[11534] = 1
      "000001" when "0010110100001111", -- t[11535] = 1
      "000001" when "0010110100010000", -- t[11536] = 1
      "000001" when "0010110100010001", -- t[11537] = 1
      "000001" when "0010110100010010", -- t[11538] = 1
      "000001" when "0010110100010011", -- t[11539] = 1
      "000001" when "0010110100010100", -- t[11540] = 1
      "000001" when "0010110100010101", -- t[11541] = 1
      "000001" when "0010110100010110", -- t[11542] = 1
      "000001" when "0010110100010111", -- t[11543] = 1
      "000001" when "0010110100011000", -- t[11544] = 1
      "000001" when "0010110100011001", -- t[11545] = 1
      "000001" when "0010110100011010", -- t[11546] = 1
      "000001" when "0010110100011011", -- t[11547] = 1
      "000001" when "0010110100011100", -- t[11548] = 1
      "000001" when "0010110100011101", -- t[11549] = 1
      "000001" when "0010110100011110", -- t[11550] = 1
      "000001" when "0010110100011111", -- t[11551] = 1
      "000001" when "0010110100100000", -- t[11552] = 1
      "000001" when "0010110100100001", -- t[11553] = 1
      "000001" when "0010110100100010", -- t[11554] = 1
      "000001" when "0010110100100011", -- t[11555] = 1
      "000001" when "0010110100100100", -- t[11556] = 1
      "000001" when "0010110100100101", -- t[11557] = 1
      "000001" when "0010110100100110", -- t[11558] = 1
      "000001" when "0010110100100111", -- t[11559] = 1
      "000001" when "0010110100101000", -- t[11560] = 1
      "000001" when "0010110100101001", -- t[11561] = 1
      "000001" when "0010110100101010", -- t[11562] = 1
      "000001" when "0010110100101011", -- t[11563] = 1
      "000001" when "0010110100101100", -- t[11564] = 1
      "000001" when "0010110100101101", -- t[11565] = 1
      "000001" when "0010110100101110", -- t[11566] = 1
      "000001" when "0010110100101111", -- t[11567] = 1
      "000001" when "0010110100110000", -- t[11568] = 1
      "000001" when "0010110100110001", -- t[11569] = 1
      "000001" when "0010110100110010", -- t[11570] = 1
      "000001" when "0010110100110011", -- t[11571] = 1
      "000001" when "0010110100110100", -- t[11572] = 1
      "000001" when "0010110100110101", -- t[11573] = 1
      "000001" when "0010110100110110", -- t[11574] = 1
      "000001" when "0010110100110111", -- t[11575] = 1
      "000001" when "0010110100111000", -- t[11576] = 1
      "000001" when "0010110100111001", -- t[11577] = 1
      "000001" when "0010110100111010", -- t[11578] = 1
      "000001" when "0010110100111011", -- t[11579] = 1
      "000001" when "0010110100111100", -- t[11580] = 1
      "000001" when "0010110100111101", -- t[11581] = 1
      "000001" when "0010110100111110", -- t[11582] = 1
      "000001" when "0010110100111111", -- t[11583] = 1
      "000001" when "0010110101000000", -- t[11584] = 1
      "000001" when "0010110101000001", -- t[11585] = 1
      "000001" when "0010110101000010", -- t[11586] = 1
      "000001" when "0010110101000011", -- t[11587] = 1
      "000001" when "0010110101000100", -- t[11588] = 1
      "000001" when "0010110101000101", -- t[11589] = 1
      "000001" when "0010110101000110", -- t[11590] = 1
      "000001" when "0010110101000111", -- t[11591] = 1
      "000001" when "0010110101001000", -- t[11592] = 1
      "000001" when "0010110101001001", -- t[11593] = 1
      "000001" when "0010110101001010", -- t[11594] = 1
      "000001" when "0010110101001011", -- t[11595] = 1
      "000001" when "0010110101001100", -- t[11596] = 1
      "000001" when "0010110101001101", -- t[11597] = 1
      "000001" when "0010110101001110", -- t[11598] = 1
      "000001" when "0010110101001111", -- t[11599] = 1
      "000001" when "0010110101010000", -- t[11600] = 1
      "000001" when "0010110101010001", -- t[11601] = 1
      "000001" when "0010110101010010", -- t[11602] = 1
      "000001" when "0010110101010011", -- t[11603] = 1
      "000001" when "0010110101010100", -- t[11604] = 1
      "000001" when "0010110101010101", -- t[11605] = 1
      "000001" when "0010110101010110", -- t[11606] = 1
      "000001" when "0010110101010111", -- t[11607] = 1
      "000001" when "0010110101011000", -- t[11608] = 1
      "000001" when "0010110101011001", -- t[11609] = 1
      "000001" when "0010110101011010", -- t[11610] = 1
      "000001" when "0010110101011011", -- t[11611] = 1
      "000001" when "0010110101011100", -- t[11612] = 1
      "000001" when "0010110101011101", -- t[11613] = 1
      "000001" when "0010110101011110", -- t[11614] = 1
      "000001" when "0010110101011111", -- t[11615] = 1
      "000001" when "0010110101100000", -- t[11616] = 1
      "000001" when "0010110101100001", -- t[11617] = 1
      "000001" when "0010110101100010", -- t[11618] = 1
      "000001" when "0010110101100011", -- t[11619] = 1
      "000001" when "0010110101100100", -- t[11620] = 1
      "000001" when "0010110101100101", -- t[11621] = 1
      "000001" when "0010110101100110", -- t[11622] = 1
      "000001" when "0010110101100111", -- t[11623] = 1
      "000001" when "0010110101101000", -- t[11624] = 1
      "000001" when "0010110101101001", -- t[11625] = 1
      "000001" when "0010110101101010", -- t[11626] = 1
      "000001" when "0010110101101011", -- t[11627] = 1
      "000001" when "0010110101101100", -- t[11628] = 1
      "000001" when "0010110101101101", -- t[11629] = 1
      "000001" when "0010110101101110", -- t[11630] = 1
      "000001" when "0010110101101111", -- t[11631] = 1
      "000001" when "0010110101110000", -- t[11632] = 1
      "000001" when "0010110101110001", -- t[11633] = 1
      "000001" when "0010110101110010", -- t[11634] = 1
      "000001" when "0010110101110011", -- t[11635] = 1
      "000001" when "0010110101110100", -- t[11636] = 1
      "000001" when "0010110101110101", -- t[11637] = 1
      "000001" when "0010110101110110", -- t[11638] = 1
      "000001" when "0010110101110111", -- t[11639] = 1
      "000001" when "0010110101111000", -- t[11640] = 1
      "000001" when "0010110101111001", -- t[11641] = 1
      "000001" when "0010110101111010", -- t[11642] = 1
      "000001" when "0010110101111011", -- t[11643] = 1
      "000001" when "0010110101111100", -- t[11644] = 1
      "000001" when "0010110101111101", -- t[11645] = 1
      "000001" when "0010110101111110", -- t[11646] = 1
      "000001" when "0010110101111111", -- t[11647] = 1
      "000001" when "0010110110000000", -- t[11648] = 1
      "000001" when "0010110110000001", -- t[11649] = 1
      "000001" when "0010110110000010", -- t[11650] = 1
      "000001" when "0010110110000011", -- t[11651] = 1
      "000001" when "0010110110000100", -- t[11652] = 1
      "000001" when "0010110110000101", -- t[11653] = 1
      "000001" when "0010110110000110", -- t[11654] = 1
      "000001" when "0010110110000111", -- t[11655] = 1
      "000001" when "0010110110001000", -- t[11656] = 1
      "000001" when "0010110110001001", -- t[11657] = 1
      "000001" when "0010110110001010", -- t[11658] = 1
      "000001" when "0010110110001011", -- t[11659] = 1
      "000001" when "0010110110001100", -- t[11660] = 1
      "000001" when "0010110110001101", -- t[11661] = 1
      "000001" when "0010110110001110", -- t[11662] = 1
      "000001" when "0010110110001111", -- t[11663] = 1
      "000001" when "0010110110010000", -- t[11664] = 1
      "000001" when "0010110110010001", -- t[11665] = 1
      "000001" when "0010110110010010", -- t[11666] = 1
      "000001" when "0010110110010011", -- t[11667] = 1
      "000001" when "0010110110010100", -- t[11668] = 1
      "000001" when "0010110110010101", -- t[11669] = 1
      "000001" when "0010110110010110", -- t[11670] = 1
      "000001" when "0010110110010111", -- t[11671] = 1
      "000001" when "0010110110011000", -- t[11672] = 1
      "000001" when "0010110110011001", -- t[11673] = 1
      "000001" when "0010110110011010", -- t[11674] = 1
      "000001" when "0010110110011011", -- t[11675] = 1
      "000001" when "0010110110011100", -- t[11676] = 1
      "000001" when "0010110110011101", -- t[11677] = 1
      "000001" when "0010110110011110", -- t[11678] = 1
      "000001" when "0010110110011111", -- t[11679] = 1
      "000001" when "0010110110100000", -- t[11680] = 1
      "000001" when "0010110110100001", -- t[11681] = 1
      "000001" when "0010110110100010", -- t[11682] = 1
      "000001" when "0010110110100011", -- t[11683] = 1
      "000001" when "0010110110100100", -- t[11684] = 1
      "000001" when "0010110110100101", -- t[11685] = 1
      "000001" when "0010110110100110", -- t[11686] = 1
      "000001" when "0010110110100111", -- t[11687] = 1
      "000001" when "0010110110101000", -- t[11688] = 1
      "000001" when "0010110110101001", -- t[11689] = 1
      "000001" when "0010110110101010", -- t[11690] = 1
      "000001" when "0010110110101011", -- t[11691] = 1
      "000001" when "0010110110101100", -- t[11692] = 1
      "000001" when "0010110110101101", -- t[11693] = 1
      "000001" when "0010110110101110", -- t[11694] = 1
      "000001" when "0010110110101111", -- t[11695] = 1
      "000001" when "0010110110110000", -- t[11696] = 1
      "000001" when "0010110110110001", -- t[11697] = 1
      "000001" when "0010110110110010", -- t[11698] = 1
      "000001" when "0010110110110011", -- t[11699] = 1
      "000001" when "0010110110110100", -- t[11700] = 1
      "000001" when "0010110110110101", -- t[11701] = 1
      "000001" when "0010110110110110", -- t[11702] = 1
      "000001" when "0010110110110111", -- t[11703] = 1
      "000001" when "0010110110111000", -- t[11704] = 1
      "000001" when "0010110110111001", -- t[11705] = 1
      "000001" when "0010110110111010", -- t[11706] = 1
      "000001" when "0010110110111011", -- t[11707] = 1
      "000001" when "0010110110111100", -- t[11708] = 1
      "000001" when "0010110110111101", -- t[11709] = 1
      "000001" when "0010110110111110", -- t[11710] = 1
      "000001" when "0010110110111111", -- t[11711] = 1
      "000001" when "0010110111000000", -- t[11712] = 1
      "000001" when "0010110111000001", -- t[11713] = 1
      "000001" when "0010110111000010", -- t[11714] = 1
      "000001" when "0010110111000011", -- t[11715] = 1
      "000001" when "0010110111000100", -- t[11716] = 1
      "000001" when "0010110111000101", -- t[11717] = 1
      "000001" when "0010110111000110", -- t[11718] = 1
      "000001" when "0010110111000111", -- t[11719] = 1
      "000001" when "0010110111001000", -- t[11720] = 1
      "000001" when "0010110111001001", -- t[11721] = 1
      "000001" when "0010110111001010", -- t[11722] = 1
      "000001" when "0010110111001011", -- t[11723] = 1
      "000001" when "0010110111001100", -- t[11724] = 1
      "000001" when "0010110111001101", -- t[11725] = 1
      "000001" when "0010110111001110", -- t[11726] = 1
      "000001" when "0010110111001111", -- t[11727] = 1
      "000001" when "0010110111010000", -- t[11728] = 1
      "000001" when "0010110111010001", -- t[11729] = 1
      "000001" when "0010110111010010", -- t[11730] = 1
      "000001" when "0010110111010011", -- t[11731] = 1
      "000001" when "0010110111010100", -- t[11732] = 1
      "000001" when "0010110111010101", -- t[11733] = 1
      "000001" when "0010110111010110", -- t[11734] = 1
      "000001" when "0010110111010111", -- t[11735] = 1
      "000001" when "0010110111011000", -- t[11736] = 1
      "000001" when "0010110111011001", -- t[11737] = 1
      "000001" when "0010110111011010", -- t[11738] = 1
      "000001" when "0010110111011011", -- t[11739] = 1
      "000001" when "0010110111011100", -- t[11740] = 1
      "000001" when "0010110111011101", -- t[11741] = 1
      "000001" when "0010110111011110", -- t[11742] = 1
      "000001" when "0010110111011111", -- t[11743] = 1
      "000001" when "0010110111100000", -- t[11744] = 1
      "000001" when "0010110111100001", -- t[11745] = 1
      "000001" when "0010110111100010", -- t[11746] = 1
      "000001" when "0010110111100011", -- t[11747] = 1
      "000001" when "0010110111100100", -- t[11748] = 1
      "000001" when "0010110111100101", -- t[11749] = 1
      "000001" when "0010110111100110", -- t[11750] = 1
      "000001" when "0010110111100111", -- t[11751] = 1
      "000001" when "0010110111101000", -- t[11752] = 1
      "000001" when "0010110111101001", -- t[11753] = 1
      "000001" when "0010110111101010", -- t[11754] = 1
      "000001" when "0010110111101011", -- t[11755] = 1
      "000001" when "0010110111101100", -- t[11756] = 1
      "000001" when "0010110111101101", -- t[11757] = 1
      "000001" when "0010110111101110", -- t[11758] = 1
      "000001" when "0010110111101111", -- t[11759] = 1
      "000001" when "0010110111110000", -- t[11760] = 1
      "000001" when "0010110111110001", -- t[11761] = 1
      "000001" when "0010110111110010", -- t[11762] = 1
      "000001" when "0010110111110011", -- t[11763] = 1
      "000001" when "0010110111110100", -- t[11764] = 1
      "000001" when "0010110111110101", -- t[11765] = 1
      "000001" when "0010110111110110", -- t[11766] = 1
      "000001" when "0010110111110111", -- t[11767] = 1
      "000001" when "0010110111111000", -- t[11768] = 1
      "000001" when "0010110111111001", -- t[11769] = 1
      "000001" when "0010110111111010", -- t[11770] = 1
      "000001" when "0010110111111011", -- t[11771] = 1
      "000001" when "0010110111111100", -- t[11772] = 1
      "000001" when "0010110111111101", -- t[11773] = 1
      "000001" when "0010110111111110", -- t[11774] = 1
      "000001" when "0010110111111111", -- t[11775] = 1
      "000001" when "0010111000000000", -- t[11776] = 1
      "000001" when "0010111000000001", -- t[11777] = 1
      "000001" when "0010111000000010", -- t[11778] = 1
      "000001" when "0010111000000011", -- t[11779] = 1
      "000001" when "0010111000000100", -- t[11780] = 1
      "000001" when "0010111000000101", -- t[11781] = 1
      "000001" when "0010111000000110", -- t[11782] = 1
      "000001" when "0010111000000111", -- t[11783] = 1
      "000001" when "0010111000001000", -- t[11784] = 1
      "000001" when "0010111000001001", -- t[11785] = 1
      "000001" when "0010111000001010", -- t[11786] = 1
      "000001" when "0010111000001011", -- t[11787] = 1
      "000001" when "0010111000001100", -- t[11788] = 1
      "000001" when "0010111000001101", -- t[11789] = 1
      "000001" when "0010111000001110", -- t[11790] = 1
      "000001" when "0010111000001111", -- t[11791] = 1
      "000001" when "0010111000010000", -- t[11792] = 1
      "000001" when "0010111000010001", -- t[11793] = 1
      "000001" when "0010111000010010", -- t[11794] = 1
      "000001" when "0010111000010011", -- t[11795] = 1
      "000001" when "0010111000010100", -- t[11796] = 1
      "000001" when "0010111000010101", -- t[11797] = 1
      "000001" when "0010111000010110", -- t[11798] = 1
      "000001" when "0010111000010111", -- t[11799] = 1
      "000001" when "0010111000011000", -- t[11800] = 1
      "000001" when "0010111000011001", -- t[11801] = 1
      "000001" when "0010111000011010", -- t[11802] = 1
      "000001" when "0010111000011011", -- t[11803] = 1
      "000001" when "0010111000011100", -- t[11804] = 1
      "000001" when "0010111000011101", -- t[11805] = 1
      "000001" when "0010111000011110", -- t[11806] = 1
      "000001" when "0010111000011111", -- t[11807] = 1
      "000001" when "0010111000100000", -- t[11808] = 1
      "000001" when "0010111000100001", -- t[11809] = 1
      "000001" when "0010111000100010", -- t[11810] = 1
      "000001" when "0010111000100011", -- t[11811] = 1
      "000001" when "0010111000100100", -- t[11812] = 1
      "000001" when "0010111000100101", -- t[11813] = 1
      "000001" when "0010111000100110", -- t[11814] = 1
      "000001" when "0010111000100111", -- t[11815] = 1
      "000001" when "0010111000101000", -- t[11816] = 1
      "000001" when "0010111000101001", -- t[11817] = 1
      "000001" when "0010111000101010", -- t[11818] = 1
      "000001" when "0010111000101011", -- t[11819] = 1
      "000001" when "0010111000101100", -- t[11820] = 1
      "000001" when "0010111000101101", -- t[11821] = 1
      "000001" when "0010111000101110", -- t[11822] = 1
      "000001" when "0010111000101111", -- t[11823] = 1
      "000001" when "0010111000110000", -- t[11824] = 1
      "000001" when "0010111000110001", -- t[11825] = 1
      "000001" when "0010111000110010", -- t[11826] = 1
      "000001" when "0010111000110011", -- t[11827] = 1
      "000001" when "0010111000110100", -- t[11828] = 1
      "000001" when "0010111000110101", -- t[11829] = 1
      "000001" when "0010111000110110", -- t[11830] = 1
      "000001" when "0010111000110111", -- t[11831] = 1
      "000001" when "0010111000111000", -- t[11832] = 1
      "000001" when "0010111000111001", -- t[11833] = 1
      "000001" when "0010111000111010", -- t[11834] = 1
      "000001" when "0010111000111011", -- t[11835] = 1
      "000001" when "0010111000111100", -- t[11836] = 1
      "000001" when "0010111000111101", -- t[11837] = 1
      "000001" when "0010111000111110", -- t[11838] = 1
      "000001" when "0010111000111111", -- t[11839] = 1
      "000001" when "0010111001000000", -- t[11840] = 1
      "000001" when "0010111001000001", -- t[11841] = 1
      "000001" when "0010111001000010", -- t[11842] = 1
      "000001" when "0010111001000011", -- t[11843] = 1
      "000001" when "0010111001000100", -- t[11844] = 1
      "000001" when "0010111001000101", -- t[11845] = 1
      "000001" when "0010111001000110", -- t[11846] = 1
      "000001" when "0010111001000111", -- t[11847] = 1
      "000001" when "0010111001001000", -- t[11848] = 1
      "000001" when "0010111001001001", -- t[11849] = 1
      "000001" when "0010111001001010", -- t[11850] = 1
      "000001" when "0010111001001011", -- t[11851] = 1
      "000001" when "0010111001001100", -- t[11852] = 1
      "000001" when "0010111001001101", -- t[11853] = 1
      "000001" when "0010111001001110", -- t[11854] = 1
      "000001" when "0010111001001111", -- t[11855] = 1
      "000001" when "0010111001010000", -- t[11856] = 1
      "000001" when "0010111001010001", -- t[11857] = 1
      "000001" when "0010111001010010", -- t[11858] = 1
      "000001" when "0010111001010011", -- t[11859] = 1
      "000001" when "0010111001010100", -- t[11860] = 1
      "000001" when "0010111001010101", -- t[11861] = 1
      "000001" when "0010111001010110", -- t[11862] = 1
      "000001" when "0010111001010111", -- t[11863] = 1
      "000001" when "0010111001011000", -- t[11864] = 1
      "000001" when "0010111001011001", -- t[11865] = 1
      "000001" when "0010111001011010", -- t[11866] = 1
      "000001" when "0010111001011011", -- t[11867] = 1
      "000001" when "0010111001011100", -- t[11868] = 1
      "000001" when "0010111001011101", -- t[11869] = 1
      "000001" when "0010111001011110", -- t[11870] = 1
      "000001" when "0010111001011111", -- t[11871] = 1
      "000001" when "0010111001100000", -- t[11872] = 1
      "000001" when "0010111001100001", -- t[11873] = 1
      "000001" when "0010111001100010", -- t[11874] = 1
      "000001" when "0010111001100011", -- t[11875] = 1
      "000001" when "0010111001100100", -- t[11876] = 1
      "000001" when "0010111001100101", -- t[11877] = 1
      "000001" when "0010111001100110", -- t[11878] = 1
      "000001" when "0010111001100111", -- t[11879] = 1
      "000001" when "0010111001101000", -- t[11880] = 1
      "000001" when "0010111001101001", -- t[11881] = 1
      "000001" when "0010111001101010", -- t[11882] = 1
      "000001" when "0010111001101011", -- t[11883] = 1
      "000001" when "0010111001101100", -- t[11884] = 1
      "000001" when "0010111001101101", -- t[11885] = 1
      "000001" when "0010111001101110", -- t[11886] = 1
      "000001" when "0010111001101111", -- t[11887] = 1
      "000001" when "0010111001110000", -- t[11888] = 1
      "000001" when "0010111001110001", -- t[11889] = 1
      "000001" when "0010111001110010", -- t[11890] = 1
      "000001" when "0010111001110011", -- t[11891] = 1
      "000001" when "0010111001110100", -- t[11892] = 1
      "000001" when "0010111001110101", -- t[11893] = 1
      "000001" when "0010111001110110", -- t[11894] = 1
      "000001" when "0010111001110111", -- t[11895] = 1
      "000001" when "0010111001111000", -- t[11896] = 1
      "000001" when "0010111001111001", -- t[11897] = 1
      "000001" when "0010111001111010", -- t[11898] = 1
      "000001" when "0010111001111011", -- t[11899] = 1
      "000001" when "0010111001111100", -- t[11900] = 1
      "000001" when "0010111001111101", -- t[11901] = 1
      "000001" when "0010111001111110", -- t[11902] = 1
      "000001" when "0010111001111111", -- t[11903] = 1
      "000001" when "0010111010000000", -- t[11904] = 1
      "000001" when "0010111010000001", -- t[11905] = 1
      "000001" when "0010111010000010", -- t[11906] = 1
      "000001" when "0010111010000011", -- t[11907] = 1
      "000001" when "0010111010000100", -- t[11908] = 1
      "000001" when "0010111010000101", -- t[11909] = 1
      "000001" when "0010111010000110", -- t[11910] = 1
      "000001" when "0010111010000111", -- t[11911] = 1
      "000001" when "0010111010001000", -- t[11912] = 1
      "000001" when "0010111010001001", -- t[11913] = 1
      "000001" when "0010111010001010", -- t[11914] = 1
      "000001" when "0010111010001011", -- t[11915] = 1
      "000001" when "0010111010001100", -- t[11916] = 1
      "000001" when "0010111010001101", -- t[11917] = 1
      "000001" when "0010111010001110", -- t[11918] = 1
      "000001" when "0010111010001111", -- t[11919] = 1
      "000001" when "0010111010010000", -- t[11920] = 1
      "000001" when "0010111010010001", -- t[11921] = 1
      "000001" when "0010111010010010", -- t[11922] = 1
      "000001" when "0010111010010011", -- t[11923] = 1
      "000001" when "0010111010010100", -- t[11924] = 1
      "000001" when "0010111010010101", -- t[11925] = 1
      "000001" when "0010111010010110", -- t[11926] = 1
      "000001" when "0010111010010111", -- t[11927] = 1
      "000001" when "0010111010011000", -- t[11928] = 1
      "000001" when "0010111010011001", -- t[11929] = 1
      "000001" when "0010111010011010", -- t[11930] = 1
      "000001" when "0010111010011011", -- t[11931] = 1
      "000001" when "0010111010011100", -- t[11932] = 1
      "000001" when "0010111010011101", -- t[11933] = 1
      "000001" when "0010111010011110", -- t[11934] = 1
      "000001" when "0010111010011111", -- t[11935] = 1
      "000001" when "0010111010100000", -- t[11936] = 1
      "000001" when "0010111010100001", -- t[11937] = 1
      "000001" when "0010111010100010", -- t[11938] = 1
      "000001" when "0010111010100011", -- t[11939] = 1
      "000001" when "0010111010100100", -- t[11940] = 1
      "000001" when "0010111010100101", -- t[11941] = 1
      "000001" when "0010111010100110", -- t[11942] = 1
      "000001" when "0010111010100111", -- t[11943] = 1
      "000001" when "0010111010101000", -- t[11944] = 1
      "000001" when "0010111010101001", -- t[11945] = 1
      "000001" when "0010111010101010", -- t[11946] = 1
      "000001" when "0010111010101011", -- t[11947] = 1
      "000001" when "0010111010101100", -- t[11948] = 1
      "000001" when "0010111010101101", -- t[11949] = 1
      "000001" when "0010111010101110", -- t[11950] = 1
      "000001" when "0010111010101111", -- t[11951] = 1
      "000001" when "0010111010110000", -- t[11952] = 1
      "000001" when "0010111010110001", -- t[11953] = 1
      "000001" when "0010111010110010", -- t[11954] = 1
      "000001" when "0010111010110011", -- t[11955] = 1
      "000001" when "0010111010110100", -- t[11956] = 1
      "000001" when "0010111010110101", -- t[11957] = 1
      "000001" when "0010111010110110", -- t[11958] = 1
      "000001" when "0010111010110111", -- t[11959] = 1
      "000001" when "0010111010111000", -- t[11960] = 1
      "000001" when "0010111010111001", -- t[11961] = 1
      "000001" when "0010111010111010", -- t[11962] = 1
      "000001" when "0010111010111011", -- t[11963] = 1
      "000001" when "0010111010111100", -- t[11964] = 1
      "000001" when "0010111010111101", -- t[11965] = 1
      "000001" when "0010111010111110", -- t[11966] = 1
      "000001" when "0010111010111111", -- t[11967] = 1
      "000001" when "0010111011000000", -- t[11968] = 1
      "000001" when "0010111011000001", -- t[11969] = 1
      "000001" when "0010111011000010", -- t[11970] = 1
      "000001" when "0010111011000011", -- t[11971] = 1
      "000001" when "0010111011000100", -- t[11972] = 1
      "000001" when "0010111011000101", -- t[11973] = 1
      "000001" when "0010111011000110", -- t[11974] = 1
      "000001" when "0010111011000111", -- t[11975] = 1
      "000001" when "0010111011001000", -- t[11976] = 1
      "000001" when "0010111011001001", -- t[11977] = 1
      "000001" when "0010111011001010", -- t[11978] = 1
      "000001" when "0010111011001011", -- t[11979] = 1
      "000001" when "0010111011001100", -- t[11980] = 1
      "000001" when "0010111011001101", -- t[11981] = 1
      "000001" when "0010111011001110", -- t[11982] = 1
      "000001" when "0010111011001111", -- t[11983] = 1
      "000001" when "0010111011010000", -- t[11984] = 1
      "000001" when "0010111011010001", -- t[11985] = 1
      "000001" when "0010111011010010", -- t[11986] = 1
      "000001" when "0010111011010011", -- t[11987] = 1
      "000001" when "0010111011010100", -- t[11988] = 1
      "000001" when "0010111011010101", -- t[11989] = 1
      "000001" when "0010111011010110", -- t[11990] = 1
      "000001" when "0010111011010111", -- t[11991] = 1
      "000001" when "0010111011011000", -- t[11992] = 1
      "000001" when "0010111011011001", -- t[11993] = 1
      "000001" when "0010111011011010", -- t[11994] = 1
      "000001" when "0010111011011011", -- t[11995] = 1
      "000001" when "0010111011011100", -- t[11996] = 1
      "000001" when "0010111011011101", -- t[11997] = 1
      "000001" when "0010111011011110", -- t[11998] = 1
      "000001" when "0010111011011111", -- t[11999] = 1
      "000001" when "0010111011100000", -- t[12000] = 1
      "000001" when "0010111011100001", -- t[12001] = 1
      "000001" when "0010111011100010", -- t[12002] = 1
      "000001" when "0010111011100011", -- t[12003] = 1
      "000001" when "0010111011100100", -- t[12004] = 1
      "000001" when "0010111011100101", -- t[12005] = 1
      "000001" when "0010111011100110", -- t[12006] = 1
      "000001" when "0010111011100111", -- t[12007] = 1
      "000001" when "0010111011101000", -- t[12008] = 1
      "000001" when "0010111011101001", -- t[12009] = 1
      "000001" when "0010111011101010", -- t[12010] = 1
      "000001" when "0010111011101011", -- t[12011] = 1
      "000001" when "0010111011101100", -- t[12012] = 1
      "000001" when "0010111011101101", -- t[12013] = 1
      "000001" when "0010111011101110", -- t[12014] = 1
      "000001" when "0010111011101111", -- t[12015] = 1
      "000001" when "0010111011110000", -- t[12016] = 1
      "000001" when "0010111011110001", -- t[12017] = 1
      "000001" when "0010111011110010", -- t[12018] = 1
      "000001" when "0010111011110011", -- t[12019] = 1
      "000001" when "0010111011110100", -- t[12020] = 1
      "000001" when "0010111011110101", -- t[12021] = 1
      "000001" when "0010111011110110", -- t[12022] = 1
      "000001" when "0010111011110111", -- t[12023] = 1
      "000001" when "0010111011111000", -- t[12024] = 1
      "000001" when "0010111011111001", -- t[12025] = 1
      "000001" when "0010111011111010", -- t[12026] = 1
      "000001" when "0010111011111011", -- t[12027] = 1
      "000001" when "0010111011111100", -- t[12028] = 1
      "000001" when "0010111011111101", -- t[12029] = 1
      "000001" when "0010111011111110", -- t[12030] = 1
      "000001" when "0010111011111111", -- t[12031] = 1
      "000001" when "0010111100000000", -- t[12032] = 1
      "000001" when "0010111100000001", -- t[12033] = 1
      "000001" when "0010111100000010", -- t[12034] = 1
      "000001" when "0010111100000011", -- t[12035] = 1
      "000001" when "0010111100000100", -- t[12036] = 1
      "000001" when "0010111100000101", -- t[12037] = 1
      "000001" when "0010111100000110", -- t[12038] = 1
      "000001" when "0010111100000111", -- t[12039] = 1
      "000001" when "0010111100001000", -- t[12040] = 1
      "000001" when "0010111100001001", -- t[12041] = 1
      "000001" when "0010111100001010", -- t[12042] = 1
      "000001" when "0010111100001011", -- t[12043] = 1
      "000001" when "0010111100001100", -- t[12044] = 1
      "000001" when "0010111100001101", -- t[12045] = 1
      "000001" when "0010111100001110", -- t[12046] = 1
      "000001" when "0010111100001111", -- t[12047] = 1
      "000001" when "0010111100010000", -- t[12048] = 1
      "000001" when "0010111100010001", -- t[12049] = 1
      "000001" when "0010111100010010", -- t[12050] = 1
      "000001" when "0010111100010011", -- t[12051] = 1
      "000001" when "0010111100010100", -- t[12052] = 1
      "000001" when "0010111100010101", -- t[12053] = 1
      "000001" when "0010111100010110", -- t[12054] = 1
      "000001" when "0010111100010111", -- t[12055] = 1
      "000001" when "0010111100011000", -- t[12056] = 1
      "000001" when "0010111100011001", -- t[12057] = 1
      "000001" when "0010111100011010", -- t[12058] = 1
      "000001" when "0010111100011011", -- t[12059] = 1
      "000001" when "0010111100011100", -- t[12060] = 1
      "000001" when "0010111100011101", -- t[12061] = 1
      "000001" when "0010111100011110", -- t[12062] = 1
      "000001" when "0010111100011111", -- t[12063] = 1
      "000001" when "0010111100100000", -- t[12064] = 1
      "000001" when "0010111100100001", -- t[12065] = 1
      "000001" when "0010111100100010", -- t[12066] = 1
      "000001" when "0010111100100011", -- t[12067] = 1
      "000001" when "0010111100100100", -- t[12068] = 1
      "000001" when "0010111100100101", -- t[12069] = 1
      "000001" when "0010111100100110", -- t[12070] = 1
      "000001" when "0010111100100111", -- t[12071] = 1
      "000001" when "0010111100101000", -- t[12072] = 1
      "000001" when "0010111100101001", -- t[12073] = 1
      "000001" when "0010111100101010", -- t[12074] = 1
      "000001" when "0010111100101011", -- t[12075] = 1
      "000001" when "0010111100101100", -- t[12076] = 1
      "000001" when "0010111100101101", -- t[12077] = 1
      "000001" when "0010111100101110", -- t[12078] = 1
      "000001" when "0010111100101111", -- t[12079] = 1
      "000001" when "0010111100110000", -- t[12080] = 1
      "000001" when "0010111100110001", -- t[12081] = 1
      "000001" when "0010111100110010", -- t[12082] = 1
      "000001" when "0010111100110011", -- t[12083] = 1
      "000001" when "0010111100110100", -- t[12084] = 1
      "000001" when "0010111100110101", -- t[12085] = 1
      "000001" when "0010111100110110", -- t[12086] = 1
      "000001" when "0010111100110111", -- t[12087] = 1
      "000001" when "0010111100111000", -- t[12088] = 1
      "000001" when "0010111100111001", -- t[12089] = 1
      "000001" when "0010111100111010", -- t[12090] = 1
      "000001" when "0010111100111011", -- t[12091] = 1
      "000001" when "0010111100111100", -- t[12092] = 1
      "000001" when "0010111100111101", -- t[12093] = 1
      "000001" when "0010111100111110", -- t[12094] = 1
      "000001" when "0010111100111111", -- t[12095] = 1
      "000001" when "0010111101000000", -- t[12096] = 1
      "000001" when "0010111101000001", -- t[12097] = 1
      "000001" when "0010111101000010", -- t[12098] = 1
      "000001" when "0010111101000011", -- t[12099] = 1
      "000001" when "0010111101000100", -- t[12100] = 1
      "000001" when "0010111101000101", -- t[12101] = 1
      "000001" when "0010111101000110", -- t[12102] = 1
      "000001" when "0010111101000111", -- t[12103] = 1
      "000001" when "0010111101001000", -- t[12104] = 1
      "000001" when "0010111101001001", -- t[12105] = 1
      "000001" when "0010111101001010", -- t[12106] = 1
      "000001" when "0010111101001011", -- t[12107] = 1
      "000001" when "0010111101001100", -- t[12108] = 1
      "000001" when "0010111101001101", -- t[12109] = 1
      "000001" when "0010111101001110", -- t[12110] = 1
      "000001" when "0010111101001111", -- t[12111] = 1
      "000001" when "0010111101010000", -- t[12112] = 1
      "000001" when "0010111101010001", -- t[12113] = 1
      "000001" when "0010111101010010", -- t[12114] = 1
      "000001" when "0010111101010011", -- t[12115] = 1
      "000001" when "0010111101010100", -- t[12116] = 1
      "000001" when "0010111101010101", -- t[12117] = 1
      "000001" when "0010111101010110", -- t[12118] = 1
      "000001" when "0010111101010111", -- t[12119] = 1
      "000001" when "0010111101011000", -- t[12120] = 1
      "000001" when "0010111101011001", -- t[12121] = 1
      "000001" when "0010111101011010", -- t[12122] = 1
      "000001" when "0010111101011011", -- t[12123] = 1
      "000001" when "0010111101011100", -- t[12124] = 1
      "000001" when "0010111101011101", -- t[12125] = 1
      "000001" when "0010111101011110", -- t[12126] = 1
      "000001" when "0010111101011111", -- t[12127] = 1
      "000001" when "0010111101100000", -- t[12128] = 1
      "000001" when "0010111101100001", -- t[12129] = 1
      "000001" when "0010111101100010", -- t[12130] = 1
      "000001" when "0010111101100011", -- t[12131] = 1
      "000001" when "0010111101100100", -- t[12132] = 1
      "000001" when "0010111101100101", -- t[12133] = 1
      "000001" when "0010111101100110", -- t[12134] = 1
      "000001" when "0010111101100111", -- t[12135] = 1
      "000001" when "0010111101101000", -- t[12136] = 1
      "000001" when "0010111101101001", -- t[12137] = 1
      "000001" when "0010111101101010", -- t[12138] = 1
      "000001" when "0010111101101011", -- t[12139] = 1
      "000001" when "0010111101101100", -- t[12140] = 1
      "000001" when "0010111101101101", -- t[12141] = 1
      "000001" when "0010111101101110", -- t[12142] = 1
      "000001" when "0010111101101111", -- t[12143] = 1
      "000001" when "0010111101110000", -- t[12144] = 1
      "000001" when "0010111101110001", -- t[12145] = 1
      "000001" when "0010111101110010", -- t[12146] = 1
      "000001" when "0010111101110011", -- t[12147] = 1
      "000001" when "0010111101110100", -- t[12148] = 1
      "000001" when "0010111101110101", -- t[12149] = 1
      "000001" when "0010111101110110", -- t[12150] = 1
      "000001" when "0010111101110111", -- t[12151] = 1
      "000001" when "0010111101111000", -- t[12152] = 1
      "000001" when "0010111101111001", -- t[12153] = 1
      "000001" when "0010111101111010", -- t[12154] = 1
      "000001" when "0010111101111011", -- t[12155] = 1
      "000001" when "0010111101111100", -- t[12156] = 1
      "000001" when "0010111101111101", -- t[12157] = 1
      "000001" when "0010111101111110", -- t[12158] = 1
      "000001" when "0010111101111111", -- t[12159] = 1
      "000001" when "0010111110000000", -- t[12160] = 1
      "000001" when "0010111110000001", -- t[12161] = 1
      "000001" when "0010111110000010", -- t[12162] = 1
      "000001" when "0010111110000011", -- t[12163] = 1
      "000001" when "0010111110000100", -- t[12164] = 1
      "000001" when "0010111110000101", -- t[12165] = 1
      "000001" when "0010111110000110", -- t[12166] = 1
      "000001" when "0010111110000111", -- t[12167] = 1
      "000001" when "0010111110001000", -- t[12168] = 1
      "000001" when "0010111110001001", -- t[12169] = 1
      "000001" when "0010111110001010", -- t[12170] = 1
      "000001" when "0010111110001011", -- t[12171] = 1
      "000001" when "0010111110001100", -- t[12172] = 1
      "000001" when "0010111110001101", -- t[12173] = 1
      "000001" when "0010111110001110", -- t[12174] = 1
      "000001" when "0010111110001111", -- t[12175] = 1
      "000001" when "0010111110010000", -- t[12176] = 1
      "000001" when "0010111110010001", -- t[12177] = 1
      "000001" when "0010111110010010", -- t[12178] = 1
      "000001" when "0010111110010011", -- t[12179] = 1
      "000001" when "0010111110010100", -- t[12180] = 1
      "000001" when "0010111110010101", -- t[12181] = 1
      "000001" when "0010111110010110", -- t[12182] = 1
      "000001" when "0010111110010111", -- t[12183] = 1
      "000001" when "0010111110011000", -- t[12184] = 1
      "000001" when "0010111110011001", -- t[12185] = 1
      "000001" when "0010111110011010", -- t[12186] = 1
      "000001" when "0010111110011011", -- t[12187] = 1
      "000001" when "0010111110011100", -- t[12188] = 1
      "000001" when "0010111110011101", -- t[12189] = 1
      "000001" when "0010111110011110", -- t[12190] = 1
      "000001" when "0010111110011111", -- t[12191] = 1
      "000001" when "0010111110100000", -- t[12192] = 1
      "000001" when "0010111110100001", -- t[12193] = 1
      "000001" when "0010111110100010", -- t[12194] = 1
      "000001" when "0010111110100011", -- t[12195] = 1
      "000001" when "0010111110100100", -- t[12196] = 1
      "000001" when "0010111110100101", -- t[12197] = 1
      "000001" when "0010111110100110", -- t[12198] = 1
      "000001" when "0010111110100111", -- t[12199] = 1
      "000001" when "0010111110101000", -- t[12200] = 1
      "000001" when "0010111110101001", -- t[12201] = 1
      "000001" when "0010111110101010", -- t[12202] = 1
      "000001" when "0010111110101011", -- t[12203] = 1
      "000001" when "0010111110101100", -- t[12204] = 1
      "000001" when "0010111110101101", -- t[12205] = 1
      "000001" when "0010111110101110", -- t[12206] = 1
      "000001" when "0010111110101111", -- t[12207] = 1
      "000001" when "0010111110110000", -- t[12208] = 1
      "000001" when "0010111110110001", -- t[12209] = 1
      "000001" when "0010111110110010", -- t[12210] = 1
      "000001" when "0010111110110011", -- t[12211] = 1
      "000001" when "0010111110110100", -- t[12212] = 1
      "000001" when "0010111110110101", -- t[12213] = 1
      "000001" when "0010111110110110", -- t[12214] = 1
      "000001" when "0010111110110111", -- t[12215] = 1
      "000001" when "0010111110111000", -- t[12216] = 1
      "000001" when "0010111110111001", -- t[12217] = 1
      "000001" when "0010111110111010", -- t[12218] = 1
      "000001" when "0010111110111011", -- t[12219] = 1
      "000001" when "0010111110111100", -- t[12220] = 1
      "000001" when "0010111110111101", -- t[12221] = 1
      "000001" when "0010111110111110", -- t[12222] = 1
      "000001" when "0010111110111111", -- t[12223] = 1
      "000001" when "0010111111000000", -- t[12224] = 1
      "000001" when "0010111111000001", -- t[12225] = 1
      "000001" when "0010111111000010", -- t[12226] = 1
      "000001" when "0010111111000011", -- t[12227] = 1
      "000001" when "0010111111000100", -- t[12228] = 1
      "000001" when "0010111111000101", -- t[12229] = 1
      "000001" when "0010111111000110", -- t[12230] = 1
      "000001" when "0010111111000111", -- t[12231] = 1
      "000001" when "0010111111001000", -- t[12232] = 1
      "000001" when "0010111111001001", -- t[12233] = 1
      "000001" when "0010111111001010", -- t[12234] = 1
      "000001" when "0010111111001011", -- t[12235] = 1
      "000001" when "0010111111001100", -- t[12236] = 1
      "000001" when "0010111111001101", -- t[12237] = 1
      "000001" when "0010111111001110", -- t[12238] = 1
      "000001" when "0010111111001111", -- t[12239] = 1
      "000001" when "0010111111010000", -- t[12240] = 1
      "000001" when "0010111111010001", -- t[12241] = 1
      "000001" when "0010111111010010", -- t[12242] = 1
      "000001" when "0010111111010011", -- t[12243] = 1
      "000001" when "0010111111010100", -- t[12244] = 1
      "000001" when "0010111111010101", -- t[12245] = 1
      "000001" when "0010111111010110", -- t[12246] = 1
      "000001" when "0010111111010111", -- t[12247] = 1
      "000001" when "0010111111011000", -- t[12248] = 1
      "000001" when "0010111111011001", -- t[12249] = 1
      "000001" when "0010111111011010", -- t[12250] = 1
      "000001" when "0010111111011011", -- t[12251] = 1
      "000001" when "0010111111011100", -- t[12252] = 1
      "000001" when "0010111111011101", -- t[12253] = 1
      "000001" when "0010111111011110", -- t[12254] = 1
      "000001" when "0010111111011111", -- t[12255] = 1
      "000001" when "0010111111100000", -- t[12256] = 1
      "000001" when "0010111111100001", -- t[12257] = 1
      "000001" when "0010111111100010", -- t[12258] = 1
      "000001" when "0010111111100011", -- t[12259] = 1
      "000001" when "0010111111100100", -- t[12260] = 1
      "000001" when "0010111111100101", -- t[12261] = 1
      "000001" when "0010111111100110", -- t[12262] = 1
      "000001" when "0010111111100111", -- t[12263] = 1
      "000001" when "0010111111101000", -- t[12264] = 1
      "000001" when "0010111111101001", -- t[12265] = 1
      "000001" when "0010111111101010", -- t[12266] = 1
      "000001" when "0010111111101011", -- t[12267] = 1
      "000001" when "0010111111101100", -- t[12268] = 1
      "000001" when "0010111111101101", -- t[12269] = 1
      "000001" when "0010111111101110", -- t[12270] = 1
      "000001" when "0010111111101111", -- t[12271] = 1
      "000001" when "0010111111110000", -- t[12272] = 1
      "000001" when "0010111111110001", -- t[12273] = 1
      "000001" when "0010111111110010", -- t[12274] = 1
      "000001" when "0010111111110011", -- t[12275] = 1
      "000001" when "0010111111110100", -- t[12276] = 1
      "000001" when "0010111111110101", -- t[12277] = 1
      "000001" when "0010111111110110", -- t[12278] = 1
      "000001" when "0010111111110111", -- t[12279] = 1
      "000001" when "0010111111111000", -- t[12280] = 1
      "000001" when "0010111111111001", -- t[12281] = 1
      "000001" when "0010111111111010", -- t[12282] = 1
      "000001" when "0010111111111011", -- t[12283] = 1
      "000001" when "0010111111111100", -- t[12284] = 1
      "000001" when "0010111111111101", -- t[12285] = 1
      "000001" when "0010111111111110", -- t[12286] = 1
      "000001" when "0010111111111111", -- t[12287] = 1
      "000001" when "0011000000000000", -- t[12288] = 1
      "000001" when "0011000000000001", -- t[12289] = 1
      "000001" when "0011000000000010", -- t[12290] = 1
      "000001" when "0011000000000011", -- t[12291] = 1
      "000001" when "0011000000000100", -- t[12292] = 1
      "000001" when "0011000000000101", -- t[12293] = 1
      "000001" when "0011000000000110", -- t[12294] = 1
      "000001" when "0011000000000111", -- t[12295] = 1
      "000001" when "0011000000001000", -- t[12296] = 1
      "000001" when "0011000000001001", -- t[12297] = 1
      "000001" when "0011000000001010", -- t[12298] = 1
      "000001" when "0011000000001011", -- t[12299] = 1
      "000001" when "0011000000001100", -- t[12300] = 1
      "000001" when "0011000000001101", -- t[12301] = 1
      "000001" when "0011000000001110", -- t[12302] = 1
      "000001" when "0011000000001111", -- t[12303] = 1
      "000001" when "0011000000010000", -- t[12304] = 1
      "000001" when "0011000000010001", -- t[12305] = 1
      "000001" when "0011000000010010", -- t[12306] = 1
      "000001" when "0011000000010011", -- t[12307] = 1
      "000001" when "0011000000010100", -- t[12308] = 1
      "000001" when "0011000000010101", -- t[12309] = 1
      "000001" when "0011000000010110", -- t[12310] = 1
      "000001" when "0011000000010111", -- t[12311] = 1
      "000001" when "0011000000011000", -- t[12312] = 1
      "000001" when "0011000000011001", -- t[12313] = 1
      "000001" when "0011000000011010", -- t[12314] = 1
      "000001" when "0011000000011011", -- t[12315] = 1
      "000001" when "0011000000011100", -- t[12316] = 1
      "000001" when "0011000000011101", -- t[12317] = 1
      "000001" when "0011000000011110", -- t[12318] = 1
      "000001" when "0011000000011111", -- t[12319] = 1
      "000001" when "0011000000100000", -- t[12320] = 1
      "000001" when "0011000000100001", -- t[12321] = 1
      "000001" when "0011000000100010", -- t[12322] = 1
      "000001" when "0011000000100011", -- t[12323] = 1
      "000001" when "0011000000100100", -- t[12324] = 1
      "000001" when "0011000000100101", -- t[12325] = 1
      "000001" when "0011000000100110", -- t[12326] = 1
      "000001" when "0011000000100111", -- t[12327] = 1
      "000001" when "0011000000101000", -- t[12328] = 1
      "000001" when "0011000000101001", -- t[12329] = 1
      "000001" when "0011000000101010", -- t[12330] = 1
      "000001" when "0011000000101011", -- t[12331] = 1
      "000001" when "0011000000101100", -- t[12332] = 1
      "000001" when "0011000000101101", -- t[12333] = 1
      "000001" when "0011000000101110", -- t[12334] = 1
      "000001" when "0011000000101111", -- t[12335] = 1
      "000001" when "0011000000110000", -- t[12336] = 1
      "000001" when "0011000000110001", -- t[12337] = 1
      "000001" when "0011000000110010", -- t[12338] = 1
      "000001" when "0011000000110011", -- t[12339] = 1
      "000001" when "0011000000110100", -- t[12340] = 1
      "000001" when "0011000000110101", -- t[12341] = 1
      "000001" when "0011000000110110", -- t[12342] = 1
      "000001" when "0011000000110111", -- t[12343] = 1
      "000001" when "0011000000111000", -- t[12344] = 1
      "000001" when "0011000000111001", -- t[12345] = 1
      "000001" when "0011000000111010", -- t[12346] = 1
      "000001" when "0011000000111011", -- t[12347] = 1
      "000001" when "0011000000111100", -- t[12348] = 1
      "000001" when "0011000000111101", -- t[12349] = 1
      "000001" when "0011000000111110", -- t[12350] = 1
      "000001" when "0011000000111111", -- t[12351] = 1
      "000001" when "0011000001000000", -- t[12352] = 1
      "000001" when "0011000001000001", -- t[12353] = 1
      "000001" when "0011000001000010", -- t[12354] = 1
      "000001" when "0011000001000011", -- t[12355] = 1
      "000001" when "0011000001000100", -- t[12356] = 1
      "000001" when "0011000001000101", -- t[12357] = 1
      "000001" when "0011000001000110", -- t[12358] = 1
      "000001" when "0011000001000111", -- t[12359] = 1
      "000001" when "0011000001001000", -- t[12360] = 1
      "000001" when "0011000001001001", -- t[12361] = 1
      "000001" when "0011000001001010", -- t[12362] = 1
      "000001" when "0011000001001011", -- t[12363] = 1
      "000001" when "0011000001001100", -- t[12364] = 1
      "000001" when "0011000001001101", -- t[12365] = 1
      "000001" when "0011000001001110", -- t[12366] = 1
      "000001" when "0011000001001111", -- t[12367] = 1
      "000001" when "0011000001010000", -- t[12368] = 1
      "000001" when "0011000001010001", -- t[12369] = 1
      "000001" when "0011000001010010", -- t[12370] = 1
      "000001" when "0011000001010011", -- t[12371] = 1
      "000001" when "0011000001010100", -- t[12372] = 1
      "000001" when "0011000001010101", -- t[12373] = 1
      "000001" when "0011000001010110", -- t[12374] = 1
      "000001" when "0011000001010111", -- t[12375] = 1
      "000001" when "0011000001011000", -- t[12376] = 1
      "000001" when "0011000001011001", -- t[12377] = 1
      "000001" when "0011000001011010", -- t[12378] = 1
      "000001" when "0011000001011011", -- t[12379] = 1
      "000001" when "0011000001011100", -- t[12380] = 1
      "000001" when "0011000001011101", -- t[12381] = 1
      "000001" when "0011000001011110", -- t[12382] = 1
      "000001" when "0011000001011111", -- t[12383] = 1
      "000001" when "0011000001100000", -- t[12384] = 1
      "000001" when "0011000001100001", -- t[12385] = 1
      "000001" when "0011000001100010", -- t[12386] = 1
      "000001" when "0011000001100011", -- t[12387] = 1
      "000001" when "0011000001100100", -- t[12388] = 1
      "000001" when "0011000001100101", -- t[12389] = 1
      "000001" when "0011000001100110", -- t[12390] = 1
      "000001" when "0011000001100111", -- t[12391] = 1
      "000001" when "0011000001101000", -- t[12392] = 1
      "000001" when "0011000001101001", -- t[12393] = 1
      "000001" when "0011000001101010", -- t[12394] = 1
      "000001" when "0011000001101011", -- t[12395] = 1
      "000001" when "0011000001101100", -- t[12396] = 1
      "000001" when "0011000001101101", -- t[12397] = 1
      "000001" when "0011000001101110", -- t[12398] = 1
      "000001" when "0011000001101111", -- t[12399] = 1
      "000001" when "0011000001110000", -- t[12400] = 1
      "000001" when "0011000001110001", -- t[12401] = 1
      "000001" when "0011000001110010", -- t[12402] = 1
      "000001" when "0011000001110011", -- t[12403] = 1
      "000001" when "0011000001110100", -- t[12404] = 1
      "000001" when "0011000001110101", -- t[12405] = 1
      "000001" when "0011000001110110", -- t[12406] = 1
      "000001" when "0011000001110111", -- t[12407] = 1
      "000001" when "0011000001111000", -- t[12408] = 1
      "000001" when "0011000001111001", -- t[12409] = 1
      "000001" when "0011000001111010", -- t[12410] = 1
      "000001" when "0011000001111011", -- t[12411] = 1
      "000001" when "0011000001111100", -- t[12412] = 1
      "000001" when "0011000001111101", -- t[12413] = 1
      "000001" when "0011000001111110", -- t[12414] = 1
      "000001" when "0011000001111111", -- t[12415] = 1
      "000001" when "0011000010000000", -- t[12416] = 1
      "000001" when "0011000010000001", -- t[12417] = 1
      "000001" when "0011000010000010", -- t[12418] = 1
      "000001" when "0011000010000011", -- t[12419] = 1
      "000001" when "0011000010000100", -- t[12420] = 1
      "000001" when "0011000010000101", -- t[12421] = 1
      "000001" when "0011000010000110", -- t[12422] = 1
      "000001" when "0011000010000111", -- t[12423] = 1
      "000001" when "0011000010001000", -- t[12424] = 1
      "000001" when "0011000010001001", -- t[12425] = 1
      "000001" when "0011000010001010", -- t[12426] = 1
      "000001" when "0011000010001011", -- t[12427] = 1
      "000001" when "0011000010001100", -- t[12428] = 1
      "000001" when "0011000010001101", -- t[12429] = 1
      "000001" when "0011000010001110", -- t[12430] = 1
      "000001" when "0011000010001111", -- t[12431] = 1
      "000001" when "0011000010010000", -- t[12432] = 1
      "000001" when "0011000010010001", -- t[12433] = 1
      "000001" when "0011000010010010", -- t[12434] = 1
      "000001" when "0011000010010011", -- t[12435] = 1
      "000001" when "0011000010010100", -- t[12436] = 1
      "000001" when "0011000010010101", -- t[12437] = 1
      "000001" when "0011000010010110", -- t[12438] = 1
      "000001" when "0011000010010111", -- t[12439] = 1
      "000001" when "0011000010011000", -- t[12440] = 1
      "000001" when "0011000010011001", -- t[12441] = 1
      "000001" when "0011000010011010", -- t[12442] = 1
      "000001" when "0011000010011011", -- t[12443] = 1
      "000001" when "0011000010011100", -- t[12444] = 1
      "000001" when "0011000010011101", -- t[12445] = 1
      "000001" when "0011000010011110", -- t[12446] = 1
      "000001" when "0011000010011111", -- t[12447] = 1
      "000001" when "0011000010100000", -- t[12448] = 1
      "000001" when "0011000010100001", -- t[12449] = 1
      "000001" when "0011000010100010", -- t[12450] = 1
      "000001" when "0011000010100011", -- t[12451] = 1
      "000001" when "0011000010100100", -- t[12452] = 1
      "000001" when "0011000010100101", -- t[12453] = 1
      "000001" when "0011000010100110", -- t[12454] = 1
      "000001" when "0011000010100111", -- t[12455] = 1
      "000001" when "0011000010101000", -- t[12456] = 1
      "000001" when "0011000010101001", -- t[12457] = 1
      "000001" when "0011000010101010", -- t[12458] = 1
      "000001" when "0011000010101011", -- t[12459] = 1
      "000001" when "0011000010101100", -- t[12460] = 1
      "000001" when "0011000010101101", -- t[12461] = 1
      "000001" when "0011000010101110", -- t[12462] = 1
      "000001" when "0011000010101111", -- t[12463] = 1
      "000001" when "0011000010110000", -- t[12464] = 1
      "000001" when "0011000010110001", -- t[12465] = 1
      "000001" when "0011000010110010", -- t[12466] = 1
      "000001" when "0011000010110011", -- t[12467] = 1
      "000001" when "0011000010110100", -- t[12468] = 1
      "000001" when "0011000010110101", -- t[12469] = 1
      "000001" when "0011000010110110", -- t[12470] = 1
      "000001" when "0011000010110111", -- t[12471] = 1
      "000001" when "0011000010111000", -- t[12472] = 1
      "000001" when "0011000010111001", -- t[12473] = 1
      "000001" when "0011000010111010", -- t[12474] = 1
      "000001" when "0011000010111011", -- t[12475] = 1
      "000001" when "0011000010111100", -- t[12476] = 1
      "000001" when "0011000010111101", -- t[12477] = 1
      "000001" when "0011000010111110", -- t[12478] = 1
      "000001" when "0011000010111111", -- t[12479] = 1
      "000001" when "0011000011000000", -- t[12480] = 1
      "000001" when "0011000011000001", -- t[12481] = 1
      "000001" when "0011000011000010", -- t[12482] = 1
      "000001" when "0011000011000011", -- t[12483] = 1
      "000001" when "0011000011000100", -- t[12484] = 1
      "000001" when "0011000011000101", -- t[12485] = 1
      "000001" when "0011000011000110", -- t[12486] = 1
      "000001" when "0011000011000111", -- t[12487] = 1
      "000001" when "0011000011001000", -- t[12488] = 1
      "000001" when "0011000011001001", -- t[12489] = 1
      "000001" when "0011000011001010", -- t[12490] = 1
      "000001" when "0011000011001011", -- t[12491] = 1
      "000001" when "0011000011001100", -- t[12492] = 1
      "000001" when "0011000011001101", -- t[12493] = 1
      "000001" when "0011000011001110", -- t[12494] = 1
      "000001" when "0011000011001111", -- t[12495] = 1
      "000001" when "0011000011010000", -- t[12496] = 1
      "000001" when "0011000011010001", -- t[12497] = 1
      "000001" when "0011000011010010", -- t[12498] = 1
      "000001" when "0011000011010011", -- t[12499] = 1
      "000001" when "0011000011010100", -- t[12500] = 1
      "000001" when "0011000011010101", -- t[12501] = 1
      "000001" when "0011000011010110", -- t[12502] = 1
      "000001" when "0011000011010111", -- t[12503] = 1
      "000001" when "0011000011011000", -- t[12504] = 1
      "000001" when "0011000011011001", -- t[12505] = 1
      "000001" when "0011000011011010", -- t[12506] = 1
      "000001" when "0011000011011011", -- t[12507] = 1
      "000001" when "0011000011011100", -- t[12508] = 1
      "000001" when "0011000011011101", -- t[12509] = 1
      "000001" when "0011000011011110", -- t[12510] = 1
      "000001" when "0011000011011111", -- t[12511] = 1
      "000001" when "0011000011100000", -- t[12512] = 1
      "000001" when "0011000011100001", -- t[12513] = 1
      "000001" when "0011000011100010", -- t[12514] = 1
      "000001" when "0011000011100011", -- t[12515] = 1
      "000001" when "0011000011100100", -- t[12516] = 1
      "000001" when "0011000011100101", -- t[12517] = 1
      "000001" when "0011000011100110", -- t[12518] = 1
      "000001" when "0011000011100111", -- t[12519] = 1
      "000001" when "0011000011101000", -- t[12520] = 1
      "000001" when "0011000011101001", -- t[12521] = 1
      "000001" when "0011000011101010", -- t[12522] = 1
      "000001" when "0011000011101011", -- t[12523] = 1
      "000001" when "0011000011101100", -- t[12524] = 1
      "000001" when "0011000011101101", -- t[12525] = 1
      "000001" when "0011000011101110", -- t[12526] = 1
      "000001" when "0011000011101111", -- t[12527] = 1
      "000001" when "0011000011110000", -- t[12528] = 1
      "000001" when "0011000011110001", -- t[12529] = 1
      "000001" when "0011000011110010", -- t[12530] = 1
      "000001" when "0011000011110011", -- t[12531] = 1
      "000001" when "0011000011110100", -- t[12532] = 1
      "000001" when "0011000011110101", -- t[12533] = 1
      "000001" when "0011000011110110", -- t[12534] = 1
      "000001" when "0011000011110111", -- t[12535] = 1
      "000001" when "0011000011111000", -- t[12536] = 1
      "000001" when "0011000011111001", -- t[12537] = 1
      "000001" when "0011000011111010", -- t[12538] = 1
      "000001" when "0011000011111011", -- t[12539] = 1
      "000001" when "0011000011111100", -- t[12540] = 1
      "000001" when "0011000011111101", -- t[12541] = 1
      "000001" when "0011000011111110", -- t[12542] = 1
      "000001" when "0011000011111111", -- t[12543] = 1
      "000001" when "0011000100000000", -- t[12544] = 1
      "000001" when "0011000100000001", -- t[12545] = 1
      "000001" when "0011000100000010", -- t[12546] = 1
      "000001" when "0011000100000011", -- t[12547] = 1
      "000001" when "0011000100000100", -- t[12548] = 1
      "000001" when "0011000100000101", -- t[12549] = 1
      "000001" when "0011000100000110", -- t[12550] = 1
      "000001" when "0011000100000111", -- t[12551] = 1
      "000001" when "0011000100001000", -- t[12552] = 1
      "000001" when "0011000100001001", -- t[12553] = 1
      "000001" when "0011000100001010", -- t[12554] = 1
      "000001" when "0011000100001011", -- t[12555] = 1
      "000001" when "0011000100001100", -- t[12556] = 1
      "000001" when "0011000100001101", -- t[12557] = 1
      "000001" when "0011000100001110", -- t[12558] = 1
      "000001" when "0011000100001111", -- t[12559] = 1
      "000001" when "0011000100010000", -- t[12560] = 1
      "000001" when "0011000100010001", -- t[12561] = 1
      "000001" when "0011000100010010", -- t[12562] = 1
      "000001" when "0011000100010011", -- t[12563] = 1
      "000001" when "0011000100010100", -- t[12564] = 1
      "000001" when "0011000100010101", -- t[12565] = 1
      "000001" when "0011000100010110", -- t[12566] = 1
      "000001" when "0011000100010111", -- t[12567] = 1
      "000001" when "0011000100011000", -- t[12568] = 1
      "000001" when "0011000100011001", -- t[12569] = 1
      "000001" when "0011000100011010", -- t[12570] = 1
      "000001" when "0011000100011011", -- t[12571] = 1
      "000001" when "0011000100011100", -- t[12572] = 1
      "000001" when "0011000100011101", -- t[12573] = 1
      "000001" when "0011000100011110", -- t[12574] = 1
      "000001" when "0011000100011111", -- t[12575] = 1
      "000001" when "0011000100100000", -- t[12576] = 1
      "000001" when "0011000100100001", -- t[12577] = 1
      "000001" when "0011000100100010", -- t[12578] = 1
      "000001" when "0011000100100011", -- t[12579] = 1
      "000001" when "0011000100100100", -- t[12580] = 1
      "000001" when "0011000100100101", -- t[12581] = 1
      "000001" when "0011000100100110", -- t[12582] = 1
      "000001" when "0011000100100111", -- t[12583] = 1
      "000001" when "0011000100101000", -- t[12584] = 1
      "000001" when "0011000100101001", -- t[12585] = 1
      "000001" when "0011000100101010", -- t[12586] = 1
      "000001" when "0011000100101011", -- t[12587] = 1
      "000001" when "0011000100101100", -- t[12588] = 1
      "000001" when "0011000100101101", -- t[12589] = 1
      "000001" when "0011000100101110", -- t[12590] = 1
      "000001" when "0011000100101111", -- t[12591] = 1
      "000001" when "0011000100110000", -- t[12592] = 1
      "000001" when "0011000100110001", -- t[12593] = 1
      "000001" when "0011000100110010", -- t[12594] = 1
      "000001" when "0011000100110011", -- t[12595] = 1
      "000001" when "0011000100110100", -- t[12596] = 1
      "000001" when "0011000100110101", -- t[12597] = 1
      "000001" when "0011000100110110", -- t[12598] = 1
      "000001" when "0011000100110111", -- t[12599] = 1
      "000001" when "0011000100111000", -- t[12600] = 1
      "000001" when "0011000100111001", -- t[12601] = 1
      "000001" when "0011000100111010", -- t[12602] = 1
      "000001" when "0011000100111011", -- t[12603] = 1
      "000001" when "0011000100111100", -- t[12604] = 1
      "000001" when "0011000100111101", -- t[12605] = 1
      "000001" when "0011000100111110", -- t[12606] = 1
      "000001" when "0011000100111111", -- t[12607] = 1
      "000001" when "0011000101000000", -- t[12608] = 1
      "000001" when "0011000101000001", -- t[12609] = 1
      "000001" when "0011000101000010", -- t[12610] = 1
      "000001" when "0011000101000011", -- t[12611] = 1
      "000001" when "0011000101000100", -- t[12612] = 1
      "000001" when "0011000101000101", -- t[12613] = 1
      "000001" when "0011000101000110", -- t[12614] = 1
      "000001" when "0011000101000111", -- t[12615] = 1
      "000001" when "0011000101001000", -- t[12616] = 1
      "000001" when "0011000101001001", -- t[12617] = 1
      "000001" when "0011000101001010", -- t[12618] = 1
      "000001" when "0011000101001011", -- t[12619] = 1
      "000001" when "0011000101001100", -- t[12620] = 1
      "000001" when "0011000101001101", -- t[12621] = 1
      "000001" when "0011000101001110", -- t[12622] = 1
      "000001" when "0011000101001111", -- t[12623] = 1
      "000001" when "0011000101010000", -- t[12624] = 1
      "000001" when "0011000101010001", -- t[12625] = 1
      "000001" when "0011000101010010", -- t[12626] = 1
      "000001" when "0011000101010011", -- t[12627] = 1
      "000001" when "0011000101010100", -- t[12628] = 1
      "000001" when "0011000101010101", -- t[12629] = 1
      "000001" when "0011000101010110", -- t[12630] = 1
      "000001" when "0011000101010111", -- t[12631] = 1
      "000001" when "0011000101011000", -- t[12632] = 1
      "000001" when "0011000101011001", -- t[12633] = 1
      "000001" when "0011000101011010", -- t[12634] = 1
      "000001" when "0011000101011011", -- t[12635] = 1
      "000001" when "0011000101011100", -- t[12636] = 1
      "000001" when "0011000101011101", -- t[12637] = 1
      "000001" when "0011000101011110", -- t[12638] = 1
      "000001" when "0011000101011111", -- t[12639] = 1
      "000001" when "0011000101100000", -- t[12640] = 1
      "000001" when "0011000101100001", -- t[12641] = 1
      "000001" when "0011000101100010", -- t[12642] = 1
      "000001" when "0011000101100011", -- t[12643] = 1
      "000001" when "0011000101100100", -- t[12644] = 1
      "000001" when "0011000101100101", -- t[12645] = 1
      "000001" when "0011000101100110", -- t[12646] = 1
      "000001" when "0011000101100111", -- t[12647] = 1
      "000001" when "0011000101101000", -- t[12648] = 1
      "000001" when "0011000101101001", -- t[12649] = 1
      "000001" when "0011000101101010", -- t[12650] = 1
      "000001" when "0011000101101011", -- t[12651] = 1
      "000001" when "0011000101101100", -- t[12652] = 1
      "000001" when "0011000101101101", -- t[12653] = 1
      "000001" when "0011000101101110", -- t[12654] = 1
      "000001" when "0011000101101111", -- t[12655] = 1
      "000001" when "0011000101110000", -- t[12656] = 1
      "000001" when "0011000101110001", -- t[12657] = 1
      "000001" when "0011000101110010", -- t[12658] = 1
      "000001" when "0011000101110011", -- t[12659] = 1
      "000001" when "0011000101110100", -- t[12660] = 1
      "000001" when "0011000101110101", -- t[12661] = 1
      "000001" when "0011000101110110", -- t[12662] = 1
      "000001" when "0011000101110111", -- t[12663] = 1
      "000001" when "0011000101111000", -- t[12664] = 1
      "000001" when "0011000101111001", -- t[12665] = 1
      "000001" when "0011000101111010", -- t[12666] = 1
      "000001" when "0011000101111011", -- t[12667] = 1
      "000001" when "0011000101111100", -- t[12668] = 1
      "000001" when "0011000101111101", -- t[12669] = 1
      "000001" when "0011000101111110", -- t[12670] = 1
      "000001" when "0011000101111111", -- t[12671] = 1
      "000001" when "0011000110000000", -- t[12672] = 1
      "000001" when "0011000110000001", -- t[12673] = 1
      "000001" when "0011000110000010", -- t[12674] = 1
      "000001" when "0011000110000011", -- t[12675] = 1
      "000001" when "0011000110000100", -- t[12676] = 1
      "000001" when "0011000110000101", -- t[12677] = 1
      "000001" when "0011000110000110", -- t[12678] = 1
      "000001" when "0011000110000111", -- t[12679] = 1
      "000001" when "0011000110001000", -- t[12680] = 1
      "000001" when "0011000110001001", -- t[12681] = 1
      "000001" when "0011000110001010", -- t[12682] = 1
      "000001" when "0011000110001011", -- t[12683] = 1
      "000001" when "0011000110001100", -- t[12684] = 1
      "000001" when "0011000110001101", -- t[12685] = 1
      "000001" when "0011000110001110", -- t[12686] = 1
      "000001" when "0011000110001111", -- t[12687] = 1
      "000001" when "0011000110010000", -- t[12688] = 1
      "000001" when "0011000110010001", -- t[12689] = 1
      "000001" when "0011000110010010", -- t[12690] = 1
      "000001" when "0011000110010011", -- t[12691] = 1
      "000001" when "0011000110010100", -- t[12692] = 1
      "000001" when "0011000110010101", -- t[12693] = 1
      "000001" when "0011000110010110", -- t[12694] = 1
      "000001" when "0011000110010111", -- t[12695] = 1
      "000001" when "0011000110011000", -- t[12696] = 1
      "000001" when "0011000110011001", -- t[12697] = 1
      "000001" when "0011000110011010", -- t[12698] = 1
      "000001" when "0011000110011011", -- t[12699] = 1
      "000001" when "0011000110011100", -- t[12700] = 1
      "000001" when "0011000110011101", -- t[12701] = 1
      "000001" when "0011000110011110", -- t[12702] = 1
      "000001" when "0011000110011111", -- t[12703] = 1
      "000001" when "0011000110100000", -- t[12704] = 1
      "000001" when "0011000110100001", -- t[12705] = 1
      "000001" when "0011000110100010", -- t[12706] = 1
      "000001" when "0011000110100011", -- t[12707] = 1
      "000001" when "0011000110100100", -- t[12708] = 1
      "000001" when "0011000110100101", -- t[12709] = 1
      "000001" when "0011000110100110", -- t[12710] = 1
      "000001" when "0011000110100111", -- t[12711] = 1
      "000001" when "0011000110101000", -- t[12712] = 1
      "000001" when "0011000110101001", -- t[12713] = 1
      "000001" when "0011000110101010", -- t[12714] = 1
      "000001" when "0011000110101011", -- t[12715] = 1
      "000001" when "0011000110101100", -- t[12716] = 1
      "000001" when "0011000110101101", -- t[12717] = 1
      "000001" when "0011000110101110", -- t[12718] = 1
      "000001" when "0011000110101111", -- t[12719] = 1
      "000001" when "0011000110110000", -- t[12720] = 1
      "000001" when "0011000110110001", -- t[12721] = 1
      "000001" when "0011000110110010", -- t[12722] = 1
      "000001" when "0011000110110011", -- t[12723] = 1
      "000001" when "0011000110110100", -- t[12724] = 1
      "000001" when "0011000110110101", -- t[12725] = 1
      "000001" when "0011000110110110", -- t[12726] = 1
      "000001" when "0011000110110111", -- t[12727] = 1
      "000001" when "0011000110111000", -- t[12728] = 1
      "000001" when "0011000110111001", -- t[12729] = 1
      "000001" when "0011000110111010", -- t[12730] = 1
      "000001" when "0011000110111011", -- t[12731] = 1
      "000001" when "0011000110111100", -- t[12732] = 1
      "000001" when "0011000110111101", -- t[12733] = 1
      "000001" when "0011000110111110", -- t[12734] = 1
      "000001" when "0011000110111111", -- t[12735] = 1
      "000001" when "0011000111000000", -- t[12736] = 1
      "000001" when "0011000111000001", -- t[12737] = 1
      "000001" when "0011000111000010", -- t[12738] = 1
      "000001" when "0011000111000011", -- t[12739] = 1
      "000001" when "0011000111000100", -- t[12740] = 1
      "000001" when "0011000111000101", -- t[12741] = 1
      "000001" when "0011000111000110", -- t[12742] = 1
      "000001" when "0011000111000111", -- t[12743] = 1
      "000001" when "0011000111001000", -- t[12744] = 1
      "000001" when "0011000111001001", -- t[12745] = 1
      "000001" when "0011000111001010", -- t[12746] = 1
      "000001" when "0011000111001011", -- t[12747] = 1
      "000001" when "0011000111001100", -- t[12748] = 1
      "000001" when "0011000111001101", -- t[12749] = 1
      "000001" when "0011000111001110", -- t[12750] = 1
      "000001" when "0011000111001111", -- t[12751] = 1
      "000001" when "0011000111010000", -- t[12752] = 1
      "000001" when "0011000111010001", -- t[12753] = 1
      "000001" when "0011000111010010", -- t[12754] = 1
      "000001" when "0011000111010011", -- t[12755] = 1
      "000001" when "0011000111010100", -- t[12756] = 1
      "000001" when "0011000111010101", -- t[12757] = 1
      "000001" when "0011000111010110", -- t[12758] = 1
      "000001" when "0011000111010111", -- t[12759] = 1
      "000001" when "0011000111011000", -- t[12760] = 1
      "000001" when "0011000111011001", -- t[12761] = 1
      "000001" when "0011000111011010", -- t[12762] = 1
      "000001" when "0011000111011011", -- t[12763] = 1
      "000001" when "0011000111011100", -- t[12764] = 1
      "000001" when "0011000111011101", -- t[12765] = 1
      "000001" when "0011000111011110", -- t[12766] = 1
      "000001" when "0011000111011111", -- t[12767] = 1
      "000001" when "0011000111100000", -- t[12768] = 1
      "000001" when "0011000111100001", -- t[12769] = 1
      "000001" when "0011000111100010", -- t[12770] = 1
      "000001" when "0011000111100011", -- t[12771] = 1
      "000001" when "0011000111100100", -- t[12772] = 1
      "000001" when "0011000111100101", -- t[12773] = 1
      "000001" when "0011000111100110", -- t[12774] = 1
      "000001" when "0011000111100111", -- t[12775] = 1
      "000001" when "0011000111101000", -- t[12776] = 1
      "000001" when "0011000111101001", -- t[12777] = 1
      "000001" when "0011000111101010", -- t[12778] = 1
      "000001" when "0011000111101011", -- t[12779] = 1
      "000001" when "0011000111101100", -- t[12780] = 1
      "000001" when "0011000111101101", -- t[12781] = 1
      "000001" when "0011000111101110", -- t[12782] = 1
      "000001" when "0011000111101111", -- t[12783] = 1
      "000001" when "0011000111110000", -- t[12784] = 1
      "000001" when "0011000111110001", -- t[12785] = 1
      "000001" when "0011000111110010", -- t[12786] = 1
      "000001" when "0011000111110011", -- t[12787] = 1
      "000001" when "0011000111110100", -- t[12788] = 1
      "000001" when "0011000111110101", -- t[12789] = 1
      "000001" when "0011000111110110", -- t[12790] = 1
      "000001" when "0011000111110111", -- t[12791] = 1
      "000001" when "0011000111111000", -- t[12792] = 1
      "000001" when "0011000111111001", -- t[12793] = 1
      "000001" when "0011000111111010", -- t[12794] = 1
      "000001" when "0011000111111011", -- t[12795] = 1
      "000001" when "0011000111111100", -- t[12796] = 1
      "000001" when "0011000111111101", -- t[12797] = 1
      "000001" when "0011000111111110", -- t[12798] = 1
      "000001" when "0011000111111111", -- t[12799] = 1
      "000001" when "0011001000000000", -- t[12800] = 1
      "000001" when "0011001000000001", -- t[12801] = 1
      "000001" when "0011001000000010", -- t[12802] = 1
      "000001" when "0011001000000011", -- t[12803] = 1
      "000001" when "0011001000000100", -- t[12804] = 1
      "000001" when "0011001000000101", -- t[12805] = 1
      "000001" when "0011001000000110", -- t[12806] = 1
      "000001" when "0011001000000111", -- t[12807] = 1
      "000001" when "0011001000001000", -- t[12808] = 1
      "000001" when "0011001000001001", -- t[12809] = 1
      "000001" when "0011001000001010", -- t[12810] = 1
      "000001" when "0011001000001011", -- t[12811] = 1
      "000001" when "0011001000001100", -- t[12812] = 1
      "000001" when "0011001000001101", -- t[12813] = 1
      "000001" when "0011001000001110", -- t[12814] = 1
      "000001" when "0011001000001111", -- t[12815] = 1
      "000001" when "0011001000010000", -- t[12816] = 1
      "000001" when "0011001000010001", -- t[12817] = 1
      "000001" when "0011001000010010", -- t[12818] = 1
      "000001" when "0011001000010011", -- t[12819] = 1
      "000001" when "0011001000010100", -- t[12820] = 1
      "000001" when "0011001000010101", -- t[12821] = 1
      "000001" when "0011001000010110", -- t[12822] = 1
      "000001" when "0011001000010111", -- t[12823] = 1
      "000001" when "0011001000011000", -- t[12824] = 1
      "000001" when "0011001000011001", -- t[12825] = 1
      "000001" when "0011001000011010", -- t[12826] = 1
      "000001" when "0011001000011011", -- t[12827] = 1
      "000001" when "0011001000011100", -- t[12828] = 1
      "000001" when "0011001000011101", -- t[12829] = 1
      "000001" when "0011001000011110", -- t[12830] = 1
      "000001" when "0011001000011111", -- t[12831] = 1
      "000001" when "0011001000100000", -- t[12832] = 1
      "000001" when "0011001000100001", -- t[12833] = 1
      "000001" when "0011001000100010", -- t[12834] = 1
      "000001" when "0011001000100011", -- t[12835] = 1
      "000001" when "0011001000100100", -- t[12836] = 1
      "000001" when "0011001000100101", -- t[12837] = 1
      "000001" when "0011001000100110", -- t[12838] = 1
      "000001" when "0011001000100111", -- t[12839] = 1
      "000001" when "0011001000101000", -- t[12840] = 1
      "000001" when "0011001000101001", -- t[12841] = 1
      "000001" when "0011001000101010", -- t[12842] = 1
      "000001" when "0011001000101011", -- t[12843] = 1
      "000001" when "0011001000101100", -- t[12844] = 1
      "000001" when "0011001000101101", -- t[12845] = 1
      "000001" when "0011001000101110", -- t[12846] = 1
      "000001" when "0011001000101111", -- t[12847] = 1
      "000001" when "0011001000110000", -- t[12848] = 1
      "000001" when "0011001000110001", -- t[12849] = 1
      "000001" when "0011001000110010", -- t[12850] = 1
      "000001" when "0011001000110011", -- t[12851] = 1
      "000001" when "0011001000110100", -- t[12852] = 1
      "000001" when "0011001000110101", -- t[12853] = 1
      "000001" when "0011001000110110", -- t[12854] = 1
      "000001" when "0011001000110111", -- t[12855] = 1
      "000001" when "0011001000111000", -- t[12856] = 1
      "000001" when "0011001000111001", -- t[12857] = 1
      "000001" when "0011001000111010", -- t[12858] = 1
      "000001" when "0011001000111011", -- t[12859] = 1
      "000001" when "0011001000111100", -- t[12860] = 1
      "000001" when "0011001000111101", -- t[12861] = 1
      "000001" when "0011001000111110", -- t[12862] = 1
      "000001" when "0011001000111111", -- t[12863] = 1
      "000001" when "0011001001000000", -- t[12864] = 1
      "000001" when "0011001001000001", -- t[12865] = 1
      "000001" when "0011001001000010", -- t[12866] = 1
      "000001" when "0011001001000011", -- t[12867] = 1
      "000001" when "0011001001000100", -- t[12868] = 1
      "000001" when "0011001001000101", -- t[12869] = 1
      "000001" when "0011001001000110", -- t[12870] = 1
      "000001" when "0011001001000111", -- t[12871] = 1
      "000001" when "0011001001001000", -- t[12872] = 1
      "000001" when "0011001001001001", -- t[12873] = 1
      "000001" when "0011001001001010", -- t[12874] = 1
      "000001" when "0011001001001011", -- t[12875] = 1
      "000001" when "0011001001001100", -- t[12876] = 1
      "000001" when "0011001001001101", -- t[12877] = 1
      "000001" when "0011001001001110", -- t[12878] = 1
      "000001" when "0011001001001111", -- t[12879] = 1
      "000001" when "0011001001010000", -- t[12880] = 1
      "000001" when "0011001001010001", -- t[12881] = 1
      "000001" when "0011001001010010", -- t[12882] = 1
      "000001" when "0011001001010011", -- t[12883] = 1
      "000001" when "0011001001010100", -- t[12884] = 1
      "000001" when "0011001001010101", -- t[12885] = 1
      "000001" when "0011001001010110", -- t[12886] = 1
      "000001" when "0011001001010111", -- t[12887] = 1
      "000001" when "0011001001011000", -- t[12888] = 1
      "000001" when "0011001001011001", -- t[12889] = 1
      "000001" when "0011001001011010", -- t[12890] = 1
      "000001" when "0011001001011011", -- t[12891] = 1
      "000001" when "0011001001011100", -- t[12892] = 1
      "000001" when "0011001001011101", -- t[12893] = 1
      "000001" when "0011001001011110", -- t[12894] = 1
      "000001" when "0011001001011111", -- t[12895] = 1
      "000001" when "0011001001100000", -- t[12896] = 1
      "000001" when "0011001001100001", -- t[12897] = 1
      "000001" when "0011001001100010", -- t[12898] = 1
      "000001" when "0011001001100011", -- t[12899] = 1
      "000001" when "0011001001100100", -- t[12900] = 1
      "000001" when "0011001001100101", -- t[12901] = 1
      "000001" when "0011001001100110", -- t[12902] = 1
      "000001" when "0011001001100111", -- t[12903] = 1
      "000001" when "0011001001101000", -- t[12904] = 1
      "000001" when "0011001001101001", -- t[12905] = 1
      "000001" when "0011001001101010", -- t[12906] = 1
      "000001" when "0011001001101011", -- t[12907] = 1
      "000001" when "0011001001101100", -- t[12908] = 1
      "000001" when "0011001001101101", -- t[12909] = 1
      "000001" when "0011001001101110", -- t[12910] = 1
      "000001" when "0011001001101111", -- t[12911] = 1
      "000001" when "0011001001110000", -- t[12912] = 1
      "000001" when "0011001001110001", -- t[12913] = 1
      "000001" when "0011001001110010", -- t[12914] = 1
      "000001" when "0011001001110011", -- t[12915] = 1
      "000001" when "0011001001110100", -- t[12916] = 1
      "000001" when "0011001001110101", -- t[12917] = 1
      "000001" when "0011001001110110", -- t[12918] = 1
      "000001" when "0011001001110111", -- t[12919] = 1
      "000001" when "0011001001111000", -- t[12920] = 1
      "000001" when "0011001001111001", -- t[12921] = 1
      "000001" when "0011001001111010", -- t[12922] = 1
      "000001" when "0011001001111011", -- t[12923] = 1
      "000001" when "0011001001111100", -- t[12924] = 1
      "000001" when "0011001001111101", -- t[12925] = 1
      "000001" when "0011001001111110", -- t[12926] = 1
      "000001" when "0011001001111111", -- t[12927] = 1
      "000001" when "0011001010000000", -- t[12928] = 1
      "000001" when "0011001010000001", -- t[12929] = 1
      "000001" when "0011001010000010", -- t[12930] = 1
      "000001" when "0011001010000011", -- t[12931] = 1
      "000001" when "0011001010000100", -- t[12932] = 1
      "000001" when "0011001010000101", -- t[12933] = 1
      "000001" when "0011001010000110", -- t[12934] = 1
      "000001" when "0011001010000111", -- t[12935] = 1
      "000001" when "0011001010001000", -- t[12936] = 1
      "000001" when "0011001010001001", -- t[12937] = 1
      "000001" when "0011001010001010", -- t[12938] = 1
      "000001" when "0011001010001011", -- t[12939] = 1
      "000001" when "0011001010001100", -- t[12940] = 1
      "000001" when "0011001010001101", -- t[12941] = 1
      "000001" when "0011001010001110", -- t[12942] = 1
      "000001" when "0011001010001111", -- t[12943] = 1
      "000001" when "0011001010010000", -- t[12944] = 1
      "000001" when "0011001010010001", -- t[12945] = 1
      "000001" when "0011001010010010", -- t[12946] = 1
      "000001" when "0011001010010011", -- t[12947] = 1
      "000001" when "0011001010010100", -- t[12948] = 1
      "000001" when "0011001010010101", -- t[12949] = 1
      "000001" when "0011001010010110", -- t[12950] = 1
      "000001" when "0011001010010111", -- t[12951] = 1
      "000001" when "0011001010011000", -- t[12952] = 1
      "000001" when "0011001010011001", -- t[12953] = 1
      "000001" when "0011001010011010", -- t[12954] = 1
      "000001" when "0011001010011011", -- t[12955] = 1
      "000001" when "0011001010011100", -- t[12956] = 1
      "000001" when "0011001010011101", -- t[12957] = 1
      "000001" when "0011001010011110", -- t[12958] = 1
      "000001" when "0011001010011111", -- t[12959] = 1
      "000001" when "0011001010100000", -- t[12960] = 1
      "000001" when "0011001010100001", -- t[12961] = 1
      "000001" when "0011001010100010", -- t[12962] = 1
      "000001" when "0011001010100011", -- t[12963] = 1
      "000001" when "0011001010100100", -- t[12964] = 1
      "000001" when "0011001010100101", -- t[12965] = 1
      "000001" when "0011001010100110", -- t[12966] = 1
      "000001" when "0011001010100111", -- t[12967] = 1
      "000001" when "0011001010101000", -- t[12968] = 1
      "000001" when "0011001010101001", -- t[12969] = 1
      "000001" when "0011001010101010", -- t[12970] = 1
      "000001" when "0011001010101011", -- t[12971] = 1
      "000001" when "0011001010101100", -- t[12972] = 1
      "000001" when "0011001010101101", -- t[12973] = 1
      "000001" when "0011001010101110", -- t[12974] = 1
      "000001" when "0011001010101111", -- t[12975] = 1
      "000001" when "0011001010110000", -- t[12976] = 1
      "000001" when "0011001010110001", -- t[12977] = 1
      "000001" when "0011001010110010", -- t[12978] = 1
      "000001" when "0011001010110011", -- t[12979] = 1
      "000001" when "0011001010110100", -- t[12980] = 1
      "000001" when "0011001010110101", -- t[12981] = 1
      "000001" when "0011001010110110", -- t[12982] = 1
      "000001" when "0011001010110111", -- t[12983] = 1
      "000001" when "0011001010111000", -- t[12984] = 1
      "000001" when "0011001010111001", -- t[12985] = 1
      "000001" when "0011001010111010", -- t[12986] = 1
      "000001" when "0011001010111011", -- t[12987] = 1
      "000001" when "0011001010111100", -- t[12988] = 1
      "000001" when "0011001010111101", -- t[12989] = 1
      "000001" when "0011001010111110", -- t[12990] = 1
      "000001" when "0011001010111111", -- t[12991] = 1
      "000001" when "0011001011000000", -- t[12992] = 1
      "000001" when "0011001011000001", -- t[12993] = 1
      "000001" when "0011001011000010", -- t[12994] = 1
      "000001" when "0011001011000011", -- t[12995] = 1
      "000001" when "0011001011000100", -- t[12996] = 1
      "000001" when "0011001011000101", -- t[12997] = 1
      "000001" when "0011001011000110", -- t[12998] = 1
      "000001" when "0011001011000111", -- t[12999] = 1
      "000001" when "0011001011001000", -- t[13000] = 1
      "000001" when "0011001011001001", -- t[13001] = 1
      "000001" when "0011001011001010", -- t[13002] = 1
      "000001" when "0011001011001011", -- t[13003] = 1
      "000001" when "0011001011001100", -- t[13004] = 1
      "000001" when "0011001011001101", -- t[13005] = 1
      "000001" when "0011001011001110", -- t[13006] = 1
      "000001" when "0011001011001111", -- t[13007] = 1
      "000001" when "0011001011010000", -- t[13008] = 1
      "000001" when "0011001011010001", -- t[13009] = 1
      "000001" when "0011001011010010", -- t[13010] = 1
      "000001" when "0011001011010011", -- t[13011] = 1
      "000001" when "0011001011010100", -- t[13012] = 1
      "000001" when "0011001011010101", -- t[13013] = 1
      "000001" when "0011001011010110", -- t[13014] = 1
      "000001" when "0011001011010111", -- t[13015] = 1
      "000001" when "0011001011011000", -- t[13016] = 1
      "000001" when "0011001011011001", -- t[13017] = 1
      "000001" when "0011001011011010", -- t[13018] = 1
      "000001" when "0011001011011011", -- t[13019] = 1
      "000001" when "0011001011011100", -- t[13020] = 1
      "000001" when "0011001011011101", -- t[13021] = 1
      "000001" when "0011001011011110", -- t[13022] = 1
      "000001" when "0011001011011111", -- t[13023] = 1
      "000001" when "0011001011100000", -- t[13024] = 1
      "000001" when "0011001011100001", -- t[13025] = 1
      "000001" when "0011001011100010", -- t[13026] = 1
      "000001" when "0011001011100011", -- t[13027] = 1
      "000001" when "0011001011100100", -- t[13028] = 1
      "000001" when "0011001011100101", -- t[13029] = 1
      "000001" when "0011001011100110", -- t[13030] = 1
      "000001" when "0011001011100111", -- t[13031] = 1
      "000001" when "0011001011101000", -- t[13032] = 1
      "000001" when "0011001011101001", -- t[13033] = 1
      "000001" when "0011001011101010", -- t[13034] = 1
      "000001" when "0011001011101011", -- t[13035] = 1
      "000001" when "0011001011101100", -- t[13036] = 1
      "000001" when "0011001011101101", -- t[13037] = 1
      "000001" when "0011001011101110", -- t[13038] = 1
      "000001" when "0011001011101111", -- t[13039] = 1
      "000001" when "0011001011110000", -- t[13040] = 1
      "000001" when "0011001011110001", -- t[13041] = 1
      "000001" when "0011001011110010", -- t[13042] = 1
      "000001" when "0011001011110011", -- t[13043] = 1
      "000001" when "0011001011110100", -- t[13044] = 1
      "000001" when "0011001011110101", -- t[13045] = 1
      "000001" when "0011001011110110", -- t[13046] = 1
      "000001" when "0011001011110111", -- t[13047] = 1
      "000001" when "0011001011111000", -- t[13048] = 1
      "000001" when "0011001011111001", -- t[13049] = 1
      "000001" when "0011001011111010", -- t[13050] = 1
      "000001" when "0011001011111011", -- t[13051] = 1
      "000001" when "0011001011111100", -- t[13052] = 1
      "000001" when "0011001011111101", -- t[13053] = 1
      "000001" when "0011001011111110", -- t[13054] = 1
      "000001" when "0011001011111111", -- t[13055] = 1
      "000001" when "0011001100000000", -- t[13056] = 1
      "000001" when "0011001100000001", -- t[13057] = 1
      "000001" when "0011001100000010", -- t[13058] = 1
      "000001" when "0011001100000011", -- t[13059] = 1
      "000001" when "0011001100000100", -- t[13060] = 1
      "000001" when "0011001100000101", -- t[13061] = 1
      "000001" when "0011001100000110", -- t[13062] = 1
      "000001" when "0011001100000111", -- t[13063] = 1
      "000001" when "0011001100001000", -- t[13064] = 1
      "000001" when "0011001100001001", -- t[13065] = 1
      "000001" when "0011001100001010", -- t[13066] = 1
      "000001" when "0011001100001011", -- t[13067] = 1
      "000001" when "0011001100001100", -- t[13068] = 1
      "000001" when "0011001100001101", -- t[13069] = 1
      "000001" when "0011001100001110", -- t[13070] = 1
      "000001" when "0011001100001111", -- t[13071] = 1
      "000001" when "0011001100010000", -- t[13072] = 1
      "000001" when "0011001100010001", -- t[13073] = 1
      "000001" when "0011001100010010", -- t[13074] = 1
      "000001" when "0011001100010011", -- t[13075] = 1
      "000001" when "0011001100010100", -- t[13076] = 1
      "000001" when "0011001100010101", -- t[13077] = 1
      "000001" when "0011001100010110", -- t[13078] = 1
      "000001" when "0011001100010111", -- t[13079] = 1
      "000001" when "0011001100011000", -- t[13080] = 1
      "000001" when "0011001100011001", -- t[13081] = 1
      "000001" when "0011001100011010", -- t[13082] = 1
      "000001" when "0011001100011011", -- t[13083] = 1
      "000001" when "0011001100011100", -- t[13084] = 1
      "000001" when "0011001100011101", -- t[13085] = 1
      "000001" when "0011001100011110", -- t[13086] = 1
      "000001" when "0011001100011111", -- t[13087] = 1
      "000001" when "0011001100100000", -- t[13088] = 1
      "000001" when "0011001100100001", -- t[13089] = 1
      "000001" when "0011001100100010", -- t[13090] = 1
      "000001" when "0011001100100011", -- t[13091] = 1
      "000001" when "0011001100100100", -- t[13092] = 1
      "000001" when "0011001100100101", -- t[13093] = 1
      "000001" when "0011001100100110", -- t[13094] = 1
      "000001" when "0011001100100111", -- t[13095] = 1
      "000001" when "0011001100101000", -- t[13096] = 1
      "000001" when "0011001100101001", -- t[13097] = 1
      "000001" when "0011001100101010", -- t[13098] = 1
      "000001" when "0011001100101011", -- t[13099] = 1
      "000001" when "0011001100101100", -- t[13100] = 1
      "000001" when "0011001100101101", -- t[13101] = 1
      "000001" when "0011001100101110", -- t[13102] = 1
      "000001" when "0011001100101111", -- t[13103] = 1
      "000001" when "0011001100110000", -- t[13104] = 1
      "000001" when "0011001100110001", -- t[13105] = 1
      "000001" when "0011001100110010", -- t[13106] = 1
      "000001" when "0011001100110011", -- t[13107] = 1
      "000001" when "0011001100110100", -- t[13108] = 1
      "000001" when "0011001100110101", -- t[13109] = 1
      "000001" when "0011001100110110", -- t[13110] = 1
      "000001" when "0011001100110111", -- t[13111] = 1
      "000001" when "0011001100111000", -- t[13112] = 1
      "000001" when "0011001100111001", -- t[13113] = 1
      "000001" when "0011001100111010", -- t[13114] = 1
      "000001" when "0011001100111011", -- t[13115] = 1
      "000001" when "0011001100111100", -- t[13116] = 1
      "000001" when "0011001100111101", -- t[13117] = 1
      "000001" when "0011001100111110", -- t[13118] = 1
      "000001" when "0011001100111111", -- t[13119] = 1
      "000001" when "0011001101000000", -- t[13120] = 1
      "000001" when "0011001101000001", -- t[13121] = 1
      "000001" when "0011001101000010", -- t[13122] = 1
      "000001" when "0011001101000011", -- t[13123] = 1
      "000001" when "0011001101000100", -- t[13124] = 1
      "000001" when "0011001101000101", -- t[13125] = 1
      "000001" when "0011001101000110", -- t[13126] = 1
      "000001" when "0011001101000111", -- t[13127] = 1
      "000001" when "0011001101001000", -- t[13128] = 1
      "000001" when "0011001101001001", -- t[13129] = 1
      "000001" when "0011001101001010", -- t[13130] = 1
      "000001" when "0011001101001011", -- t[13131] = 1
      "000001" when "0011001101001100", -- t[13132] = 1
      "000001" when "0011001101001101", -- t[13133] = 1
      "000001" when "0011001101001110", -- t[13134] = 1
      "000001" when "0011001101001111", -- t[13135] = 1
      "000001" when "0011001101010000", -- t[13136] = 1
      "000001" when "0011001101010001", -- t[13137] = 1
      "000001" when "0011001101010010", -- t[13138] = 1
      "000001" when "0011001101010011", -- t[13139] = 1
      "000001" when "0011001101010100", -- t[13140] = 1
      "000001" when "0011001101010101", -- t[13141] = 1
      "000001" when "0011001101010110", -- t[13142] = 1
      "000001" when "0011001101010111", -- t[13143] = 1
      "000001" when "0011001101011000", -- t[13144] = 1
      "000001" when "0011001101011001", -- t[13145] = 1
      "000001" when "0011001101011010", -- t[13146] = 1
      "000001" when "0011001101011011", -- t[13147] = 1
      "000001" when "0011001101011100", -- t[13148] = 1
      "000001" when "0011001101011101", -- t[13149] = 1
      "000001" when "0011001101011110", -- t[13150] = 1
      "000001" when "0011001101011111", -- t[13151] = 1
      "000001" when "0011001101100000", -- t[13152] = 1
      "000001" when "0011001101100001", -- t[13153] = 1
      "000001" when "0011001101100010", -- t[13154] = 1
      "000001" when "0011001101100011", -- t[13155] = 1
      "000001" when "0011001101100100", -- t[13156] = 1
      "000001" when "0011001101100101", -- t[13157] = 1
      "000001" when "0011001101100110", -- t[13158] = 1
      "000001" when "0011001101100111", -- t[13159] = 1
      "000001" when "0011001101101000", -- t[13160] = 1
      "000001" when "0011001101101001", -- t[13161] = 1
      "000001" when "0011001101101010", -- t[13162] = 1
      "000001" when "0011001101101011", -- t[13163] = 1
      "000001" when "0011001101101100", -- t[13164] = 1
      "000001" when "0011001101101101", -- t[13165] = 1
      "000001" when "0011001101101110", -- t[13166] = 1
      "000001" when "0011001101101111", -- t[13167] = 1
      "000001" when "0011001101110000", -- t[13168] = 1
      "000001" when "0011001101110001", -- t[13169] = 1
      "000001" when "0011001101110010", -- t[13170] = 1
      "000001" when "0011001101110011", -- t[13171] = 1
      "000001" when "0011001101110100", -- t[13172] = 1
      "000001" when "0011001101110101", -- t[13173] = 1
      "000001" when "0011001101110110", -- t[13174] = 1
      "000001" when "0011001101110111", -- t[13175] = 1
      "000001" when "0011001101111000", -- t[13176] = 1
      "000001" when "0011001101111001", -- t[13177] = 1
      "000001" when "0011001101111010", -- t[13178] = 1
      "000001" when "0011001101111011", -- t[13179] = 1
      "000001" when "0011001101111100", -- t[13180] = 1
      "000001" when "0011001101111101", -- t[13181] = 1
      "000001" when "0011001101111110", -- t[13182] = 1
      "000001" when "0011001101111111", -- t[13183] = 1
      "000001" when "0011001110000000", -- t[13184] = 1
      "000001" when "0011001110000001", -- t[13185] = 1
      "000001" when "0011001110000010", -- t[13186] = 1
      "000001" when "0011001110000011", -- t[13187] = 1
      "000001" when "0011001110000100", -- t[13188] = 1
      "000001" when "0011001110000101", -- t[13189] = 1
      "000001" when "0011001110000110", -- t[13190] = 1
      "000001" when "0011001110000111", -- t[13191] = 1
      "000001" when "0011001110001000", -- t[13192] = 1
      "000001" when "0011001110001001", -- t[13193] = 1
      "000001" when "0011001110001010", -- t[13194] = 1
      "000001" when "0011001110001011", -- t[13195] = 1
      "000001" when "0011001110001100", -- t[13196] = 1
      "000001" when "0011001110001101", -- t[13197] = 1
      "000001" when "0011001110001110", -- t[13198] = 1
      "000001" when "0011001110001111", -- t[13199] = 1
      "000001" when "0011001110010000", -- t[13200] = 1
      "000001" when "0011001110010001", -- t[13201] = 1
      "000001" when "0011001110010010", -- t[13202] = 1
      "000001" when "0011001110010011", -- t[13203] = 1
      "000001" when "0011001110010100", -- t[13204] = 1
      "000001" when "0011001110010101", -- t[13205] = 1
      "000001" when "0011001110010110", -- t[13206] = 1
      "000001" when "0011001110010111", -- t[13207] = 1
      "000001" when "0011001110011000", -- t[13208] = 1
      "000001" when "0011001110011001", -- t[13209] = 1
      "000001" when "0011001110011010", -- t[13210] = 1
      "000001" when "0011001110011011", -- t[13211] = 1
      "000001" when "0011001110011100", -- t[13212] = 1
      "000001" when "0011001110011101", -- t[13213] = 1
      "000001" when "0011001110011110", -- t[13214] = 1
      "000001" when "0011001110011111", -- t[13215] = 1
      "000001" when "0011001110100000", -- t[13216] = 1
      "000001" when "0011001110100001", -- t[13217] = 1
      "000001" when "0011001110100010", -- t[13218] = 1
      "000001" when "0011001110100011", -- t[13219] = 1
      "000001" when "0011001110100100", -- t[13220] = 1
      "000001" when "0011001110100101", -- t[13221] = 1
      "000001" when "0011001110100110", -- t[13222] = 1
      "000001" when "0011001110100111", -- t[13223] = 1
      "000001" when "0011001110101000", -- t[13224] = 1
      "000001" when "0011001110101001", -- t[13225] = 1
      "000001" when "0011001110101010", -- t[13226] = 1
      "000001" when "0011001110101011", -- t[13227] = 1
      "000001" when "0011001110101100", -- t[13228] = 1
      "000001" when "0011001110101101", -- t[13229] = 1
      "000001" when "0011001110101110", -- t[13230] = 1
      "000001" when "0011001110101111", -- t[13231] = 1
      "000001" when "0011001110110000", -- t[13232] = 1
      "000001" when "0011001110110001", -- t[13233] = 1
      "000001" when "0011001110110010", -- t[13234] = 1
      "000001" when "0011001110110011", -- t[13235] = 1
      "000001" when "0011001110110100", -- t[13236] = 1
      "000001" when "0011001110110101", -- t[13237] = 1
      "000001" when "0011001110110110", -- t[13238] = 1
      "000001" when "0011001110110111", -- t[13239] = 1
      "000001" when "0011001110111000", -- t[13240] = 1
      "000001" when "0011001110111001", -- t[13241] = 1
      "000001" when "0011001110111010", -- t[13242] = 1
      "000001" when "0011001110111011", -- t[13243] = 1
      "000001" when "0011001110111100", -- t[13244] = 1
      "000001" when "0011001110111101", -- t[13245] = 1
      "000001" when "0011001110111110", -- t[13246] = 1
      "000001" when "0011001110111111", -- t[13247] = 1
      "000001" when "0011001111000000", -- t[13248] = 1
      "000001" when "0011001111000001", -- t[13249] = 1
      "000001" when "0011001111000010", -- t[13250] = 1
      "000001" when "0011001111000011", -- t[13251] = 1
      "000001" when "0011001111000100", -- t[13252] = 1
      "000001" when "0011001111000101", -- t[13253] = 1
      "000001" when "0011001111000110", -- t[13254] = 1
      "000001" when "0011001111000111", -- t[13255] = 1
      "000001" when "0011001111001000", -- t[13256] = 1
      "000001" when "0011001111001001", -- t[13257] = 1
      "000001" when "0011001111001010", -- t[13258] = 1
      "000001" when "0011001111001011", -- t[13259] = 1
      "000001" when "0011001111001100", -- t[13260] = 1
      "000001" when "0011001111001101", -- t[13261] = 1
      "000001" when "0011001111001110", -- t[13262] = 1
      "000001" when "0011001111001111", -- t[13263] = 1
      "000001" when "0011001111010000", -- t[13264] = 1
      "000001" when "0011001111010001", -- t[13265] = 1
      "000001" when "0011001111010010", -- t[13266] = 1
      "000001" when "0011001111010011", -- t[13267] = 1
      "000001" when "0011001111010100", -- t[13268] = 1
      "000001" when "0011001111010101", -- t[13269] = 1
      "000001" when "0011001111010110", -- t[13270] = 1
      "000001" when "0011001111010111", -- t[13271] = 1
      "000001" when "0011001111011000", -- t[13272] = 1
      "000001" when "0011001111011001", -- t[13273] = 1
      "000001" when "0011001111011010", -- t[13274] = 1
      "000001" when "0011001111011011", -- t[13275] = 1
      "000001" when "0011001111011100", -- t[13276] = 1
      "000001" when "0011001111011101", -- t[13277] = 1
      "000001" when "0011001111011110", -- t[13278] = 1
      "000001" when "0011001111011111", -- t[13279] = 1
      "000001" when "0011001111100000", -- t[13280] = 1
      "000001" when "0011001111100001", -- t[13281] = 1
      "000001" when "0011001111100010", -- t[13282] = 1
      "000001" when "0011001111100011", -- t[13283] = 1
      "000001" when "0011001111100100", -- t[13284] = 1
      "000001" when "0011001111100101", -- t[13285] = 1
      "000001" when "0011001111100110", -- t[13286] = 1
      "000001" when "0011001111100111", -- t[13287] = 1
      "000001" when "0011001111101000", -- t[13288] = 1
      "000001" when "0011001111101001", -- t[13289] = 1
      "000001" when "0011001111101010", -- t[13290] = 1
      "000001" when "0011001111101011", -- t[13291] = 1
      "000001" when "0011001111101100", -- t[13292] = 1
      "000001" when "0011001111101101", -- t[13293] = 1
      "000001" when "0011001111101110", -- t[13294] = 1
      "000001" when "0011001111101111", -- t[13295] = 1
      "000001" when "0011001111110000", -- t[13296] = 1
      "000001" when "0011001111110001", -- t[13297] = 1
      "000001" when "0011001111110010", -- t[13298] = 1
      "000001" when "0011001111110011", -- t[13299] = 1
      "000001" when "0011001111110100", -- t[13300] = 1
      "000001" when "0011001111110101", -- t[13301] = 1
      "000001" when "0011001111110110", -- t[13302] = 1
      "000001" when "0011001111110111", -- t[13303] = 1
      "000001" when "0011001111111000", -- t[13304] = 1
      "000001" when "0011001111111001", -- t[13305] = 1
      "000001" when "0011001111111010", -- t[13306] = 1
      "000001" when "0011001111111011", -- t[13307] = 1
      "000001" when "0011001111111100", -- t[13308] = 1
      "000001" when "0011001111111101", -- t[13309] = 1
      "000001" when "0011001111111110", -- t[13310] = 1
      "000001" when "0011001111111111", -- t[13311] = 1
      "000001" when "0011010000000000", -- t[13312] = 1
      "000001" when "0011010000000001", -- t[13313] = 1
      "000001" when "0011010000000010", -- t[13314] = 1
      "000001" when "0011010000000011", -- t[13315] = 1
      "000001" when "0011010000000100", -- t[13316] = 1
      "000001" when "0011010000000101", -- t[13317] = 1
      "000001" when "0011010000000110", -- t[13318] = 1
      "000001" when "0011010000000111", -- t[13319] = 1
      "000001" when "0011010000001000", -- t[13320] = 1
      "000001" when "0011010000001001", -- t[13321] = 1
      "000001" when "0011010000001010", -- t[13322] = 1
      "000001" when "0011010000001011", -- t[13323] = 1
      "000001" when "0011010000001100", -- t[13324] = 1
      "000001" when "0011010000001101", -- t[13325] = 1
      "000001" when "0011010000001110", -- t[13326] = 1
      "000001" when "0011010000001111", -- t[13327] = 1
      "000001" when "0011010000010000", -- t[13328] = 1
      "000001" when "0011010000010001", -- t[13329] = 1
      "000001" when "0011010000010010", -- t[13330] = 1
      "000001" when "0011010000010011", -- t[13331] = 1
      "000001" when "0011010000010100", -- t[13332] = 1
      "000001" when "0011010000010101", -- t[13333] = 1
      "000001" when "0011010000010110", -- t[13334] = 1
      "000001" when "0011010000010111", -- t[13335] = 1
      "000001" when "0011010000011000", -- t[13336] = 1
      "000001" when "0011010000011001", -- t[13337] = 1
      "000001" when "0011010000011010", -- t[13338] = 1
      "000001" when "0011010000011011", -- t[13339] = 1
      "000001" when "0011010000011100", -- t[13340] = 1
      "000001" when "0011010000011101", -- t[13341] = 1
      "000001" when "0011010000011110", -- t[13342] = 1
      "000001" when "0011010000011111", -- t[13343] = 1
      "000001" when "0011010000100000", -- t[13344] = 1
      "000001" when "0011010000100001", -- t[13345] = 1
      "000001" when "0011010000100010", -- t[13346] = 1
      "000001" when "0011010000100011", -- t[13347] = 1
      "000001" when "0011010000100100", -- t[13348] = 1
      "000001" when "0011010000100101", -- t[13349] = 1
      "000001" when "0011010000100110", -- t[13350] = 1
      "000001" when "0011010000100111", -- t[13351] = 1
      "000001" when "0011010000101000", -- t[13352] = 1
      "000001" when "0011010000101001", -- t[13353] = 1
      "000001" when "0011010000101010", -- t[13354] = 1
      "000001" when "0011010000101011", -- t[13355] = 1
      "000001" when "0011010000101100", -- t[13356] = 1
      "000001" when "0011010000101101", -- t[13357] = 1
      "000001" when "0011010000101110", -- t[13358] = 1
      "000001" when "0011010000101111", -- t[13359] = 1
      "000001" when "0011010000110000", -- t[13360] = 1
      "000001" when "0011010000110001", -- t[13361] = 1
      "000001" when "0011010000110010", -- t[13362] = 1
      "000001" when "0011010000110011", -- t[13363] = 1
      "000001" when "0011010000110100", -- t[13364] = 1
      "000001" when "0011010000110101", -- t[13365] = 1
      "000001" when "0011010000110110", -- t[13366] = 1
      "000001" when "0011010000110111", -- t[13367] = 1
      "000001" when "0011010000111000", -- t[13368] = 1
      "000001" when "0011010000111001", -- t[13369] = 1
      "000001" when "0011010000111010", -- t[13370] = 1
      "000001" when "0011010000111011", -- t[13371] = 1
      "000001" when "0011010000111100", -- t[13372] = 1
      "000001" when "0011010000111101", -- t[13373] = 1
      "000001" when "0011010000111110", -- t[13374] = 1
      "000001" when "0011010000111111", -- t[13375] = 1
      "000001" when "0011010001000000", -- t[13376] = 1
      "000001" when "0011010001000001", -- t[13377] = 1
      "000001" when "0011010001000010", -- t[13378] = 1
      "000001" when "0011010001000011", -- t[13379] = 1
      "000001" when "0011010001000100", -- t[13380] = 1
      "000001" when "0011010001000101", -- t[13381] = 1
      "000001" when "0011010001000110", -- t[13382] = 1
      "000001" when "0011010001000111", -- t[13383] = 1
      "000001" when "0011010001001000", -- t[13384] = 1
      "000001" when "0011010001001001", -- t[13385] = 1
      "000001" when "0011010001001010", -- t[13386] = 1
      "000001" when "0011010001001011", -- t[13387] = 1
      "000001" when "0011010001001100", -- t[13388] = 1
      "000001" when "0011010001001101", -- t[13389] = 1
      "000001" when "0011010001001110", -- t[13390] = 1
      "000001" when "0011010001001111", -- t[13391] = 1
      "000001" when "0011010001010000", -- t[13392] = 1
      "000001" when "0011010001010001", -- t[13393] = 1
      "000001" when "0011010001010010", -- t[13394] = 1
      "000001" when "0011010001010011", -- t[13395] = 1
      "000001" when "0011010001010100", -- t[13396] = 1
      "000001" when "0011010001010101", -- t[13397] = 1
      "000001" when "0011010001010110", -- t[13398] = 1
      "000001" when "0011010001010111", -- t[13399] = 1
      "000001" when "0011010001011000", -- t[13400] = 1
      "000001" when "0011010001011001", -- t[13401] = 1
      "000001" when "0011010001011010", -- t[13402] = 1
      "000001" when "0011010001011011", -- t[13403] = 1
      "000001" when "0011010001011100", -- t[13404] = 1
      "000001" when "0011010001011101", -- t[13405] = 1
      "000001" when "0011010001011110", -- t[13406] = 1
      "000001" when "0011010001011111", -- t[13407] = 1
      "000001" when "0011010001100000", -- t[13408] = 1
      "000001" when "0011010001100001", -- t[13409] = 1
      "000001" when "0011010001100010", -- t[13410] = 1
      "000001" when "0011010001100011", -- t[13411] = 1
      "000001" when "0011010001100100", -- t[13412] = 1
      "000001" when "0011010001100101", -- t[13413] = 1
      "000001" when "0011010001100110", -- t[13414] = 1
      "000001" when "0011010001100111", -- t[13415] = 1
      "000001" when "0011010001101000", -- t[13416] = 1
      "000001" when "0011010001101001", -- t[13417] = 1
      "000001" when "0011010001101010", -- t[13418] = 1
      "000001" when "0011010001101011", -- t[13419] = 1
      "000001" when "0011010001101100", -- t[13420] = 1
      "000001" when "0011010001101101", -- t[13421] = 1
      "000001" when "0011010001101110", -- t[13422] = 1
      "000001" when "0011010001101111", -- t[13423] = 1
      "000001" when "0011010001110000", -- t[13424] = 1
      "000001" when "0011010001110001", -- t[13425] = 1
      "000001" when "0011010001110010", -- t[13426] = 1
      "000001" when "0011010001110011", -- t[13427] = 1
      "000001" when "0011010001110100", -- t[13428] = 1
      "000001" when "0011010001110101", -- t[13429] = 1
      "000001" when "0011010001110110", -- t[13430] = 1
      "000001" when "0011010001110111", -- t[13431] = 1
      "000001" when "0011010001111000", -- t[13432] = 1
      "000001" when "0011010001111001", -- t[13433] = 1
      "000001" when "0011010001111010", -- t[13434] = 1
      "000001" when "0011010001111011", -- t[13435] = 1
      "000001" when "0011010001111100", -- t[13436] = 1
      "000001" when "0011010001111101", -- t[13437] = 1
      "000001" when "0011010001111110", -- t[13438] = 1
      "000001" when "0011010001111111", -- t[13439] = 1
      "000001" when "0011010010000000", -- t[13440] = 1
      "000001" when "0011010010000001", -- t[13441] = 1
      "000001" when "0011010010000010", -- t[13442] = 1
      "000001" when "0011010010000011", -- t[13443] = 1
      "000001" when "0011010010000100", -- t[13444] = 1
      "000001" when "0011010010000101", -- t[13445] = 1
      "000001" when "0011010010000110", -- t[13446] = 1
      "000001" when "0011010010000111", -- t[13447] = 1
      "000001" when "0011010010001000", -- t[13448] = 1
      "000001" when "0011010010001001", -- t[13449] = 1
      "000001" when "0011010010001010", -- t[13450] = 1
      "000001" when "0011010010001011", -- t[13451] = 1
      "000001" when "0011010010001100", -- t[13452] = 1
      "000001" when "0011010010001101", -- t[13453] = 1
      "000001" when "0011010010001110", -- t[13454] = 1
      "000001" when "0011010010001111", -- t[13455] = 1
      "000001" when "0011010010010000", -- t[13456] = 1
      "000001" when "0011010010010001", -- t[13457] = 1
      "000001" when "0011010010010010", -- t[13458] = 1
      "000001" when "0011010010010011", -- t[13459] = 1
      "000001" when "0011010010010100", -- t[13460] = 1
      "000001" when "0011010010010101", -- t[13461] = 1
      "000001" when "0011010010010110", -- t[13462] = 1
      "000001" when "0011010010010111", -- t[13463] = 1
      "000001" when "0011010010011000", -- t[13464] = 1
      "000001" when "0011010010011001", -- t[13465] = 1
      "000001" when "0011010010011010", -- t[13466] = 1
      "000001" when "0011010010011011", -- t[13467] = 1
      "000001" when "0011010010011100", -- t[13468] = 1
      "000001" when "0011010010011101", -- t[13469] = 1
      "000001" when "0011010010011110", -- t[13470] = 1
      "000001" when "0011010010011111", -- t[13471] = 1
      "000001" when "0011010010100000", -- t[13472] = 1
      "000001" when "0011010010100001", -- t[13473] = 1
      "000001" when "0011010010100010", -- t[13474] = 1
      "000001" when "0011010010100011", -- t[13475] = 1
      "000001" when "0011010010100100", -- t[13476] = 1
      "000001" when "0011010010100101", -- t[13477] = 1
      "000001" when "0011010010100110", -- t[13478] = 1
      "000001" when "0011010010100111", -- t[13479] = 1
      "000001" when "0011010010101000", -- t[13480] = 1
      "000001" when "0011010010101001", -- t[13481] = 1
      "000001" when "0011010010101010", -- t[13482] = 1
      "000001" when "0011010010101011", -- t[13483] = 1
      "000001" when "0011010010101100", -- t[13484] = 1
      "000001" when "0011010010101101", -- t[13485] = 1
      "000001" when "0011010010101110", -- t[13486] = 1
      "000001" when "0011010010101111", -- t[13487] = 1
      "000001" when "0011010010110000", -- t[13488] = 1
      "000001" when "0011010010110001", -- t[13489] = 1
      "000001" when "0011010010110010", -- t[13490] = 1
      "000001" when "0011010010110011", -- t[13491] = 1
      "000001" when "0011010010110100", -- t[13492] = 1
      "000001" when "0011010010110101", -- t[13493] = 1
      "000001" when "0011010010110110", -- t[13494] = 1
      "000001" when "0011010010110111", -- t[13495] = 1
      "000001" when "0011010010111000", -- t[13496] = 1
      "000001" when "0011010010111001", -- t[13497] = 1
      "000001" when "0011010010111010", -- t[13498] = 1
      "000001" when "0011010010111011", -- t[13499] = 1
      "000001" when "0011010010111100", -- t[13500] = 1
      "000001" when "0011010010111101", -- t[13501] = 1
      "000001" when "0011010010111110", -- t[13502] = 1
      "000001" when "0011010010111111", -- t[13503] = 1
      "000001" when "0011010011000000", -- t[13504] = 1
      "000001" when "0011010011000001", -- t[13505] = 1
      "000001" when "0011010011000010", -- t[13506] = 1
      "000001" when "0011010011000011", -- t[13507] = 1
      "000001" when "0011010011000100", -- t[13508] = 1
      "000001" when "0011010011000101", -- t[13509] = 1
      "000001" when "0011010011000110", -- t[13510] = 1
      "000001" when "0011010011000111", -- t[13511] = 1
      "000001" when "0011010011001000", -- t[13512] = 1
      "000001" when "0011010011001001", -- t[13513] = 1
      "000001" when "0011010011001010", -- t[13514] = 1
      "000001" when "0011010011001011", -- t[13515] = 1
      "000001" when "0011010011001100", -- t[13516] = 1
      "000001" when "0011010011001101", -- t[13517] = 1
      "000001" when "0011010011001110", -- t[13518] = 1
      "000001" when "0011010011001111", -- t[13519] = 1
      "000001" when "0011010011010000", -- t[13520] = 1
      "000001" when "0011010011010001", -- t[13521] = 1
      "000001" when "0011010011010010", -- t[13522] = 1
      "000001" when "0011010011010011", -- t[13523] = 1
      "000001" when "0011010011010100", -- t[13524] = 1
      "000001" when "0011010011010101", -- t[13525] = 1
      "000001" when "0011010011010110", -- t[13526] = 1
      "000001" when "0011010011010111", -- t[13527] = 1
      "000001" when "0011010011011000", -- t[13528] = 1
      "000001" when "0011010011011001", -- t[13529] = 1
      "000001" when "0011010011011010", -- t[13530] = 1
      "000001" when "0011010011011011", -- t[13531] = 1
      "000001" when "0011010011011100", -- t[13532] = 1
      "000001" when "0011010011011101", -- t[13533] = 1
      "000001" when "0011010011011110", -- t[13534] = 1
      "000001" when "0011010011011111", -- t[13535] = 1
      "000001" when "0011010011100000", -- t[13536] = 1
      "000001" when "0011010011100001", -- t[13537] = 1
      "000001" when "0011010011100010", -- t[13538] = 1
      "000001" when "0011010011100011", -- t[13539] = 1
      "000001" when "0011010011100100", -- t[13540] = 1
      "000001" when "0011010011100101", -- t[13541] = 1
      "000001" when "0011010011100110", -- t[13542] = 1
      "000001" when "0011010011100111", -- t[13543] = 1
      "000001" when "0011010011101000", -- t[13544] = 1
      "000001" when "0011010011101001", -- t[13545] = 1
      "000001" when "0011010011101010", -- t[13546] = 1
      "000001" when "0011010011101011", -- t[13547] = 1
      "000001" when "0011010011101100", -- t[13548] = 1
      "000001" when "0011010011101101", -- t[13549] = 1
      "000001" when "0011010011101110", -- t[13550] = 1
      "000001" when "0011010011101111", -- t[13551] = 1
      "000001" when "0011010011110000", -- t[13552] = 1
      "000001" when "0011010011110001", -- t[13553] = 1
      "000001" when "0011010011110010", -- t[13554] = 1
      "000001" when "0011010011110011", -- t[13555] = 1
      "000001" when "0011010011110100", -- t[13556] = 1
      "000001" when "0011010011110101", -- t[13557] = 1
      "000001" when "0011010011110110", -- t[13558] = 1
      "000001" when "0011010011110111", -- t[13559] = 1
      "000001" when "0011010011111000", -- t[13560] = 1
      "000001" when "0011010011111001", -- t[13561] = 1
      "000001" when "0011010011111010", -- t[13562] = 1
      "000001" when "0011010011111011", -- t[13563] = 1
      "000001" when "0011010011111100", -- t[13564] = 1
      "000001" when "0011010011111101", -- t[13565] = 1
      "000001" when "0011010011111110", -- t[13566] = 1
      "000001" when "0011010011111111", -- t[13567] = 1
      "000001" when "0011010100000000", -- t[13568] = 1
      "000001" when "0011010100000001", -- t[13569] = 1
      "000001" when "0011010100000010", -- t[13570] = 1
      "000001" when "0011010100000011", -- t[13571] = 1
      "000001" when "0011010100000100", -- t[13572] = 1
      "000001" when "0011010100000101", -- t[13573] = 1
      "000001" when "0011010100000110", -- t[13574] = 1
      "000001" when "0011010100000111", -- t[13575] = 1
      "000001" when "0011010100001000", -- t[13576] = 1
      "000001" when "0011010100001001", -- t[13577] = 1
      "000001" when "0011010100001010", -- t[13578] = 1
      "000001" when "0011010100001011", -- t[13579] = 1
      "000001" when "0011010100001100", -- t[13580] = 1
      "000001" when "0011010100001101", -- t[13581] = 1
      "000001" when "0011010100001110", -- t[13582] = 1
      "000001" when "0011010100001111", -- t[13583] = 1
      "000001" when "0011010100010000", -- t[13584] = 1
      "000001" when "0011010100010001", -- t[13585] = 1
      "000001" when "0011010100010010", -- t[13586] = 1
      "000001" when "0011010100010011", -- t[13587] = 1
      "000001" when "0011010100010100", -- t[13588] = 1
      "000001" when "0011010100010101", -- t[13589] = 1
      "000001" when "0011010100010110", -- t[13590] = 1
      "000001" when "0011010100010111", -- t[13591] = 1
      "000001" when "0011010100011000", -- t[13592] = 1
      "000001" when "0011010100011001", -- t[13593] = 1
      "000001" when "0011010100011010", -- t[13594] = 1
      "000001" when "0011010100011011", -- t[13595] = 1
      "000001" when "0011010100011100", -- t[13596] = 1
      "000001" when "0011010100011101", -- t[13597] = 1
      "000001" when "0011010100011110", -- t[13598] = 1
      "000001" when "0011010100011111", -- t[13599] = 1
      "000001" when "0011010100100000", -- t[13600] = 1
      "000001" when "0011010100100001", -- t[13601] = 1
      "000001" when "0011010100100010", -- t[13602] = 1
      "000001" when "0011010100100011", -- t[13603] = 1
      "000001" when "0011010100100100", -- t[13604] = 1
      "000001" when "0011010100100101", -- t[13605] = 1
      "000001" when "0011010100100110", -- t[13606] = 1
      "000001" when "0011010100100111", -- t[13607] = 1
      "000001" when "0011010100101000", -- t[13608] = 1
      "000001" when "0011010100101001", -- t[13609] = 1
      "000001" when "0011010100101010", -- t[13610] = 1
      "000001" when "0011010100101011", -- t[13611] = 1
      "000001" when "0011010100101100", -- t[13612] = 1
      "000001" when "0011010100101101", -- t[13613] = 1
      "000001" when "0011010100101110", -- t[13614] = 1
      "000001" when "0011010100101111", -- t[13615] = 1
      "000001" when "0011010100110000", -- t[13616] = 1
      "000001" when "0011010100110001", -- t[13617] = 1
      "000001" when "0011010100110010", -- t[13618] = 1
      "000001" when "0011010100110011", -- t[13619] = 1
      "000001" when "0011010100110100", -- t[13620] = 1
      "000001" when "0011010100110101", -- t[13621] = 1
      "000001" when "0011010100110110", -- t[13622] = 1
      "000001" when "0011010100110111", -- t[13623] = 1
      "000001" when "0011010100111000", -- t[13624] = 1
      "000001" when "0011010100111001", -- t[13625] = 1
      "000001" when "0011010100111010", -- t[13626] = 1
      "000001" when "0011010100111011", -- t[13627] = 1
      "000001" when "0011010100111100", -- t[13628] = 1
      "000001" when "0011010100111101", -- t[13629] = 1
      "000001" when "0011010100111110", -- t[13630] = 1
      "000001" when "0011010100111111", -- t[13631] = 1
      "000001" when "0011010101000000", -- t[13632] = 1
      "000001" when "0011010101000001", -- t[13633] = 1
      "000001" when "0011010101000010", -- t[13634] = 1
      "000001" when "0011010101000011", -- t[13635] = 1
      "000001" when "0011010101000100", -- t[13636] = 1
      "000001" when "0011010101000101", -- t[13637] = 1
      "000001" when "0011010101000110", -- t[13638] = 1
      "000001" when "0011010101000111", -- t[13639] = 1
      "000001" when "0011010101001000", -- t[13640] = 1
      "000001" when "0011010101001001", -- t[13641] = 1
      "000001" when "0011010101001010", -- t[13642] = 1
      "000001" when "0011010101001011", -- t[13643] = 1
      "000001" when "0011010101001100", -- t[13644] = 1
      "000001" when "0011010101001101", -- t[13645] = 1
      "000001" when "0011010101001110", -- t[13646] = 1
      "000001" when "0011010101001111", -- t[13647] = 1
      "000001" when "0011010101010000", -- t[13648] = 1
      "000001" when "0011010101010001", -- t[13649] = 1
      "000001" when "0011010101010010", -- t[13650] = 1
      "000001" when "0011010101010011", -- t[13651] = 1
      "000001" when "0011010101010100", -- t[13652] = 1
      "000001" when "0011010101010101", -- t[13653] = 1
      "000001" when "0011010101010110", -- t[13654] = 1
      "000001" when "0011010101010111", -- t[13655] = 1
      "000001" when "0011010101011000", -- t[13656] = 1
      "000001" when "0011010101011001", -- t[13657] = 1
      "000001" when "0011010101011010", -- t[13658] = 1
      "000001" when "0011010101011011", -- t[13659] = 1
      "000001" when "0011010101011100", -- t[13660] = 1
      "000001" when "0011010101011101", -- t[13661] = 1
      "000001" when "0011010101011110", -- t[13662] = 1
      "000001" when "0011010101011111", -- t[13663] = 1
      "000001" when "0011010101100000", -- t[13664] = 1
      "000001" when "0011010101100001", -- t[13665] = 1
      "000001" when "0011010101100010", -- t[13666] = 1
      "000001" when "0011010101100011", -- t[13667] = 1
      "000001" when "0011010101100100", -- t[13668] = 1
      "000001" when "0011010101100101", -- t[13669] = 1
      "000001" when "0011010101100110", -- t[13670] = 1
      "000001" when "0011010101100111", -- t[13671] = 1
      "000001" when "0011010101101000", -- t[13672] = 1
      "000001" when "0011010101101001", -- t[13673] = 1
      "000001" when "0011010101101010", -- t[13674] = 1
      "000001" when "0011010101101011", -- t[13675] = 1
      "000001" when "0011010101101100", -- t[13676] = 1
      "000001" when "0011010101101101", -- t[13677] = 1
      "000001" when "0011010101101110", -- t[13678] = 1
      "000001" when "0011010101101111", -- t[13679] = 1
      "000001" when "0011010101110000", -- t[13680] = 1
      "000001" when "0011010101110001", -- t[13681] = 1
      "000001" when "0011010101110010", -- t[13682] = 1
      "000001" when "0011010101110011", -- t[13683] = 1
      "000001" when "0011010101110100", -- t[13684] = 1
      "000001" when "0011010101110101", -- t[13685] = 1
      "000001" when "0011010101110110", -- t[13686] = 1
      "000001" when "0011010101110111", -- t[13687] = 1
      "000001" when "0011010101111000", -- t[13688] = 1
      "000001" when "0011010101111001", -- t[13689] = 1
      "000001" when "0011010101111010", -- t[13690] = 1
      "000001" when "0011010101111011", -- t[13691] = 1
      "000001" when "0011010101111100", -- t[13692] = 1
      "000001" when "0011010101111101", -- t[13693] = 1
      "000001" when "0011010101111110", -- t[13694] = 1
      "000001" when "0011010101111111", -- t[13695] = 1
      "000001" when "0011010110000000", -- t[13696] = 1
      "000001" when "0011010110000001", -- t[13697] = 1
      "000001" when "0011010110000010", -- t[13698] = 1
      "000001" when "0011010110000011", -- t[13699] = 1
      "000001" when "0011010110000100", -- t[13700] = 1
      "000001" when "0011010110000101", -- t[13701] = 1
      "000001" when "0011010110000110", -- t[13702] = 1
      "000001" when "0011010110000111", -- t[13703] = 1
      "000001" when "0011010110001000", -- t[13704] = 1
      "000001" when "0011010110001001", -- t[13705] = 1
      "000001" when "0011010110001010", -- t[13706] = 1
      "000001" when "0011010110001011", -- t[13707] = 1
      "000001" when "0011010110001100", -- t[13708] = 1
      "000001" when "0011010110001101", -- t[13709] = 1
      "000001" when "0011010110001110", -- t[13710] = 1
      "000001" when "0011010110001111", -- t[13711] = 1
      "000001" when "0011010110010000", -- t[13712] = 1
      "000001" when "0011010110010001", -- t[13713] = 1
      "000001" when "0011010110010010", -- t[13714] = 1
      "000001" when "0011010110010011", -- t[13715] = 1
      "000001" when "0011010110010100", -- t[13716] = 1
      "000001" when "0011010110010101", -- t[13717] = 1
      "000001" when "0011010110010110", -- t[13718] = 1
      "000001" when "0011010110010111", -- t[13719] = 1
      "000001" when "0011010110011000", -- t[13720] = 1
      "000001" when "0011010110011001", -- t[13721] = 1
      "000001" when "0011010110011010", -- t[13722] = 1
      "000001" when "0011010110011011", -- t[13723] = 1
      "000001" when "0011010110011100", -- t[13724] = 1
      "000001" when "0011010110011101", -- t[13725] = 1
      "000001" when "0011010110011110", -- t[13726] = 1
      "000001" when "0011010110011111", -- t[13727] = 1
      "000001" when "0011010110100000", -- t[13728] = 1
      "000001" when "0011010110100001", -- t[13729] = 1
      "000001" when "0011010110100010", -- t[13730] = 1
      "000001" when "0011010110100011", -- t[13731] = 1
      "000001" when "0011010110100100", -- t[13732] = 1
      "000001" when "0011010110100101", -- t[13733] = 1
      "000001" when "0011010110100110", -- t[13734] = 1
      "000001" when "0011010110100111", -- t[13735] = 1
      "000001" when "0011010110101000", -- t[13736] = 1
      "000001" when "0011010110101001", -- t[13737] = 1
      "000001" when "0011010110101010", -- t[13738] = 1
      "000001" when "0011010110101011", -- t[13739] = 1
      "000001" when "0011010110101100", -- t[13740] = 1
      "000001" when "0011010110101101", -- t[13741] = 1
      "000001" when "0011010110101110", -- t[13742] = 1
      "000001" when "0011010110101111", -- t[13743] = 1
      "000001" when "0011010110110000", -- t[13744] = 1
      "000001" when "0011010110110001", -- t[13745] = 1
      "000001" when "0011010110110010", -- t[13746] = 1
      "000001" when "0011010110110011", -- t[13747] = 1
      "000001" when "0011010110110100", -- t[13748] = 1
      "000001" when "0011010110110101", -- t[13749] = 1
      "000001" when "0011010110110110", -- t[13750] = 1
      "000001" when "0011010110110111", -- t[13751] = 1
      "000001" when "0011010110111000", -- t[13752] = 1
      "000001" when "0011010110111001", -- t[13753] = 1
      "000001" when "0011010110111010", -- t[13754] = 1
      "000001" when "0011010110111011", -- t[13755] = 1
      "000001" when "0011010110111100", -- t[13756] = 1
      "000001" when "0011010110111101", -- t[13757] = 1
      "000001" when "0011010110111110", -- t[13758] = 1
      "000001" when "0011010110111111", -- t[13759] = 1
      "000001" when "0011010111000000", -- t[13760] = 1
      "000001" when "0011010111000001", -- t[13761] = 1
      "000001" when "0011010111000010", -- t[13762] = 1
      "000001" when "0011010111000011", -- t[13763] = 1
      "000001" when "0011010111000100", -- t[13764] = 1
      "000001" when "0011010111000101", -- t[13765] = 1
      "000001" when "0011010111000110", -- t[13766] = 1
      "000001" when "0011010111000111", -- t[13767] = 1
      "000001" when "0011010111001000", -- t[13768] = 1
      "000001" when "0011010111001001", -- t[13769] = 1
      "000001" when "0011010111001010", -- t[13770] = 1
      "000001" when "0011010111001011", -- t[13771] = 1
      "000001" when "0011010111001100", -- t[13772] = 1
      "000001" when "0011010111001101", -- t[13773] = 1
      "000001" when "0011010111001110", -- t[13774] = 1
      "000001" when "0011010111001111", -- t[13775] = 1
      "000001" when "0011010111010000", -- t[13776] = 1
      "000001" when "0011010111010001", -- t[13777] = 1
      "000001" when "0011010111010010", -- t[13778] = 1
      "000001" when "0011010111010011", -- t[13779] = 1
      "000001" when "0011010111010100", -- t[13780] = 1
      "000001" when "0011010111010101", -- t[13781] = 1
      "000001" when "0011010111010110", -- t[13782] = 1
      "000001" when "0011010111010111", -- t[13783] = 1
      "000001" when "0011010111011000", -- t[13784] = 1
      "000001" when "0011010111011001", -- t[13785] = 1
      "000001" when "0011010111011010", -- t[13786] = 1
      "000001" when "0011010111011011", -- t[13787] = 1
      "000001" when "0011010111011100", -- t[13788] = 1
      "000001" when "0011010111011101", -- t[13789] = 1
      "000001" when "0011010111011110", -- t[13790] = 1
      "000001" when "0011010111011111", -- t[13791] = 1
      "000001" when "0011010111100000", -- t[13792] = 1
      "000001" when "0011010111100001", -- t[13793] = 1
      "000001" when "0011010111100010", -- t[13794] = 1
      "000001" when "0011010111100011", -- t[13795] = 1
      "000001" when "0011010111100100", -- t[13796] = 1
      "000001" when "0011010111100101", -- t[13797] = 1
      "000001" when "0011010111100110", -- t[13798] = 1
      "000001" when "0011010111100111", -- t[13799] = 1
      "000001" when "0011010111101000", -- t[13800] = 1
      "000001" when "0011010111101001", -- t[13801] = 1
      "000001" when "0011010111101010", -- t[13802] = 1
      "000001" when "0011010111101011", -- t[13803] = 1
      "000001" when "0011010111101100", -- t[13804] = 1
      "000001" when "0011010111101101", -- t[13805] = 1
      "000001" when "0011010111101110", -- t[13806] = 1
      "000001" when "0011010111101111", -- t[13807] = 1
      "000001" when "0011010111110000", -- t[13808] = 1
      "000001" when "0011010111110001", -- t[13809] = 1
      "000001" when "0011010111110010", -- t[13810] = 1
      "000001" when "0011010111110011", -- t[13811] = 1
      "000001" when "0011010111110100", -- t[13812] = 1
      "000001" when "0011010111110101", -- t[13813] = 1
      "000001" when "0011010111110110", -- t[13814] = 1
      "000001" when "0011010111110111", -- t[13815] = 1
      "000001" when "0011010111111000", -- t[13816] = 1
      "000001" when "0011010111111001", -- t[13817] = 1
      "000001" when "0011010111111010", -- t[13818] = 1
      "000001" when "0011010111111011", -- t[13819] = 1
      "000001" when "0011010111111100", -- t[13820] = 1
      "000001" when "0011010111111101", -- t[13821] = 1
      "000001" when "0011010111111110", -- t[13822] = 1
      "000001" when "0011010111111111", -- t[13823] = 1
      "000001" when "0011011000000000", -- t[13824] = 1
      "000001" when "0011011000000001", -- t[13825] = 1
      "000001" when "0011011000000010", -- t[13826] = 1
      "000001" when "0011011000000011", -- t[13827] = 1
      "000001" when "0011011000000100", -- t[13828] = 1
      "000001" when "0011011000000101", -- t[13829] = 1
      "000001" when "0011011000000110", -- t[13830] = 1
      "000001" when "0011011000000111", -- t[13831] = 1
      "000001" when "0011011000001000", -- t[13832] = 1
      "000001" when "0011011000001001", -- t[13833] = 1
      "000001" when "0011011000001010", -- t[13834] = 1
      "000001" when "0011011000001011", -- t[13835] = 1
      "000001" when "0011011000001100", -- t[13836] = 1
      "000001" when "0011011000001101", -- t[13837] = 1
      "000001" when "0011011000001110", -- t[13838] = 1
      "000001" when "0011011000001111", -- t[13839] = 1
      "000001" when "0011011000010000", -- t[13840] = 1
      "000001" when "0011011000010001", -- t[13841] = 1
      "000001" when "0011011000010010", -- t[13842] = 1
      "000001" when "0011011000010011", -- t[13843] = 1
      "000001" when "0011011000010100", -- t[13844] = 1
      "000001" when "0011011000010101", -- t[13845] = 1
      "000001" when "0011011000010110", -- t[13846] = 1
      "000001" when "0011011000010111", -- t[13847] = 1
      "000001" when "0011011000011000", -- t[13848] = 1
      "000001" when "0011011000011001", -- t[13849] = 1
      "000001" when "0011011000011010", -- t[13850] = 1
      "000001" when "0011011000011011", -- t[13851] = 1
      "000001" when "0011011000011100", -- t[13852] = 1
      "000001" when "0011011000011101", -- t[13853] = 1
      "000001" when "0011011000011110", -- t[13854] = 1
      "000001" when "0011011000011111", -- t[13855] = 1
      "000001" when "0011011000100000", -- t[13856] = 1
      "000001" when "0011011000100001", -- t[13857] = 1
      "000001" when "0011011000100010", -- t[13858] = 1
      "000001" when "0011011000100011", -- t[13859] = 1
      "000001" when "0011011000100100", -- t[13860] = 1
      "000001" when "0011011000100101", -- t[13861] = 1
      "000001" when "0011011000100110", -- t[13862] = 1
      "000001" when "0011011000100111", -- t[13863] = 1
      "000001" when "0011011000101000", -- t[13864] = 1
      "000001" when "0011011000101001", -- t[13865] = 1
      "000001" when "0011011000101010", -- t[13866] = 1
      "000001" when "0011011000101011", -- t[13867] = 1
      "000001" when "0011011000101100", -- t[13868] = 1
      "000001" when "0011011000101101", -- t[13869] = 1
      "000001" when "0011011000101110", -- t[13870] = 1
      "000001" when "0011011000101111", -- t[13871] = 1
      "000001" when "0011011000110000", -- t[13872] = 1
      "000001" when "0011011000110001", -- t[13873] = 1
      "000001" when "0011011000110010", -- t[13874] = 1
      "000001" when "0011011000110011", -- t[13875] = 1
      "000001" when "0011011000110100", -- t[13876] = 1
      "000001" when "0011011000110101", -- t[13877] = 1
      "000001" when "0011011000110110", -- t[13878] = 1
      "000001" when "0011011000110111", -- t[13879] = 1
      "000001" when "0011011000111000", -- t[13880] = 1
      "000001" when "0011011000111001", -- t[13881] = 1
      "000001" when "0011011000111010", -- t[13882] = 1
      "000001" when "0011011000111011", -- t[13883] = 1
      "000001" when "0011011000111100", -- t[13884] = 1
      "000001" when "0011011000111101", -- t[13885] = 1
      "000001" when "0011011000111110", -- t[13886] = 1
      "000001" when "0011011000111111", -- t[13887] = 1
      "000001" when "0011011001000000", -- t[13888] = 1
      "000001" when "0011011001000001", -- t[13889] = 1
      "000001" when "0011011001000010", -- t[13890] = 1
      "000001" when "0011011001000011", -- t[13891] = 1
      "000001" when "0011011001000100", -- t[13892] = 1
      "000001" when "0011011001000101", -- t[13893] = 1
      "000001" when "0011011001000110", -- t[13894] = 1
      "000001" when "0011011001000111", -- t[13895] = 1
      "000001" when "0011011001001000", -- t[13896] = 1
      "000001" when "0011011001001001", -- t[13897] = 1
      "000001" when "0011011001001010", -- t[13898] = 1
      "000001" when "0011011001001011", -- t[13899] = 1
      "000001" when "0011011001001100", -- t[13900] = 1
      "000001" when "0011011001001101", -- t[13901] = 1
      "000001" when "0011011001001110", -- t[13902] = 1
      "000001" when "0011011001001111", -- t[13903] = 1
      "000001" when "0011011001010000", -- t[13904] = 1
      "000001" when "0011011001010001", -- t[13905] = 1
      "000001" when "0011011001010010", -- t[13906] = 1
      "000001" when "0011011001010011", -- t[13907] = 1
      "000001" when "0011011001010100", -- t[13908] = 1
      "000001" when "0011011001010101", -- t[13909] = 1
      "000001" when "0011011001010110", -- t[13910] = 1
      "000001" when "0011011001010111", -- t[13911] = 1
      "000001" when "0011011001011000", -- t[13912] = 1
      "000001" when "0011011001011001", -- t[13913] = 1
      "000001" when "0011011001011010", -- t[13914] = 1
      "000001" when "0011011001011011", -- t[13915] = 1
      "000001" when "0011011001011100", -- t[13916] = 1
      "000001" when "0011011001011101", -- t[13917] = 1
      "000001" when "0011011001011110", -- t[13918] = 1
      "000001" when "0011011001011111", -- t[13919] = 1
      "000001" when "0011011001100000", -- t[13920] = 1
      "000001" when "0011011001100001", -- t[13921] = 1
      "000001" when "0011011001100010", -- t[13922] = 1
      "000001" when "0011011001100011", -- t[13923] = 1
      "000001" when "0011011001100100", -- t[13924] = 1
      "000001" when "0011011001100101", -- t[13925] = 1
      "000001" when "0011011001100110", -- t[13926] = 1
      "000001" when "0011011001100111", -- t[13927] = 1
      "000001" when "0011011001101000", -- t[13928] = 1
      "000001" when "0011011001101001", -- t[13929] = 1
      "000001" when "0011011001101010", -- t[13930] = 1
      "000001" when "0011011001101011", -- t[13931] = 1
      "000001" when "0011011001101100", -- t[13932] = 1
      "000001" when "0011011001101101", -- t[13933] = 1
      "000001" when "0011011001101110", -- t[13934] = 1
      "000001" when "0011011001101111", -- t[13935] = 1
      "000001" when "0011011001110000", -- t[13936] = 1
      "000001" when "0011011001110001", -- t[13937] = 1
      "000001" when "0011011001110010", -- t[13938] = 1
      "000001" when "0011011001110011", -- t[13939] = 1
      "000001" when "0011011001110100", -- t[13940] = 1
      "000001" when "0011011001110101", -- t[13941] = 1
      "000001" when "0011011001110110", -- t[13942] = 1
      "000001" when "0011011001110111", -- t[13943] = 1
      "000001" when "0011011001111000", -- t[13944] = 1
      "000001" when "0011011001111001", -- t[13945] = 1
      "000001" when "0011011001111010", -- t[13946] = 1
      "000001" when "0011011001111011", -- t[13947] = 1
      "000001" when "0011011001111100", -- t[13948] = 1
      "000001" when "0011011001111101", -- t[13949] = 1
      "000001" when "0011011001111110", -- t[13950] = 1
      "000001" when "0011011001111111", -- t[13951] = 1
      "000001" when "0011011010000000", -- t[13952] = 1
      "000001" when "0011011010000001", -- t[13953] = 1
      "000001" when "0011011010000010", -- t[13954] = 1
      "000001" when "0011011010000011", -- t[13955] = 1
      "000001" when "0011011010000100", -- t[13956] = 1
      "000001" when "0011011010000101", -- t[13957] = 1
      "000001" when "0011011010000110", -- t[13958] = 1
      "000001" when "0011011010000111", -- t[13959] = 1
      "000001" when "0011011010001000", -- t[13960] = 1
      "000001" when "0011011010001001", -- t[13961] = 1
      "000001" when "0011011010001010", -- t[13962] = 1
      "000001" when "0011011010001011", -- t[13963] = 1
      "000001" when "0011011010001100", -- t[13964] = 1
      "000001" when "0011011010001101", -- t[13965] = 1
      "000001" when "0011011010001110", -- t[13966] = 1
      "000001" when "0011011010001111", -- t[13967] = 1
      "000001" when "0011011010010000", -- t[13968] = 1
      "000001" when "0011011010010001", -- t[13969] = 1
      "000001" when "0011011010010010", -- t[13970] = 1
      "000001" when "0011011010010011", -- t[13971] = 1
      "000001" when "0011011010010100", -- t[13972] = 1
      "000001" when "0011011010010101", -- t[13973] = 1
      "000001" when "0011011010010110", -- t[13974] = 1
      "000001" when "0011011010010111", -- t[13975] = 1
      "000001" when "0011011010011000", -- t[13976] = 1
      "000001" when "0011011010011001", -- t[13977] = 1
      "000001" when "0011011010011010", -- t[13978] = 1
      "000001" when "0011011010011011", -- t[13979] = 1
      "000001" when "0011011010011100", -- t[13980] = 1
      "000001" when "0011011010011101", -- t[13981] = 1
      "000001" when "0011011010011110", -- t[13982] = 1
      "000001" when "0011011010011111", -- t[13983] = 1
      "000001" when "0011011010100000", -- t[13984] = 1
      "000001" when "0011011010100001", -- t[13985] = 1
      "000001" when "0011011010100010", -- t[13986] = 1
      "000001" when "0011011010100011", -- t[13987] = 1
      "000001" when "0011011010100100", -- t[13988] = 1
      "000001" when "0011011010100101", -- t[13989] = 1
      "000001" when "0011011010100110", -- t[13990] = 1
      "000001" when "0011011010100111", -- t[13991] = 1
      "000001" when "0011011010101000", -- t[13992] = 1
      "000001" when "0011011010101001", -- t[13993] = 1
      "000001" when "0011011010101010", -- t[13994] = 1
      "000001" when "0011011010101011", -- t[13995] = 1
      "000001" when "0011011010101100", -- t[13996] = 1
      "000001" when "0011011010101101", -- t[13997] = 1
      "000001" when "0011011010101110", -- t[13998] = 1
      "000001" when "0011011010101111", -- t[13999] = 1
      "000001" when "0011011010110000", -- t[14000] = 1
      "000001" when "0011011010110001", -- t[14001] = 1
      "000001" when "0011011010110010", -- t[14002] = 1
      "000001" when "0011011010110011", -- t[14003] = 1
      "000001" when "0011011010110100", -- t[14004] = 1
      "000001" when "0011011010110101", -- t[14005] = 1
      "000001" when "0011011010110110", -- t[14006] = 1
      "000001" when "0011011010110111", -- t[14007] = 1
      "000001" when "0011011010111000", -- t[14008] = 1
      "000001" when "0011011010111001", -- t[14009] = 1
      "000001" when "0011011010111010", -- t[14010] = 1
      "000001" when "0011011010111011", -- t[14011] = 1
      "000001" when "0011011010111100", -- t[14012] = 1
      "000001" when "0011011010111101", -- t[14013] = 1
      "000001" when "0011011010111110", -- t[14014] = 1
      "000001" when "0011011010111111", -- t[14015] = 1
      "000001" when "0011011011000000", -- t[14016] = 1
      "000001" when "0011011011000001", -- t[14017] = 1
      "000001" when "0011011011000010", -- t[14018] = 1
      "000001" when "0011011011000011", -- t[14019] = 1
      "000001" when "0011011011000100", -- t[14020] = 1
      "000001" when "0011011011000101", -- t[14021] = 1
      "000001" when "0011011011000110", -- t[14022] = 1
      "000001" when "0011011011000111", -- t[14023] = 1
      "000001" when "0011011011001000", -- t[14024] = 1
      "000001" when "0011011011001001", -- t[14025] = 1
      "000001" when "0011011011001010", -- t[14026] = 1
      "000001" when "0011011011001011", -- t[14027] = 1
      "000001" when "0011011011001100", -- t[14028] = 1
      "000001" when "0011011011001101", -- t[14029] = 1
      "000001" when "0011011011001110", -- t[14030] = 1
      "000001" when "0011011011001111", -- t[14031] = 1
      "000001" when "0011011011010000", -- t[14032] = 1
      "000001" when "0011011011010001", -- t[14033] = 1
      "000001" when "0011011011010010", -- t[14034] = 1
      "000001" when "0011011011010011", -- t[14035] = 1
      "000001" when "0011011011010100", -- t[14036] = 1
      "000001" when "0011011011010101", -- t[14037] = 1
      "000001" when "0011011011010110", -- t[14038] = 1
      "000001" when "0011011011010111", -- t[14039] = 1
      "000001" when "0011011011011000", -- t[14040] = 1
      "000001" when "0011011011011001", -- t[14041] = 1
      "000001" when "0011011011011010", -- t[14042] = 1
      "000001" when "0011011011011011", -- t[14043] = 1
      "000001" when "0011011011011100", -- t[14044] = 1
      "000001" when "0011011011011101", -- t[14045] = 1
      "000001" when "0011011011011110", -- t[14046] = 1
      "000001" when "0011011011011111", -- t[14047] = 1
      "000001" when "0011011011100000", -- t[14048] = 1
      "000001" when "0011011011100001", -- t[14049] = 1
      "000001" when "0011011011100010", -- t[14050] = 1
      "000001" when "0011011011100011", -- t[14051] = 1
      "000001" when "0011011011100100", -- t[14052] = 1
      "000001" when "0011011011100101", -- t[14053] = 1
      "000001" when "0011011011100110", -- t[14054] = 1
      "000001" when "0011011011100111", -- t[14055] = 1
      "000001" when "0011011011101000", -- t[14056] = 1
      "000001" when "0011011011101001", -- t[14057] = 1
      "000001" when "0011011011101010", -- t[14058] = 1
      "000001" when "0011011011101011", -- t[14059] = 1
      "000001" when "0011011011101100", -- t[14060] = 1
      "000001" when "0011011011101101", -- t[14061] = 1
      "000001" when "0011011011101110", -- t[14062] = 1
      "000001" when "0011011011101111", -- t[14063] = 1
      "000001" when "0011011011110000", -- t[14064] = 1
      "000001" when "0011011011110001", -- t[14065] = 1
      "000001" when "0011011011110010", -- t[14066] = 1
      "000001" when "0011011011110011", -- t[14067] = 1
      "000001" when "0011011011110100", -- t[14068] = 1
      "000001" when "0011011011110101", -- t[14069] = 1
      "000001" when "0011011011110110", -- t[14070] = 1
      "000001" when "0011011011110111", -- t[14071] = 1
      "000001" when "0011011011111000", -- t[14072] = 1
      "000001" when "0011011011111001", -- t[14073] = 1
      "000001" when "0011011011111010", -- t[14074] = 1
      "000001" when "0011011011111011", -- t[14075] = 1
      "000001" when "0011011011111100", -- t[14076] = 1
      "000001" when "0011011011111101", -- t[14077] = 1
      "000001" when "0011011011111110", -- t[14078] = 1
      "000001" when "0011011011111111", -- t[14079] = 1
      "000001" when "0011011100000000", -- t[14080] = 1
      "000001" when "0011011100000001", -- t[14081] = 1
      "000001" when "0011011100000010", -- t[14082] = 1
      "000001" when "0011011100000011", -- t[14083] = 1
      "000001" when "0011011100000100", -- t[14084] = 1
      "000001" when "0011011100000101", -- t[14085] = 1
      "000001" when "0011011100000110", -- t[14086] = 1
      "000001" when "0011011100000111", -- t[14087] = 1
      "000001" when "0011011100001000", -- t[14088] = 1
      "000001" when "0011011100001001", -- t[14089] = 1
      "000001" when "0011011100001010", -- t[14090] = 1
      "000001" when "0011011100001011", -- t[14091] = 1
      "000001" when "0011011100001100", -- t[14092] = 1
      "000001" when "0011011100001101", -- t[14093] = 1
      "000001" when "0011011100001110", -- t[14094] = 1
      "000001" when "0011011100001111", -- t[14095] = 1
      "000001" when "0011011100010000", -- t[14096] = 1
      "000001" when "0011011100010001", -- t[14097] = 1
      "000001" when "0011011100010010", -- t[14098] = 1
      "000001" when "0011011100010011", -- t[14099] = 1
      "000001" when "0011011100010100", -- t[14100] = 1
      "000001" when "0011011100010101", -- t[14101] = 1
      "000001" when "0011011100010110", -- t[14102] = 1
      "000001" when "0011011100010111", -- t[14103] = 1
      "000001" when "0011011100011000", -- t[14104] = 1
      "000001" when "0011011100011001", -- t[14105] = 1
      "000001" when "0011011100011010", -- t[14106] = 1
      "000001" when "0011011100011011", -- t[14107] = 1
      "000001" when "0011011100011100", -- t[14108] = 1
      "000001" when "0011011100011101", -- t[14109] = 1
      "000001" when "0011011100011110", -- t[14110] = 1
      "000001" when "0011011100011111", -- t[14111] = 1
      "000001" when "0011011100100000", -- t[14112] = 1
      "000001" when "0011011100100001", -- t[14113] = 1
      "000001" when "0011011100100010", -- t[14114] = 1
      "000001" when "0011011100100011", -- t[14115] = 1
      "000001" when "0011011100100100", -- t[14116] = 1
      "000001" when "0011011100100101", -- t[14117] = 1
      "000001" when "0011011100100110", -- t[14118] = 1
      "000001" when "0011011100100111", -- t[14119] = 1
      "000001" when "0011011100101000", -- t[14120] = 1
      "000001" when "0011011100101001", -- t[14121] = 1
      "000001" when "0011011100101010", -- t[14122] = 1
      "000001" when "0011011100101011", -- t[14123] = 1
      "000001" when "0011011100101100", -- t[14124] = 1
      "000001" when "0011011100101101", -- t[14125] = 1
      "000001" when "0011011100101110", -- t[14126] = 1
      "000001" when "0011011100101111", -- t[14127] = 1
      "000001" when "0011011100110000", -- t[14128] = 1
      "000001" when "0011011100110001", -- t[14129] = 1
      "000001" when "0011011100110010", -- t[14130] = 1
      "000001" when "0011011100110011", -- t[14131] = 1
      "000001" when "0011011100110100", -- t[14132] = 1
      "000001" when "0011011100110101", -- t[14133] = 1
      "000001" when "0011011100110110", -- t[14134] = 1
      "000001" when "0011011100110111", -- t[14135] = 1
      "000001" when "0011011100111000", -- t[14136] = 1
      "000001" when "0011011100111001", -- t[14137] = 1
      "000001" when "0011011100111010", -- t[14138] = 1
      "000001" when "0011011100111011", -- t[14139] = 1
      "000001" when "0011011100111100", -- t[14140] = 1
      "000001" when "0011011100111101", -- t[14141] = 1
      "000001" when "0011011100111110", -- t[14142] = 1
      "000001" when "0011011100111111", -- t[14143] = 1
      "000001" when "0011011101000000", -- t[14144] = 1
      "000001" when "0011011101000001", -- t[14145] = 1
      "000001" when "0011011101000010", -- t[14146] = 1
      "000001" when "0011011101000011", -- t[14147] = 1
      "000001" when "0011011101000100", -- t[14148] = 1
      "000001" when "0011011101000101", -- t[14149] = 1
      "000001" when "0011011101000110", -- t[14150] = 1
      "000001" when "0011011101000111", -- t[14151] = 1
      "000001" when "0011011101001000", -- t[14152] = 1
      "000001" when "0011011101001001", -- t[14153] = 1
      "000001" when "0011011101001010", -- t[14154] = 1
      "000001" when "0011011101001011", -- t[14155] = 1
      "000001" when "0011011101001100", -- t[14156] = 1
      "000001" when "0011011101001101", -- t[14157] = 1
      "000001" when "0011011101001110", -- t[14158] = 1
      "000001" when "0011011101001111", -- t[14159] = 1
      "000001" when "0011011101010000", -- t[14160] = 1
      "000001" when "0011011101010001", -- t[14161] = 1
      "000001" when "0011011101010010", -- t[14162] = 1
      "000001" when "0011011101010011", -- t[14163] = 1
      "000001" when "0011011101010100", -- t[14164] = 1
      "000001" when "0011011101010101", -- t[14165] = 1
      "000001" when "0011011101010110", -- t[14166] = 1
      "000001" when "0011011101010111", -- t[14167] = 1
      "000001" when "0011011101011000", -- t[14168] = 1
      "000001" when "0011011101011001", -- t[14169] = 1
      "000001" when "0011011101011010", -- t[14170] = 1
      "000001" when "0011011101011011", -- t[14171] = 1
      "000001" when "0011011101011100", -- t[14172] = 1
      "000001" when "0011011101011101", -- t[14173] = 1
      "000001" when "0011011101011110", -- t[14174] = 1
      "000001" when "0011011101011111", -- t[14175] = 1
      "000001" when "0011011101100000", -- t[14176] = 1
      "000001" when "0011011101100001", -- t[14177] = 1
      "000001" when "0011011101100010", -- t[14178] = 1
      "000001" when "0011011101100011", -- t[14179] = 1
      "000001" when "0011011101100100", -- t[14180] = 1
      "000001" when "0011011101100101", -- t[14181] = 1
      "000001" when "0011011101100110", -- t[14182] = 1
      "000001" when "0011011101100111", -- t[14183] = 1
      "000001" when "0011011101101000", -- t[14184] = 1
      "000001" when "0011011101101001", -- t[14185] = 1
      "000001" when "0011011101101010", -- t[14186] = 1
      "000001" when "0011011101101011", -- t[14187] = 1
      "000001" when "0011011101101100", -- t[14188] = 1
      "000001" when "0011011101101101", -- t[14189] = 1
      "000001" when "0011011101101110", -- t[14190] = 1
      "000001" when "0011011101101111", -- t[14191] = 1
      "000001" when "0011011101110000", -- t[14192] = 1
      "000001" when "0011011101110001", -- t[14193] = 1
      "000001" when "0011011101110010", -- t[14194] = 1
      "000001" when "0011011101110011", -- t[14195] = 1
      "000001" when "0011011101110100", -- t[14196] = 1
      "000001" when "0011011101110101", -- t[14197] = 1
      "000001" when "0011011101110110", -- t[14198] = 1
      "000001" when "0011011101110111", -- t[14199] = 1
      "000001" when "0011011101111000", -- t[14200] = 1
      "000001" when "0011011101111001", -- t[14201] = 1
      "000001" when "0011011101111010", -- t[14202] = 1
      "000001" when "0011011101111011", -- t[14203] = 1
      "000001" when "0011011101111100", -- t[14204] = 1
      "000001" when "0011011101111101", -- t[14205] = 1
      "000001" when "0011011101111110", -- t[14206] = 1
      "000001" when "0011011101111111", -- t[14207] = 1
      "000001" when "0011011110000000", -- t[14208] = 1
      "000001" when "0011011110000001", -- t[14209] = 1
      "000001" when "0011011110000010", -- t[14210] = 1
      "000001" when "0011011110000011", -- t[14211] = 1
      "000001" when "0011011110000100", -- t[14212] = 1
      "000001" when "0011011110000101", -- t[14213] = 1
      "000001" when "0011011110000110", -- t[14214] = 1
      "000001" when "0011011110000111", -- t[14215] = 1
      "000001" when "0011011110001000", -- t[14216] = 1
      "000001" when "0011011110001001", -- t[14217] = 1
      "000001" when "0011011110001010", -- t[14218] = 1
      "000001" when "0011011110001011", -- t[14219] = 1
      "000001" when "0011011110001100", -- t[14220] = 1
      "000001" when "0011011110001101", -- t[14221] = 1
      "000001" when "0011011110001110", -- t[14222] = 1
      "000001" when "0011011110001111", -- t[14223] = 1
      "000001" when "0011011110010000", -- t[14224] = 1
      "000001" when "0011011110010001", -- t[14225] = 1
      "000001" when "0011011110010010", -- t[14226] = 1
      "000001" when "0011011110010011", -- t[14227] = 1
      "000001" when "0011011110010100", -- t[14228] = 1
      "000001" when "0011011110010101", -- t[14229] = 1
      "000001" when "0011011110010110", -- t[14230] = 1
      "000001" when "0011011110010111", -- t[14231] = 1
      "000001" when "0011011110011000", -- t[14232] = 1
      "000001" when "0011011110011001", -- t[14233] = 1
      "000001" when "0011011110011010", -- t[14234] = 1
      "000001" when "0011011110011011", -- t[14235] = 1
      "000001" when "0011011110011100", -- t[14236] = 1
      "000001" when "0011011110011101", -- t[14237] = 1
      "000001" when "0011011110011110", -- t[14238] = 1
      "000001" when "0011011110011111", -- t[14239] = 1
      "000001" when "0011011110100000", -- t[14240] = 1
      "000001" when "0011011110100001", -- t[14241] = 1
      "000001" when "0011011110100010", -- t[14242] = 1
      "000001" when "0011011110100011", -- t[14243] = 1
      "000001" when "0011011110100100", -- t[14244] = 1
      "000001" when "0011011110100101", -- t[14245] = 1
      "000001" when "0011011110100110", -- t[14246] = 1
      "000001" when "0011011110100111", -- t[14247] = 1
      "000001" when "0011011110101000", -- t[14248] = 1
      "000001" when "0011011110101001", -- t[14249] = 1
      "000001" when "0011011110101010", -- t[14250] = 1
      "000001" when "0011011110101011", -- t[14251] = 1
      "000001" when "0011011110101100", -- t[14252] = 1
      "000001" when "0011011110101101", -- t[14253] = 1
      "000001" when "0011011110101110", -- t[14254] = 1
      "000001" when "0011011110101111", -- t[14255] = 1
      "000001" when "0011011110110000", -- t[14256] = 1
      "000001" when "0011011110110001", -- t[14257] = 1
      "000001" when "0011011110110010", -- t[14258] = 1
      "000001" when "0011011110110011", -- t[14259] = 1
      "000001" when "0011011110110100", -- t[14260] = 1
      "000001" when "0011011110110101", -- t[14261] = 1
      "000001" when "0011011110110110", -- t[14262] = 1
      "000001" when "0011011110110111", -- t[14263] = 1
      "000001" when "0011011110111000", -- t[14264] = 1
      "000001" when "0011011110111001", -- t[14265] = 1
      "000001" when "0011011110111010", -- t[14266] = 1
      "000001" when "0011011110111011", -- t[14267] = 1
      "000001" when "0011011110111100", -- t[14268] = 1
      "000001" when "0011011110111101", -- t[14269] = 1
      "000001" when "0011011110111110", -- t[14270] = 1
      "000001" when "0011011110111111", -- t[14271] = 1
      "000001" when "0011011111000000", -- t[14272] = 1
      "000001" when "0011011111000001", -- t[14273] = 1
      "000001" when "0011011111000010", -- t[14274] = 1
      "000001" when "0011011111000011", -- t[14275] = 1
      "000001" when "0011011111000100", -- t[14276] = 1
      "000001" when "0011011111000101", -- t[14277] = 1
      "000001" when "0011011111000110", -- t[14278] = 1
      "000001" when "0011011111000111", -- t[14279] = 1
      "000001" when "0011011111001000", -- t[14280] = 1
      "000001" when "0011011111001001", -- t[14281] = 1
      "000001" when "0011011111001010", -- t[14282] = 1
      "000001" when "0011011111001011", -- t[14283] = 1
      "000001" when "0011011111001100", -- t[14284] = 1
      "000001" when "0011011111001101", -- t[14285] = 1
      "000001" when "0011011111001110", -- t[14286] = 1
      "000001" when "0011011111001111", -- t[14287] = 1
      "000001" when "0011011111010000", -- t[14288] = 1
      "000001" when "0011011111010001", -- t[14289] = 1
      "000001" when "0011011111010010", -- t[14290] = 1
      "000001" when "0011011111010011", -- t[14291] = 1
      "000001" when "0011011111010100", -- t[14292] = 1
      "000001" when "0011011111010101", -- t[14293] = 1
      "000001" when "0011011111010110", -- t[14294] = 1
      "000001" when "0011011111010111", -- t[14295] = 1
      "000001" when "0011011111011000", -- t[14296] = 1
      "000001" when "0011011111011001", -- t[14297] = 1
      "000001" when "0011011111011010", -- t[14298] = 1
      "000001" when "0011011111011011", -- t[14299] = 1
      "000001" when "0011011111011100", -- t[14300] = 1
      "000001" when "0011011111011101", -- t[14301] = 1
      "000001" when "0011011111011110", -- t[14302] = 1
      "000001" when "0011011111011111", -- t[14303] = 1
      "000001" when "0011011111100000", -- t[14304] = 1
      "000001" when "0011011111100001", -- t[14305] = 1
      "000001" when "0011011111100010", -- t[14306] = 1
      "000001" when "0011011111100011", -- t[14307] = 1
      "000001" when "0011011111100100", -- t[14308] = 1
      "000001" when "0011011111100101", -- t[14309] = 1
      "000001" when "0011011111100110", -- t[14310] = 1
      "000001" when "0011011111100111", -- t[14311] = 1
      "000001" when "0011011111101000", -- t[14312] = 1
      "000001" when "0011011111101001", -- t[14313] = 1
      "000001" when "0011011111101010", -- t[14314] = 1
      "000001" when "0011011111101011", -- t[14315] = 1
      "000001" when "0011011111101100", -- t[14316] = 1
      "000001" when "0011011111101101", -- t[14317] = 1
      "000001" when "0011011111101110", -- t[14318] = 1
      "000001" when "0011011111101111", -- t[14319] = 1
      "000001" when "0011011111110000", -- t[14320] = 1
      "000001" when "0011011111110001", -- t[14321] = 1
      "000001" when "0011011111110010", -- t[14322] = 1
      "000001" when "0011011111110011", -- t[14323] = 1
      "000001" when "0011011111110100", -- t[14324] = 1
      "000001" when "0011011111110101", -- t[14325] = 1
      "000001" when "0011011111110110", -- t[14326] = 1
      "000001" when "0011011111110111", -- t[14327] = 1
      "000001" when "0011011111111000", -- t[14328] = 1
      "000001" when "0011011111111001", -- t[14329] = 1
      "000001" when "0011011111111010", -- t[14330] = 1
      "000001" when "0011011111111011", -- t[14331] = 1
      "000001" when "0011011111111100", -- t[14332] = 1
      "000001" when "0011011111111101", -- t[14333] = 1
      "000001" when "0011011111111110", -- t[14334] = 1
      "000001" when "0011011111111111", -- t[14335] = 1
      "000001" when "0011100000000000", -- t[14336] = 1
      "000001" when "0011100000000001", -- t[14337] = 1
      "000001" when "0011100000000010", -- t[14338] = 1
      "000001" when "0011100000000011", -- t[14339] = 1
      "000001" when "0011100000000100", -- t[14340] = 1
      "000001" when "0011100000000101", -- t[14341] = 1
      "000001" when "0011100000000110", -- t[14342] = 1
      "000001" when "0011100000000111", -- t[14343] = 1
      "000001" when "0011100000001000", -- t[14344] = 1
      "000001" when "0011100000001001", -- t[14345] = 1
      "000001" when "0011100000001010", -- t[14346] = 1
      "000001" when "0011100000001011", -- t[14347] = 1
      "000001" when "0011100000001100", -- t[14348] = 1
      "000001" when "0011100000001101", -- t[14349] = 1
      "000001" when "0011100000001110", -- t[14350] = 1
      "000001" when "0011100000001111", -- t[14351] = 1
      "000001" when "0011100000010000", -- t[14352] = 1
      "000001" when "0011100000010001", -- t[14353] = 1
      "000001" when "0011100000010010", -- t[14354] = 1
      "000001" when "0011100000010011", -- t[14355] = 1
      "000001" when "0011100000010100", -- t[14356] = 1
      "000001" when "0011100000010101", -- t[14357] = 1
      "000001" when "0011100000010110", -- t[14358] = 1
      "000001" when "0011100000010111", -- t[14359] = 1
      "000001" when "0011100000011000", -- t[14360] = 1
      "000001" when "0011100000011001", -- t[14361] = 1
      "000001" when "0011100000011010", -- t[14362] = 1
      "000001" when "0011100000011011", -- t[14363] = 1
      "000001" when "0011100000011100", -- t[14364] = 1
      "000001" when "0011100000011101", -- t[14365] = 1
      "000001" when "0011100000011110", -- t[14366] = 1
      "000001" when "0011100000011111", -- t[14367] = 1
      "000001" when "0011100000100000", -- t[14368] = 1
      "000001" when "0011100000100001", -- t[14369] = 1
      "000001" when "0011100000100010", -- t[14370] = 1
      "000001" when "0011100000100011", -- t[14371] = 1
      "000001" when "0011100000100100", -- t[14372] = 1
      "000001" when "0011100000100101", -- t[14373] = 1
      "000001" when "0011100000100110", -- t[14374] = 1
      "000001" when "0011100000100111", -- t[14375] = 1
      "000001" when "0011100000101000", -- t[14376] = 1
      "000001" when "0011100000101001", -- t[14377] = 1
      "000001" when "0011100000101010", -- t[14378] = 1
      "000001" when "0011100000101011", -- t[14379] = 1
      "000001" when "0011100000101100", -- t[14380] = 1
      "000001" when "0011100000101101", -- t[14381] = 1
      "000001" when "0011100000101110", -- t[14382] = 1
      "000001" when "0011100000101111", -- t[14383] = 1
      "000001" when "0011100000110000", -- t[14384] = 1
      "000001" when "0011100000110001", -- t[14385] = 1
      "000001" when "0011100000110010", -- t[14386] = 1
      "000001" when "0011100000110011", -- t[14387] = 1
      "000001" when "0011100000110100", -- t[14388] = 1
      "000001" when "0011100000110101", -- t[14389] = 1
      "000001" when "0011100000110110", -- t[14390] = 1
      "000001" when "0011100000110111", -- t[14391] = 1
      "000001" when "0011100000111000", -- t[14392] = 1
      "000001" when "0011100000111001", -- t[14393] = 1
      "000001" when "0011100000111010", -- t[14394] = 1
      "000001" when "0011100000111011", -- t[14395] = 1
      "000001" when "0011100000111100", -- t[14396] = 1
      "000001" when "0011100000111101", -- t[14397] = 1
      "000001" when "0011100000111110", -- t[14398] = 1
      "000001" when "0011100000111111", -- t[14399] = 1
      "000001" when "0011100001000000", -- t[14400] = 1
      "000001" when "0011100001000001", -- t[14401] = 1
      "000001" when "0011100001000010", -- t[14402] = 1
      "000001" when "0011100001000011", -- t[14403] = 1
      "000001" when "0011100001000100", -- t[14404] = 1
      "000001" when "0011100001000101", -- t[14405] = 1
      "000001" when "0011100001000110", -- t[14406] = 1
      "000001" when "0011100001000111", -- t[14407] = 1
      "000001" when "0011100001001000", -- t[14408] = 1
      "000001" when "0011100001001001", -- t[14409] = 1
      "000001" when "0011100001001010", -- t[14410] = 1
      "000001" when "0011100001001011", -- t[14411] = 1
      "000001" when "0011100001001100", -- t[14412] = 1
      "000001" when "0011100001001101", -- t[14413] = 1
      "000001" when "0011100001001110", -- t[14414] = 1
      "000001" when "0011100001001111", -- t[14415] = 1
      "000001" when "0011100001010000", -- t[14416] = 1
      "000001" when "0011100001010001", -- t[14417] = 1
      "000001" when "0011100001010010", -- t[14418] = 1
      "000001" when "0011100001010011", -- t[14419] = 1
      "000001" when "0011100001010100", -- t[14420] = 1
      "000001" when "0011100001010101", -- t[14421] = 1
      "000001" when "0011100001010110", -- t[14422] = 1
      "000001" when "0011100001010111", -- t[14423] = 1
      "000001" when "0011100001011000", -- t[14424] = 1
      "000001" when "0011100001011001", -- t[14425] = 1
      "000001" when "0011100001011010", -- t[14426] = 1
      "000001" when "0011100001011011", -- t[14427] = 1
      "000001" when "0011100001011100", -- t[14428] = 1
      "000001" when "0011100001011101", -- t[14429] = 1
      "000001" when "0011100001011110", -- t[14430] = 1
      "000001" when "0011100001011111", -- t[14431] = 1
      "000001" when "0011100001100000", -- t[14432] = 1
      "000001" when "0011100001100001", -- t[14433] = 1
      "000001" when "0011100001100010", -- t[14434] = 1
      "000001" when "0011100001100011", -- t[14435] = 1
      "000001" when "0011100001100100", -- t[14436] = 1
      "000001" when "0011100001100101", -- t[14437] = 1
      "000001" when "0011100001100110", -- t[14438] = 1
      "000001" when "0011100001100111", -- t[14439] = 1
      "000001" when "0011100001101000", -- t[14440] = 1
      "000001" when "0011100001101001", -- t[14441] = 1
      "000001" when "0011100001101010", -- t[14442] = 1
      "000001" when "0011100001101011", -- t[14443] = 1
      "000001" when "0011100001101100", -- t[14444] = 1
      "000001" when "0011100001101101", -- t[14445] = 1
      "000001" when "0011100001101110", -- t[14446] = 1
      "000001" when "0011100001101111", -- t[14447] = 1
      "000001" when "0011100001110000", -- t[14448] = 1
      "000001" when "0011100001110001", -- t[14449] = 1
      "000001" when "0011100001110010", -- t[14450] = 1
      "000001" when "0011100001110011", -- t[14451] = 1
      "000001" when "0011100001110100", -- t[14452] = 1
      "000001" when "0011100001110101", -- t[14453] = 1
      "000001" when "0011100001110110", -- t[14454] = 1
      "000001" when "0011100001110111", -- t[14455] = 1
      "000001" when "0011100001111000", -- t[14456] = 1
      "000001" when "0011100001111001", -- t[14457] = 1
      "000001" when "0011100001111010", -- t[14458] = 1
      "000001" when "0011100001111011", -- t[14459] = 1
      "000001" when "0011100001111100", -- t[14460] = 1
      "000001" when "0011100001111101", -- t[14461] = 1
      "000001" when "0011100001111110", -- t[14462] = 1
      "000001" when "0011100001111111", -- t[14463] = 1
      "000001" when "0011100010000000", -- t[14464] = 1
      "000001" when "0011100010000001", -- t[14465] = 1
      "000001" when "0011100010000010", -- t[14466] = 1
      "000001" when "0011100010000011", -- t[14467] = 1
      "000001" when "0011100010000100", -- t[14468] = 1
      "000001" when "0011100010000101", -- t[14469] = 1
      "000001" when "0011100010000110", -- t[14470] = 1
      "000001" when "0011100010000111", -- t[14471] = 1
      "000001" when "0011100010001000", -- t[14472] = 1
      "000001" when "0011100010001001", -- t[14473] = 1
      "000001" when "0011100010001010", -- t[14474] = 1
      "000001" when "0011100010001011", -- t[14475] = 1
      "000001" when "0011100010001100", -- t[14476] = 1
      "000001" when "0011100010001101", -- t[14477] = 1
      "000001" when "0011100010001110", -- t[14478] = 1
      "000001" when "0011100010001111", -- t[14479] = 1
      "000001" when "0011100010010000", -- t[14480] = 1
      "000001" when "0011100010010001", -- t[14481] = 1
      "000001" when "0011100010010010", -- t[14482] = 1
      "000001" when "0011100010010011", -- t[14483] = 1
      "000001" when "0011100010010100", -- t[14484] = 1
      "000001" when "0011100010010101", -- t[14485] = 1
      "000001" when "0011100010010110", -- t[14486] = 1
      "000001" when "0011100010010111", -- t[14487] = 1
      "000001" when "0011100010011000", -- t[14488] = 1
      "000001" when "0011100010011001", -- t[14489] = 1
      "000001" when "0011100010011010", -- t[14490] = 1
      "000001" when "0011100010011011", -- t[14491] = 1
      "000001" when "0011100010011100", -- t[14492] = 1
      "000001" when "0011100010011101", -- t[14493] = 1
      "000001" when "0011100010011110", -- t[14494] = 1
      "000001" when "0011100010011111", -- t[14495] = 1
      "000001" when "0011100010100000", -- t[14496] = 1
      "000001" when "0011100010100001", -- t[14497] = 1
      "000001" when "0011100010100010", -- t[14498] = 1
      "000001" when "0011100010100011", -- t[14499] = 1
      "000001" when "0011100010100100", -- t[14500] = 1
      "000001" when "0011100010100101", -- t[14501] = 1
      "000001" when "0011100010100110", -- t[14502] = 1
      "000001" when "0011100010100111", -- t[14503] = 1
      "000001" when "0011100010101000", -- t[14504] = 1
      "000001" when "0011100010101001", -- t[14505] = 1
      "000001" when "0011100010101010", -- t[14506] = 1
      "000001" when "0011100010101011", -- t[14507] = 1
      "000001" when "0011100010101100", -- t[14508] = 1
      "000001" when "0011100010101101", -- t[14509] = 1
      "000001" when "0011100010101110", -- t[14510] = 1
      "000001" when "0011100010101111", -- t[14511] = 1
      "000001" when "0011100010110000", -- t[14512] = 1
      "000001" when "0011100010110001", -- t[14513] = 1
      "000001" when "0011100010110010", -- t[14514] = 1
      "000001" when "0011100010110011", -- t[14515] = 1
      "000001" when "0011100010110100", -- t[14516] = 1
      "000001" when "0011100010110101", -- t[14517] = 1
      "000001" when "0011100010110110", -- t[14518] = 1
      "000001" when "0011100010110111", -- t[14519] = 1
      "000001" when "0011100010111000", -- t[14520] = 1
      "000001" when "0011100010111001", -- t[14521] = 1
      "000001" when "0011100010111010", -- t[14522] = 1
      "000001" when "0011100010111011", -- t[14523] = 1
      "000001" when "0011100010111100", -- t[14524] = 1
      "000001" when "0011100010111101", -- t[14525] = 1
      "000001" when "0011100010111110", -- t[14526] = 1
      "000001" when "0011100010111111", -- t[14527] = 1
      "000001" when "0011100011000000", -- t[14528] = 1
      "000001" when "0011100011000001", -- t[14529] = 1
      "000001" when "0011100011000010", -- t[14530] = 1
      "000001" when "0011100011000011", -- t[14531] = 1
      "000001" when "0011100011000100", -- t[14532] = 1
      "000001" when "0011100011000101", -- t[14533] = 1
      "000001" when "0011100011000110", -- t[14534] = 1
      "000001" when "0011100011000111", -- t[14535] = 1
      "000001" when "0011100011001000", -- t[14536] = 1
      "000001" when "0011100011001001", -- t[14537] = 1
      "000001" when "0011100011001010", -- t[14538] = 1
      "000001" when "0011100011001011", -- t[14539] = 1
      "000001" when "0011100011001100", -- t[14540] = 1
      "000001" when "0011100011001101", -- t[14541] = 1
      "000001" when "0011100011001110", -- t[14542] = 1
      "000001" when "0011100011001111", -- t[14543] = 1
      "000001" when "0011100011010000", -- t[14544] = 1
      "000001" when "0011100011010001", -- t[14545] = 1
      "000001" when "0011100011010010", -- t[14546] = 1
      "000001" when "0011100011010011", -- t[14547] = 1
      "000001" when "0011100011010100", -- t[14548] = 1
      "000001" when "0011100011010101", -- t[14549] = 1
      "000001" when "0011100011010110", -- t[14550] = 1
      "000001" when "0011100011010111", -- t[14551] = 1
      "000001" when "0011100011011000", -- t[14552] = 1
      "000001" when "0011100011011001", -- t[14553] = 1
      "000001" when "0011100011011010", -- t[14554] = 1
      "000001" when "0011100011011011", -- t[14555] = 1
      "000001" when "0011100011011100", -- t[14556] = 1
      "000001" when "0011100011011101", -- t[14557] = 1
      "000001" when "0011100011011110", -- t[14558] = 1
      "000001" when "0011100011011111", -- t[14559] = 1
      "000001" when "0011100011100000", -- t[14560] = 1
      "000001" when "0011100011100001", -- t[14561] = 1
      "000001" when "0011100011100010", -- t[14562] = 1
      "000001" when "0011100011100011", -- t[14563] = 1
      "000001" when "0011100011100100", -- t[14564] = 1
      "000001" when "0011100011100101", -- t[14565] = 1
      "000001" when "0011100011100110", -- t[14566] = 1
      "000001" when "0011100011100111", -- t[14567] = 1
      "000001" when "0011100011101000", -- t[14568] = 1
      "000001" when "0011100011101001", -- t[14569] = 1
      "000001" when "0011100011101010", -- t[14570] = 1
      "000001" when "0011100011101011", -- t[14571] = 1
      "000001" when "0011100011101100", -- t[14572] = 1
      "000001" when "0011100011101101", -- t[14573] = 1
      "000001" when "0011100011101110", -- t[14574] = 1
      "000001" when "0011100011101111", -- t[14575] = 1
      "000001" when "0011100011110000", -- t[14576] = 1
      "000001" when "0011100011110001", -- t[14577] = 1
      "000001" when "0011100011110010", -- t[14578] = 1
      "000001" when "0011100011110011", -- t[14579] = 1
      "000001" when "0011100011110100", -- t[14580] = 1
      "000001" when "0011100011110101", -- t[14581] = 1
      "000001" when "0011100011110110", -- t[14582] = 1
      "000001" when "0011100011110111", -- t[14583] = 1
      "000001" when "0011100011111000", -- t[14584] = 1
      "000001" when "0011100011111001", -- t[14585] = 1
      "000001" when "0011100011111010", -- t[14586] = 1
      "000001" when "0011100011111011", -- t[14587] = 1
      "000001" when "0011100011111100", -- t[14588] = 1
      "000001" when "0011100011111101", -- t[14589] = 1
      "000001" when "0011100011111110", -- t[14590] = 1
      "000001" when "0011100011111111", -- t[14591] = 1
      "000001" when "0011100100000000", -- t[14592] = 1
      "000001" when "0011100100000001", -- t[14593] = 1
      "000001" when "0011100100000010", -- t[14594] = 1
      "000001" when "0011100100000011", -- t[14595] = 1
      "000001" when "0011100100000100", -- t[14596] = 1
      "000001" when "0011100100000101", -- t[14597] = 1
      "000001" when "0011100100000110", -- t[14598] = 1
      "000001" when "0011100100000111", -- t[14599] = 1
      "000001" when "0011100100001000", -- t[14600] = 1
      "000001" when "0011100100001001", -- t[14601] = 1
      "000001" when "0011100100001010", -- t[14602] = 1
      "000001" when "0011100100001011", -- t[14603] = 1
      "000001" when "0011100100001100", -- t[14604] = 1
      "000001" when "0011100100001101", -- t[14605] = 1
      "000001" when "0011100100001110", -- t[14606] = 1
      "000001" when "0011100100001111", -- t[14607] = 1
      "000001" when "0011100100010000", -- t[14608] = 1
      "000001" when "0011100100010001", -- t[14609] = 1
      "000001" when "0011100100010010", -- t[14610] = 1
      "000001" when "0011100100010011", -- t[14611] = 1
      "000001" when "0011100100010100", -- t[14612] = 1
      "000001" when "0011100100010101", -- t[14613] = 1
      "000001" when "0011100100010110", -- t[14614] = 1
      "000001" when "0011100100010111", -- t[14615] = 1
      "000001" when "0011100100011000", -- t[14616] = 1
      "000001" when "0011100100011001", -- t[14617] = 1
      "000001" when "0011100100011010", -- t[14618] = 1
      "000001" when "0011100100011011", -- t[14619] = 1
      "000001" when "0011100100011100", -- t[14620] = 1
      "000001" when "0011100100011101", -- t[14621] = 1
      "000001" when "0011100100011110", -- t[14622] = 1
      "000001" when "0011100100011111", -- t[14623] = 1
      "000001" when "0011100100100000", -- t[14624] = 1
      "000001" when "0011100100100001", -- t[14625] = 1
      "000001" when "0011100100100010", -- t[14626] = 1
      "000001" when "0011100100100011", -- t[14627] = 1
      "000001" when "0011100100100100", -- t[14628] = 1
      "000001" when "0011100100100101", -- t[14629] = 1
      "000001" when "0011100100100110", -- t[14630] = 1
      "000001" when "0011100100100111", -- t[14631] = 1
      "000001" when "0011100100101000", -- t[14632] = 1
      "000001" when "0011100100101001", -- t[14633] = 1
      "000001" when "0011100100101010", -- t[14634] = 1
      "000001" when "0011100100101011", -- t[14635] = 1
      "000001" when "0011100100101100", -- t[14636] = 1
      "000001" when "0011100100101101", -- t[14637] = 1
      "000001" when "0011100100101110", -- t[14638] = 1
      "000001" when "0011100100101111", -- t[14639] = 1
      "000001" when "0011100100110000", -- t[14640] = 1
      "000001" when "0011100100110001", -- t[14641] = 1
      "000001" when "0011100100110010", -- t[14642] = 1
      "000001" when "0011100100110011", -- t[14643] = 1
      "000001" when "0011100100110100", -- t[14644] = 1
      "000001" when "0011100100110101", -- t[14645] = 1
      "000001" when "0011100100110110", -- t[14646] = 1
      "000001" when "0011100100110111", -- t[14647] = 1
      "000001" when "0011100100111000", -- t[14648] = 1
      "000001" when "0011100100111001", -- t[14649] = 1
      "000001" when "0011100100111010", -- t[14650] = 1
      "000001" when "0011100100111011", -- t[14651] = 1
      "000001" when "0011100100111100", -- t[14652] = 1
      "000001" when "0011100100111101", -- t[14653] = 1
      "000001" when "0011100100111110", -- t[14654] = 1
      "000001" when "0011100100111111", -- t[14655] = 1
      "000001" when "0011100101000000", -- t[14656] = 1
      "000001" when "0011100101000001", -- t[14657] = 1
      "000001" when "0011100101000010", -- t[14658] = 1
      "000001" when "0011100101000011", -- t[14659] = 1
      "000001" when "0011100101000100", -- t[14660] = 1
      "000001" when "0011100101000101", -- t[14661] = 1
      "000001" when "0011100101000110", -- t[14662] = 1
      "000001" when "0011100101000111", -- t[14663] = 1
      "000001" when "0011100101001000", -- t[14664] = 1
      "000001" when "0011100101001001", -- t[14665] = 1
      "000001" when "0011100101001010", -- t[14666] = 1
      "000001" when "0011100101001011", -- t[14667] = 1
      "000001" when "0011100101001100", -- t[14668] = 1
      "000001" when "0011100101001101", -- t[14669] = 1
      "000001" when "0011100101001110", -- t[14670] = 1
      "000001" when "0011100101001111", -- t[14671] = 1
      "000001" when "0011100101010000", -- t[14672] = 1
      "000001" when "0011100101010001", -- t[14673] = 1
      "000001" when "0011100101010010", -- t[14674] = 1
      "000001" when "0011100101010011", -- t[14675] = 1
      "000001" when "0011100101010100", -- t[14676] = 1
      "000001" when "0011100101010101", -- t[14677] = 1
      "000001" when "0011100101010110", -- t[14678] = 1
      "000001" when "0011100101010111", -- t[14679] = 1
      "000001" when "0011100101011000", -- t[14680] = 1
      "000001" when "0011100101011001", -- t[14681] = 1
      "000001" when "0011100101011010", -- t[14682] = 1
      "000001" when "0011100101011011", -- t[14683] = 1
      "000001" when "0011100101011100", -- t[14684] = 1
      "000001" when "0011100101011101", -- t[14685] = 1
      "000001" when "0011100101011110", -- t[14686] = 1
      "000001" when "0011100101011111", -- t[14687] = 1
      "000001" when "0011100101100000", -- t[14688] = 1
      "000001" when "0011100101100001", -- t[14689] = 1
      "000001" when "0011100101100010", -- t[14690] = 1
      "000001" when "0011100101100011", -- t[14691] = 1
      "000001" when "0011100101100100", -- t[14692] = 1
      "000001" when "0011100101100101", -- t[14693] = 1
      "000001" when "0011100101100110", -- t[14694] = 1
      "000001" when "0011100101100111", -- t[14695] = 1
      "000001" when "0011100101101000", -- t[14696] = 1
      "000001" when "0011100101101001", -- t[14697] = 1
      "000001" when "0011100101101010", -- t[14698] = 1
      "000001" when "0011100101101011", -- t[14699] = 1
      "000001" when "0011100101101100", -- t[14700] = 1
      "000001" when "0011100101101101", -- t[14701] = 1
      "000001" when "0011100101101110", -- t[14702] = 1
      "000001" when "0011100101101111", -- t[14703] = 1
      "000001" when "0011100101110000", -- t[14704] = 1
      "000001" when "0011100101110001", -- t[14705] = 1
      "000001" when "0011100101110010", -- t[14706] = 1
      "000001" when "0011100101110011", -- t[14707] = 1
      "000001" when "0011100101110100", -- t[14708] = 1
      "000001" when "0011100101110101", -- t[14709] = 1
      "000001" when "0011100101110110", -- t[14710] = 1
      "000001" when "0011100101110111", -- t[14711] = 1
      "000001" when "0011100101111000", -- t[14712] = 1
      "000001" when "0011100101111001", -- t[14713] = 1
      "000001" when "0011100101111010", -- t[14714] = 1
      "000001" when "0011100101111011", -- t[14715] = 1
      "000001" when "0011100101111100", -- t[14716] = 1
      "000001" when "0011100101111101", -- t[14717] = 1
      "000001" when "0011100101111110", -- t[14718] = 1
      "000001" when "0011100101111111", -- t[14719] = 1
      "000001" when "0011100110000000", -- t[14720] = 1
      "000001" when "0011100110000001", -- t[14721] = 1
      "000001" when "0011100110000010", -- t[14722] = 1
      "000001" when "0011100110000011", -- t[14723] = 1
      "000001" when "0011100110000100", -- t[14724] = 1
      "000001" when "0011100110000101", -- t[14725] = 1
      "000001" when "0011100110000110", -- t[14726] = 1
      "000001" when "0011100110000111", -- t[14727] = 1
      "000001" when "0011100110001000", -- t[14728] = 1
      "000001" when "0011100110001001", -- t[14729] = 1
      "000001" when "0011100110001010", -- t[14730] = 1
      "000001" when "0011100110001011", -- t[14731] = 1
      "000001" when "0011100110001100", -- t[14732] = 1
      "000001" when "0011100110001101", -- t[14733] = 1
      "000001" when "0011100110001110", -- t[14734] = 1
      "000001" when "0011100110001111", -- t[14735] = 1
      "000001" when "0011100110010000", -- t[14736] = 1
      "000001" when "0011100110010001", -- t[14737] = 1
      "000001" when "0011100110010010", -- t[14738] = 1
      "000001" when "0011100110010011", -- t[14739] = 1
      "000001" when "0011100110010100", -- t[14740] = 1
      "000001" when "0011100110010101", -- t[14741] = 1
      "000001" when "0011100110010110", -- t[14742] = 1
      "000001" when "0011100110010111", -- t[14743] = 1
      "000001" when "0011100110011000", -- t[14744] = 1
      "000001" when "0011100110011001", -- t[14745] = 1
      "000001" when "0011100110011010", -- t[14746] = 1
      "000001" when "0011100110011011", -- t[14747] = 1
      "000001" when "0011100110011100", -- t[14748] = 1
      "000001" when "0011100110011101", -- t[14749] = 1
      "000001" when "0011100110011110", -- t[14750] = 1
      "000001" when "0011100110011111", -- t[14751] = 1
      "000001" when "0011100110100000", -- t[14752] = 1
      "000001" when "0011100110100001", -- t[14753] = 1
      "000001" when "0011100110100010", -- t[14754] = 1
      "000001" when "0011100110100011", -- t[14755] = 1
      "000001" when "0011100110100100", -- t[14756] = 1
      "000001" when "0011100110100101", -- t[14757] = 1
      "000001" when "0011100110100110", -- t[14758] = 1
      "000001" when "0011100110100111", -- t[14759] = 1
      "000001" when "0011100110101000", -- t[14760] = 1
      "000001" when "0011100110101001", -- t[14761] = 1
      "000001" when "0011100110101010", -- t[14762] = 1
      "000001" when "0011100110101011", -- t[14763] = 1
      "000001" when "0011100110101100", -- t[14764] = 1
      "000001" when "0011100110101101", -- t[14765] = 1
      "000001" when "0011100110101110", -- t[14766] = 1
      "000001" when "0011100110101111", -- t[14767] = 1
      "000001" when "0011100110110000", -- t[14768] = 1
      "000001" when "0011100110110001", -- t[14769] = 1
      "000001" when "0011100110110010", -- t[14770] = 1
      "000001" when "0011100110110011", -- t[14771] = 1
      "000001" when "0011100110110100", -- t[14772] = 1
      "000001" when "0011100110110101", -- t[14773] = 1
      "000001" when "0011100110110110", -- t[14774] = 1
      "000001" when "0011100110110111", -- t[14775] = 1
      "000001" when "0011100110111000", -- t[14776] = 1
      "000001" when "0011100110111001", -- t[14777] = 1
      "000001" when "0011100110111010", -- t[14778] = 1
      "000001" when "0011100110111011", -- t[14779] = 1
      "000001" when "0011100110111100", -- t[14780] = 1
      "000001" when "0011100110111101", -- t[14781] = 1
      "000001" when "0011100110111110", -- t[14782] = 1
      "000001" when "0011100110111111", -- t[14783] = 1
      "000001" when "0011100111000000", -- t[14784] = 1
      "000001" when "0011100111000001", -- t[14785] = 1
      "000001" when "0011100111000010", -- t[14786] = 1
      "000001" when "0011100111000011", -- t[14787] = 1
      "000001" when "0011100111000100", -- t[14788] = 1
      "000001" when "0011100111000101", -- t[14789] = 1
      "000001" when "0011100111000110", -- t[14790] = 1
      "000001" when "0011100111000111", -- t[14791] = 1
      "000001" when "0011100111001000", -- t[14792] = 1
      "000001" when "0011100111001001", -- t[14793] = 1
      "000001" when "0011100111001010", -- t[14794] = 1
      "000001" when "0011100111001011", -- t[14795] = 1
      "000001" when "0011100111001100", -- t[14796] = 1
      "000001" when "0011100111001101", -- t[14797] = 1
      "000001" when "0011100111001110", -- t[14798] = 1
      "000001" when "0011100111001111", -- t[14799] = 1
      "000001" when "0011100111010000", -- t[14800] = 1
      "000001" when "0011100111010001", -- t[14801] = 1
      "000001" when "0011100111010010", -- t[14802] = 1
      "000001" when "0011100111010011", -- t[14803] = 1
      "000001" when "0011100111010100", -- t[14804] = 1
      "000001" when "0011100111010101", -- t[14805] = 1
      "000001" when "0011100111010110", -- t[14806] = 1
      "000001" when "0011100111010111", -- t[14807] = 1
      "000001" when "0011100111011000", -- t[14808] = 1
      "000001" when "0011100111011001", -- t[14809] = 1
      "000001" when "0011100111011010", -- t[14810] = 1
      "000001" when "0011100111011011", -- t[14811] = 1
      "000001" when "0011100111011100", -- t[14812] = 1
      "000001" when "0011100111011101", -- t[14813] = 1
      "000001" when "0011100111011110", -- t[14814] = 1
      "000001" when "0011100111011111", -- t[14815] = 1
      "000001" when "0011100111100000", -- t[14816] = 1
      "000001" when "0011100111100001", -- t[14817] = 1
      "000001" when "0011100111100010", -- t[14818] = 1
      "000001" when "0011100111100011", -- t[14819] = 1
      "000001" when "0011100111100100", -- t[14820] = 1
      "000001" when "0011100111100101", -- t[14821] = 1
      "000001" when "0011100111100110", -- t[14822] = 1
      "000001" when "0011100111100111", -- t[14823] = 1
      "000001" when "0011100111101000", -- t[14824] = 1
      "000001" when "0011100111101001", -- t[14825] = 1
      "000001" when "0011100111101010", -- t[14826] = 1
      "000001" when "0011100111101011", -- t[14827] = 1
      "000001" when "0011100111101100", -- t[14828] = 1
      "000001" when "0011100111101101", -- t[14829] = 1
      "000001" when "0011100111101110", -- t[14830] = 1
      "000001" when "0011100111101111", -- t[14831] = 1
      "000001" when "0011100111110000", -- t[14832] = 1
      "000001" when "0011100111110001", -- t[14833] = 1
      "000001" when "0011100111110010", -- t[14834] = 1
      "000001" when "0011100111110011", -- t[14835] = 1
      "000001" when "0011100111110100", -- t[14836] = 1
      "000001" when "0011100111110101", -- t[14837] = 1
      "000001" when "0011100111110110", -- t[14838] = 1
      "000001" when "0011100111110111", -- t[14839] = 1
      "000001" when "0011100111111000", -- t[14840] = 1
      "000001" when "0011100111111001", -- t[14841] = 1
      "000001" when "0011100111111010", -- t[14842] = 1
      "000001" when "0011100111111011", -- t[14843] = 1
      "000001" when "0011100111111100", -- t[14844] = 1
      "000001" when "0011100111111101", -- t[14845] = 1
      "000001" when "0011100111111110", -- t[14846] = 1
      "000001" when "0011100111111111", -- t[14847] = 1
      "000001" when "0011101000000000", -- t[14848] = 1
      "000001" when "0011101000000001", -- t[14849] = 1
      "000001" when "0011101000000010", -- t[14850] = 1
      "000001" when "0011101000000011", -- t[14851] = 1
      "000001" when "0011101000000100", -- t[14852] = 1
      "000001" when "0011101000000101", -- t[14853] = 1
      "000001" when "0011101000000110", -- t[14854] = 1
      "000001" when "0011101000000111", -- t[14855] = 1
      "000001" when "0011101000001000", -- t[14856] = 1
      "000001" when "0011101000001001", -- t[14857] = 1
      "000001" when "0011101000001010", -- t[14858] = 1
      "000001" when "0011101000001011", -- t[14859] = 1
      "000001" when "0011101000001100", -- t[14860] = 1
      "000001" when "0011101000001101", -- t[14861] = 1
      "000001" when "0011101000001110", -- t[14862] = 1
      "000001" when "0011101000001111", -- t[14863] = 1
      "000001" when "0011101000010000", -- t[14864] = 1
      "000001" when "0011101000010001", -- t[14865] = 1
      "000001" when "0011101000010010", -- t[14866] = 1
      "000001" when "0011101000010011", -- t[14867] = 1
      "000001" when "0011101000010100", -- t[14868] = 1
      "000001" when "0011101000010101", -- t[14869] = 1
      "000001" when "0011101000010110", -- t[14870] = 1
      "000001" when "0011101000010111", -- t[14871] = 1
      "000001" when "0011101000011000", -- t[14872] = 1
      "000001" when "0011101000011001", -- t[14873] = 1
      "000001" when "0011101000011010", -- t[14874] = 1
      "000001" when "0011101000011011", -- t[14875] = 1
      "000001" when "0011101000011100", -- t[14876] = 1
      "000001" when "0011101000011101", -- t[14877] = 1
      "000001" when "0011101000011110", -- t[14878] = 1
      "000001" when "0011101000011111", -- t[14879] = 1
      "000001" when "0011101000100000", -- t[14880] = 1
      "000001" when "0011101000100001", -- t[14881] = 1
      "000001" when "0011101000100010", -- t[14882] = 1
      "000001" when "0011101000100011", -- t[14883] = 1
      "000001" when "0011101000100100", -- t[14884] = 1
      "000001" when "0011101000100101", -- t[14885] = 1
      "000001" when "0011101000100110", -- t[14886] = 1
      "000001" when "0011101000100111", -- t[14887] = 1
      "000001" when "0011101000101000", -- t[14888] = 1
      "000001" when "0011101000101001", -- t[14889] = 1
      "000001" when "0011101000101010", -- t[14890] = 1
      "000001" when "0011101000101011", -- t[14891] = 1
      "000001" when "0011101000101100", -- t[14892] = 1
      "000001" when "0011101000101101", -- t[14893] = 1
      "000001" when "0011101000101110", -- t[14894] = 1
      "000001" when "0011101000101111", -- t[14895] = 1
      "000001" when "0011101000110000", -- t[14896] = 1
      "000001" when "0011101000110001", -- t[14897] = 1
      "000001" when "0011101000110010", -- t[14898] = 1
      "000001" when "0011101000110011", -- t[14899] = 1
      "000001" when "0011101000110100", -- t[14900] = 1
      "000001" when "0011101000110101", -- t[14901] = 1
      "000001" when "0011101000110110", -- t[14902] = 1
      "000001" when "0011101000110111", -- t[14903] = 1
      "000001" when "0011101000111000", -- t[14904] = 1
      "000001" when "0011101000111001", -- t[14905] = 1
      "000001" when "0011101000111010", -- t[14906] = 1
      "000001" when "0011101000111011", -- t[14907] = 1
      "000001" when "0011101000111100", -- t[14908] = 1
      "000001" when "0011101000111101", -- t[14909] = 1
      "000001" when "0011101000111110", -- t[14910] = 1
      "000001" when "0011101000111111", -- t[14911] = 1
      "000001" when "0011101001000000", -- t[14912] = 1
      "000001" when "0011101001000001", -- t[14913] = 1
      "000001" when "0011101001000010", -- t[14914] = 1
      "000001" when "0011101001000011", -- t[14915] = 1
      "000001" when "0011101001000100", -- t[14916] = 1
      "000001" when "0011101001000101", -- t[14917] = 1
      "000001" when "0011101001000110", -- t[14918] = 1
      "000001" when "0011101001000111", -- t[14919] = 1
      "000001" when "0011101001001000", -- t[14920] = 1
      "000001" when "0011101001001001", -- t[14921] = 1
      "000001" when "0011101001001010", -- t[14922] = 1
      "000001" when "0011101001001011", -- t[14923] = 1
      "000001" when "0011101001001100", -- t[14924] = 1
      "000001" when "0011101001001101", -- t[14925] = 1
      "000001" when "0011101001001110", -- t[14926] = 1
      "000001" when "0011101001001111", -- t[14927] = 1
      "000001" when "0011101001010000", -- t[14928] = 1
      "000001" when "0011101001010001", -- t[14929] = 1
      "000001" when "0011101001010010", -- t[14930] = 1
      "000001" when "0011101001010011", -- t[14931] = 1
      "000001" when "0011101001010100", -- t[14932] = 1
      "000001" when "0011101001010101", -- t[14933] = 1
      "000001" when "0011101001010110", -- t[14934] = 1
      "000001" when "0011101001010111", -- t[14935] = 1
      "000001" when "0011101001011000", -- t[14936] = 1
      "000001" when "0011101001011001", -- t[14937] = 1
      "000001" when "0011101001011010", -- t[14938] = 1
      "000001" when "0011101001011011", -- t[14939] = 1
      "000001" when "0011101001011100", -- t[14940] = 1
      "000001" when "0011101001011101", -- t[14941] = 1
      "000001" when "0011101001011110", -- t[14942] = 1
      "000001" when "0011101001011111", -- t[14943] = 1
      "000001" when "0011101001100000", -- t[14944] = 1
      "000001" when "0011101001100001", -- t[14945] = 1
      "000001" when "0011101001100010", -- t[14946] = 1
      "000001" when "0011101001100011", -- t[14947] = 1
      "000001" when "0011101001100100", -- t[14948] = 1
      "000001" when "0011101001100101", -- t[14949] = 1
      "000001" when "0011101001100110", -- t[14950] = 1
      "000001" when "0011101001100111", -- t[14951] = 1
      "000001" when "0011101001101000", -- t[14952] = 1
      "000001" when "0011101001101001", -- t[14953] = 1
      "000001" when "0011101001101010", -- t[14954] = 1
      "000001" when "0011101001101011", -- t[14955] = 1
      "000001" when "0011101001101100", -- t[14956] = 1
      "000001" when "0011101001101101", -- t[14957] = 1
      "000001" when "0011101001101110", -- t[14958] = 1
      "000001" when "0011101001101111", -- t[14959] = 1
      "000001" when "0011101001110000", -- t[14960] = 1
      "000001" when "0011101001110001", -- t[14961] = 1
      "000001" when "0011101001110010", -- t[14962] = 1
      "000001" when "0011101001110011", -- t[14963] = 1
      "000001" when "0011101001110100", -- t[14964] = 1
      "000001" when "0011101001110101", -- t[14965] = 1
      "000001" when "0011101001110110", -- t[14966] = 1
      "000001" when "0011101001110111", -- t[14967] = 1
      "000001" when "0011101001111000", -- t[14968] = 1
      "000001" when "0011101001111001", -- t[14969] = 1
      "000001" when "0011101001111010", -- t[14970] = 1
      "000001" when "0011101001111011", -- t[14971] = 1
      "000001" when "0011101001111100", -- t[14972] = 1
      "000001" when "0011101001111101", -- t[14973] = 1
      "000001" when "0011101001111110", -- t[14974] = 1
      "000001" when "0011101001111111", -- t[14975] = 1
      "000001" when "0011101010000000", -- t[14976] = 1
      "000001" when "0011101010000001", -- t[14977] = 1
      "000001" when "0011101010000010", -- t[14978] = 1
      "000001" when "0011101010000011", -- t[14979] = 1
      "000001" when "0011101010000100", -- t[14980] = 1
      "000001" when "0011101010000101", -- t[14981] = 1
      "000001" when "0011101010000110", -- t[14982] = 1
      "000001" when "0011101010000111", -- t[14983] = 1
      "000001" when "0011101010001000", -- t[14984] = 1
      "000001" when "0011101010001001", -- t[14985] = 1
      "000001" when "0011101010001010", -- t[14986] = 1
      "000001" when "0011101010001011", -- t[14987] = 1
      "000001" when "0011101010001100", -- t[14988] = 1
      "000001" when "0011101010001101", -- t[14989] = 1
      "000001" when "0011101010001110", -- t[14990] = 1
      "000001" when "0011101010001111", -- t[14991] = 1
      "000001" when "0011101010010000", -- t[14992] = 1
      "000001" when "0011101010010001", -- t[14993] = 1
      "000001" when "0011101010010010", -- t[14994] = 1
      "000001" when "0011101010010011", -- t[14995] = 1
      "000001" when "0011101010010100", -- t[14996] = 1
      "000001" when "0011101010010101", -- t[14997] = 1
      "000001" when "0011101010010110", -- t[14998] = 1
      "000001" when "0011101010010111", -- t[14999] = 1
      "000001" when "0011101010011000", -- t[15000] = 1
      "000001" when "0011101010011001", -- t[15001] = 1
      "000001" when "0011101010011010", -- t[15002] = 1
      "000001" when "0011101010011011", -- t[15003] = 1
      "000001" when "0011101010011100", -- t[15004] = 1
      "000001" when "0011101010011101", -- t[15005] = 1
      "000001" when "0011101010011110", -- t[15006] = 1
      "000001" when "0011101010011111", -- t[15007] = 1
      "000001" when "0011101010100000", -- t[15008] = 1
      "000001" when "0011101010100001", -- t[15009] = 1
      "000001" when "0011101010100010", -- t[15010] = 1
      "000001" when "0011101010100011", -- t[15011] = 1
      "000001" when "0011101010100100", -- t[15012] = 1
      "000001" when "0011101010100101", -- t[15013] = 1
      "000001" when "0011101010100110", -- t[15014] = 1
      "000001" when "0011101010100111", -- t[15015] = 1
      "000001" when "0011101010101000", -- t[15016] = 1
      "000001" when "0011101010101001", -- t[15017] = 1
      "000001" when "0011101010101010", -- t[15018] = 1
      "000001" when "0011101010101011", -- t[15019] = 1
      "000001" when "0011101010101100", -- t[15020] = 1
      "000001" when "0011101010101101", -- t[15021] = 1
      "000001" when "0011101010101110", -- t[15022] = 1
      "000001" when "0011101010101111", -- t[15023] = 1
      "000001" when "0011101010110000", -- t[15024] = 1
      "000001" when "0011101010110001", -- t[15025] = 1
      "000001" when "0011101010110010", -- t[15026] = 1
      "000001" when "0011101010110011", -- t[15027] = 1
      "000001" when "0011101010110100", -- t[15028] = 1
      "000001" when "0011101010110101", -- t[15029] = 1
      "000001" when "0011101010110110", -- t[15030] = 1
      "000001" when "0011101010110111", -- t[15031] = 1
      "000001" when "0011101010111000", -- t[15032] = 1
      "000001" when "0011101010111001", -- t[15033] = 1
      "000001" when "0011101010111010", -- t[15034] = 1
      "000001" when "0011101010111011", -- t[15035] = 1
      "000001" when "0011101010111100", -- t[15036] = 1
      "000001" when "0011101010111101", -- t[15037] = 1
      "000001" when "0011101010111110", -- t[15038] = 1
      "000001" when "0011101010111111", -- t[15039] = 1
      "000001" when "0011101011000000", -- t[15040] = 1
      "000001" when "0011101011000001", -- t[15041] = 1
      "000001" when "0011101011000010", -- t[15042] = 1
      "000001" when "0011101011000011", -- t[15043] = 1
      "000001" when "0011101011000100", -- t[15044] = 1
      "000001" when "0011101011000101", -- t[15045] = 1
      "000001" when "0011101011000110", -- t[15046] = 1
      "000001" when "0011101011000111", -- t[15047] = 1
      "000001" when "0011101011001000", -- t[15048] = 1
      "000001" when "0011101011001001", -- t[15049] = 1
      "000001" when "0011101011001010", -- t[15050] = 1
      "000001" when "0011101011001011", -- t[15051] = 1
      "000001" when "0011101011001100", -- t[15052] = 1
      "000001" when "0011101011001101", -- t[15053] = 1
      "000001" when "0011101011001110", -- t[15054] = 1
      "000001" when "0011101011001111", -- t[15055] = 1
      "000001" when "0011101011010000", -- t[15056] = 1
      "000001" when "0011101011010001", -- t[15057] = 1
      "000001" when "0011101011010010", -- t[15058] = 1
      "000001" when "0011101011010011", -- t[15059] = 1
      "000001" when "0011101011010100", -- t[15060] = 1
      "000001" when "0011101011010101", -- t[15061] = 1
      "000001" when "0011101011010110", -- t[15062] = 1
      "000001" when "0011101011010111", -- t[15063] = 1
      "000001" when "0011101011011000", -- t[15064] = 1
      "000001" when "0011101011011001", -- t[15065] = 1
      "000001" when "0011101011011010", -- t[15066] = 1
      "000001" when "0011101011011011", -- t[15067] = 1
      "000001" when "0011101011011100", -- t[15068] = 1
      "000001" when "0011101011011101", -- t[15069] = 1
      "000001" when "0011101011011110", -- t[15070] = 1
      "000001" when "0011101011011111", -- t[15071] = 1
      "000001" when "0011101011100000", -- t[15072] = 1
      "000001" when "0011101011100001", -- t[15073] = 1
      "000001" when "0011101011100010", -- t[15074] = 1
      "000001" when "0011101011100011", -- t[15075] = 1
      "000001" when "0011101011100100", -- t[15076] = 1
      "000001" when "0011101011100101", -- t[15077] = 1
      "000001" when "0011101011100110", -- t[15078] = 1
      "000001" when "0011101011100111", -- t[15079] = 1
      "000001" when "0011101011101000", -- t[15080] = 1
      "000001" when "0011101011101001", -- t[15081] = 1
      "000001" when "0011101011101010", -- t[15082] = 1
      "000001" when "0011101011101011", -- t[15083] = 1
      "000001" when "0011101011101100", -- t[15084] = 1
      "000001" when "0011101011101101", -- t[15085] = 1
      "000001" when "0011101011101110", -- t[15086] = 1
      "000001" when "0011101011101111", -- t[15087] = 1
      "000001" when "0011101011110000", -- t[15088] = 1
      "000001" when "0011101011110001", -- t[15089] = 1
      "000001" when "0011101011110010", -- t[15090] = 1
      "000001" when "0011101011110011", -- t[15091] = 1
      "000001" when "0011101011110100", -- t[15092] = 1
      "000001" when "0011101011110101", -- t[15093] = 1
      "000001" when "0011101011110110", -- t[15094] = 1
      "000001" when "0011101011110111", -- t[15095] = 1
      "000001" when "0011101011111000", -- t[15096] = 1
      "000001" when "0011101011111001", -- t[15097] = 1
      "000001" when "0011101011111010", -- t[15098] = 1
      "000001" when "0011101011111011", -- t[15099] = 1
      "000001" when "0011101011111100", -- t[15100] = 1
      "000001" when "0011101011111101", -- t[15101] = 1
      "000001" when "0011101011111110", -- t[15102] = 1
      "000001" when "0011101011111111", -- t[15103] = 1
      "000001" when "0011101100000000", -- t[15104] = 1
      "000001" when "0011101100000001", -- t[15105] = 1
      "000001" when "0011101100000010", -- t[15106] = 1
      "000001" when "0011101100000011", -- t[15107] = 1
      "000001" when "0011101100000100", -- t[15108] = 1
      "000001" when "0011101100000101", -- t[15109] = 1
      "000001" when "0011101100000110", -- t[15110] = 1
      "000001" when "0011101100000111", -- t[15111] = 1
      "000001" when "0011101100001000", -- t[15112] = 1
      "000001" when "0011101100001001", -- t[15113] = 1
      "000001" when "0011101100001010", -- t[15114] = 1
      "000001" when "0011101100001011", -- t[15115] = 1
      "000001" when "0011101100001100", -- t[15116] = 1
      "000001" when "0011101100001101", -- t[15117] = 1
      "000001" when "0011101100001110", -- t[15118] = 1
      "000001" when "0011101100001111", -- t[15119] = 1
      "000001" when "0011101100010000", -- t[15120] = 1
      "000001" when "0011101100010001", -- t[15121] = 1
      "000001" when "0011101100010010", -- t[15122] = 1
      "000001" when "0011101100010011", -- t[15123] = 1
      "000001" when "0011101100010100", -- t[15124] = 1
      "000001" when "0011101100010101", -- t[15125] = 1
      "000001" when "0011101100010110", -- t[15126] = 1
      "000001" when "0011101100010111", -- t[15127] = 1
      "000001" when "0011101100011000", -- t[15128] = 1
      "000001" when "0011101100011001", -- t[15129] = 1
      "000001" when "0011101100011010", -- t[15130] = 1
      "000001" when "0011101100011011", -- t[15131] = 1
      "000001" when "0011101100011100", -- t[15132] = 1
      "000001" when "0011101100011101", -- t[15133] = 1
      "000001" when "0011101100011110", -- t[15134] = 1
      "000001" when "0011101100011111", -- t[15135] = 1
      "000001" when "0011101100100000", -- t[15136] = 1
      "000001" when "0011101100100001", -- t[15137] = 1
      "000001" when "0011101100100010", -- t[15138] = 1
      "000001" when "0011101100100011", -- t[15139] = 1
      "000001" when "0011101100100100", -- t[15140] = 1
      "000001" when "0011101100100101", -- t[15141] = 1
      "000001" when "0011101100100110", -- t[15142] = 1
      "000001" when "0011101100100111", -- t[15143] = 1
      "000001" when "0011101100101000", -- t[15144] = 1
      "000001" when "0011101100101001", -- t[15145] = 1
      "000001" when "0011101100101010", -- t[15146] = 1
      "000001" when "0011101100101011", -- t[15147] = 1
      "000001" when "0011101100101100", -- t[15148] = 1
      "000001" when "0011101100101101", -- t[15149] = 1
      "000001" when "0011101100101110", -- t[15150] = 1
      "000001" when "0011101100101111", -- t[15151] = 1
      "000001" when "0011101100110000", -- t[15152] = 1
      "000001" when "0011101100110001", -- t[15153] = 1
      "000001" when "0011101100110010", -- t[15154] = 1
      "000001" when "0011101100110011", -- t[15155] = 1
      "000001" when "0011101100110100", -- t[15156] = 1
      "000001" when "0011101100110101", -- t[15157] = 1
      "000001" when "0011101100110110", -- t[15158] = 1
      "000001" when "0011101100110111", -- t[15159] = 1
      "000001" when "0011101100111000", -- t[15160] = 1
      "000001" when "0011101100111001", -- t[15161] = 1
      "000001" when "0011101100111010", -- t[15162] = 1
      "000001" when "0011101100111011", -- t[15163] = 1
      "000001" when "0011101100111100", -- t[15164] = 1
      "000001" when "0011101100111101", -- t[15165] = 1
      "000001" when "0011101100111110", -- t[15166] = 1
      "000001" when "0011101100111111", -- t[15167] = 1
      "000001" when "0011101101000000", -- t[15168] = 1
      "000001" when "0011101101000001", -- t[15169] = 1
      "000001" when "0011101101000010", -- t[15170] = 1
      "000001" when "0011101101000011", -- t[15171] = 1
      "000001" when "0011101101000100", -- t[15172] = 1
      "000001" when "0011101101000101", -- t[15173] = 1
      "000001" when "0011101101000110", -- t[15174] = 1
      "000001" when "0011101101000111", -- t[15175] = 1
      "000001" when "0011101101001000", -- t[15176] = 1
      "000001" when "0011101101001001", -- t[15177] = 1
      "000001" when "0011101101001010", -- t[15178] = 1
      "000001" when "0011101101001011", -- t[15179] = 1
      "000001" when "0011101101001100", -- t[15180] = 1
      "000001" when "0011101101001101", -- t[15181] = 1
      "000001" when "0011101101001110", -- t[15182] = 1
      "000001" when "0011101101001111", -- t[15183] = 1
      "000001" when "0011101101010000", -- t[15184] = 1
      "000001" when "0011101101010001", -- t[15185] = 1
      "000001" when "0011101101010010", -- t[15186] = 1
      "000001" when "0011101101010011", -- t[15187] = 1
      "000001" when "0011101101010100", -- t[15188] = 1
      "000001" when "0011101101010101", -- t[15189] = 1
      "000001" when "0011101101010110", -- t[15190] = 1
      "000001" when "0011101101010111", -- t[15191] = 1
      "000001" when "0011101101011000", -- t[15192] = 1
      "000001" when "0011101101011001", -- t[15193] = 1
      "000001" when "0011101101011010", -- t[15194] = 1
      "000001" when "0011101101011011", -- t[15195] = 1
      "000001" when "0011101101011100", -- t[15196] = 1
      "000001" when "0011101101011101", -- t[15197] = 1
      "000001" when "0011101101011110", -- t[15198] = 1
      "000001" when "0011101101011111", -- t[15199] = 1
      "000001" when "0011101101100000", -- t[15200] = 1
      "000001" when "0011101101100001", -- t[15201] = 1
      "000001" when "0011101101100010", -- t[15202] = 1
      "000001" when "0011101101100011", -- t[15203] = 1
      "000001" when "0011101101100100", -- t[15204] = 1
      "000001" when "0011101101100101", -- t[15205] = 1
      "000001" when "0011101101100110", -- t[15206] = 1
      "000001" when "0011101101100111", -- t[15207] = 1
      "000001" when "0011101101101000", -- t[15208] = 1
      "000001" when "0011101101101001", -- t[15209] = 1
      "000001" when "0011101101101010", -- t[15210] = 1
      "000001" when "0011101101101011", -- t[15211] = 1
      "000001" when "0011101101101100", -- t[15212] = 1
      "000001" when "0011101101101101", -- t[15213] = 1
      "000001" when "0011101101101110", -- t[15214] = 1
      "000001" when "0011101101101111", -- t[15215] = 1
      "000001" when "0011101101110000", -- t[15216] = 1
      "000001" when "0011101101110001", -- t[15217] = 1
      "000001" when "0011101101110010", -- t[15218] = 1
      "000001" when "0011101101110011", -- t[15219] = 1
      "000001" when "0011101101110100", -- t[15220] = 1
      "000001" when "0011101101110101", -- t[15221] = 1
      "000001" when "0011101101110110", -- t[15222] = 1
      "000001" when "0011101101110111", -- t[15223] = 1
      "000001" when "0011101101111000", -- t[15224] = 1
      "000001" when "0011101101111001", -- t[15225] = 1
      "000001" when "0011101101111010", -- t[15226] = 1
      "000001" when "0011101101111011", -- t[15227] = 1
      "000001" when "0011101101111100", -- t[15228] = 1
      "000001" when "0011101101111101", -- t[15229] = 1
      "000001" when "0011101101111110", -- t[15230] = 1
      "000001" when "0011101101111111", -- t[15231] = 1
      "000001" when "0011101110000000", -- t[15232] = 1
      "000001" when "0011101110000001", -- t[15233] = 1
      "000001" when "0011101110000010", -- t[15234] = 1
      "000001" when "0011101110000011", -- t[15235] = 1
      "000001" when "0011101110000100", -- t[15236] = 1
      "000001" when "0011101110000101", -- t[15237] = 1
      "000001" when "0011101110000110", -- t[15238] = 1
      "000001" when "0011101110000111", -- t[15239] = 1
      "000001" when "0011101110001000", -- t[15240] = 1
      "000001" when "0011101110001001", -- t[15241] = 1
      "000001" when "0011101110001010", -- t[15242] = 1
      "000001" when "0011101110001011", -- t[15243] = 1
      "000001" when "0011101110001100", -- t[15244] = 1
      "000001" when "0011101110001101", -- t[15245] = 1
      "000001" when "0011101110001110", -- t[15246] = 1
      "000001" when "0011101110001111", -- t[15247] = 1
      "000001" when "0011101110010000", -- t[15248] = 1
      "000001" when "0011101110010001", -- t[15249] = 1
      "000001" when "0011101110010010", -- t[15250] = 1
      "000001" when "0011101110010011", -- t[15251] = 1
      "000001" when "0011101110010100", -- t[15252] = 1
      "000001" when "0011101110010101", -- t[15253] = 1
      "000001" when "0011101110010110", -- t[15254] = 1
      "000001" when "0011101110010111", -- t[15255] = 1
      "000001" when "0011101110011000", -- t[15256] = 1
      "000001" when "0011101110011001", -- t[15257] = 1
      "000001" when "0011101110011010", -- t[15258] = 1
      "000001" when "0011101110011011", -- t[15259] = 1
      "000001" when "0011101110011100", -- t[15260] = 1
      "000001" when "0011101110011101", -- t[15261] = 1
      "000001" when "0011101110011110", -- t[15262] = 1
      "000001" when "0011101110011111", -- t[15263] = 1
      "000001" when "0011101110100000", -- t[15264] = 1
      "000001" when "0011101110100001", -- t[15265] = 1
      "000001" when "0011101110100010", -- t[15266] = 1
      "000001" when "0011101110100011", -- t[15267] = 1
      "000001" when "0011101110100100", -- t[15268] = 1
      "000001" when "0011101110100101", -- t[15269] = 1
      "000001" when "0011101110100110", -- t[15270] = 1
      "000001" when "0011101110100111", -- t[15271] = 1
      "000001" when "0011101110101000", -- t[15272] = 1
      "000001" when "0011101110101001", -- t[15273] = 1
      "000001" when "0011101110101010", -- t[15274] = 1
      "000001" when "0011101110101011", -- t[15275] = 1
      "000001" when "0011101110101100", -- t[15276] = 1
      "000001" when "0011101110101101", -- t[15277] = 1
      "000001" when "0011101110101110", -- t[15278] = 1
      "000001" when "0011101110101111", -- t[15279] = 1
      "000001" when "0011101110110000", -- t[15280] = 1
      "000001" when "0011101110110001", -- t[15281] = 1
      "000001" when "0011101110110010", -- t[15282] = 1
      "000001" when "0011101110110011", -- t[15283] = 1
      "000001" when "0011101110110100", -- t[15284] = 1
      "000001" when "0011101110110101", -- t[15285] = 1
      "000001" when "0011101110110110", -- t[15286] = 1
      "000001" when "0011101110110111", -- t[15287] = 1
      "000001" when "0011101110111000", -- t[15288] = 1
      "000001" when "0011101110111001", -- t[15289] = 1
      "000001" when "0011101110111010", -- t[15290] = 1
      "000001" when "0011101110111011", -- t[15291] = 1
      "000001" when "0011101110111100", -- t[15292] = 1
      "000001" when "0011101110111101", -- t[15293] = 1
      "000001" when "0011101110111110", -- t[15294] = 1
      "000001" when "0011101110111111", -- t[15295] = 1
      "000001" when "0011101111000000", -- t[15296] = 1
      "000001" when "0011101111000001", -- t[15297] = 1
      "000001" when "0011101111000010", -- t[15298] = 1
      "000001" when "0011101111000011", -- t[15299] = 1
      "000001" when "0011101111000100", -- t[15300] = 1
      "000001" when "0011101111000101", -- t[15301] = 1
      "000001" when "0011101111000110", -- t[15302] = 1
      "000001" when "0011101111000111", -- t[15303] = 1
      "000001" when "0011101111001000", -- t[15304] = 1
      "000001" when "0011101111001001", -- t[15305] = 1
      "000001" when "0011101111001010", -- t[15306] = 1
      "000001" when "0011101111001011", -- t[15307] = 1
      "000001" when "0011101111001100", -- t[15308] = 1
      "000001" when "0011101111001101", -- t[15309] = 1
      "000001" when "0011101111001110", -- t[15310] = 1
      "000001" when "0011101111001111", -- t[15311] = 1
      "000001" when "0011101111010000", -- t[15312] = 1
      "000001" when "0011101111010001", -- t[15313] = 1
      "000001" when "0011101111010010", -- t[15314] = 1
      "000001" when "0011101111010011", -- t[15315] = 1
      "000001" when "0011101111010100", -- t[15316] = 1
      "000001" when "0011101111010101", -- t[15317] = 1
      "000001" when "0011101111010110", -- t[15318] = 1
      "000001" when "0011101111010111", -- t[15319] = 1
      "000001" when "0011101111011000", -- t[15320] = 1
      "000001" when "0011101111011001", -- t[15321] = 1
      "000001" when "0011101111011010", -- t[15322] = 1
      "000001" when "0011101111011011", -- t[15323] = 1
      "000001" when "0011101111011100", -- t[15324] = 1
      "000001" when "0011101111011101", -- t[15325] = 1
      "000001" when "0011101111011110", -- t[15326] = 1
      "000001" when "0011101111011111", -- t[15327] = 1
      "000001" when "0011101111100000", -- t[15328] = 1
      "000001" when "0011101111100001", -- t[15329] = 1
      "000001" when "0011101111100010", -- t[15330] = 1
      "000001" when "0011101111100011", -- t[15331] = 1
      "000001" when "0011101111100100", -- t[15332] = 1
      "000001" when "0011101111100101", -- t[15333] = 1
      "000001" when "0011101111100110", -- t[15334] = 1
      "000001" when "0011101111100111", -- t[15335] = 1
      "000001" when "0011101111101000", -- t[15336] = 1
      "000001" when "0011101111101001", -- t[15337] = 1
      "000001" when "0011101111101010", -- t[15338] = 1
      "000001" when "0011101111101011", -- t[15339] = 1
      "000001" when "0011101111101100", -- t[15340] = 1
      "000001" when "0011101111101101", -- t[15341] = 1
      "000001" when "0011101111101110", -- t[15342] = 1
      "000001" when "0011101111101111", -- t[15343] = 1
      "000001" when "0011101111110000", -- t[15344] = 1
      "000001" when "0011101111110001", -- t[15345] = 1
      "000001" when "0011101111110010", -- t[15346] = 1
      "000001" when "0011101111110011", -- t[15347] = 1
      "000001" when "0011101111110100", -- t[15348] = 1
      "000001" when "0011101111110101", -- t[15349] = 1
      "000001" when "0011101111110110", -- t[15350] = 1
      "000001" when "0011101111110111", -- t[15351] = 1
      "000001" when "0011101111111000", -- t[15352] = 1
      "000001" when "0011101111111001", -- t[15353] = 1
      "000001" when "0011101111111010", -- t[15354] = 1
      "000001" when "0011101111111011", -- t[15355] = 1
      "000001" when "0011101111111100", -- t[15356] = 1
      "000001" when "0011101111111101", -- t[15357] = 1
      "000001" when "0011101111111110", -- t[15358] = 1
      "000001" when "0011101111111111", -- t[15359] = 1
      "000001" when "0011110000000000", -- t[15360] = 1
      "000001" when "0011110000000001", -- t[15361] = 1
      "000001" when "0011110000000010", -- t[15362] = 1
      "000001" when "0011110000000011", -- t[15363] = 1
      "000001" when "0011110000000100", -- t[15364] = 1
      "000001" when "0011110000000101", -- t[15365] = 1
      "000001" when "0011110000000110", -- t[15366] = 1
      "000001" when "0011110000000111", -- t[15367] = 1
      "000001" when "0011110000001000", -- t[15368] = 1
      "000001" when "0011110000001001", -- t[15369] = 1
      "000001" when "0011110000001010", -- t[15370] = 1
      "000001" when "0011110000001011", -- t[15371] = 1
      "000001" when "0011110000001100", -- t[15372] = 1
      "000001" when "0011110000001101", -- t[15373] = 1
      "000001" when "0011110000001110", -- t[15374] = 1
      "000001" when "0011110000001111", -- t[15375] = 1
      "000001" when "0011110000010000", -- t[15376] = 1
      "000001" when "0011110000010001", -- t[15377] = 1
      "000001" when "0011110000010010", -- t[15378] = 1
      "000001" when "0011110000010011", -- t[15379] = 1
      "000001" when "0011110000010100", -- t[15380] = 1
      "000001" when "0011110000010101", -- t[15381] = 1
      "000001" when "0011110000010110", -- t[15382] = 1
      "000001" when "0011110000010111", -- t[15383] = 1
      "000001" when "0011110000011000", -- t[15384] = 1
      "000001" when "0011110000011001", -- t[15385] = 1
      "000001" when "0011110000011010", -- t[15386] = 1
      "000001" when "0011110000011011", -- t[15387] = 1
      "000001" when "0011110000011100", -- t[15388] = 1
      "000001" when "0011110000011101", -- t[15389] = 1
      "000001" when "0011110000011110", -- t[15390] = 1
      "000001" when "0011110000011111", -- t[15391] = 1
      "000001" when "0011110000100000", -- t[15392] = 1
      "000001" when "0011110000100001", -- t[15393] = 1
      "000001" when "0011110000100010", -- t[15394] = 1
      "000001" when "0011110000100011", -- t[15395] = 1
      "000001" when "0011110000100100", -- t[15396] = 1
      "000001" when "0011110000100101", -- t[15397] = 1
      "000001" when "0011110000100110", -- t[15398] = 1
      "000001" when "0011110000100111", -- t[15399] = 1
      "000001" when "0011110000101000", -- t[15400] = 1
      "000001" when "0011110000101001", -- t[15401] = 1
      "000001" when "0011110000101010", -- t[15402] = 1
      "000001" when "0011110000101011", -- t[15403] = 1
      "000001" when "0011110000101100", -- t[15404] = 1
      "000001" when "0011110000101101", -- t[15405] = 1
      "000001" when "0011110000101110", -- t[15406] = 1
      "000001" when "0011110000101111", -- t[15407] = 1
      "000001" when "0011110000110000", -- t[15408] = 1
      "000001" when "0011110000110001", -- t[15409] = 1
      "000001" when "0011110000110010", -- t[15410] = 1
      "000001" when "0011110000110011", -- t[15411] = 1
      "000001" when "0011110000110100", -- t[15412] = 1
      "000001" when "0011110000110101", -- t[15413] = 1
      "000001" when "0011110000110110", -- t[15414] = 1
      "000001" when "0011110000110111", -- t[15415] = 1
      "000001" when "0011110000111000", -- t[15416] = 1
      "000001" when "0011110000111001", -- t[15417] = 1
      "000001" when "0011110000111010", -- t[15418] = 1
      "000001" when "0011110000111011", -- t[15419] = 1
      "000001" when "0011110000111100", -- t[15420] = 1
      "000001" when "0011110000111101", -- t[15421] = 1
      "000001" when "0011110000111110", -- t[15422] = 1
      "000001" when "0011110000111111", -- t[15423] = 1
      "000001" when "0011110001000000", -- t[15424] = 1
      "000001" when "0011110001000001", -- t[15425] = 1
      "000001" when "0011110001000010", -- t[15426] = 1
      "000001" when "0011110001000011", -- t[15427] = 1
      "000001" when "0011110001000100", -- t[15428] = 1
      "000001" when "0011110001000101", -- t[15429] = 1
      "000001" when "0011110001000110", -- t[15430] = 1
      "000001" when "0011110001000111", -- t[15431] = 1
      "000001" when "0011110001001000", -- t[15432] = 1
      "000001" when "0011110001001001", -- t[15433] = 1
      "000001" when "0011110001001010", -- t[15434] = 1
      "000001" when "0011110001001011", -- t[15435] = 1
      "000001" when "0011110001001100", -- t[15436] = 1
      "000001" when "0011110001001101", -- t[15437] = 1
      "000001" when "0011110001001110", -- t[15438] = 1
      "000001" when "0011110001001111", -- t[15439] = 1
      "000001" when "0011110001010000", -- t[15440] = 1
      "000001" when "0011110001010001", -- t[15441] = 1
      "000001" when "0011110001010010", -- t[15442] = 1
      "000001" when "0011110001010011", -- t[15443] = 1
      "000001" when "0011110001010100", -- t[15444] = 1
      "000001" when "0011110001010101", -- t[15445] = 1
      "000001" when "0011110001010110", -- t[15446] = 1
      "000001" when "0011110001010111", -- t[15447] = 1
      "000001" when "0011110001011000", -- t[15448] = 1
      "000001" when "0011110001011001", -- t[15449] = 1
      "000001" when "0011110001011010", -- t[15450] = 1
      "000001" when "0011110001011011", -- t[15451] = 1
      "000001" when "0011110001011100", -- t[15452] = 1
      "000001" when "0011110001011101", -- t[15453] = 1
      "000001" when "0011110001011110", -- t[15454] = 1
      "000001" when "0011110001011111", -- t[15455] = 1
      "000001" when "0011110001100000", -- t[15456] = 1
      "000001" when "0011110001100001", -- t[15457] = 1
      "000001" when "0011110001100010", -- t[15458] = 1
      "000001" when "0011110001100011", -- t[15459] = 1
      "000001" when "0011110001100100", -- t[15460] = 1
      "000001" when "0011110001100101", -- t[15461] = 1
      "000001" when "0011110001100110", -- t[15462] = 1
      "000001" when "0011110001100111", -- t[15463] = 1
      "000001" when "0011110001101000", -- t[15464] = 1
      "000001" when "0011110001101001", -- t[15465] = 1
      "000001" when "0011110001101010", -- t[15466] = 1
      "000001" when "0011110001101011", -- t[15467] = 1
      "000001" when "0011110001101100", -- t[15468] = 1
      "000001" when "0011110001101101", -- t[15469] = 1
      "000001" when "0011110001101110", -- t[15470] = 1
      "000001" when "0011110001101111", -- t[15471] = 1
      "000001" when "0011110001110000", -- t[15472] = 1
      "000001" when "0011110001110001", -- t[15473] = 1
      "000001" when "0011110001110010", -- t[15474] = 1
      "000001" when "0011110001110011", -- t[15475] = 1
      "000001" when "0011110001110100", -- t[15476] = 1
      "000001" when "0011110001110101", -- t[15477] = 1
      "000001" when "0011110001110110", -- t[15478] = 1
      "000001" when "0011110001110111", -- t[15479] = 1
      "000001" when "0011110001111000", -- t[15480] = 1
      "000001" when "0011110001111001", -- t[15481] = 1
      "000001" when "0011110001111010", -- t[15482] = 1
      "000001" when "0011110001111011", -- t[15483] = 1
      "000001" when "0011110001111100", -- t[15484] = 1
      "000001" when "0011110001111101", -- t[15485] = 1
      "000001" when "0011110001111110", -- t[15486] = 1
      "000001" when "0011110001111111", -- t[15487] = 1
      "000001" when "0011110010000000", -- t[15488] = 1
      "000001" when "0011110010000001", -- t[15489] = 1
      "000001" when "0011110010000010", -- t[15490] = 1
      "000001" when "0011110010000011", -- t[15491] = 1
      "000001" when "0011110010000100", -- t[15492] = 1
      "000001" when "0011110010000101", -- t[15493] = 1
      "000001" when "0011110010000110", -- t[15494] = 1
      "000001" when "0011110010000111", -- t[15495] = 1
      "000001" when "0011110010001000", -- t[15496] = 1
      "000001" when "0011110010001001", -- t[15497] = 1
      "000001" when "0011110010001010", -- t[15498] = 1
      "000001" when "0011110010001011", -- t[15499] = 1
      "000001" when "0011110010001100", -- t[15500] = 1
      "000001" when "0011110010001101", -- t[15501] = 1
      "000001" when "0011110010001110", -- t[15502] = 1
      "000001" when "0011110010001111", -- t[15503] = 1
      "000001" when "0011110010010000", -- t[15504] = 1
      "000001" when "0011110010010001", -- t[15505] = 1
      "000001" when "0011110010010010", -- t[15506] = 1
      "000001" when "0011110010010011", -- t[15507] = 1
      "000001" when "0011110010010100", -- t[15508] = 1
      "000001" when "0011110010010101", -- t[15509] = 1
      "000001" when "0011110010010110", -- t[15510] = 1
      "000001" when "0011110010010111", -- t[15511] = 1
      "000001" when "0011110010011000", -- t[15512] = 1
      "000001" when "0011110010011001", -- t[15513] = 1
      "000001" when "0011110010011010", -- t[15514] = 1
      "000001" when "0011110010011011", -- t[15515] = 1
      "000001" when "0011110010011100", -- t[15516] = 1
      "000001" when "0011110010011101", -- t[15517] = 1
      "000001" when "0011110010011110", -- t[15518] = 1
      "000001" when "0011110010011111", -- t[15519] = 1
      "000001" when "0011110010100000", -- t[15520] = 1
      "000001" when "0011110010100001", -- t[15521] = 1
      "000001" when "0011110010100010", -- t[15522] = 1
      "000001" when "0011110010100011", -- t[15523] = 1
      "000001" when "0011110010100100", -- t[15524] = 1
      "000001" when "0011110010100101", -- t[15525] = 1
      "000001" when "0011110010100110", -- t[15526] = 1
      "000001" when "0011110010100111", -- t[15527] = 1
      "000001" when "0011110010101000", -- t[15528] = 1
      "000001" when "0011110010101001", -- t[15529] = 1
      "000001" when "0011110010101010", -- t[15530] = 1
      "000001" when "0011110010101011", -- t[15531] = 1
      "000001" when "0011110010101100", -- t[15532] = 1
      "000001" when "0011110010101101", -- t[15533] = 1
      "000001" when "0011110010101110", -- t[15534] = 1
      "000001" when "0011110010101111", -- t[15535] = 1
      "000001" when "0011110010110000", -- t[15536] = 1
      "000001" when "0011110010110001", -- t[15537] = 1
      "000001" when "0011110010110010", -- t[15538] = 1
      "000001" when "0011110010110011", -- t[15539] = 1
      "000001" when "0011110010110100", -- t[15540] = 1
      "000001" when "0011110010110101", -- t[15541] = 1
      "000001" when "0011110010110110", -- t[15542] = 1
      "000001" when "0011110010110111", -- t[15543] = 1
      "000001" when "0011110010111000", -- t[15544] = 1
      "000001" when "0011110010111001", -- t[15545] = 1
      "000001" when "0011110010111010", -- t[15546] = 1
      "000001" when "0011110010111011", -- t[15547] = 1
      "000001" when "0011110010111100", -- t[15548] = 1
      "000001" when "0011110010111101", -- t[15549] = 1
      "000001" when "0011110010111110", -- t[15550] = 1
      "000001" when "0011110010111111", -- t[15551] = 1
      "000001" when "0011110011000000", -- t[15552] = 1
      "000001" when "0011110011000001", -- t[15553] = 1
      "000001" when "0011110011000010", -- t[15554] = 1
      "000001" when "0011110011000011", -- t[15555] = 1
      "000001" when "0011110011000100", -- t[15556] = 1
      "000001" when "0011110011000101", -- t[15557] = 1
      "000001" when "0011110011000110", -- t[15558] = 1
      "000001" when "0011110011000111", -- t[15559] = 1
      "000001" when "0011110011001000", -- t[15560] = 1
      "000001" when "0011110011001001", -- t[15561] = 1
      "000001" when "0011110011001010", -- t[15562] = 1
      "000001" when "0011110011001011", -- t[15563] = 1
      "000001" when "0011110011001100", -- t[15564] = 1
      "000001" when "0011110011001101", -- t[15565] = 1
      "000001" when "0011110011001110", -- t[15566] = 1
      "000001" when "0011110011001111", -- t[15567] = 1
      "000001" when "0011110011010000", -- t[15568] = 1
      "000001" when "0011110011010001", -- t[15569] = 1
      "000001" when "0011110011010010", -- t[15570] = 1
      "000001" when "0011110011010011", -- t[15571] = 1
      "000001" when "0011110011010100", -- t[15572] = 1
      "000001" when "0011110011010101", -- t[15573] = 1
      "000001" when "0011110011010110", -- t[15574] = 1
      "000001" when "0011110011010111", -- t[15575] = 1
      "000001" when "0011110011011000", -- t[15576] = 1
      "000001" when "0011110011011001", -- t[15577] = 1
      "000001" when "0011110011011010", -- t[15578] = 1
      "000001" when "0011110011011011", -- t[15579] = 1
      "000001" when "0011110011011100", -- t[15580] = 1
      "000001" when "0011110011011101", -- t[15581] = 1
      "000001" when "0011110011011110", -- t[15582] = 1
      "000001" when "0011110011011111", -- t[15583] = 1
      "000001" when "0011110011100000", -- t[15584] = 1
      "000001" when "0011110011100001", -- t[15585] = 1
      "000001" when "0011110011100010", -- t[15586] = 1
      "000001" when "0011110011100011", -- t[15587] = 1
      "000001" when "0011110011100100", -- t[15588] = 1
      "000001" when "0011110011100101", -- t[15589] = 1
      "000001" when "0011110011100110", -- t[15590] = 1
      "000001" when "0011110011100111", -- t[15591] = 1
      "000001" when "0011110011101000", -- t[15592] = 1
      "000001" when "0011110011101001", -- t[15593] = 1
      "000001" when "0011110011101010", -- t[15594] = 1
      "000001" when "0011110011101011", -- t[15595] = 1
      "000001" when "0011110011101100", -- t[15596] = 1
      "000001" when "0011110011101101", -- t[15597] = 1
      "000001" when "0011110011101110", -- t[15598] = 1
      "000001" when "0011110011101111", -- t[15599] = 1
      "000001" when "0011110011110000", -- t[15600] = 1
      "000001" when "0011110011110001", -- t[15601] = 1
      "000001" when "0011110011110010", -- t[15602] = 1
      "000001" when "0011110011110011", -- t[15603] = 1
      "000001" when "0011110011110100", -- t[15604] = 1
      "000001" when "0011110011110101", -- t[15605] = 1
      "000001" when "0011110011110110", -- t[15606] = 1
      "000001" when "0011110011110111", -- t[15607] = 1
      "000001" when "0011110011111000", -- t[15608] = 1
      "000001" when "0011110011111001", -- t[15609] = 1
      "000001" when "0011110011111010", -- t[15610] = 1
      "000001" when "0011110011111011", -- t[15611] = 1
      "000001" when "0011110011111100", -- t[15612] = 1
      "000001" when "0011110011111101", -- t[15613] = 1
      "000001" when "0011110011111110", -- t[15614] = 1
      "000001" when "0011110011111111", -- t[15615] = 1
      "000001" when "0011110100000000", -- t[15616] = 1
      "000001" when "0011110100000001", -- t[15617] = 1
      "000001" when "0011110100000010", -- t[15618] = 1
      "000001" when "0011110100000011", -- t[15619] = 1
      "000001" when "0011110100000100", -- t[15620] = 1
      "000001" when "0011110100000101", -- t[15621] = 1
      "000001" when "0011110100000110", -- t[15622] = 1
      "000001" when "0011110100000111", -- t[15623] = 1
      "000001" when "0011110100001000", -- t[15624] = 1
      "000001" when "0011110100001001", -- t[15625] = 1
      "000001" when "0011110100001010", -- t[15626] = 1
      "000001" when "0011110100001011", -- t[15627] = 1
      "000001" when "0011110100001100", -- t[15628] = 1
      "000001" when "0011110100001101", -- t[15629] = 1
      "000001" when "0011110100001110", -- t[15630] = 1
      "000001" when "0011110100001111", -- t[15631] = 1
      "000001" when "0011110100010000", -- t[15632] = 1
      "000001" when "0011110100010001", -- t[15633] = 1
      "000001" when "0011110100010010", -- t[15634] = 1
      "000001" when "0011110100010011", -- t[15635] = 1
      "000001" when "0011110100010100", -- t[15636] = 1
      "000001" when "0011110100010101", -- t[15637] = 1
      "000001" when "0011110100010110", -- t[15638] = 1
      "000001" when "0011110100010111", -- t[15639] = 1
      "000001" when "0011110100011000", -- t[15640] = 1
      "000001" when "0011110100011001", -- t[15641] = 1
      "000001" when "0011110100011010", -- t[15642] = 1
      "000001" when "0011110100011011", -- t[15643] = 1
      "000001" when "0011110100011100", -- t[15644] = 1
      "000001" when "0011110100011101", -- t[15645] = 1
      "000001" when "0011110100011110", -- t[15646] = 1
      "000001" when "0011110100011111", -- t[15647] = 1
      "000001" when "0011110100100000", -- t[15648] = 1
      "000001" when "0011110100100001", -- t[15649] = 1
      "000001" when "0011110100100010", -- t[15650] = 1
      "000001" when "0011110100100011", -- t[15651] = 1
      "000001" when "0011110100100100", -- t[15652] = 1
      "000001" when "0011110100100101", -- t[15653] = 1
      "000001" when "0011110100100110", -- t[15654] = 1
      "000001" when "0011110100100111", -- t[15655] = 1
      "000001" when "0011110100101000", -- t[15656] = 1
      "000001" when "0011110100101001", -- t[15657] = 1
      "000001" when "0011110100101010", -- t[15658] = 1
      "000001" when "0011110100101011", -- t[15659] = 1
      "000001" when "0011110100101100", -- t[15660] = 1
      "000001" when "0011110100101101", -- t[15661] = 1
      "000001" when "0011110100101110", -- t[15662] = 1
      "000001" when "0011110100101111", -- t[15663] = 1
      "000001" when "0011110100110000", -- t[15664] = 1
      "000001" when "0011110100110001", -- t[15665] = 1
      "000001" when "0011110100110010", -- t[15666] = 1
      "000001" when "0011110100110011", -- t[15667] = 1
      "000001" when "0011110100110100", -- t[15668] = 1
      "000001" when "0011110100110101", -- t[15669] = 1
      "000001" when "0011110100110110", -- t[15670] = 1
      "000001" when "0011110100110111", -- t[15671] = 1
      "000001" when "0011110100111000", -- t[15672] = 1
      "000001" when "0011110100111001", -- t[15673] = 1
      "000001" when "0011110100111010", -- t[15674] = 1
      "000001" when "0011110100111011", -- t[15675] = 1
      "000001" when "0011110100111100", -- t[15676] = 1
      "000001" when "0011110100111101", -- t[15677] = 1
      "000001" when "0011110100111110", -- t[15678] = 1
      "000001" when "0011110100111111", -- t[15679] = 1
      "000001" when "0011110101000000", -- t[15680] = 1
      "000001" when "0011110101000001", -- t[15681] = 1
      "000001" when "0011110101000010", -- t[15682] = 1
      "000001" when "0011110101000011", -- t[15683] = 1
      "000001" when "0011110101000100", -- t[15684] = 1
      "000001" when "0011110101000101", -- t[15685] = 1
      "000001" when "0011110101000110", -- t[15686] = 1
      "000001" when "0011110101000111", -- t[15687] = 1
      "000001" when "0011110101001000", -- t[15688] = 1
      "000001" when "0011110101001001", -- t[15689] = 1
      "000001" when "0011110101001010", -- t[15690] = 1
      "000001" when "0011110101001011", -- t[15691] = 1
      "000001" when "0011110101001100", -- t[15692] = 1
      "000001" when "0011110101001101", -- t[15693] = 1
      "000001" when "0011110101001110", -- t[15694] = 1
      "000001" when "0011110101001111", -- t[15695] = 1
      "000001" when "0011110101010000", -- t[15696] = 1
      "000001" when "0011110101010001", -- t[15697] = 1
      "000001" when "0011110101010010", -- t[15698] = 1
      "000001" when "0011110101010011", -- t[15699] = 1
      "000001" when "0011110101010100", -- t[15700] = 1
      "000001" when "0011110101010101", -- t[15701] = 1
      "000001" when "0011110101010110", -- t[15702] = 1
      "000001" when "0011110101010111", -- t[15703] = 1
      "000001" when "0011110101011000", -- t[15704] = 1
      "000001" when "0011110101011001", -- t[15705] = 1
      "000001" when "0011110101011010", -- t[15706] = 1
      "000001" when "0011110101011011", -- t[15707] = 1
      "000001" when "0011110101011100", -- t[15708] = 1
      "000001" when "0011110101011101", -- t[15709] = 1
      "000001" when "0011110101011110", -- t[15710] = 1
      "000001" when "0011110101011111", -- t[15711] = 1
      "000001" when "0011110101100000", -- t[15712] = 1
      "000001" when "0011110101100001", -- t[15713] = 1
      "000001" when "0011110101100010", -- t[15714] = 1
      "000001" when "0011110101100011", -- t[15715] = 1
      "000001" when "0011110101100100", -- t[15716] = 1
      "000001" when "0011110101100101", -- t[15717] = 1
      "000001" when "0011110101100110", -- t[15718] = 1
      "000001" when "0011110101100111", -- t[15719] = 1
      "000001" when "0011110101101000", -- t[15720] = 1
      "000001" when "0011110101101001", -- t[15721] = 1
      "000001" when "0011110101101010", -- t[15722] = 1
      "000001" when "0011110101101011", -- t[15723] = 1
      "000001" when "0011110101101100", -- t[15724] = 1
      "000001" when "0011110101101101", -- t[15725] = 1
      "000001" when "0011110101101110", -- t[15726] = 1
      "000001" when "0011110101101111", -- t[15727] = 1
      "000001" when "0011110101110000", -- t[15728] = 1
      "000001" when "0011110101110001", -- t[15729] = 1
      "000001" when "0011110101110010", -- t[15730] = 1
      "000001" when "0011110101110011", -- t[15731] = 1
      "000001" when "0011110101110100", -- t[15732] = 1
      "000001" when "0011110101110101", -- t[15733] = 1
      "000001" when "0011110101110110", -- t[15734] = 1
      "000001" when "0011110101110111", -- t[15735] = 1
      "000001" when "0011110101111000", -- t[15736] = 1
      "000001" when "0011110101111001", -- t[15737] = 1
      "000001" when "0011110101111010", -- t[15738] = 1
      "000001" when "0011110101111011", -- t[15739] = 1
      "000001" when "0011110101111100", -- t[15740] = 1
      "000001" when "0011110101111101", -- t[15741] = 1
      "000001" when "0011110101111110", -- t[15742] = 1
      "000001" when "0011110101111111", -- t[15743] = 1
      "000001" when "0011110110000000", -- t[15744] = 1
      "000001" when "0011110110000001", -- t[15745] = 1
      "000001" when "0011110110000010", -- t[15746] = 1
      "000001" when "0011110110000011", -- t[15747] = 1
      "000001" when "0011110110000100", -- t[15748] = 1
      "000001" when "0011110110000101", -- t[15749] = 1
      "000001" when "0011110110000110", -- t[15750] = 1
      "000001" when "0011110110000111", -- t[15751] = 1
      "000001" when "0011110110001000", -- t[15752] = 1
      "000001" when "0011110110001001", -- t[15753] = 1
      "000001" when "0011110110001010", -- t[15754] = 1
      "000001" when "0011110110001011", -- t[15755] = 1
      "000001" when "0011110110001100", -- t[15756] = 1
      "000001" when "0011110110001101", -- t[15757] = 1
      "000001" when "0011110110001110", -- t[15758] = 1
      "000001" when "0011110110001111", -- t[15759] = 1
      "000001" when "0011110110010000", -- t[15760] = 1
      "000001" when "0011110110010001", -- t[15761] = 1
      "000001" when "0011110110010010", -- t[15762] = 1
      "000001" when "0011110110010011", -- t[15763] = 1
      "000001" when "0011110110010100", -- t[15764] = 1
      "000001" when "0011110110010101", -- t[15765] = 1
      "000001" when "0011110110010110", -- t[15766] = 1
      "000001" when "0011110110010111", -- t[15767] = 1
      "000001" when "0011110110011000", -- t[15768] = 1
      "000001" when "0011110110011001", -- t[15769] = 1
      "000001" when "0011110110011010", -- t[15770] = 1
      "000001" when "0011110110011011", -- t[15771] = 1
      "000001" when "0011110110011100", -- t[15772] = 1
      "000001" when "0011110110011101", -- t[15773] = 1
      "000001" when "0011110110011110", -- t[15774] = 1
      "000001" when "0011110110011111", -- t[15775] = 1
      "000001" when "0011110110100000", -- t[15776] = 1
      "000001" when "0011110110100001", -- t[15777] = 1
      "000001" when "0011110110100010", -- t[15778] = 1
      "000001" when "0011110110100011", -- t[15779] = 1
      "000001" when "0011110110100100", -- t[15780] = 1
      "000001" when "0011110110100101", -- t[15781] = 1
      "000001" when "0011110110100110", -- t[15782] = 1
      "000001" when "0011110110100111", -- t[15783] = 1
      "000001" when "0011110110101000", -- t[15784] = 1
      "000001" when "0011110110101001", -- t[15785] = 1
      "000001" when "0011110110101010", -- t[15786] = 1
      "000001" when "0011110110101011", -- t[15787] = 1
      "000001" when "0011110110101100", -- t[15788] = 1
      "000001" when "0011110110101101", -- t[15789] = 1
      "000001" when "0011110110101110", -- t[15790] = 1
      "000001" when "0011110110101111", -- t[15791] = 1
      "000001" when "0011110110110000", -- t[15792] = 1
      "000001" when "0011110110110001", -- t[15793] = 1
      "000001" when "0011110110110010", -- t[15794] = 1
      "000001" when "0011110110110011", -- t[15795] = 1
      "000001" when "0011110110110100", -- t[15796] = 1
      "000001" when "0011110110110101", -- t[15797] = 1
      "000001" when "0011110110110110", -- t[15798] = 1
      "000001" when "0011110110110111", -- t[15799] = 1
      "000001" when "0011110110111000", -- t[15800] = 1
      "000001" when "0011110110111001", -- t[15801] = 1
      "000001" when "0011110110111010", -- t[15802] = 1
      "000001" when "0011110110111011", -- t[15803] = 1
      "000001" when "0011110110111100", -- t[15804] = 1
      "000001" when "0011110110111101", -- t[15805] = 1
      "000001" when "0011110110111110", -- t[15806] = 1
      "000001" when "0011110110111111", -- t[15807] = 1
      "000001" when "0011110111000000", -- t[15808] = 1
      "000001" when "0011110111000001", -- t[15809] = 1
      "000001" when "0011110111000010", -- t[15810] = 1
      "000001" when "0011110111000011", -- t[15811] = 1
      "000001" when "0011110111000100", -- t[15812] = 1
      "000001" when "0011110111000101", -- t[15813] = 1
      "000001" when "0011110111000110", -- t[15814] = 1
      "000001" when "0011110111000111", -- t[15815] = 1
      "000001" when "0011110111001000", -- t[15816] = 1
      "000001" when "0011110111001001", -- t[15817] = 1
      "000001" when "0011110111001010", -- t[15818] = 1
      "000001" when "0011110111001011", -- t[15819] = 1
      "000001" when "0011110111001100", -- t[15820] = 1
      "000001" when "0011110111001101", -- t[15821] = 1
      "000001" when "0011110111001110", -- t[15822] = 1
      "000001" when "0011110111001111", -- t[15823] = 1
      "000001" when "0011110111010000", -- t[15824] = 1
      "000001" when "0011110111010001", -- t[15825] = 1
      "000001" when "0011110111010010", -- t[15826] = 1
      "000001" when "0011110111010011", -- t[15827] = 1
      "000001" when "0011110111010100", -- t[15828] = 1
      "000001" when "0011110111010101", -- t[15829] = 1
      "000001" when "0011110111010110", -- t[15830] = 1
      "000001" when "0011110111010111", -- t[15831] = 1
      "000001" when "0011110111011000", -- t[15832] = 1
      "000001" when "0011110111011001", -- t[15833] = 1
      "000001" when "0011110111011010", -- t[15834] = 1
      "000001" when "0011110111011011", -- t[15835] = 1
      "000001" when "0011110111011100", -- t[15836] = 1
      "000001" when "0011110111011101", -- t[15837] = 1
      "000001" when "0011110111011110", -- t[15838] = 1
      "000001" when "0011110111011111", -- t[15839] = 1
      "000001" when "0011110111100000", -- t[15840] = 1
      "000001" when "0011110111100001", -- t[15841] = 1
      "000001" when "0011110111100010", -- t[15842] = 1
      "000001" when "0011110111100011", -- t[15843] = 1
      "000001" when "0011110111100100", -- t[15844] = 1
      "000001" when "0011110111100101", -- t[15845] = 1
      "000001" when "0011110111100110", -- t[15846] = 1
      "000001" when "0011110111100111", -- t[15847] = 1
      "000001" when "0011110111101000", -- t[15848] = 1
      "000001" when "0011110111101001", -- t[15849] = 1
      "000001" when "0011110111101010", -- t[15850] = 1
      "000001" when "0011110111101011", -- t[15851] = 1
      "000001" when "0011110111101100", -- t[15852] = 1
      "000001" when "0011110111101101", -- t[15853] = 1
      "000001" when "0011110111101110", -- t[15854] = 1
      "000001" when "0011110111101111", -- t[15855] = 1
      "000001" when "0011110111110000", -- t[15856] = 1
      "000001" when "0011110111110001", -- t[15857] = 1
      "000001" when "0011110111110010", -- t[15858] = 1
      "000001" when "0011110111110011", -- t[15859] = 1
      "000001" when "0011110111110100", -- t[15860] = 1
      "000001" when "0011110111110101", -- t[15861] = 1
      "000001" when "0011110111110110", -- t[15862] = 1
      "000001" when "0011110111110111", -- t[15863] = 1
      "000001" when "0011110111111000", -- t[15864] = 1
      "000001" when "0011110111111001", -- t[15865] = 1
      "000001" when "0011110111111010", -- t[15866] = 1
      "000001" when "0011110111111011", -- t[15867] = 1
      "000001" when "0011110111111100", -- t[15868] = 1
      "000001" when "0011110111111101", -- t[15869] = 1
      "000001" when "0011110111111110", -- t[15870] = 1
      "000001" when "0011110111111111", -- t[15871] = 1
      "000001" when "0011111000000000", -- t[15872] = 1
      "000001" when "0011111000000001", -- t[15873] = 1
      "000001" when "0011111000000010", -- t[15874] = 1
      "000001" when "0011111000000011", -- t[15875] = 1
      "000001" when "0011111000000100", -- t[15876] = 1
      "000001" when "0011111000000101", -- t[15877] = 1
      "000001" when "0011111000000110", -- t[15878] = 1
      "000001" when "0011111000000111", -- t[15879] = 1
      "000001" when "0011111000001000", -- t[15880] = 1
      "000001" when "0011111000001001", -- t[15881] = 1
      "000001" when "0011111000001010", -- t[15882] = 1
      "000001" when "0011111000001011", -- t[15883] = 1
      "000001" when "0011111000001100", -- t[15884] = 1
      "000001" when "0011111000001101", -- t[15885] = 1
      "000001" when "0011111000001110", -- t[15886] = 1
      "000001" when "0011111000001111", -- t[15887] = 1
      "000001" when "0011111000010000", -- t[15888] = 1
      "000001" when "0011111000010001", -- t[15889] = 1
      "000001" when "0011111000010010", -- t[15890] = 1
      "000001" when "0011111000010011", -- t[15891] = 1
      "000001" when "0011111000010100", -- t[15892] = 1
      "000001" when "0011111000010101", -- t[15893] = 1
      "000001" when "0011111000010110", -- t[15894] = 1
      "000001" when "0011111000010111", -- t[15895] = 1
      "000001" when "0011111000011000", -- t[15896] = 1
      "000001" when "0011111000011001", -- t[15897] = 1
      "000001" when "0011111000011010", -- t[15898] = 1
      "000001" when "0011111000011011", -- t[15899] = 1
      "000001" when "0011111000011100", -- t[15900] = 1
      "000001" when "0011111000011101", -- t[15901] = 1
      "000001" when "0011111000011110", -- t[15902] = 1
      "000001" when "0011111000011111", -- t[15903] = 1
      "000001" when "0011111000100000", -- t[15904] = 1
      "000001" when "0011111000100001", -- t[15905] = 1
      "000001" when "0011111000100010", -- t[15906] = 1
      "000001" when "0011111000100011", -- t[15907] = 1
      "000001" when "0011111000100100", -- t[15908] = 1
      "000001" when "0011111000100101", -- t[15909] = 1
      "000001" when "0011111000100110", -- t[15910] = 1
      "000001" when "0011111000100111", -- t[15911] = 1
      "000001" when "0011111000101000", -- t[15912] = 1
      "000001" when "0011111000101001", -- t[15913] = 1
      "000001" when "0011111000101010", -- t[15914] = 1
      "000001" when "0011111000101011", -- t[15915] = 1
      "000001" when "0011111000101100", -- t[15916] = 1
      "000001" when "0011111000101101", -- t[15917] = 1
      "000001" when "0011111000101110", -- t[15918] = 1
      "000001" when "0011111000101111", -- t[15919] = 1
      "000001" when "0011111000110000", -- t[15920] = 1
      "000001" when "0011111000110001", -- t[15921] = 1
      "000001" when "0011111000110010", -- t[15922] = 1
      "000001" when "0011111000110011", -- t[15923] = 1
      "000001" when "0011111000110100", -- t[15924] = 1
      "000001" when "0011111000110101", -- t[15925] = 1
      "000001" when "0011111000110110", -- t[15926] = 1
      "000001" when "0011111000110111", -- t[15927] = 1
      "000001" when "0011111000111000", -- t[15928] = 1
      "000001" when "0011111000111001", -- t[15929] = 1
      "000001" when "0011111000111010", -- t[15930] = 1
      "000001" when "0011111000111011", -- t[15931] = 1
      "000001" when "0011111000111100", -- t[15932] = 1
      "000001" when "0011111000111101", -- t[15933] = 1
      "000001" when "0011111000111110", -- t[15934] = 1
      "000001" when "0011111000111111", -- t[15935] = 1
      "000001" when "0011111001000000", -- t[15936] = 1
      "000001" when "0011111001000001", -- t[15937] = 1
      "000001" when "0011111001000010", -- t[15938] = 1
      "000001" when "0011111001000011", -- t[15939] = 1
      "000001" when "0011111001000100", -- t[15940] = 1
      "000001" when "0011111001000101", -- t[15941] = 1
      "000001" when "0011111001000110", -- t[15942] = 1
      "000001" when "0011111001000111", -- t[15943] = 1
      "000001" when "0011111001001000", -- t[15944] = 1
      "000001" when "0011111001001001", -- t[15945] = 1
      "000001" when "0011111001001010", -- t[15946] = 1
      "000001" when "0011111001001011", -- t[15947] = 1
      "000001" when "0011111001001100", -- t[15948] = 1
      "000001" when "0011111001001101", -- t[15949] = 1
      "000001" when "0011111001001110", -- t[15950] = 1
      "000001" when "0011111001001111", -- t[15951] = 1
      "000001" when "0011111001010000", -- t[15952] = 1
      "000001" when "0011111001010001", -- t[15953] = 1
      "000001" when "0011111001010010", -- t[15954] = 1
      "000001" when "0011111001010011", -- t[15955] = 1
      "000001" when "0011111001010100", -- t[15956] = 1
      "000001" when "0011111001010101", -- t[15957] = 1
      "000001" when "0011111001010110", -- t[15958] = 1
      "000001" when "0011111001010111", -- t[15959] = 1
      "000001" when "0011111001011000", -- t[15960] = 1
      "000001" when "0011111001011001", -- t[15961] = 1
      "000001" when "0011111001011010", -- t[15962] = 1
      "000001" when "0011111001011011", -- t[15963] = 1
      "000001" when "0011111001011100", -- t[15964] = 1
      "000001" when "0011111001011101", -- t[15965] = 1
      "000001" when "0011111001011110", -- t[15966] = 1
      "000001" when "0011111001011111", -- t[15967] = 1
      "000001" when "0011111001100000", -- t[15968] = 1
      "000001" when "0011111001100001", -- t[15969] = 1
      "000001" when "0011111001100010", -- t[15970] = 1
      "000001" when "0011111001100011", -- t[15971] = 1
      "000001" when "0011111001100100", -- t[15972] = 1
      "000001" when "0011111001100101", -- t[15973] = 1
      "000001" when "0011111001100110", -- t[15974] = 1
      "000001" when "0011111001100111", -- t[15975] = 1
      "000001" when "0011111001101000", -- t[15976] = 1
      "000001" when "0011111001101001", -- t[15977] = 1
      "000001" when "0011111001101010", -- t[15978] = 1
      "000001" when "0011111001101011", -- t[15979] = 1
      "000001" when "0011111001101100", -- t[15980] = 1
      "000001" when "0011111001101101", -- t[15981] = 1
      "000001" when "0011111001101110", -- t[15982] = 1
      "000001" when "0011111001101111", -- t[15983] = 1
      "000001" when "0011111001110000", -- t[15984] = 1
      "000001" when "0011111001110001", -- t[15985] = 1
      "000001" when "0011111001110010", -- t[15986] = 1
      "000001" when "0011111001110011", -- t[15987] = 1
      "000001" when "0011111001110100", -- t[15988] = 1
      "000001" when "0011111001110101", -- t[15989] = 1
      "000001" when "0011111001110110", -- t[15990] = 1
      "000001" when "0011111001110111", -- t[15991] = 1
      "000001" when "0011111001111000", -- t[15992] = 1
      "000001" when "0011111001111001", -- t[15993] = 1
      "000001" when "0011111001111010", -- t[15994] = 1
      "000001" when "0011111001111011", -- t[15995] = 1
      "000001" when "0011111001111100", -- t[15996] = 1
      "000001" when "0011111001111101", -- t[15997] = 1
      "000001" when "0011111001111110", -- t[15998] = 1
      "000001" when "0011111001111111", -- t[15999] = 1
      "000001" when "0011111010000000", -- t[16000] = 1
      "000001" when "0011111010000001", -- t[16001] = 1
      "000001" when "0011111010000010", -- t[16002] = 1
      "000001" when "0011111010000011", -- t[16003] = 1
      "000001" when "0011111010000100", -- t[16004] = 1
      "000001" when "0011111010000101", -- t[16005] = 1
      "000001" when "0011111010000110", -- t[16006] = 1
      "000001" when "0011111010000111", -- t[16007] = 1
      "000001" when "0011111010001000", -- t[16008] = 1
      "000001" when "0011111010001001", -- t[16009] = 1
      "000001" when "0011111010001010", -- t[16010] = 1
      "000001" when "0011111010001011", -- t[16011] = 1
      "000001" when "0011111010001100", -- t[16012] = 1
      "000001" when "0011111010001101", -- t[16013] = 1
      "000001" when "0011111010001110", -- t[16014] = 1
      "000001" when "0011111010001111", -- t[16015] = 1
      "000001" when "0011111010010000", -- t[16016] = 1
      "000001" when "0011111010010001", -- t[16017] = 1
      "000001" when "0011111010010010", -- t[16018] = 1
      "000001" when "0011111010010011", -- t[16019] = 1
      "000001" when "0011111010010100", -- t[16020] = 1
      "000001" when "0011111010010101", -- t[16021] = 1
      "000001" when "0011111010010110", -- t[16022] = 1
      "000001" when "0011111010010111", -- t[16023] = 1
      "000001" when "0011111010011000", -- t[16024] = 1
      "000001" when "0011111010011001", -- t[16025] = 1
      "000001" when "0011111010011010", -- t[16026] = 1
      "000001" when "0011111010011011", -- t[16027] = 1
      "000001" when "0011111010011100", -- t[16028] = 1
      "000001" when "0011111010011101", -- t[16029] = 1
      "000001" when "0011111010011110", -- t[16030] = 1
      "000001" when "0011111010011111", -- t[16031] = 1
      "000001" when "0011111010100000", -- t[16032] = 1
      "000001" when "0011111010100001", -- t[16033] = 1
      "000001" when "0011111010100010", -- t[16034] = 1
      "000001" when "0011111010100011", -- t[16035] = 1
      "000001" when "0011111010100100", -- t[16036] = 1
      "000001" when "0011111010100101", -- t[16037] = 1
      "000001" when "0011111010100110", -- t[16038] = 1
      "000001" when "0011111010100111", -- t[16039] = 1
      "000001" when "0011111010101000", -- t[16040] = 1
      "000001" when "0011111010101001", -- t[16041] = 1
      "000001" when "0011111010101010", -- t[16042] = 1
      "000001" when "0011111010101011", -- t[16043] = 1
      "000001" when "0011111010101100", -- t[16044] = 1
      "000001" when "0011111010101101", -- t[16045] = 1
      "000001" when "0011111010101110", -- t[16046] = 1
      "000001" when "0011111010101111", -- t[16047] = 1
      "000001" when "0011111010110000", -- t[16048] = 1
      "000001" when "0011111010110001", -- t[16049] = 1
      "000001" when "0011111010110010", -- t[16050] = 1
      "000001" when "0011111010110011", -- t[16051] = 1
      "000001" when "0011111010110100", -- t[16052] = 1
      "000001" when "0011111010110101", -- t[16053] = 1
      "000001" when "0011111010110110", -- t[16054] = 1
      "000001" when "0011111010110111", -- t[16055] = 1
      "000001" when "0011111010111000", -- t[16056] = 1
      "000001" when "0011111010111001", -- t[16057] = 1
      "000001" when "0011111010111010", -- t[16058] = 1
      "000001" when "0011111010111011", -- t[16059] = 1
      "000001" when "0011111010111100", -- t[16060] = 1
      "000001" when "0011111010111101", -- t[16061] = 1
      "000001" when "0011111010111110", -- t[16062] = 1
      "000001" when "0011111010111111", -- t[16063] = 1
      "000001" when "0011111011000000", -- t[16064] = 1
      "000001" when "0011111011000001", -- t[16065] = 1
      "000001" when "0011111011000010", -- t[16066] = 1
      "000001" when "0011111011000011", -- t[16067] = 1
      "000001" when "0011111011000100", -- t[16068] = 1
      "000001" when "0011111011000101", -- t[16069] = 1
      "000001" when "0011111011000110", -- t[16070] = 1
      "000001" when "0011111011000111", -- t[16071] = 1
      "000001" when "0011111011001000", -- t[16072] = 1
      "000001" when "0011111011001001", -- t[16073] = 1
      "000001" when "0011111011001010", -- t[16074] = 1
      "000001" when "0011111011001011", -- t[16075] = 1
      "000001" when "0011111011001100", -- t[16076] = 1
      "000001" when "0011111011001101", -- t[16077] = 1
      "000001" when "0011111011001110", -- t[16078] = 1
      "000001" when "0011111011001111", -- t[16079] = 1
      "000001" when "0011111011010000", -- t[16080] = 1
      "000001" when "0011111011010001", -- t[16081] = 1
      "000001" when "0011111011010010", -- t[16082] = 1
      "000001" when "0011111011010011", -- t[16083] = 1
      "000001" when "0011111011010100", -- t[16084] = 1
      "000001" when "0011111011010101", -- t[16085] = 1
      "000001" when "0011111011010110", -- t[16086] = 1
      "000001" when "0011111011010111", -- t[16087] = 1
      "000001" when "0011111011011000", -- t[16088] = 1
      "000001" when "0011111011011001", -- t[16089] = 1
      "000001" when "0011111011011010", -- t[16090] = 1
      "000001" when "0011111011011011", -- t[16091] = 1
      "000001" when "0011111011011100", -- t[16092] = 1
      "000001" when "0011111011011101", -- t[16093] = 1
      "000001" when "0011111011011110", -- t[16094] = 1
      "000001" when "0011111011011111", -- t[16095] = 1
      "000001" when "0011111011100000", -- t[16096] = 1
      "000001" when "0011111011100001", -- t[16097] = 1
      "000001" when "0011111011100010", -- t[16098] = 1
      "000001" when "0011111011100011", -- t[16099] = 1
      "000001" when "0011111011100100", -- t[16100] = 1
      "000001" when "0011111011100101", -- t[16101] = 1
      "000001" when "0011111011100110", -- t[16102] = 1
      "000001" when "0011111011100111", -- t[16103] = 1
      "000001" when "0011111011101000", -- t[16104] = 1
      "000001" when "0011111011101001", -- t[16105] = 1
      "000001" when "0011111011101010", -- t[16106] = 1
      "000001" when "0011111011101011", -- t[16107] = 1
      "000001" when "0011111011101100", -- t[16108] = 1
      "000001" when "0011111011101101", -- t[16109] = 1
      "000001" when "0011111011101110", -- t[16110] = 1
      "000001" when "0011111011101111", -- t[16111] = 1
      "000001" when "0011111011110000", -- t[16112] = 1
      "000001" when "0011111011110001", -- t[16113] = 1
      "000001" when "0011111011110010", -- t[16114] = 1
      "000001" when "0011111011110011", -- t[16115] = 1
      "000001" when "0011111011110100", -- t[16116] = 1
      "000001" when "0011111011110101", -- t[16117] = 1
      "000001" when "0011111011110110", -- t[16118] = 1
      "000001" when "0011111011110111", -- t[16119] = 1
      "000001" when "0011111011111000", -- t[16120] = 1
      "000001" when "0011111011111001", -- t[16121] = 1
      "000001" when "0011111011111010", -- t[16122] = 1
      "000001" when "0011111011111011", -- t[16123] = 1
      "000001" when "0011111011111100", -- t[16124] = 1
      "000001" when "0011111011111101", -- t[16125] = 1
      "000001" when "0011111011111110", -- t[16126] = 1
      "000001" when "0011111011111111", -- t[16127] = 1
      "000001" when "0011111100000000", -- t[16128] = 1
      "000001" when "0011111100000001", -- t[16129] = 1
      "000001" when "0011111100000010", -- t[16130] = 1
      "000001" when "0011111100000011", -- t[16131] = 1
      "000001" when "0011111100000100", -- t[16132] = 1
      "000001" when "0011111100000101", -- t[16133] = 1
      "000001" when "0011111100000110", -- t[16134] = 1
      "000001" when "0011111100000111", -- t[16135] = 1
      "000001" when "0011111100001000", -- t[16136] = 1
      "000001" when "0011111100001001", -- t[16137] = 1
      "000001" when "0011111100001010", -- t[16138] = 1
      "000001" when "0011111100001011", -- t[16139] = 1
      "000001" when "0011111100001100", -- t[16140] = 1
      "000001" when "0011111100001101", -- t[16141] = 1
      "000001" when "0011111100001110", -- t[16142] = 1
      "000001" when "0011111100001111", -- t[16143] = 1
      "000001" when "0011111100010000", -- t[16144] = 1
      "000001" when "0011111100010001", -- t[16145] = 1
      "000001" when "0011111100010010", -- t[16146] = 1
      "000001" when "0011111100010011", -- t[16147] = 1
      "000001" when "0011111100010100", -- t[16148] = 1
      "000001" when "0011111100010101", -- t[16149] = 1
      "000001" when "0011111100010110", -- t[16150] = 1
      "000001" when "0011111100010111", -- t[16151] = 1
      "000001" when "0011111100011000", -- t[16152] = 1
      "000001" when "0011111100011001", -- t[16153] = 1
      "000001" when "0011111100011010", -- t[16154] = 1
      "000001" when "0011111100011011", -- t[16155] = 1
      "000001" when "0011111100011100", -- t[16156] = 1
      "000001" when "0011111100011101", -- t[16157] = 1
      "000001" when "0011111100011110", -- t[16158] = 1
      "000001" when "0011111100011111", -- t[16159] = 1
      "000001" when "0011111100100000", -- t[16160] = 1
      "000001" when "0011111100100001", -- t[16161] = 1
      "000001" when "0011111100100010", -- t[16162] = 1
      "000001" when "0011111100100011", -- t[16163] = 1
      "000001" when "0011111100100100", -- t[16164] = 1
      "000001" when "0011111100100101", -- t[16165] = 1
      "000001" when "0011111100100110", -- t[16166] = 1
      "000001" when "0011111100100111", -- t[16167] = 1
      "000001" when "0011111100101000", -- t[16168] = 1
      "000001" when "0011111100101001", -- t[16169] = 1
      "000001" when "0011111100101010", -- t[16170] = 1
      "000001" when "0011111100101011", -- t[16171] = 1
      "000001" when "0011111100101100", -- t[16172] = 1
      "000001" when "0011111100101101", -- t[16173] = 1
      "000001" when "0011111100101110", -- t[16174] = 1
      "000001" when "0011111100101111", -- t[16175] = 1
      "000001" when "0011111100110000", -- t[16176] = 1
      "000001" when "0011111100110001", -- t[16177] = 1
      "000001" when "0011111100110010", -- t[16178] = 1
      "000001" when "0011111100110011", -- t[16179] = 1
      "000001" when "0011111100110100", -- t[16180] = 1
      "000001" when "0011111100110101", -- t[16181] = 1
      "000001" when "0011111100110110", -- t[16182] = 1
      "000001" when "0011111100110111", -- t[16183] = 1
      "000001" when "0011111100111000", -- t[16184] = 1
      "000001" when "0011111100111001", -- t[16185] = 1
      "000001" when "0011111100111010", -- t[16186] = 1
      "000001" when "0011111100111011", -- t[16187] = 1
      "000001" when "0011111100111100", -- t[16188] = 1
      "000001" when "0011111100111101", -- t[16189] = 1
      "000001" when "0011111100111110", -- t[16190] = 1
      "000001" when "0011111100111111", -- t[16191] = 1
      "000001" when "0011111101000000", -- t[16192] = 1
      "000001" when "0011111101000001", -- t[16193] = 1
      "000001" when "0011111101000010", -- t[16194] = 1
      "000001" when "0011111101000011", -- t[16195] = 1
      "000001" when "0011111101000100", -- t[16196] = 1
      "000001" when "0011111101000101", -- t[16197] = 1
      "000001" when "0011111101000110", -- t[16198] = 1
      "000001" when "0011111101000111", -- t[16199] = 1
      "000001" when "0011111101001000", -- t[16200] = 1
      "000001" when "0011111101001001", -- t[16201] = 1
      "000001" when "0011111101001010", -- t[16202] = 1
      "000001" when "0011111101001011", -- t[16203] = 1
      "000001" when "0011111101001100", -- t[16204] = 1
      "000001" when "0011111101001101", -- t[16205] = 1
      "000001" when "0011111101001110", -- t[16206] = 1
      "000001" when "0011111101001111", -- t[16207] = 1
      "000001" when "0011111101010000", -- t[16208] = 1
      "000001" when "0011111101010001", -- t[16209] = 1
      "000001" when "0011111101010010", -- t[16210] = 1
      "000001" when "0011111101010011", -- t[16211] = 1
      "000001" when "0011111101010100", -- t[16212] = 1
      "000001" when "0011111101010101", -- t[16213] = 1
      "000001" when "0011111101010110", -- t[16214] = 1
      "000001" when "0011111101010111", -- t[16215] = 1
      "000001" when "0011111101011000", -- t[16216] = 1
      "000001" when "0011111101011001", -- t[16217] = 1
      "000001" when "0011111101011010", -- t[16218] = 1
      "000001" when "0011111101011011", -- t[16219] = 1
      "000001" when "0011111101011100", -- t[16220] = 1
      "000001" when "0011111101011101", -- t[16221] = 1
      "000001" when "0011111101011110", -- t[16222] = 1
      "000001" when "0011111101011111", -- t[16223] = 1
      "000001" when "0011111101100000", -- t[16224] = 1
      "000001" when "0011111101100001", -- t[16225] = 1
      "000001" when "0011111101100010", -- t[16226] = 1
      "000001" when "0011111101100011", -- t[16227] = 1
      "000001" when "0011111101100100", -- t[16228] = 1
      "000001" when "0011111101100101", -- t[16229] = 1
      "000001" when "0011111101100110", -- t[16230] = 1
      "000001" when "0011111101100111", -- t[16231] = 1
      "000001" when "0011111101101000", -- t[16232] = 1
      "000001" when "0011111101101001", -- t[16233] = 1
      "000001" when "0011111101101010", -- t[16234] = 1
      "000001" when "0011111101101011", -- t[16235] = 1
      "000001" when "0011111101101100", -- t[16236] = 1
      "000001" when "0011111101101101", -- t[16237] = 1
      "000001" when "0011111101101110", -- t[16238] = 1
      "000001" when "0011111101101111", -- t[16239] = 1
      "000001" when "0011111101110000", -- t[16240] = 1
      "000001" when "0011111101110001", -- t[16241] = 1
      "000001" when "0011111101110010", -- t[16242] = 1
      "000001" when "0011111101110011", -- t[16243] = 1
      "000001" when "0011111101110100", -- t[16244] = 1
      "000001" when "0011111101110101", -- t[16245] = 1
      "000001" when "0011111101110110", -- t[16246] = 1
      "000001" when "0011111101110111", -- t[16247] = 1
      "000001" when "0011111101111000", -- t[16248] = 1
      "000001" when "0011111101111001", -- t[16249] = 1
      "000001" when "0011111101111010", -- t[16250] = 1
      "000001" when "0011111101111011", -- t[16251] = 1
      "000001" when "0011111101111100", -- t[16252] = 1
      "000001" when "0011111101111101", -- t[16253] = 1
      "000001" when "0011111101111110", -- t[16254] = 1
      "000001" when "0011111101111111", -- t[16255] = 1
      "000001" when "0011111110000000", -- t[16256] = 1
      "000001" when "0011111110000001", -- t[16257] = 1
      "000001" when "0011111110000010", -- t[16258] = 1
      "000001" when "0011111110000011", -- t[16259] = 1
      "000001" when "0011111110000100", -- t[16260] = 1
      "000001" when "0011111110000101", -- t[16261] = 1
      "000001" when "0011111110000110", -- t[16262] = 1
      "000001" when "0011111110000111", -- t[16263] = 1
      "000001" when "0011111110001000", -- t[16264] = 1
      "000001" when "0011111110001001", -- t[16265] = 1
      "000001" when "0011111110001010", -- t[16266] = 1
      "000001" when "0011111110001011", -- t[16267] = 1
      "000001" when "0011111110001100", -- t[16268] = 1
      "000001" when "0011111110001101", -- t[16269] = 1
      "000001" when "0011111110001110", -- t[16270] = 1
      "000001" when "0011111110001111", -- t[16271] = 1
      "000001" when "0011111110010000", -- t[16272] = 1
      "000001" when "0011111110010001", -- t[16273] = 1
      "000001" when "0011111110010010", -- t[16274] = 1
      "000001" when "0011111110010011", -- t[16275] = 1
      "000001" when "0011111110010100", -- t[16276] = 1
      "000001" when "0011111110010101", -- t[16277] = 1
      "000001" when "0011111110010110", -- t[16278] = 1
      "000001" when "0011111110010111", -- t[16279] = 1
      "000001" when "0011111110011000", -- t[16280] = 1
      "000001" when "0011111110011001", -- t[16281] = 1
      "000001" when "0011111110011010", -- t[16282] = 1
      "000001" when "0011111110011011", -- t[16283] = 1
      "000001" when "0011111110011100", -- t[16284] = 1
      "000001" when "0011111110011101", -- t[16285] = 1
      "000001" when "0011111110011110", -- t[16286] = 1
      "000001" when "0011111110011111", -- t[16287] = 1
      "000001" when "0011111110100000", -- t[16288] = 1
      "000001" when "0011111110100001", -- t[16289] = 1
      "000001" when "0011111110100010", -- t[16290] = 1
      "000001" when "0011111110100011", -- t[16291] = 1
      "000001" when "0011111110100100", -- t[16292] = 1
      "000001" when "0011111110100101", -- t[16293] = 1
      "000001" when "0011111110100110", -- t[16294] = 1
      "000001" when "0011111110100111", -- t[16295] = 1
      "000001" when "0011111110101000", -- t[16296] = 1
      "000001" when "0011111110101001", -- t[16297] = 1
      "000001" when "0011111110101010", -- t[16298] = 1
      "000001" when "0011111110101011", -- t[16299] = 1
      "000001" when "0011111110101100", -- t[16300] = 1
      "000001" when "0011111110101101", -- t[16301] = 1
      "000001" when "0011111110101110", -- t[16302] = 1
      "000001" when "0011111110101111", -- t[16303] = 1
      "000001" when "0011111110110000", -- t[16304] = 1
      "000001" when "0011111110110001", -- t[16305] = 1
      "000001" when "0011111110110010", -- t[16306] = 1
      "000001" when "0011111110110011", -- t[16307] = 1
      "000001" when "0011111110110100", -- t[16308] = 1
      "000001" when "0011111110110101", -- t[16309] = 1
      "000001" when "0011111110110110", -- t[16310] = 1
      "000001" when "0011111110110111", -- t[16311] = 1
      "000001" when "0011111110111000", -- t[16312] = 1
      "000001" when "0011111110111001", -- t[16313] = 1
      "000001" when "0011111110111010", -- t[16314] = 1
      "000001" when "0011111110111011", -- t[16315] = 1
      "000001" when "0011111110111100", -- t[16316] = 1
      "000001" when "0011111110111101", -- t[16317] = 1
      "000001" when "0011111110111110", -- t[16318] = 1
      "000001" when "0011111110111111", -- t[16319] = 1
      "000001" when "0011111111000000", -- t[16320] = 1
      "000001" when "0011111111000001", -- t[16321] = 1
      "000001" when "0011111111000010", -- t[16322] = 1
      "000001" when "0011111111000011", -- t[16323] = 1
      "000001" when "0011111111000100", -- t[16324] = 1
      "000001" when "0011111111000101", -- t[16325] = 1
      "000001" when "0011111111000110", -- t[16326] = 1
      "000001" when "0011111111000111", -- t[16327] = 1
      "000001" when "0011111111001000", -- t[16328] = 1
      "000001" when "0011111111001001", -- t[16329] = 1
      "000001" when "0011111111001010", -- t[16330] = 1
      "000001" when "0011111111001011", -- t[16331] = 1
      "000001" when "0011111111001100", -- t[16332] = 1
      "000001" when "0011111111001101", -- t[16333] = 1
      "000001" when "0011111111001110", -- t[16334] = 1
      "000001" when "0011111111001111", -- t[16335] = 1
      "000001" when "0011111111010000", -- t[16336] = 1
      "000001" when "0011111111010001", -- t[16337] = 1
      "000001" when "0011111111010010", -- t[16338] = 1
      "000001" when "0011111111010011", -- t[16339] = 1
      "000001" when "0011111111010100", -- t[16340] = 1
      "000001" when "0011111111010101", -- t[16341] = 1
      "000001" when "0011111111010110", -- t[16342] = 1
      "000001" when "0011111111010111", -- t[16343] = 1
      "000001" when "0011111111011000", -- t[16344] = 1
      "000001" when "0011111111011001", -- t[16345] = 1
      "000001" when "0011111111011010", -- t[16346] = 1
      "000001" when "0011111111011011", -- t[16347] = 1
      "000001" when "0011111111011100", -- t[16348] = 1
      "000001" when "0011111111011101", -- t[16349] = 1
      "000001" when "0011111111011110", -- t[16350] = 1
      "000001" when "0011111111011111", -- t[16351] = 1
      "000001" when "0011111111100000", -- t[16352] = 1
      "000001" when "0011111111100001", -- t[16353] = 1
      "000001" when "0011111111100010", -- t[16354] = 1
      "000001" when "0011111111100011", -- t[16355] = 1
      "000001" when "0011111111100100", -- t[16356] = 1
      "000001" when "0011111111100101", -- t[16357] = 1
      "000001" when "0011111111100110", -- t[16358] = 1
      "000001" when "0011111111100111", -- t[16359] = 1
      "000001" when "0011111111101000", -- t[16360] = 1
      "000001" when "0011111111101001", -- t[16361] = 1
      "000001" when "0011111111101010", -- t[16362] = 1
      "000001" when "0011111111101011", -- t[16363] = 1
      "000001" when "0011111111101100", -- t[16364] = 1
      "000001" when "0011111111101101", -- t[16365] = 1
      "000001" when "0011111111101110", -- t[16366] = 1
      "000001" when "0011111111101111", -- t[16367] = 1
      "000001" when "0011111111110000", -- t[16368] = 1
      "000001" when "0011111111110001", -- t[16369] = 1
      "000001" when "0011111111110010", -- t[16370] = 1
      "000001" when "0011111111110011", -- t[16371] = 1
      "000001" when "0011111111110100", -- t[16372] = 1
      "000001" when "0011111111110101", -- t[16373] = 1
      "000001" when "0011111111110110", -- t[16374] = 1
      "000001" when "0011111111110111", -- t[16375] = 1
      "000001" when "0011111111111000", -- t[16376] = 1
      "000001" when "0011111111111001", -- t[16377] = 1
      "000001" when "0011111111111010", -- t[16378] = 1
      "000001" when "0011111111111011", -- t[16379] = 1
      "000001" when "0011111111111100", -- t[16380] = 1
      "000001" when "0011111111111101", -- t[16381] = 1
      "000001" when "0011111111111110", -- t[16382] = 1
      "000001" when "0011111111111111", -- t[16383] = 1
      "000001" when "0100000000000000", -- t[16384] = 1
      "000001" when "0100000000000001", -- t[16385] = 1
      "000001" when "0100000000000010", -- t[16386] = 1
      "000001" when "0100000000000011", -- t[16387] = 1
      "000001" when "0100000000000100", -- t[16388] = 1
      "000001" when "0100000000000101", -- t[16389] = 1
      "000001" when "0100000000000110", -- t[16390] = 1
      "000001" when "0100000000000111", -- t[16391] = 1
      "000001" when "0100000000001000", -- t[16392] = 1
      "000001" when "0100000000001001", -- t[16393] = 1
      "000001" when "0100000000001010", -- t[16394] = 1
      "000001" when "0100000000001011", -- t[16395] = 1
      "000001" when "0100000000001100", -- t[16396] = 1
      "000001" when "0100000000001101", -- t[16397] = 1
      "000001" when "0100000000001110", -- t[16398] = 1
      "000001" when "0100000000001111", -- t[16399] = 1
      "000001" when "0100000000010000", -- t[16400] = 1
      "000001" when "0100000000010001", -- t[16401] = 1
      "000001" when "0100000000010010", -- t[16402] = 1
      "000001" when "0100000000010011", -- t[16403] = 1
      "000001" when "0100000000010100", -- t[16404] = 1
      "000001" when "0100000000010101", -- t[16405] = 1
      "000001" when "0100000000010110", -- t[16406] = 1
      "000001" when "0100000000010111", -- t[16407] = 1
      "000001" when "0100000000011000", -- t[16408] = 1
      "000001" when "0100000000011001", -- t[16409] = 1
      "000001" when "0100000000011010", -- t[16410] = 1
      "000001" when "0100000000011011", -- t[16411] = 1
      "000001" when "0100000000011100", -- t[16412] = 1
      "000001" when "0100000000011101", -- t[16413] = 1
      "000001" when "0100000000011110", -- t[16414] = 1
      "000001" when "0100000000011111", -- t[16415] = 1
      "000001" when "0100000000100000", -- t[16416] = 1
      "000001" when "0100000000100001", -- t[16417] = 1
      "000001" when "0100000000100010", -- t[16418] = 1
      "000001" when "0100000000100011", -- t[16419] = 1
      "000001" when "0100000000100100", -- t[16420] = 1
      "000001" when "0100000000100101", -- t[16421] = 1
      "000001" when "0100000000100110", -- t[16422] = 1
      "000001" when "0100000000100111", -- t[16423] = 1
      "000001" when "0100000000101000", -- t[16424] = 1
      "000001" when "0100000000101001", -- t[16425] = 1
      "000001" when "0100000000101010", -- t[16426] = 1
      "000001" when "0100000000101011", -- t[16427] = 1
      "000001" when "0100000000101100", -- t[16428] = 1
      "000001" when "0100000000101101", -- t[16429] = 1
      "000001" when "0100000000101110", -- t[16430] = 1
      "000001" when "0100000000101111", -- t[16431] = 1
      "000001" when "0100000000110000", -- t[16432] = 1
      "000001" when "0100000000110001", -- t[16433] = 1
      "000001" when "0100000000110010", -- t[16434] = 1
      "000001" when "0100000000110011", -- t[16435] = 1
      "000001" when "0100000000110100", -- t[16436] = 1
      "000001" when "0100000000110101", -- t[16437] = 1
      "000001" when "0100000000110110", -- t[16438] = 1
      "000001" when "0100000000110111", -- t[16439] = 1
      "000001" when "0100000000111000", -- t[16440] = 1
      "000001" when "0100000000111001", -- t[16441] = 1
      "000001" when "0100000000111010", -- t[16442] = 1
      "000001" when "0100000000111011", -- t[16443] = 1
      "000001" when "0100000000111100", -- t[16444] = 1
      "000001" when "0100000000111101", -- t[16445] = 1
      "000001" when "0100000000111110", -- t[16446] = 1
      "000001" when "0100000000111111", -- t[16447] = 1
      "000001" when "0100000001000000", -- t[16448] = 1
      "000001" when "0100000001000001", -- t[16449] = 1
      "000001" when "0100000001000010", -- t[16450] = 1
      "000001" when "0100000001000011", -- t[16451] = 1
      "000001" when "0100000001000100", -- t[16452] = 1
      "000001" when "0100000001000101", -- t[16453] = 1
      "000001" when "0100000001000110", -- t[16454] = 1
      "000001" when "0100000001000111", -- t[16455] = 1
      "000001" when "0100000001001000", -- t[16456] = 1
      "000001" when "0100000001001001", -- t[16457] = 1
      "000001" when "0100000001001010", -- t[16458] = 1
      "000001" when "0100000001001011", -- t[16459] = 1
      "000001" when "0100000001001100", -- t[16460] = 1
      "000001" when "0100000001001101", -- t[16461] = 1
      "000001" when "0100000001001110", -- t[16462] = 1
      "000001" when "0100000001001111", -- t[16463] = 1
      "000001" when "0100000001010000", -- t[16464] = 1
      "000001" when "0100000001010001", -- t[16465] = 1
      "000001" when "0100000001010010", -- t[16466] = 1
      "000001" when "0100000001010011", -- t[16467] = 1
      "000001" when "0100000001010100", -- t[16468] = 1
      "000001" when "0100000001010101", -- t[16469] = 1
      "000001" when "0100000001010110", -- t[16470] = 1
      "000001" when "0100000001010111", -- t[16471] = 1
      "000001" when "0100000001011000", -- t[16472] = 1
      "000001" when "0100000001011001", -- t[16473] = 1
      "000001" when "0100000001011010", -- t[16474] = 1
      "000001" when "0100000001011011", -- t[16475] = 1
      "000001" when "0100000001011100", -- t[16476] = 1
      "000001" when "0100000001011101", -- t[16477] = 1
      "000001" when "0100000001011110", -- t[16478] = 1
      "000001" when "0100000001011111", -- t[16479] = 1
      "000001" when "0100000001100000", -- t[16480] = 1
      "000001" when "0100000001100001", -- t[16481] = 1
      "000001" when "0100000001100010", -- t[16482] = 1
      "000001" when "0100000001100011", -- t[16483] = 1
      "000001" when "0100000001100100", -- t[16484] = 1
      "000001" when "0100000001100101", -- t[16485] = 1
      "000001" when "0100000001100110", -- t[16486] = 1
      "000001" when "0100000001100111", -- t[16487] = 1
      "000001" when "0100000001101000", -- t[16488] = 1
      "000001" when "0100000001101001", -- t[16489] = 1
      "000001" when "0100000001101010", -- t[16490] = 1
      "000001" when "0100000001101011", -- t[16491] = 1
      "000001" when "0100000001101100", -- t[16492] = 1
      "000001" when "0100000001101101", -- t[16493] = 1
      "000001" when "0100000001101110", -- t[16494] = 1
      "000001" when "0100000001101111", -- t[16495] = 1
      "000001" when "0100000001110000", -- t[16496] = 1
      "000001" when "0100000001110001", -- t[16497] = 1
      "000001" when "0100000001110010", -- t[16498] = 1
      "000001" when "0100000001110011", -- t[16499] = 1
      "000001" when "0100000001110100", -- t[16500] = 1
      "000001" when "0100000001110101", -- t[16501] = 1
      "000001" when "0100000001110110", -- t[16502] = 1
      "000001" when "0100000001110111", -- t[16503] = 1
      "000001" when "0100000001111000", -- t[16504] = 1
      "000001" when "0100000001111001", -- t[16505] = 1
      "000001" when "0100000001111010", -- t[16506] = 1
      "000001" when "0100000001111011", -- t[16507] = 1
      "000001" when "0100000001111100", -- t[16508] = 1
      "000001" when "0100000001111101", -- t[16509] = 1
      "000001" when "0100000001111110", -- t[16510] = 1
      "000001" when "0100000001111111", -- t[16511] = 1
      "000001" when "0100000010000000", -- t[16512] = 1
      "000001" when "0100000010000001", -- t[16513] = 1
      "000001" when "0100000010000010", -- t[16514] = 1
      "000001" when "0100000010000011", -- t[16515] = 1
      "000001" when "0100000010000100", -- t[16516] = 1
      "000001" when "0100000010000101", -- t[16517] = 1
      "000001" when "0100000010000110", -- t[16518] = 1
      "000001" when "0100000010000111", -- t[16519] = 1
      "000001" when "0100000010001000", -- t[16520] = 1
      "000001" when "0100000010001001", -- t[16521] = 1
      "000001" when "0100000010001010", -- t[16522] = 1
      "000001" when "0100000010001011", -- t[16523] = 1
      "000001" when "0100000010001100", -- t[16524] = 1
      "000001" when "0100000010001101", -- t[16525] = 1
      "000001" when "0100000010001110", -- t[16526] = 1
      "000001" when "0100000010001111", -- t[16527] = 1
      "000001" when "0100000010010000", -- t[16528] = 1
      "000001" when "0100000010010001", -- t[16529] = 1
      "000001" when "0100000010010010", -- t[16530] = 1
      "000001" when "0100000010010011", -- t[16531] = 1
      "000001" when "0100000010010100", -- t[16532] = 1
      "000001" when "0100000010010101", -- t[16533] = 1
      "000001" when "0100000010010110", -- t[16534] = 1
      "000001" when "0100000010010111", -- t[16535] = 1
      "000001" when "0100000010011000", -- t[16536] = 1
      "000001" when "0100000010011001", -- t[16537] = 1
      "000001" when "0100000010011010", -- t[16538] = 1
      "000001" when "0100000010011011", -- t[16539] = 1
      "000001" when "0100000010011100", -- t[16540] = 1
      "000001" when "0100000010011101", -- t[16541] = 1
      "000001" when "0100000010011110", -- t[16542] = 1
      "000001" when "0100000010011111", -- t[16543] = 1
      "000001" when "0100000010100000", -- t[16544] = 1
      "000001" when "0100000010100001", -- t[16545] = 1
      "000001" when "0100000010100010", -- t[16546] = 1
      "000001" when "0100000010100011", -- t[16547] = 1
      "000001" when "0100000010100100", -- t[16548] = 1
      "000001" when "0100000010100101", -- t[16549] = 1
      "000001" when "0100000010100110", -- t[16550] = 1
      "000001" when "0100000010100111", -- t[16551] = 1
      "000001" when "0100000010101000", -- t[16552] = 1
      "000001" when "0100000010101001", -- t[16553] = 1
      "000001" when "0100000010101010", -- t[16554] = 1
      "000001" when "0100000010101011", -- t[16555] = 1
      "000001" when "0100000010101100", -- t[16556] = 1
      "000001" when "0100000010101101", -- t[16557] = 1
      "000001" when "0100000010101110", -- t[16558] = 1
      "000001" when "0100000010101111", -- t[16559] = 1
      "000001" when "0100000010110000", -- t[16560] = 1
      "000001" when "0100000010110001", -- t[16561] = 1
      "000001" when "0100000010110010", -- t[16562] = 1
      "000001" when "0100000010110011", -- t[16563] = 1
      "000001" when "0100000010110100", -- t[16564] = 1
      "000001" when "0100000010110101", -- t[16565] = 1
      "000001" when "0100000010110110", -- t[16566] = 1
      "000001" when "0100000010110111", -- t[16567] = 1
      "000001" when "0100000010111000", -- t[16568] = 1
      "000001" when "0100000010111001", -- t[16569] = 1
      "000001" when "0100000010111010", -- t[16570] = 1
      "000001" when "0100000010111011", -- t[16571] = 1
      "000001" when "0100000010111100", -- t[16572] = 1
      "000001" when "0100000010111101", -- t[16573] = 1
      "000001" when "0100000010111110", -- t[16574] = 1
      "000001" when "0100000010111111", -- t[16575] = 1
      "000001" when "0100000011000000", -- t[16576] = 1
      "000001" when "0100000011000001", -- t[16577] = 1
      "000001" when "0100000011000010", -- t[16578] = 1
      "000001" when "0100000011000011", -- t[16579] = 1
      "000001" when "0100000011000100", -- t[16580] = 1
      "000001" when "0100000011000101", -- t[16581] = 1
      "000001" when "0100000011000110", -- t[16582] = 1
      "000001" when "0100000011000111", -- t[16583] = 1
      "000001" when "0100000011001000", -- t[16584] = 1
      "000001" when "0100000011001001", -- t[16585] = 1
      "000001" when "0100000011001010", -- t[16586] = 1
      "000001" when "0100000011001011", -- t[16587] = 1
      "000001" when "0100000011001100", -- t[16588] = 1
      "000001" when "0100000011001101", -- t[16589] = 1
      "000001" when "0100000011001110", -- t[16590] = 1
      "000001" when "0100000011001111", -- t[16591] = 1
      "000001" when "0100000011010000", -- t[16592] = 1
      "000001" when "0100000011010001", -- t[16593] = 1
      "000001" when "0100000011010010", -- t[16594] = 1
      "000001" when "0100000011010011", -- t[16595] = 1
      "000001" when "0100000011010100", -- t[16596] = 1
      "000001" when "0100000011010101", -- t[16597] = 1
      "000001" when "0100000011010110", -- t[16598] = 1
      "000001" when "0100000011010111", -- t[16599] = 1
      "000001" when "0100000011011000", -- t[16600] = 1
      "000001" when "0100000011011001", -- t[16601] = 1
      "000001" when "0100000011011010", -- t[16602] = 1
      "000001" when "0100000011011011", -- t[16603] = 1
      "000001" when "0100000011011100", -- t[16604] = 1
      "000001" when "0100000011011101", -- t[16605] = 1
      "000001" when "0100000011011110", -- t[16606] = 1
      "000001" when "0100000011011111", -- t[16607] = 1
      "000001" when "0100000011100000", -- t[16608] = 1
      "000001" when "0100000011100001", -- t[16609] = 1
      "000001" when "0100000011100010", -- t[16610] = 1
      "000001" when "0100000011100011", -- t[16611] = 1
      "000001" when "0100000011100100", -- t[16612] = 1
      "000001" when "0100000011100101", -- t[16613] = 1
      "000010" when "0100000011100110", -- t[16614] = 2
      "000010" when "0100000011100111", -- t[16615] = 2
      "000010" when "0100000011101000", -- t[16616] = 2
      "000010" when "0100000011101001", -- t[16617] = 2
      "000010" when "0100000011101010", -- t[16618] = 2
      "000010" when "0100000011101011", -- t[16619] = 2
      "000010" when "0100000011101100", -- t[16620] = 2
      "000010" when "0100000011101101", -- t[16621] = 2
      "000010" when "0100000011101110", -- t[16622] = 2
      "000010" when "0100000011101111", -- t[16623] = 2
      "000010" when "0100000011110000", -- t[16624] = 2
      "000010" when "0100000011110001", -- t[16625] = 2
      "000010" when "0100000011110010", -- t[16626] = 2
      "000010" when "0100000011110011", -- t[16627] = 2
      "000010" when "0100000011110100", -- t[16628] = 2
      "000010" when "0100000011110101", -- t[16629] = 2
      "000010" when "0100000011110110", -- t[16630] = 2
      "000010" when "0100000011110111", -- t[16631] = 2
      "000010" when "0100000011111000", -- t[16632] = 2
      "000010" when "0100000011111001", -- t[16633] = 2
      "000010" when "0100000011111010", -- t[16634] = 2
      "000010" when "0100000011111011", -- t[16635] = 2
      "000010" when "0100000011111100", -- t[16636] = 2
      "000010" when "0100000011111101", -- t[16637] = 2
      "000010" when "0100000011111110", -- t[16638] = 2
      "000010" when "0100000011111111", -- t[16639] = 2
      "000010" when "0100000100000000", -- t[16640] = 2
      "000010" when "0100000100000001", -- t[16641] = 2
      "000010" when "0100000100000010", -- t[16642] = 2
      "000010" when "0100000100000011", -- t[16643] = 2
      "000010" when "0100000100000100", -- t[16644] = 2
      "000010" when "0100000100000101", -- t[16645] = 2
      "000010" when "0100000100000110", -- t[16646] = 2
      "000010" when "0100000100000111", -- t[16647] = 2
      "000010" when "0100000100001000", -- t[16648] = 2
      "000010" when "0100000100001001", -- t[16649] = 2
      "000010" when "0100000100001010", -- t[16650] = 2
      "000010" when "0100000100001011", -- t[16651] = 2
      "000010" when "0100000100001100", -- t[16652] = 2
      "000010" when "0100000100001101", -- t[16653] = 2
      "000010" when "0100000100001110", -- t[16654] = 2
      "000010" when "0100000100001111", -- t[16655] = 2
      "000010" when "0100000100010000", -- t[16656] = 2
      "000010" when "0100000100010001", -- t[16657] = 2
      "000010" when "0100000100010010", -- t[16658] = 2
      "000010" when "0100000100010011", -- t[16659] = 2
      "000010" when "0100000100010100", -- t[16660] = 2
      "000010" when "0100000100010101", -- t[16661] = 2
      "000010" when "0100000100010110", -- t[16662] = 2
      "000010" when "0100000100010111", -- t[16663] = 2
      "000010" when "0100000100011000", -- t[16664] = 2
      "000010" when "0100000100011001", -- t[16665] = 2
      "000010" when "0100000100011010", -- t[16666] = 2
      "000010" when "0100000100011011", -- t[16667] = 2
      "000010" when "0100000100011100", -- t[16668] = 2
      "000010" when "0100000100011101", -- t[16669] = 2
      "000010" when "0100000100011110", -- t[16670] = 2
      "000010" when "0100000100011111", -- t[16671] = 2
      "000010" when "0100000100100000", -- t[16672] = 2
      "000010" when "0100000100100001", -- t[16673] = 2
      "000010" when "0100000100100010", -- t[16674] = 2
      "000010" when "0100000100100011", -- t[16675] = 2
      "000010" when "0100000100100100", -- t[16676] = 2
      "000010" when "0100000100100101", -- t[16677] = 2
      "000010" when "0100000100100110", -- t[16678] = 2
      "000010" when "0100000100100111", -- t[16679] = 2
      "000010" when "0100000100101000", -- t[16680] = 2
      "000010" when "0100000100101001", -- t[16681] = 2
      "000010" when "0100000100101010", -- t[16682] = 2
      "000010" when "0100000100101011", -- t[16683] = 2
      "000010" when "0100000100101100", -- t[16684] = 2
      "000010" when "0100000100101101", -- t[16685] = 2
      "000010" when "0100000100101110", -- t[16686] = 2
      "000010" when "0100000100101111", -- t[16687] = 2
      "000010" when "0100000100110000", -- t[16688] = 2
      "000010" when "0100000100110001", -- t[16689] = 2
      "000010" when "0100000100110010", -- t[16690] = 2
      "000010" when "0100000100110011", -- t[16691] = 2
      "000010" when "0100000100110100", -- t[16692] = 2
      "000010" when "0100000100110101", -- t[16693] = 2
      "000010" when "0100000100110110", -- t[16694] = 2
      "000010" when "0100000100110111", -- t[16695] = 2
      "000010" when "0100000100111000", -- t[16696] = 2
      "000010" when "0100000100111001", -- t[16697] = 2
      "000010" when "0100000100111010", -- t[16698] = 2
      "000010" when "0100000100111011", -- t[16699] = 2
      "000010" when "0100000100111100", -- t[16700] = 2
      "000010" when "0100000100111101", -- t[16701] = 2
      "000010" when "0100000100111110", -- t[16702] = 2
      "000010" when "0100000100111111", -- t[16703] = 2
      "000010" when "0100000101000000", -- t[16704] = 2
      "000010" when "0100000101000001", -- t[16705] = 2
      "000010" when "0100000101000010", -- t[16706] = 2
      "000010" when "0100000101000011", -- t[16707] = 2
      "000010" when "0100000101000100", -- t[16708] = 2
      "000010" when "0100000101000101", -- t[16709] = 2
      "000010" when "0100000101000110", -- t[16710] = 2
      "000010" when "0100000101000111", -- t[16711] = 2
      "000010" when "0100000101001000", -- t[16712] = 2
      "000010" when "0100000101001001", -- t[16713] = 2
      "000010" when "0100000101001010", -- t[16714] = 2
      "000010" when "0100000101001011", -- t[16715] = 2
      "000010" when "0100000101001100", -- t[16716] = 2
      "000010" when "0100000101001101", -- t[16717] = 2
      "000010" when "0100000101001110", -- t[16718] = 2
      "000010" when "0100000101001111", -- t[16719] = 2
      "000010" when "0100000101010000", -- t[16720] = 2
      "000010" when "0100000101010001", -- t[16721] = 2
      "000010" when "0100000101010010", -- t[16722] = 2
      "000010" when "0100000101010011", -- t[16723] = 2
      "000010" when "0100000101010100", -- t[16724] = 2
      "000010" when "0100000101010101", -- t[16725] = 2
      "000010" when "0100000101010110", -- t[16726] = 2
      "000010" when "0100000101010111", -- t[16727] = 2
      "000010" when "0100000101011000", -- t[16728] = 2
      "000010" when "0100000101011001", -- t[16729] = 2
      "000010" when "0100000101011010", -- t[16730] = 2
      "000010" when "0100000101011011", -- t[16731] = 2
      "000010" when "0100000101011100", -- t[16732] = 2
      "000010" when "0100000101011101", -- t[16733] = 2
      "000010" when "0100000101011110", -- t[16734] = 2
      "000010" when "0100000101011111", -- t[16735] = 2
      "000010" when "0100000101100000", -- t[16736] = 2
      "000010" when "0100000101100001", -- t[16737] = 2
      "000010" when "0100000101100010", -- t[16738] = 2
      "000010" when "0100000101100011", -- t[16739] = 2
      "000010" when "0100000101100100", -- t[16740] = 2
      "000010" when "0100000101100101", -- t[16741] = 2
      "000010" when "0100000101100110", -- t[16742] = 2
      "000010" when "0100000101100111", -- t[16743] = 2
      "000010" when "0100000101101000", -- t[16744] = 2
      "000010" when "0100000101101001", -- t[16745] = 2
      "000010" when "0100000101101010", -- t[16746] = 2
      "000010" when "0100000101101011", -- t[16747] = 2
      "000010" when "0100000101101100", -- t[16748] = 2
      "000010" when "0100000101101101", -- t[16749] = 2
      "000010" when "0100000101101110", -- t[16750] = 2
      "000010" when "0100000101101111", -- t[16751] = 2
      "000010" when "0100000101110000", -- t[16752] = 2
      "000010" when "0100000101110001", -- t[16753] = 2
      "000010" when "0100000101110010", -- t[16754] = 2
      "000010" when "0100000101110011", -- t[16755] = 2
      "000010" when "0100000101110100", -- t[16756] = 2
      "000010" when "0100000101110101", -- t[16757] = 2
      "000010" when "0100000101110110", -- t[16758] = 2
      "000010" when "0100000101110111", -- t[16759] = 2
      "000010" when "0100000101111000", -- t[16760] = 2
      "000010" when "0100000101111001", -- t[16761] = 2
      "000010" when "0100000101111010", -- t[16762] = 2
      "000010" when "0100000101111011", -- t[16763] = 2
      "000010" when "0100000101111100", -- t[16764] = 2
      "000010" when "0100000101111101", -- t[16765] = 2
      "000010" when "0100000101111110", -- t[16766] = 2
      "000010" when "0100000101111111", -- t[16767] = 2
      "000010" when "0100000110000000", -- t[16768] = 2
      "000010" when "0100000110000001", -- t[16769] = 2
      "000010" when "0100000110000010", -- t[16770] = 2
      "000010" when "0100000110000011", -- t[16771] = 2
      "000010" when "0100000110000100", -- t[16772] = 2
      "000010" when "0100000110000101", -- t[16773] = 2
      "000010" when "0100000110000110", -- t[16774] = 2
      "000010" when "0100000110000111", -- t[16775] = 2
      "000010" when "0100000110001000", -- t[16776] = 2
      "000010" when "0100000110001001", -- t[16777] = 2
      "000010" when "0100000110001010", -- t[16778] = 2
      "000010" when "0100000110001011", -- t[16779] = 2
      "000010" when "0100000110001100", -- t[16780] = 2
      "000010" when "0100000110001101", -- t[16781] = 2
      "000010" when "0100000110001110", -- t[16782] = 2
      "000010" when "0100000110001111", -- t[16783] = 2
      "000010" when "0100000110010000", -- t[16784] = 2
      "000010" when "0100000110010001", -- t[16785] = 2
      "000010" when "0100000110010010", -- t[16786] = 2
      "000010" when "0100000110010011", -- t[16787] = 2
      "000010" when "0100000110010100", -- t[16788] = 2
      "000010" when "0100000110010101", -- t[16789] = 2
      "000010" when "0100000110010110", -- t[16790] = 2
      "000010" when "0100000110010111", -- t[16791] = 2
      "000010" when "0100000110011000", -- t[16792] = 2
      "000010" when "0100000110011001", -- t[16793] = 2
      "000010" when "0100000110011010", -- t[16794] = 2
      "000010" when "0100000110011011", -- t[16795] = 2
      "000010" when "0100000110011100", -- t[16796] = 2
      "000010" when "0100000110011101", -- t[16797] = 2
      "000010" when "0100000110011110", -- t[16798] = 2
      "000010" when "0100000110011111", -- t[16799] = 2
      "000010" when "0100000110100000", -- t[16800] = 2
      "000010" when "0100000110100001", -- t[16801] = 2
      "000010" when "0100000110100010", -- t[16802] = 2
      "000010" when "0100000110100011", -- t[16803] = 2
      "000010" when "0100000110100100", -- t[16804] = 2
      "000010" when "0100000110100101", -- t[16805] = 2
      "000010" when "0100000110100110", -- t[16806] = 2
      "000010" when "0100000110100111", -- t[16807] = 2
      "000010" when "0100000110101000", -- t[16808] = 2
      "000010" when "0100000110101001", -- t[16809] = 2
      "000010" when "0100000110101010", -- t[16810] = 2
      "000010" when "0100000110101011", -- t[16811] = 2
      "000010" when "0100000110101100", -- t[16812] = 2
      "000010" when "0100000110101101", -- t[16813] = 2
      "000010" when "0100000110101110", -- t[16814] = 2
      "000010" when "0100000110101111", -- t[16815] = 2
      "000010" when "0100000110110000", -- t[16816] = 2
      "000010" when "0100000110110001", -- t[16817] = 2
      "000010" when "0100000110110010", -- t[16818] = 2
      "000010" when "0100000110110011", -- t[16819] = 2
      "000010" when "0100000110110100", -- t[16820] = 2
      "000010" when "0100000110110101", -- t[16821] = 2
      "000010" when "0100000110110110", -- t[16822] = 2
      "000010" when "0100000110110111", -- t[16823] = 2
      "000010" when "0100000110111000", -- t[16824] = 2
      "000010" when "0100000110111001", -- t[16825] = 2
      "000010" when "0100000110111010", -- t[16826] = 2
      "000010" when "0100000110111011", -- t[16827] = 2
      "000010" when "0100000110111100", -- t[16828] = 2
      "000010" when "0100000110111101", -- t[16829] = 2
      "000010" when "0100000110111110", -- t[16830] = 2
      "000010" when "0100000110111111", -- t[16831] = 2
      "000010" when "0100000111000000", -- t[16832] = 2
      "000010" when "0100000111000001", -- t[16833] = 2
      "000010" when "0100000111000010", -- t[16834] = 2
      "000010" when "0100000111000011", -- t[16835] = 2
      "000010" when "0100000111000100", -- t[16836] = 2
      "000010" when "0100000111000101", -- t[16837] = 2
      "000010" when "0100000111000110", -- t[16838] = 2
      "000010" when "0100000111000111", -- t[16839] = 2
      "000010" when "0100000111001000", -- t[16840] = 2
      "000010" when "0100000111001001", -- t[16841] = 2
      "000010" when "0100000111001010", -- t[16842] = 2
      "000010" when "0100000111001011", -- t[16843] = 2
      "000010" when "0100000111001100", -- t[16844] = 2
      "000010" when "0100000111001101", -- t[16845] = 2
      "000010" when "0100000111001110", -- t[16846] = 2
      "000010" when "0100000111001111", -- t[16847] = 2
      "000010" when "0100000111010000", -- t[16848] = 2
      "000010" when "0100000111010001", -- t[16849] = 2
      "000010" when "0100000111010010", -- t[16850] = 2
      "000010" when "0100000111010011", -- t[16851] = 2
      "000010" when "0100000111010100", -- t[16852] = 2
      "000010" when "0100000111010101", -- t[16853] = 2
      "000010" when "0100000111010110", -- t[16854] = 2
      "000010" when "0100000111010111", -- t[16855] = 2
      "000010" when "0100000111011000", -- t[16856] = 2
      "000010" when "0100000111011001", -- t[16857] = 2
      "000010" when "0100000111011010", -- t[16858] = 2
      "000010" when "0100000111011011", -- t[16859] = 2
      "000010" when "0100000111011100", -- t[16860] = 2
      "000010" when "0100000111011101", -- t[16861] = 2
      "000010" when "0100000111011110", -- t[16862] = 2
      "000010" when "0100000111011111", -- t[16863] = 2
      "000010" when "0100000111100000", -- t[16864] = 2
      "000010" when "0100000111100001", -- t[16865] = 2
      "000010" when "0100000111100010", -- t[16866] = 2
      "000010" when "0100000111100011", -- t[16867] = 2
      "000010" when "0100000111100100", -- t[16868] = 2
      "000010" when "0100000111100101", -- t[16869] = 2
      "000010" when "0100000111100110", -- t[16870] = 2
      "000010" when "0100000111100111", -- t[16871] = 2
      "000010" when "0100000111101000", -- t[16872] = 2
      "000010" when "0100000111101001", -- t[16873] = 2
      "000010" when "0100000111101010", -- t[16874] = 2
      "000010" when "0100000111101011", -- t[16875] = 2
      "000010" when "0100000111101100", -- t[16876] = 2
      "000010" when "0100000111101101", -- t[16877] = 2
      "000010" when "0100000111101110", -- t[16878] = 2
      "000010" when "0100000111101111", -- t[16879] = 2
      "000010" when "0100000111110000", -- t[16880] = 2
      "000010" when "0100000111110001", -- t[16881] = 2
      "000010" when "0100000111110010", -- t[16882] = 2
      "000010" when "0100000111110011", -- t[16883] = 2
      "000010" when "0100000111110100", -- t[16884] = 2
      "000010" when "0100000111110101", -- t[16885] = 2
      "000010" when "0100000111110110", -- t[16886] = 2
      "000010" when "0100000111110111", -- t[16887] = 2
      "000010" when "0100000111111000", -- t[16888] = 2
      "000010" when "0100000111111001", -- t[16889] = 2
      "000010" when "0100000111111010", -- t[16890] = 2
      "000010" when "0100000111111011", -- t[16891] = 2
      "000010" when "0100000111111100", -- t[16892] = 2
      "000010" when "0100000111111101", -- t[16893] = 2
      "000010" when "0100000111111110", -- t[16894] = 2
      "000010" when "0100000111111111", -- t[16895] = 2
      "000010" when "0100001000000000", -- t[16896] = 2
      "000010" when "0100001000000001", -- t[16897] = 2
      "000010" when "0100001000000010", -- t[16898] = 2
      "000010" when "0100001000000011", -- t[16899] = 2
      "000010" when "0100001000000100", -- t[16900] = 2
      "000010" when "0100001000000101", -- t[16901] = 2
      "000010" when "0100001000000110", -- t[16902] = 2
      "000010" when "0100001000000111", -- t[16903] = 2
      "000010" when "0100001000001000", -- t[16904] = 2
      "000010" when "0100001000001001", -- t[16905] = 2
      "000010" when "0100001000001010", -- t[16906] = 2
      "000010" when "0100001000001011", -- t[16907] = 2
      "000010" when "0100001000001100", -- t[16908] = 2
      "000010" when "0100001000001101", -- t[16909] = 2
      "000010" when "0100001000001110", -- t[16910] = 2
      "000010" when "0100001000001111", -- t[16911] = 2
      "000010" when "0100001000010000", -- t[16912] = 2
      "000010" when "0100001000010001", -- t[16913] = 2
      "000010" when "0100001000010010", -- t[16914] = 2
      "000010" when "0100001000010011", -- t[16915] = 2
      "000010" when "0100001000010100", -- t[16916] = 2
      "000010" when "0100001000010101", -- t[16917] = 2
      "000010" when "0100001000010110", -- t[16918] = 2
      "000010" when "0100001000010111", -- t[16919] = 2
      "000010" when "0100001000011000", -- t[16920] = 2
      "000010" when "0100001000011001", -- t[16921] = 2
      "000010" when "0100001000011010", -- t[16922] = 2
      "000010" when "0100001000011011", -- t[16923] = 2
      "000010" when "0100001000011100", -- t[16924] = 2
      "000010" when "0100001000011101", -- t[16925] = 2
      "000010" when "0100001000011110", -- t[16926] = 2
      "000010" when "0100001000011111", -- t[16927] = 2
      "000010" when "0100001000100000", -- t[16928] = 2
      "000010" when "0100001000100001", -- t[16929] = 2
      "000010" when "0100001000100010", -- t[16930] = 2
      "000010" when "0100001000100011", -- t[16931] = 2
      "000010" when "0100001000100100", -- t[16932] = 2
      "000010" when "0100001000100101", -- t[16933] = 2
      "000010" when "0100001000100110", -- t[16934] = 2
      "000010" when "0100001000100111", -- t[16935] = 2
      "000010" when "0100001000101000", -- t[16936] = 2
      "000010" when "0100001000101001", -- t[16937] = 2
      "000010" when "0100001000101010", -- t[16938] = 2
      "000010" when "0100001000101011", -- t[16939] = 2
      "000010" when "0100001000101100", -- t[16940] = 2
      "000010" when "0100001000101101", -- t[16941] = 2
      "000010" when "0100001000101110", -- t[16942] = 2
      "000010" when "0100001000101111", -- t[16943] = 2
      "000010" when "0100001000110000", -- t[16944] = 2
      "000010" when "0100001000110001", -- t[16945] = 2
      "000010" when "0100001000110010", -- t[16946] = 2
      "000010" when "0100001000110011", -- t[16947] = 2
      "000010" when "0100001000110100", -- t[16948] = 2
      "000010" when "0100001000110101", -- t[16949] = 2
      "000010" when "0100001000110110", -- t[16950] = 2
      "000010" when "0100001000110111", -- t[16951] = 2
      "000010" when "0100001000111000", -- t[16952] = 2
      "000010" when "0100001000111001", -- t[16953] = 2
      "000010" when "0100001000111010", -- t[16954] = 2
      "000010" when "0100001000111011", -- t[16955] = 2
      "000010" when "0100001000111100", -- t[16956] = 2
      "000010" when "0100001000111101", -- t[16957] = 2
      "000010" when "0100001000111110", -- t[16958] = 2
      "000010" when "0100001000111111", -- t[16959] = 2
      "000010" when "0100001001000000", -- t[16960] = 2
      "000010" when "0100001001000001", -- t[16961] = 2
      "000010" when "0100001001000010", -- t[16962] = 2
      "000010" when "0100001001000011", -- t[16963] = 2
      "000010" when "0100001001000100", -- t[16964] = 2
      "000010" when "0100001001000101", -- t[16965] = 2
      "000010" when "0100001001000110", -- t[16966] = 2
      "000010" when "0100001001000111", -- t[16967] = 2
      "000010" when "0100001001001000", -- t[16968] = 2
      "000010" when "0100001001001001", -- t[16969] = 2
      "000010" when "0100001001001010", -- t[16970] = 2
      "000010" when "0100001001001011", -- t[16971] = 2
      "000010" when "0100001001001100", -- t[16972] = 2
      "000010" when "0100001001001101", -- t[16973] = 2
      "000010" when "0100001001001110", -- t[16974] = 2
      "000010" when "0100001001001111", -- t[16975] = 2
      "000010" when "0100001001010000", -- t[16976] = 2
      "000010" when "0100001001010001", -- t[16977] = 2
      "000010" when "0100001001010010", -- t[16978] = 2
      "000010" when "0100001001010011", -- t[16979] = 2
      "000010" when "0100001001010100", -- t[16980] = 2
      "000010" when "0100001001010101", -- t[16981] = 2
      "000010" when "0100001001010110", -- t[16982] = 2
      "000010" when "0100001001010111", -- t[16983] = 2
      "000010" when "0100001001011000", -- t[16984] = 2
      "000010" when "0100001001011001", -- t[16985] = 2
      "000010" when "0100001001011010", -- t[16986] = 2
      "000010" when "0100001001011011", -- t[16987] = 2
      "000010" when "0100001001011100", -- t[16988] = 2
      "000010" when "0100001001011101", -- t[16989] = 2
      "000010" when "0100001001011110", -- t[16990] = 2
      "000010" when "0100001001011111", -- t[16991] = 2
      "000010" when "0100001001100000", -- t[16992] = 2
      "000010" when "0100001001100001", -- t[16993] = 2
      "000010" when "0100001001100010", -- t[16994] = 2
      "000010" when "0100001001100011", -- t[16995] = 2
      "000010" when "0100001001100100", -- t[16996] = 2
      "000010" when "0100001001100101", -- t[16997] = 2
      "000010" when "0100001001100110", -- t[16998] = 2
      "000010" when "0100001001100111", -- t[16999] = 2
      "000010" when "0100001001101000", -- t[17000] = 2
      "000010" when "0100001001101001", -- t[17001] = 2
      "000010" when "0100001001101010", -- t[17002] = 2
      "000010" when "0100001001101011", -- t[17003] = 2
      "000010" when "0100001001101100", -- t[17004] = 2
      "000010" when "0100001001101101", -- t[17005] = 2
      "000010" when "0100001001101110", -- t[17006] = 2
      "000010" when "0100001001101111", -- t[17007] = 2
      "000010" when "0100001001110000", -- t[17008] = 2
      "000010" when "0100001001110001", -- t[17009] = 2
      "000010" when "0100001001110010", -- t[17010] = 2
      "000010" when "0100001001110011", -- t[17011] = 2
      "000010" when "0100001001110100", -- t[17012] = 2
      "000010" when "0100001001110101", -- t[17013] = 2
      "000010" when "0100001001110110", -- t[17014] = 2
      "000010" when "0100001001110111", -- t[17015] = 2
      "000010" when "0100001001111000", -- t[17016] = 2
      "000010" when "0100001001111001", -- t[17017] = 2
      "000010" when "0100001001111010", -- t[17018] = 2
      "000010" when "0100001001111011", -- t[17019] = 2
      "000010" when "0100001001111100", -- t[17020] = 2
      "000010" when "0100001001111101", -- t[17021] = 2
      "000010" when "0100001001111110", -- t[17022] = 2
      "000010" when "0100001001111111", -- t[17023] = 2
      "000010" when "0100001010000000", -- t[17024] = 2
      "000010" when "0100001010000001", -- t[17025] = 2
      "000010" when "0100001010000010", -- t[17026] = 2
      "000010" when "0100001010000011", -- t[17027] = 2
      "000010" when "0100001010000100", -- t[17028] = 2
      "000010" when "0100001010000101", -- t[17029] = 2
      "000010" when "0100001010000110", -- t[17030] = 2
      "000010" when "0100001010000111", -- t[17031] = 2
      "000010" when "0100001010001000", -- t[17032] = 2
      "000010" when "0100001010001001", -- t[17033] = 2
      "000010" when "0100001010001010", -- t[17034] = 2
      "000010" when "0100001010001011", -- t[17035] = 2
      "000010" when "0100001010001100", -- t[17036] = 2
      "000010" when "0100001010001101", -- t[17037] = 2
      "000010" when "0100001010001110", -- t[17038] = 2
      "000010" when "0100001010001111", -- t[17039] = 2
      "000010" when "0100001010010000", -- t[17040] = 2
      "000010" when "0100001010010001", -- t[17041] = 2
      "000010" when "0100001010010010", -- t[17042] = 2
      "000010" when "0100001010010011", -- t[17043] = 2
      "000010" when "0100001010010100", -- t[17044] = 2
      "000010" when "0100001010010101", -- t[17045] = 2
      "000010" when "0100001010010110", -- t[17046] = 2
      "000010" when "0100001010010111", -- t[17047] = 2
      "000010" when "0100001010011000", -- t[17048] = 2
      "000010" when "0100001010011001", -- t[17049] = 2
      "000010" when "0100001010011010", -- t[17050] = 2
      "000010" when "0100001010011011", -- t[17051] = 2
      "000010" when "0100001010011100", -- t[17052] = 2
      "000010" when "0100001010011101", -- t[17053] = 2
      "000010" when "0100001010011110", -- t[17054] = 2
      "000010" when "0100001010011111", -- t[17055] = 2
      "000010" when "0100001010100000", -- t[17056] = 2
      "000010" when "0100001010100001", -- t[17057] = 2
      "000010" when "0100001010100010", -- t[17058] = 2
      "000010" when "0100001010100011", -- t[17059] = 2
      "000010" when "0100001010100100", -- t[17060] = 2
      "000010" when "0100001010100101", -- t[17061] = 2
      "000010" when "0100001010100110", -- t[17062] = 2
      "000010" when "0100001010100111", -- t[17063] = 2
      "000010" when "0100001010101000", -- t[17064] = 2
      "000010" when "0100001010101001", -- t[17065] = 2
      "000010" when "0100001010101010", -- t[17066] = 2
      "000010" when "0100001010101011", -- t[17067] = 2
      "000010" when "0100001010101100", -- t[17068] = 2
      "000010" when "0100001010101101", -- t[17069] = 2
      "000010" when "0100001010101110", -- t[17070] = 2
      "000010" when "0100001010101111", -- t[17071] = 2
      "000010" when "0100001010110000", -- t[17072] = 2
      "000010" when "0100001010110001", -- t[17073] = 2
      "000010" when "0100001010110010", -- t[17074] = 2
      "000010" when "0100001010110011", -- t[17075] = 2
      "000010" when "0100001010110100", -- t[17076] = 2
      "000010" when "0100001010110101", -- t[17077] = 2
      "000010" when "0100001010110110", -- t[17078] = 2
      "000010" when "0100001010110111", -- t[17079] = 2
      "000010" when "0100001010111000", -- t[17080] = 2
      "000010" when "0100001010111001", -- t[17081] = 2
      "000010" when "0100001010111010", -- t[17082] = 2
      "000010" when "0100001010111011", -- t[17083] = 2
      "000010" when "0100001010111100", -- t[17084] = 2
      "000010" when "0100001010111101", -- t[17085] = 2
      "000010" when "0100001010111110", -- t[17086] = 2
      "000010" when "0100001010111111", -- t[17087] = 2
      "000010" when "0100001011000000", -- t[17088] = 2
      "000010" when "0100001011000001", -- t[17089] = 2
      "000010" when "0100001011000010", -- t[17090] = 2
      "000010" when "0100001011000011", -- t[17091] = 2
      "000010" when "0100001011000100", -- t[17092] = 2
      "000010" when "0100001011000101", -- t[17093] = 2
      "000010" when "0100001011000110", -- t[17094] = 2
      "000010" when "0100001011000111", -- t[17095] = 2
      "000010" when "0100001011001000", -- t[17096] = 2
      "000010" when "0100001011001001", -- t[17097] = 2
      "000010" when "0100001011001010", -- t[17098] = 2
      "000010" when "0100001011001011", -- t[17099] = 2
      "000010" when "0100001011001100", -- t[17100] = 2
      "000010" when "0100001011001101", -- t[17101] = 2
      "000010" when "0100001011001110", -- t[17102] = 2
      "000010" when "0100001011001111", -- t[17103] = 2
      "000010" when "0100001011010000", -- t[17104] = 2
      "000010" when "0100001011010001", -- t[17105] = 2
      "000010" when "0100001011010010", -- t[17106] = 2
      "000010" when "0100001011010011", -- t[17107] = 2
      "000010" when "0100001011010100", -- t[17108] = 2
      "000010" when "0100001011010101", -- t[17109] = 2
      "000010" when "0100001011010110", -- t[17110] = 2
      "000010" when "0100001011010111", -- t[17111] = 2
      "000010" when "0100001011011000", -- t[17112] = 2
      "000010" when "0100001011011001", -- t[17113] = 2
      "000010" when "0100001011011010", -- t[17114] = 2
      "000010" when "0100001011011011", -- t[17115] = 2
      "000010" when "0100001011011100", -- t[17116] = 2
      "000010" when "0100001011011101", -- t[17117] = 2
      "000010" when "0100001011011110", -- t[17118] = 2
      "000010" when "0100001011011111", -- t[17119] = 2
      "000010" when "0100001011100000", -- t[17120] = 2
      "000010" when "0100001011100001", -- t[17121] = 2
      "000010" when "0100001011100010", -- t[17122] = 2
      "000010" when "0100001011100011", -- t[17123] = 2
      "000010" when "0100001011100100", -- t[17124] = 2
      "000010" when "0100001011100101", -- t[17125] = 2
      "000010" when "0100001011100110", -- t[17126] = 2
      "000010" when "0100001011100111", -- t[17127] = 2
      "000010" when "0100001011101000", -- t[17128] = 2
      "000010" when "0100001011101001", -- t[17129] = 2
      "000010" when "0100001011101010", -- t[17130] = 2
      "000010" when "0100001011101011", -- t[17131] = 2
      "000010" when "0100001011101100", -- t[17132] = 2
      "000010" when "0100001011101101", -- t[17133] = 2
      "000010" when "0100001011101110", -- t[17134] = 2
      "000010" when "0100001011101111", -- t[17135] = 2
      "000010" when "0100001011110000", -- t[17136] = 2
      "000010" when "0100001011110001", -- t[17137] = 2
      "000010" when "0100001011110010", -- t[17138] = 2
      "000010" when "0100001011110011", -- t[17139] = 2
      "000010" when "0100001011110100", -- t[17140] = 2
      "000010" when "0100001011110101", -- t[17141] = 2
      "000010" when "0100001011110110", -- t[17142] = 2
      "000010" when "0100001011110111", -- t[17143] = 2
      "000010" when "0100001011111000", -- t[17144] = 2
      "000010" when "0100001011111001", -- t[17145] = 2
      "000010" when "0100001011111010", -- t[17146] = 2
      "000010" when "0100001011111011", -- t[17147] = 2
      "000010" when "0100001011111100", -- t[17148] = 2
      "000010" when "0100001011111101", -- t[17149] = 2
      "000010" when "0100001011111110", -- t[17150] = 2
      "000010" when "0100001011111111", -- t[17151] = 2
      "000010" when "0100001100000000", -- t[17152] = 2
      "000010" when "0100001100000001", -- t[17153] = 2
      "000010" when "0100001100000010", -- t[17154] = 2
      "000010" when "0100001100000011", -- t[17155] = 2
      "000010" when "0100001100000100", -- t[17156] = 2
      "000010" when "0100001100000101", -- t[17157] = 2
      "000010" when "0100001100000110", -- t[17158] = 2
      "000010" when "0100001100000111", -- t[17159] = 2
      "000010" when "0100001100001000", -- t[17160] = 2
      "000010" when "0100001100001001", -- t[17161] = 2
      "000010" when "0100001100001010", -- t[17162] = 2
      "000010" when "0100001100001011", -- t[17163] = 2
      "000010" when "0100001100001100", -- t[17164] = 2
      "000010" when "0100001100001101", -- t[17165] = 2
      "000010" when "0100001100001110", -- t[17166] = 2
      "000010" when "0100001100001111", -- t[17167] = 2
      "000010" when "0100001100010000", -- t[17168] = 2
      "000010" when "0100001100010001", -- t[17169] = 2
      "000010" when "0100001100010010", -- t[17170] = 2
      "000010" when "0100001100010011", -- t[17171] = 2
      "000010" when "0100001100010100", -- t[17172] = 2
      "000010" when "0100001100010101", -- t[17173] = 2
      "000010" when "0100001100010110", -- t[17174] = 2
      "000010" when "0100001100010111", -- t[17175] = 2
      "000010" when "0100001100011000", -- t[17176] = 2
      "000010" when "0100001100011001", -- t[17177] = 2
      "000010" when "0100001100011010", -- t[17178] = 2
      "000010" when "0100001100011011", -- t[17179] = 2
      "000010" when "0100001100011100", -- t[17180] = 2
      "000010" when "0100001100011101", -- t[17181] = 2
      "000010" when "0100001100011110", -- t[17182] = 2
      "000010" when "0100001100011111", -- t[17183] = 2
      "000010" when "0100001100100000", -- t[17184] = 2
      "000010" when "0100001100100001", -- t[17185] = 2
      "000010" when "0100001100100010", -- t[17186] = 2
      "000010" when "0100001100100011", -- t[17187] = 2
      "000010" when "0100001100100100", -- t[17188] = 2
      "000010" when "0100001100100101", -- t[17189] = 2
      "000010" when "0100001100100110", -- t[17190] = 2
      "000010" when "0100001100100111", -- t[17191] = 2
      "000010" when "0100001100101000", -- t[17192] = 2
      "000010" when "0100001100101001", -- t[17193] = 2
      "000010" when "0100001100101010", -- t[17194] = 2
      "000010" when "0100001100101011", -- t[17195] = 2
      "000010" when "0100001100101100", -- t[17196] = 2
      "000010" when "0100001100101101", -- t[17197] = 2
      "000010" when "0100001100101110", -- t[17198] = 2
      "000010" when "0100001100101111", -- t[17199] = 2
      "000010" when "0100001100110000", -- t[17200] = 2
      "000010" when "0100001100110001", -- t[17201] = 2
      "000010" when "0100001100110010", -- t[17202] = 2
      "000010" when "0100001100110011", -- t[17203] = 2
      "000010" when "0100001100110100", -- t[17204] = 2
      "000010" when "0100001100110101", -- t[17205] = 2
      "000010" when "0100001100110110", -- t[17206] = 2
      "000010" when "0100001100110111", -- t[17207] = 2
      "000010" when "0100001100111000", -- t[17208] = 2
      "000010" when "0100001100111001", -- t[17209] = 2
      "000010" when "0100001100111010", -- t[17210] = 2
      "000010" when "0100001100111011", -- t[17211] = 2
      "000010" when "0100001100111100", -- t[17212] = 2
      "000010" when "0100001100111101", -- t[17213] = 2
      "000010" when "0100001100111110", -- t[17214] = 2
      "000010" when "0100001100111111", -- t[17215] = 2
      "000010" when "0100001101000000", -- t[17216] = 2
      "000010" when "0100001101000001", -- t[17217] = 2
      "000010" when "0100001101000010", -- t[17218] = 2
      "000010" when "0100001101000011", -- t[17219] = 2
      "000010" when "0100001101000100", -- t[17220] = 2
      "000010" when "0100001101000101", -- t[17221] = 2
      "000010" when "0100001101000110", -- t[17222] = 2
      "000010" when "0100001101000111", -- t[17223] = 2
      "000010" when "0100001101001000", -- t[17224] = 2
      "000010" when "0100001101001001", -- t[17225] = 2
      "000010" when "0100001101001010", -- t[17226] = 2
      "000010" when "0100001101001011", -- t[17227] = 2
      "000010" when "0100001101001100", -- t[17228] = 2
      "000010" when "0100001101001101", -- t[17229] = 2
      "000010" when "0100001101001110", -- t[17230] = 2
      "000010" when "0100001101001111", -- t[17231] = 2
      "000010" when "0100001101010000", -- t[17232] = 2
      "000010" when "0100001101010001", -- t[17233] = 2
      "000010" when "0100001101010010", -- t[17234] = 2
      "000010" when "0100001101010011", -- t[17235] = 2
      "000010" when "0100001101010100", -- t[17236] = 2
      "000010" when "0100001101010101", -- t[17237] = 2
      "000010" when "0100001101010110", -- t[17238] = 2
      "000010" when "0100001101010111", -- t[17239] = 2
      "000010" when "0100001101011000", -- t[17240] = 2
      "000010" when "0100001101011001", -- t[17241] = 2
      "000010" when "0100001101011010", -- t[17242] = 2
      "000010" when "0100001101011011", -- t[17243] = 2
      "000010" when "0100001101011100", -- t[17244] = 2
      "000010" when "0100001101011101", -- t[17245] = 2
      "000010" when "0100001101011110", -- t[17246] = 2
      "000010" when "0100001101011111", -- t[17247] = 2
      "000010" when "0100001101100000", -- t[17248] = 2
      "000010" when "0100001101100001", -- t[17249] = 2
      "000010" when "0100001101100010", -- t[17250] = 2
      "000010" when "0100001101100011", -- t[17251] = 2
      "000010" when "0100001101100100", -- t[17252] = 2
      "000010" when "0100001101100101", -- t[17253] = 2
      "000010" when "0100001101100110", -- t[17254] = 2
      "000010" when "0100001101100111", -- t[17255] = 2
      "000010" when "0100001101101000", -- t[17256] = 2
      "000010" when "0100001101101001", -- t[17257] = 2
      "000010" when "0100001101101010", -- t[17258] = 2
      "000010" when "0100001101101011", -- t[17259] = 2
      "000010" when "0100001101101100", -- t[17260] = 2
      "000010" when "0100001101101101", -- t[17261] = 2
      "000010" when "0100001101101110", -- t[17262] = 2
      "000010" when "0100001101101111", -- t[17263] = 2
      "000010" when "0100001101110000", -- t[17264] = 2
      "000010" when "0100001101110001", -- t[17265] = 2
      "000010" when "0100001101110010", -- t[17266] = 2
      "000010" when "0100001101110011", -- t[17267] = 2
      "000010" when "0100001101110100", -- t[17268] = 2
      "000010" when "0100001101110101", -- t[17269] = 2
      "000010" when "0100001101110110", -- t[17270] = 2
      "000010" when "0100001101110111", -- t[17271] = 2
      "000010" when "0100001101111000", -- t[17272] = 2
      "000010" when "0100001101111001", -- t[17273] = 2
      "000010" when "0100001101111010", -- t[17274] = 2
      "000010" when "0100001101111011", -- t[17275] = 2
      "000010" when "0100001101111100", -- t[17276] = 2
      "000010" when "0100001101111101", -- t[17277] = 2
      "000010" when "0100001101111110", -- t[17278] = 2
      "000010" when "0100001101111111", -- t[17279] = 2
      "000010" when "0100001110000000", -- t[17280] = 2
      "000010" when "0100001110000001", -- t[17281] = 2
      "000010" when "0100001110000010", -- t[17282] = 2
      "000010" when "0100001110000011", -- t[17283] = 2
      "000010" when "0100001110000100", -- t[17284] = 2
      "000010" when "0100001110000101", -- t[17285] = 2
      "000010" when "0100001110000110", -- t[17286] = 2
      "000010" when "0100001110000111", -- t[17287] = 2
      "000010" when "0100001110001000", -- t[17288] = 2
      "000010" when "0100001110001001", -- t[17289] = 2
      "000010" when "0100001110001010", -- t[17290] = 2
      "000010" when "0100001110001011", -- t[17291] = 2
      "000010" when "0100001110001100", -- t[17292] = 2
      "000010" when "0100001110001101", -- t[17293] = 2
      "000010" when "0100001110001110", -- t[17294] = 2
      "000010" when "0100001110001111", -- t[17295] = 2
      "000010" when "0100001110010000", -- t[17296] = 2
      "000010" when "0100001110010001", -- t[17297] = 2
      "000010" when "0100001110010010", -- t[17298] = 2
      "000010" when "0100001110010011", -- t[17299] = 2
      "000010" when "0100001110010100", -- t[17300] = 2
      "000010" when "0100001110010101", -- t[17301] = 2
      "000010" when "0100001110010110", -- t[17302] = 2
      "000010" when "0100001110010111", -- t[17303] = 2
      "000010" when "0100001110011000", -- t[17304] = 2
      "000010" when "0100001110011001", -- t[17305] = 2
      "000010" when "0100001110011010", -- t[17306] = 2
      "000010" when "0100001110011011", -- t[17307] = 2
      "000010" when "0100001110011100", -- t[17308] = 2
      "000010" when "0100001110011101", -- t[17309] = 2
      "000010" when "0100001110011110", -- t[17310] = 2
      "000010" when "0100001110011111", -- t[17311] = 2
      "000010" when "0100001110100000", -- t[17312] = 2
      "000010" when "0100001110100001", -- t[17313] = 2
      "000010" when "0100001110100010", -- t[17314] = 2
      "000010" when "0100001110100011", -- t[17315] = 2
      "000010" when "0100001110100100", -- t[17316] = 2
      "000010" when "0100001110100101", -- t[17317] = 2
      "000010" when "0100001110100110", -- t[17318] = 2
      "000010" when "0100001110100111", -- t[17319] = 2
      "000010" when "0100001110101000", -- t[17320] = 2
      "000010" when "0100001110101001", -- t[17321] = 2
      "000010" when "0100001110101010", -- t[17322] = 2
      "000010" when "0100001110101011", -- t[17323] = 2
      "000010" when "0100001110101100", -- t[17324] = 2
      "000010" when "0100001110101101", -- t[17325] = 2
      "000010" when "0100001110101110", -- t[17326] = 2
      "000010" when "0100001110101111", -- t[17327] = 2
      "000010" when "0100001110110000", -- t[17328] = 2
      "000010" when "0100001110110001", -- t[17329] = 2
      "000010" when "0100001110110010", -- t[17330] = 2
      "000010" when "0100001110110011", -- t[17331] = 2
      "000010" when "0100001110110100", -- t[17332] = 2
      "000010" when "0100001110110101", -- t[17333] = 2
      "000010" when "0100001110110110", -- t[17334] = 2
      "000010" when "0100001110110111", -- t[17335] = 2
      "000010" when "0100001110111000", -- t[17336] = 2
      "000010" when "0100001110111001", -- t[17337] = 2
      "000010" when "0100001110111010", -- t[17338] = 2
      "000010" when "0100001110111011", -- t[17339] = 2
      "000010" when "0100001110111100", -- t[17340] = 2
      "000010" when "0100001110111101", -- t[17341] = 2
      "000010" when "0100001110111110", -- t[17342] = 2
      "000010" when "0100001110111111", -- t[17343] = 2
      "000010" when "0100001111000000", -- t[17344] = 2
      "000010" when "0100001111000001", -- t[17345] = 2
      "000010" when "0100001111000010", -- t[17346] = 2
      "000010" when "0100001111000011", -- t[17347] = 2
      "000010" when "0100001111000100", -- t[17348] = 2
      "000010" when "0100001111000101", -- t[17349] = 2
      "000010" when "0100001111000110", -- t[17350] = 2
      "000010" when "0100001111000111", -- t[17351] = 2
      "000010" when "0100001111001000", -- t[17352] = 2
      "000010" when "0100001111001001", -- t[17353] = 2
      "000010" when "0100001111001010", -- t[17354] = 2
      "000010" when "0100001111001011", -- t[17355] = 2
      "000010" when "0100001111001100", -- t[17356] = 2
      "000010" when "0100001111001101", -- t[17357] = 2
      "000010" when "0100001111001110", -- t[17358] = 2
      "000010" when "0100001111001111", -- t[17359] = 2
      "000010" when "0100001111010000", -- t[17360] = 2
      "000010" when "0100001111010001", -- t[17361] = 2
      "000010" when "0100001111010010", -- t[17362] = 2
      "000010" when "0100001111010011", -- t[17363] = 2
      "000010" when "0100001111010100", -- t[17364] = 2
      "000010" when "0100001111010101", -- t[17365] = 2
      "000010" when "0100001111010110", -- t[17366] = 2
      "000010" when "0100001111010111", -- t[17367] = 2
      "000010" when "0100001111011000", -- t[17368] = 2
      "000010" when "0100001111011001", -- t[17369] = 2
      "000010" when "0100001111011010", -- t[17370] = 2
      "000010" when "0100001111011011", -- t[17371] = 2
      "000010" when "0100001111011100", -- t[17372] = 2
      "000010" when "0100001111011101", -- t[17373] = 2
      "000010" when "0100001111011110", -- t[17374] = 2
      "000010" when "0100001111011111", -- t[17375] = 2
      "000010" when "0100001111100000", -- t[17376] = 2
      "000010" when "0100001111100001", -- t[17377] = 2
      "000010" when "0100001111100010", -- t[17378] = 2
      "000010" when "0100001111100011", -- t[17379] = 2
      "000010" when "0100001111100100", -- t[17380] = 2
      "000010" when "0100001111100101", -- t[17381] = 2
      "000010" when "0100001111100110", -- t[17382] = 2
      "000010" when "0100001111100111", -- t[17383] = 2
      "000010" when "0100001111101000", -- t[17384] = 2
      "000010" when "0100001111101001", -- t[17385] = 2
      "000010" when "0100001111101010", -- t[17386] = 2
      "000010" when "0100001111101011", -- t[17387] = 2
      "000010" when "0100001111101100", -- t[17388] = 2
      "000010" when "0100001111101101", -- t[17389] = 2
      "000010" when "0100001111101110", -- t[17390] = 2
      "000010" when "0100001111101111", -- t[17391] = 2
      "000010" when "0100001111110000", -- t[17392] = 2
      "000010" when "0100001111110001", -- t[17393] = 2
      "000010" when "0100001111110010", -- t[17394] = 2
      "000010" when "0100001111110011", -- t[17395] = 2
      "000010" when "0100001111110100", -- t[17396] = 2
      "000010" when "0100001111110101", -- t[17397] = 2
      "000010" when "0100001111110110", -- t[17398] = 2
      "000010" when "0100001111110111", -- t[17399] = 2
      "000010" when "0100001111111000", -- t[17400] = 2
      "000010" when "0100001111111001", -- t[17401] = 2
      "000010" when "0100001111111010", -- t[17402] = 2
      "000010" when "0100001111111011", -- t[17403] = 2
      "000010" when "0100001111111100", -- t[17404] = 2
      "000010" when "0100001111111101", -- t[17405] = 2
      "000010" when "0100001111111110", -- t[17406] = 2
      "000010" when "0100001111111111", -- t[17407] = 2
      "000010" when "0100010000000000", -- t[17408] = 2
      "000010" when "0100010000000001", -- t[17409] = 2
      "000010" when "0100010000000010", -- t[17410] = 2
      "000010" when "0100010000000011", -- t[17411] = 2
      "000010" when "0100010000000100", -- t[17412] = 2
      "000010" when "0100010000000101", -- t[17413] = 2
      "000010" when "0100010000000110", -- t[17414] = 2
      "000010" when "0100010000000111", -- t[17415] = 2
      "000010" when "0100010000001000", -- t[17416] = 2
      "000010" when "0100010000001001", -- t[17417] = 2
      "000010" when "0100010000001010", -- t[17418] = 2
      "000010" when "0100010000001011", -- t[17419] = 2
      "000010" when "0100010000001100", -- t[17420] = 2
      "000010" when "0100010000001101", -- t[17421] = 2
      "000010" when "0100010000001110", -- t[17422] = 2
      "000010" when "0100010000001111", -- t[17423] = 2
      "000010" when "0100010000010000", -- t[17424] = 2
      "000010" when "0100010000010001", -- t[17425] = 2
      "000010" when "0100010000010010", -- t[17426] = 2
      "000010" when "0100010000010011", -- t[17427] = 2
      "000010" when "0100010000010100", -- t[17428] = 2
      "000010" when "0100010000010101", -- t[17429] = 2
      "000010" when "0100010000010110", -- t[17430] = 2
      "000010" when "0100010000010111", -- t[17431] = 2
      "000010" when "0100010000011000", -- t[17432] = 2
      "000010" when "0100010000011001", -- t[17433] = 2
      "000010" when "0100010000011010", -- t[17434] = 2
      "000010" when "0100010000011011", -- t[17435] = 2
      "000010" when "0100010000011100", -- t[17436] = 2
      "000010" when "0100010000011101", -- t[17437] = 2
      "000010" when "0100010000011110", -- t[17438] = 2
      "000010" when "0100010000011111", -- t[17439] = 2
      "000010" when "0100010000100000", -- t[17440] = 2
      "000010" when "0100010000100001", -- t[17441] = 2
      "000010" when "0100010000100010", -- t[17442] = 2
      "000010" when "0100010000100011", -- t[17443] = 2
      "000010" when "0100010000100100", -- t[17444] = 2
      "000010" when "0100010000100101", -- t[17445] = 2
      "000010" when "0100010000100110", -- t[17446] = 2
      "000010" when "0100010000100111", -- t[17447] = 2
      "000010" when "0100010000101000", -- t[17448] = 2
      "000010" when "0100010000101001", -- t[17449] = 2
      "000010" when "0100010000101010", -- t[17450] = 2
      "000010" when "0100010000101011", -- t[17451] = 2
      "000010" when "0100010000101100", -- t[17452] = 2
      "000010" when "0100010000101101", -- t[17453] = 2
      "000010" when "0100010000101110", -- t[17454] = 2
      "000010" when "0100010000101111", -- t[17455] = 2
      "000010" when "0100010000110000", -- t[17456] = 2
      "000010" when "0100010000110001", -- t[17457] = 2
      "000010" when "0100010000110010", -- t[17458] = 2
      "000010" when "0100010000110011", -- t[17459] = 2
      "000010" when "0100010000110100", -- t[17460] = 2
      "000010" when "0100010000110101", -- t[17461] = 2
      "000010" when "0100010000110110", -- t[17462] = 2
      "000010" when "0100010000110111", -- t[17463] = 2
      "000010" when "0100010000111000", -- t[17464] = 2
      "000010" when "0100010000111001", -- t[17465] = 2
      "000010" when "0100010000111010", -- t[17466] = 2
      "000010" when "0100010000111011", -- t[17467] = 2
      "000010" when "0100010000111100", -- t[17468] = 2
      "000010" when "0100010000111101", -- t[17469] = 2
      "000010" when "0100010000111110", -- t[17470] = 2
      "000010" when "0100010000111111", -- t[17471] = 2
      "000010" when "0100010001000000", -- t[17472] = 2
      "000010" when "0100010001000001", -- t[17473] = 2
      "000010" when "0100010001000010", -- t[17474] = 2
      "000010" when "0100010001000011", -- t[17475] = 2
      "000010" when "0100010001000100", -- t[17476] = 2
      "000010" when "0100010001000101", -- t[17477] = 2
      "000010" when "0100010001000110", -- t[17478] = 2
      "000010" when "0100010001000111", -- t[17479] = 2
      "000010" when "0100010001001000", -- t[17480] = 2
      "000010" when "0100010001001001", -- t[17481] = 2
      "000010" when "0100010001001010", -- t[17482] = 2
      "000010" when "0100010001001011", -- t[17483] = 2
      "000010" when "0100010001001100", -- t[17484] = 2
      "000010" when "0100010001001101", -- t[17485] = 2
      "000010" when "0100010001001110", -- t[17486] = 2
      "000010" when "0100010001001111", -- t[17487] = 2
      "000010" when "0100010001010000", -- t[17488] = 2
      "000010" when "0100010001010001", -- t[17489] = 2
      "000010" when "0100010001010010", -- t[17490] = 2
      "000010" when "0100010001010011", -- t[17491] = 2
      "000010" when "0100010001010100", -- t[17492] = 2
      "000010" when "0100010001010101", -- t[17493] = 2
      "000010" when "0100010001010110", -- t[17494] = 2
      "000010" when "0100010001010111", -- t[17495] = 2
      "000010" when "0100010001011000", -- t[17496] = 2
      "000010" when "0100010001011001", -- t[17497] = 2
      "000010" when "0100010001011010", -- t[17498] = 2
      "000010" when "0100010001011011", -- t[17499] = 2
      "000010" when "0100010001011100", -- t[17500] = 2
      "000010" when "0100010001011101", -- t[17501] = 2
      "000010" when "0100010001011110", -- t[17502] = 2
      "000010" when "0100010001011111", -- t[17503] = 2
      "000010" when "0100010001100000", -- t[17504] = 2
      "000010" when "0100010001100001", -- t[17505] = 2
      "000010" when "0100010001100010", -- t[17506] = 2
      "000010" when "0100010001100011", -- t[17507] = 2
      "000010" when "0100010001100100", -- t[17508] = 2
      "000010" when "0100010001100101", -- t[17509] = 2
      "000010" when "0100010001100110", -- t[17510] = 2
      "000010" when "0100010001100111", -- t[17511] = 2
      "000010" when "0100010001101000", -- t[17512] = 2
      "000010" when "0100010001101001", -- t[17513] = 2
      "000010" when "0100010001101010", -- t[17514] = 2
      "000010" when "0100010001101011", -- t[17515] = 2
      "000010" when "0100010001101100", -- t[17516] = 2
      "000010" when "0100010001101101", -- t[17517] = 2
      "000010" when "0100010001101110", -- t[17518] = 2
      "000010" when "0100010001101111", -- t[17519] = 2
      "000010" when "0100010001110000", -- t[17520] = 2
      "000010" when "0100010001110001", -- t[17521] = 2
      "000010" when "0100010001110010", -- t[17522] = 2
      "000010" when "0100010001110011", -- t[17523] = 2
      "000010" when "0100010001110100", -- t[17524] = 2
      "000010" when "0100010001110101", -- t[17525] = 2
      "000010" when "0100010001110110", -- t[17526] = 2
      "000010" when "0100010001110111", -- t[17527] = 2
      "000010" when "0100010001111000", -- t[17528] = 2
      "000010" when "0100010001111001", -- t[17529] = 2
      "000010" when "0100010001111010", -- t[17530] = 2
      "000010" when "0100010001111011", -- t[17531] = 2
      "000010" when "0100010001111100", -- t[17532] = 2
      "000010" when "0100010001111101", -- t[17533] = 2
      "000010" when "0100010001111110", -- t[17534] = 2
      "000010" when "0100010001111111", -- t[17535] = 2
      "000010" when "0100010010000000", -- t[17536] = 2
      "000010" when "0100010010000001", -- t[17537] = 2
      "000010" when "0100010010000010", -- t[17538] = 2
      "000010" when "0100010010000011", -- t[17539] = 2
      "000010" when "0100010010000100", -- t[17540] = 2
      "000010" when "0100010010000101", -- t[17541] = 2
      "000010" when "0100010010000110", -- t[17542] = 2
      "000010" when "0100010010000111", -- t[17543] = 2
      "000010" when "0100010010001000", -- t[17544] = 2
      "000010" when "0100010010001001", -- t[17545] = 2
      "000010" when "0100010010001010", -- t[17546] = 2
      "000010" when "0100010010001011", -- t[17547] = 2
      "000010" when "0100010010001100", -- t[17548] = 2
      "000010" when "0100010010001101", -- t[17549] = 2
      "000010" when "0100010010001110", -- t[17550] = 2
      "000010" when "0100010010001111", -- t[17551] = 2
      "000010" when "0100010010010000", -- t[17552] = 2
      "000010" when "0100010010010001", -- t[17553] = 2
      "000010" when "0100010010010010", -- t[17554] = 2
      "000010" when "0100010010010011", -- t[17555] = 2
      "000010" when "0100010010010100", -- t[17556] = 2
      "000010" when "0100010010010101", -- t[17557] = 2
      "000010" when "0100010010010110", -- t[17558] = 2
      "000010" when "0100010010010111", -- t[17559] = 2
      "000010" when "0100010010011000", -- t[17560] = 2
      "000010" when "0100010010011001", -- t[17561] = 2
      "000010" when "0100010010011010", -- t[17562] = 2
      "000010" when "0100010010011011", -- t[17563] = 2
      "000010" when "0100010010011100", -- t[17564] = 2
      "000010" when "0100010010011101", -- t[17565] = 2
      "000010" when "0100010010011110", -- t[17566] = 2
      "000010" when "0100010010011111", -- t[17567] = 2
      "000010" when "0100010010100000", -- t[17568] = 2
      "000010" when "0100010010100001", -- t[17569] = 2
      "000010" when "0100010010100010", -- t[17570] = 2
      "000010" when "0100010010100011", -- t[17571] = 2
      "000010" when "0100010010100100", -- t[17572] = 2
      "000010" when "0100010010100101", -- t[17573] = 2
      "000010" when "0100010010100110", -- t[17574] = 2
      "000010" when "0100010010100111", -- t[17575] = 2
      "000010" when "0100010010101000", -- t[17576] = 2
      "000010" when "0100010010101001", -- t[17577] = 2
      "000010" when "0100010010101010", -- t[17578] = 2
      "000010" when "0100010010101011", -- t[17579] = 2
      "000010" when "0100010010101100", -- t[17580] = 2
      "000010" when "0100010010101101", -- t[17581] = 2
      "000010" when "0100010010101110", -- t[17582] = 2
      "000010" when "0100010010101111", -- t[17583] = 2
      "000010" when "0100010010110000", -- t[17584] = 2
      "000010" when "0100010010110001", -- t[17585] = 2
      "000010" when "0100010010110010", -- t[17586] = 2
      "000010" when "0100010010110011", -- t[17587] = 2
      "000010" when "0100010010110100", -- t[17588] = 2
      "000010" when "0100010010110101", -- t[17589] = 2
      "000010" when "0100010010110110", -- t[17590] = 2
      "000010" when "0100010010110111", -- t[17591] = 2
      "000010" when "0100010010111000", -- t[17592] = 2
      "000010" when "0100010010111001", -- t[17593] = 2
      "000010" when "0100010010111010", -- t[17594] = 2
      "000010" when "0100010010111011", -- t[17595] = 2
      "000010" when "0100010010111100", -- t[17596] = 2
      "000010" when "0100010010111101", -- t[17597] = 2
      "000010" when "0100010010111110", -- t[17598] = 2
      "000010" when "0100010010111111", -- t[17599] = 2
      "000010" when "0100010011000000", -- t[17600] = 2
      "000010" when "0100010011000001", -- t[17601] = 2
      "000010" when "0100010011000010", -- t[17602] = 2
      "000010" when "0100010011000011", -- t[17603] = 2
      "000010" when "0100010011000100", -- t[17604] = 2
      "000010" when "0100010011000101", -- t[17605] = 2
      "000010" when "0100010011000110", -- t[17606] = 2
      "000010" when "0100010011000111", -- t[17607] = 2
      "000010" when "0100010011001000", -- t[17608] = 2
      "000010" when "0100010011001001", -- t[17609] = 2
      "000010" when "0100010011001010", -- t[17610] = 2
      "000010" when "0100010011001011", -- t[17611] = 2
      "000010" when "0100010011001100", -- t[17612] = 2
      "000010" when "0100010011001101", -- t[17613] = 2
      "000010" when "0100010011001110", -- t[17614] = 2
      "000010" when "0100010011001111", -- t[17615] = 2
      "000010" when "0100010011010000", -- t[17616] = 2
      "000010" when "0100010011010001", -- t[17617] = 2
      "000010" when "0100010011010010", -- t[17618] = 2
      "000010" when "0100010011010011", -- t[17619] = 2
      "000010" when "0100010011010100", -- t[17620] = 2
      "000010" when "0100010011010101", -- t[17621] = 2
      "000010" when "0100010011010110", -- t[17622] = 2
      "000010" when "0100010011010111", -- t[17623] = 2
      "000010" when "0100010011011000", -- t[17624] = 2
      "000010" when "0100010011011001", -- t[17625] = 2
      "000010" when "0100010011011010", -- t[17626] = 2
      "000010" when "0100010011011011", -- t[17627] = 2
      "000010" when "0100010011011100", -- t[17628] = 2
      "000010" when "0100010011011101", -- t[17629] = 2
      "000010" when "0100010011011110", -- t[17630] = 2
      "000010" when "0100010011011111", -- t[17631] = 2
      "000010" when "0100010011100000", -- t[17632] = 2
      "000010" when "0100010011100001", -- t[17633] = 2
      "000010" when "0100010011100010", -- t[17634] = 2
      "000010" when "0100010011100011", -- t[17635] = 2
      "000010" when "0100010011100100", -- t[17636] = 2
      "000010" when "0100010011100101", -- t[17637] = 2
      "000010" when "0100010011100110", -- t[17638] = 2
      "000010" when "0100010011100111", -- t[17639] = 2
      "000010" when "0100010011101000", -- t[17640] = 2
      "000010" when "0100010011101001", -- t[17641] = 2
      "000010" when "0100010011101010", -- t[17642] = 2
      "000010" when "0100010011101011", -- t[17643] = 2
      "000010" when "0100010011101100", -- t[17644] = 2
      "000010" when "0100010011101101", -- t[17645] = 2
      "000010" when "0100010011101110", -- t[17646] = 2
      "000010" when "0100010011101111", -- t[17647] = 2
      "000010" when "0100010011110000", -- t[17648] = 2
      "000010" when "0100010011110001", -- t[17649] = 2
      "000010" when "0100010011110010", -- t[17650] = 2
      "000010" when "0100010011110011", -- t[17651] = 2
      "000010" when "0100010011110100", -- t[17652] = 2
      "000010" when "0100010011110101", -- t[17653] = 2
      "000010" when "0100010011110110", -- t[17654] = 2
      "000010" when "0100010011110111", -- t[17655] = 2
      "000010" when "0100010011111000", -- t[17656] = 2
      "000010" when "0100010011111001", -- t[17657] = 2
      "000010" when "0100010011111010", -- t[17658] = 2
      "000010" when "0100010011111011", -- t[17659] = 2
      "000010" when "0100010011111100", -- t[17660] = 2
      "000010" when "0100010011111101", -- t[17661] = 2
      "000010" when "0100010011111110", -- t[17662] = 2
      "000010" when "0100010011111111", -- t[17663] = 2
      "000010" when "0100010100000000", -- t[17664] = 2
      "000010" when "0100010100000001", -- t[17665] = 2
      "000010" when "0100010100000010", -- t[17666] = 2
      "000010" when "0100010100000011", -- t[17667] = 2
      "000010" when "0100010100000100", -- t[17668] = 2
      "000010" when "0100010100000101", -- t[17669] = 2
      "000010" when "0100010100000110", -- t[17670] = 2
      "000010" when "0100010100000111", -- t[17671] = 2
      "000010" when "0100010100001000", -- t[17672] = 2
      "000010" when "0100010100001001", -- t[17673] = 2
      "000010" when "0100010100001010", -- t[17674] = 2
      "000010" when "0100010100001011", -- t[17675] = 2
      "000010" when "0100010100001100", -- t[17676] = 2
      "000010" when "0100010100001101", -- t[17677] = 2
      "000010" when "0100010100001110", -- t[17678] = 2
      "000010" when "0100010100001111", -- t[17679] = 2
      "000010" when "0100010100010000", -- t[17680] = 2
      "000010" when "0100010100010001", -- t[17681] = 2
      "000010" when "0100010100010010", -- t[17682] = 2
      "000010" when "0100010100010011", -- t[17683] = 2
      "000010" when "0100010100010100", -- t[17684] = 2
      "000010" when "0100010100010101", -- t[17685] = 2
      "000010" when "0100010100010110", -- t[17686] = 2
      "000010" when "0100010100010111", -- t[17687] = 2
      "000010" when "0100010100011000", -- t[17688] = 2
      "000010" when "0100010100011001", -- t[17689] = 2
      "000010" when "0100010100011010", -- t[17690] = 2
      "000010" when "0100010100011011", -- t[17691] = 2
      "000010" when "0100010100011100", -- t[17692] = 2
      "000010" when "0100010100011101", -- t[17693] = 2
      "000010" when "0100010100011110", -- t[17694] = 2
      "000010" when "0100010100011111", -- t[17695] = 2
      "000010" when "0100010100100000", -- t[17696] = 2
      "000010" when "0100010100100001", -- t[17697] = 2
      "000010" when "0100010100100010", -- t[17698] = 2
      "000010" when "0100010100100011", -- t[17699] = 2
      "000010" when "0100010100100100", -- t[17700] = 2
      "000010" when "0100010100100101", -- t[17701] = 2
      "000010" when "0100010100100110", -- t[17702] = 2
      "000010" when "0100010100100111", -- t[17703] = 2
      "000010" when "0100010100101000", -- t[17704] = 2
      "000010" when "0100010100101001", -- t[17705] = 2
      "000010" when "0100010100101010", -- t[17706] = 2
      "000010" when "0100010100101011", -- t[17707] = 2
      "000010" when "0100010100101100", -- t[17708] = 2
      "000010" when "0100010100101101", -- t[17709] = 2
      "000010" when "0100010100101110", -- t[17710] = 2
      "000010" when "0100010100101111", -- t[17711] = 2
      "000010" when "0100010100110000", -- t[17712] = 2
      "000010" when "0100010100110001", -- t[17713] = 2
      "000010" when "0100010100110010", -- t[17714] = 2
      "000010" when "0100010100110011", -- t[17715] = 2
      "000010" when "0100010100110100", -- t[17716] = 2
      "000010" when "0100010100110101", -- t[17717] = 2
      "000010" when "0100010100110110", -- t[17718] = 2
      "000010" when "0100010100110111", -- t[17719] = 2
      "000010" when "0100010100111000", -- t[17720] = 2
      "000010" when "0100010100111001", -- t[17721] = 2
      "000010" when "0100010100111010", -- t[17722] = 2
      "000010" when "0100010100111011", -- t[17723] = 2
      "000010" when "0100010100111100", -- t[17724] = 2
      "000010" when "0100010100111101", -- t[17725] = 2
      "000010" when "0100010100111110", -- t[17726] = 2
      "000010" when "0100010100111111", -- t[17727] = 2
      "000010" when "0100010101000000", -- t[17728] = 2
      "000010" when "0100010101000001", -- t[17729] = 2
      "000010" when "0100010101000010", -- t[17730] = 2
      "000010" when "0100010101000011", -- t[17731] = 2
      "000010" when "0100010101000100", -- t[17732] = 2
      "000010" when "0100010101000101", -- t[17733] = 2
      "000010" when "0100010101000110", -- t[17734] = 2
      "000010" when "0100010101000111", -- t[17735] = 2
      "000010" when "0100010101001000", -- t[17736] = 2
      "000010" when "0100010101001001", -- t[17737] = 2
      "000010" when "0100010101001010", -- t[17738] = 2
      "000010" when "0100010101001011", -- t[17739] = 2
      "000010" when "0100010101001100", -- t[17740] = 2
      "000010" when "0100010101001101", -- t[17741] = 2
      "000010" when "0100010101001110", -- t[17742] = 2
      "000010" when "0100010101001111", -- t[17743] = 2
      "000010" when "0100010101010000", -- t[17744] = 2
      "000010" when "0100010101010001", -- t[17745] = 2
      "000010" when "0100010101010010", -- t[17746] = 2
      "000010" when "0100010101010011", -- t[17747] = 2
      "000010" when "0100010101010100", -- t[17748] = 2
      "000010" when "0100010101010101", -- t[17749] = 2
      "000010" when "0100010101010110", -- t[17750] = 2
      "000010" when "0100010101010111", -- t[17751] = 2
      "000010" when "0100010101011000", -- t[17752] = 2
      "000010" when "0100010101011001", -- t[17753] = 2
      "000010" when "0100010101011010", -- t[17754] = 2
      "000010" when "0100010101011011", -- t[17755] = 2
      "000010" when "0100010101011100", -- t[17756] = 2
      "000010" when "0100010101011101", -- t[17757] = 2
      "000010" when "0100010101011110", -- t[17758] = 2
      "000010" when "0100010101011111", -- t[17759] = 2
      "000010" when "0100010101100000", -- t[17760] = 2
      "000010" when "0100010101100001", -- t[17761] = 2
      "000010" when "0100010101100010", -- t[17762] = 2
      "000010" when "0100010101100011", -- t[17763] = 2
      "000010" when "0100010101100100", -- t[17764] = 2
      "000010" when "0100010101100101", -- t[17765] = 2
      "000010" when "0100010101100110", -- t[17766] = 2
      "000010" when "0100010101100111", -- t[17767] = 2
      "000010" when "0100010101101000", -- t[17768] = 2
      "000010" when "0100010101101001", -- t[17769] = 2
      "000010" when "0100010101101010", -- t[17770] = 2
      "000010" when "0100010101101011", -- t[17771] = 2
      "000010" when "0100010101101100", -- t[17772] = 2
      "000010" when "0100010101101101", -- t[17773] = 2
      "000010" when "0100010101101110", -- t[17774] = 2
      "000010" when "0100010101101111", -- t[17775] = 2
      "000010" when "0100010101110000", -- t[17776] = 2
      "000010" when "0100010101110001", -- t[17777] = 2
      "000010" when "0100010101110010", -- t[17778] = 2
      "000010" when "0100010101110011", -- t[17779] = 2
      "000010" when "0100010101110100", -- t[17780] = 2
      "000010" when "0100010101110101", -- t[17781] = 2
      "000010" when "0100010101110110", -- t[17782] = 2
      "000010" when "0100010101110111", -- t[17783] = 2
      "000010" when "0100010101111000", -- t[17784] = 2
      "000010" when "0100010101111001", -- t[17785] = 2
      "000010" when "0100010101111010", -- t[17786] = 2
      "000010" when "0100010101111011", -- t[17787] = 2
      "000010" when "0100010101111100", -- t[17788] = 2
      "000010" when "0100010101111101", -- t[17789] = 2
      "000010" when "0100010101111110", -- t[17790] = 2
      "000010" when "0100010101111111", -- t[17791] = 2
      "000010" when "0100010110000000", -- t[17792] = 2
      "000010" when "0100010110000001", -- t[17793] = 2
      "000010" when "0100010110000010", -- t[17794] = 2
      "000010" when "0100010110000011", -- t[17795] = 2
      "000010" when "0100010110000100", -- t[17796] = 2
      "000010" when "0100010110000101", -- t[17797] = 2
      "000010" when "0100010110000110", -- t[17798] = 2
      "000010" when "0100010110000111", -- t[17799] = 2
      "000010" when "0100010110001000", -- t[17800] = 2
      "000010" when "0100010110001001", -- t[17801] = 2
      "000010" when "0100010110001010", -- t[17802] = 2
      "000010" when "0100010110001011", -- t[17803] = 2
      "000010" when "0100010110001100", -- t[17804] = 2
      "000010" when "0100010110001101", -- t[17805] = 2
      "000010" when "0100010110001110", -- t[17806] = 2
      "000010" when "0100010110001111", -- t[17807] = 2
      "000010" when "0100010110010000", -- t[17808] = 2
      "000010" when "0100010110010001", -- t[17809] = 2
      "000010" when "0100010110010010", -- t[17810] = 2
      "000010" when "0100010110010011", -- t[17811] = 2
      "000010" when "0100010110010100", -- t[17812] = 2
      "000010" when "0100010110010101", -- t[17813] = 2
      "000010" when "0100010110010110", -- t[17814] = 2
      "000010" when "0100010110010111", -- t[17815] = 2
      "000010" when "0100010110011000", -- t[17816] = 2
      "000010" when "0100010110011001", -- t[17817] = 2
      "000010" when "0100010110011010", -- t[17818] = 2
      "000010" when "0100010110011011", -- t[17819] = 2
      "000010" when "0100010110011100", -- t[17820] = 2
      "000010" when "0100010110011101", -- t[17821] = 2
      "000010" when "0100010110011110", -- t[17822] = 2
      "000010" when "0100010110011111", -- t[17823] = 2
      "000010" when "0100010110100000", -- t[17824] = 2
      "000010" when "0100010110100001", -- t[17825] = 2
      "000010" when "0100010110100010", -- t[17826] = 2
      "000010" when "0100010110100011", -- t[17827] = 2
      "000010" when "0100010110100100", -- t[17828] = 2
      "000010" when "0100010110100101", -- t[17829] = 2
      "000010" when "0100010110100110", -- t[17830] = 2
      "000010" when "0100010110100111", -- t[17831] = 2
      "000010" when "0100010110101000", -- t[17832] = 2
      "000010" when "0100010110101001", -- t[17833] = 2
      "000010" when "0100010110101010", -- t[17834] = 2
      "000010" when "0100010110101011", -- t[17835] = 2
      "000010" when "0100010110101100", -- t[17836] = 2
      "000010" when "0100010110101101", -- t[17837] = 2
      "000010" when "0100010110101110", -- t[17838] = 2
      "000010" when "0100010110101111", -- t[17839] = 2
      "000010" when "0100010110110000", -- t[17840] = 2
      "000010" when "0100010110110001", -- t[17841] = 2
      "000010" when "0100010110110010", -- t[17842] = 2
      "000010" when "0100010110110011", -- t[17843] = 2
      "000010" when "0100010110110100", -- t[17844] = 2
      "000010" when "0100010110110101", -- t[17845] = 2
      "000010" when "0100010110110110", -- t[17846] = 2
      "000010" when "0100010110110111", -- t[17847] = 2
      "000010" when "0100010110111000", -- t[17848] = 2
      "000010" when "0100010110111001", -- t[17849] = 2
      "000010" when "0100010110111010", -- t[17850] = 2
      "000010" when "0100010110111011", -- t[17851] = 2
      "000010" when "0100010110111100", -- t[17852] = 2
      "000010" when "0100010110111101", -- t[17853] = 2
      "000010" when "0100010110111110", -- t[17854] = 2
      "000010" when "0100010110111111", -- t[17855] = 2
      "000010" when "0100010111000000", -- t[17856] = 2
      "000010" when "0100010111000001", -- t[17857] = 2
      "000010" when "0100010111000010", -- t[17858] = 2
      "000010" when "0100010111000011", -- t[17859] = 2
      "000010" when "0100010111000100", -- t[17860] = 2
      "000010" when "0100010111000101", -- t[17861] = 2
      "000010" when "0100010111000110", -- t[17862] = 2
      "000010" when "0100010111000111", -- t[17863] = 2
      "000010" when "0100010111001000", -- t[17864] = 2
      "000010" when "0100010111001001", -- t[17865] = 2
      "000010" when "0100010111001010", -- t[17866] = 2
      "000010" when "0100010111001011", -- t[17867] = 2
      "000010" when "0100010111001100", -- t[17868] = 2
      "000010" when "0100010111001101", -- t[17869] = 2
      "000010" when "0100010111001110", -- t[17870] = 2
      "000010" when "0100010111001111", -- t[17871] = 2
      "000010" when "0100010111010000", -- t[17872] = 2
      "000010" when "0100010111010001", -- t[17873] = 2
      "000010" when "0100010111010010", -- t[17874] = 2
      "000010" when "0100010111010011", -- t[17875] = 2
      "000010" when "0100010111010100", -- t[17876] = 2
      "000010" when "0100010111010101", -- t[17877] = 2
      "000010" when "0100010111010110", -- t[17878] = 2
      "000010" when "0100010111010111", -- t[17879] = 2
      "000010" when "0100010111011000", -- t[17880] = 2
      "000010" when "0100010111011001", -- t[17881] = 2
      "000010" when "0100010111011010", -- t[17882] = 2
      "000010" when "0100010111011011", -- t[17883] = 2
      "000010" when "0100010111011100", -- t[17884] = 2
      "000010" when "0100010111011101", -- t[17885] = 2
      "000010" when "0100010111011110", -- t[17886] = 2
      "000010" when "0100010111011111", -- t[17887] = 2
      "000010" when "0100010111100000", -- t[17888] = 2
      "000010" when "0100010111100001", -- t[17889] = 2
      "000010" when "0100010111100010", -- t[17890] = 2
      "000010" when "0100010111100011", -- t[17891] = 2
      "000010" when "0100010111100100", -- t[17892] = 2
      "000010" when "0100010111100101", -- t[17893] = 2
      "000010" when "0100010111100110", -- t[17894] = 2
      "000010" when "0100010111100111", -- t[17895] = 2
      "000010" when "0100010111101000", -- t[17896] = 2
      "000010" when "0100010111101001", -- t[17897] = 2
      "000010" when "0100010111101010", -- t[17898] = 2
      "000010" when "0100010111101011", -- t[17899] = 2
      "000010" when "0100010111101100", -- t[17900] = 2
      "000010" when "0100010111101101", -- t[17901] = 2
      "000010" when "0100010111101110", -- t[17902] = 2
      "000010" when "0100010111101111", -- t[17903] = 2
      "000010" when "0100010111110000", -- t[17904] = 2
      "000010" when "0100010111110001", -- t[17905] = 2
      "000010" when "0100010111110010", -- t[17906] = 2
      "000010" when "0100010111110011", -- t[17907] = 2
      "000010" when "0100010111110100", -- t[17908] = 2
      "000010" when "0100010111110101", -- t[17909] = 2
      "000010" when "0100010111110110", -- t[17910] = 2
      "000010" when "0100010111110111", -- t[17911] = 2
      "000010" when "0100010111111000", -- t[17912] = 2
      "000010" when "0100010111111001", -- t[17913] = 2
      "000010" when "0100010111111010", -- t[17914] = 2
      "000010" when "0100010111111011", -- t[17915] = 2
      "000010" when "0100010111111100", -- t[17916] = 2
      "000010" when "0100010111111101", -- t[17917] = 2
      "000010" when "0100010111111110", -- t[17918] = 2
      "000010" when "0100010111111111", -- t[17919] = 2
      "000010" when "0100011000000000", -- t[17920] = 2
      "000010" when "0100011000000001", -- t[17921] = 2
      "000010" when "0100011000000010", -- t[17922] = 2
      "000010" when "0100011000000011", -- t[17923] = 2
      "000010" when "0100011000000100", -- t[17924] = 2
      "000010" when "0100011000000101", -- t[17925] = 2
      "000010" when "0100011000000110", -- t[17926] = 2
      "000010" when "0100011000000111", -- t[17927] = 2
      "000010" when "0100011000001000", -- t[17928] = 2
      "000010" when "0100011000001001", -- t[17929] = 2
      "000010" when "0100011000001010", -- t[17930] = 2
      "000010" when "0100011000001011", -- t[17931] = 2
      "000010" when "0100011000001100", -- t[17932] = 2
      "000010" when "0100011000001101", -- t[17933] = 2
      "000010" when "0100011000001110", -- t[17934] = 2
      "000010" when "0100011000001111", -- t[17935] = 2
      "000010" when "0100011000010000", -- t[17936] = 2
      "000010" when "0100011000010001", -- t[17937] = 2
      "000010" when "0100011000010010", -- t[17938] = 2
      "000010" when "0100011000010011", -- t[17939] = 2
      "000010" when "0100011000010100", -- t[17940] = 2
      "000010" when "0100011000010101", -- t[17941] = 2
      "000010" when "0100011000010110", -- t[17942] = 2
      "000010" when "0100011000010111", -- t[17943] = 2
      "000010" when "0100011000011000", -- t[17944] = 2
      "000010" when "0100011000011001", -- t[17945] = 2
      "000010" when "0100011000011010", -- t[17946] = 2
      "000010" when "0100011000011011", -- t[17947] = 2
      "000010" when "0100011000011100", -- t[17948] = 2
      "000010" when "0100011000011101", -- t[17949] = 2
      "000010" when "0100011000011110", -- t[17950] = 2
      "000010" when "0100011000011111", -- t[17951] = 2
      "000010" when "0100011000100000", -- t[17952] = 2
      "000010" when "0100011000100001", -- t[17953] = 2
      "000010" when "0100011000100010", -- t[17954] = 2
      "000010" when "0100011000100011", -- t[17955] = 2
      "000010" when "0100011000100100", -- t[17956] = 2
      "000010" when "0100011000100101", -- t[17957] = 2
      "000010" when "0100011000100110", -- t[17958] = 2
      "000010" when "0100011000100111", -- t[17959] = 2
      "000010" when "0100011000101000", -- t[17960] = 2
      "000010" when "0100011000101001", -- t[17961] = 2
      "000010" when "0100011000101010", -- t[17962] = 2
      "000010" when "0100011000101011", -- t[17963] = 2
      "000010" when "0100011000101100", -- t[17964] = 2
      "000010" when "0100011000101101", -- t[17965] = 2
      "000010" when "0100011000101110", -- t[17966] = 2
      "000010" when "0100011000101111", -- t[17967] = 2
      "000010" when "0100011000110000", -- t[17968] = 2
      "000010" when "0100011000110001", -- t[17969] = 2
      "000010" when "0100011000110010", -- t[17970] = 2
      "000010" when "0100011000110011", -- t[17971] = 2
      "000010" when "0100011000110100", -- t[17972] = 2
      "000010" when "0100011000110101", -- t[17973] = 2
      "000010" when "0100011000110110", -- t[17974] = 2
      "000010" when "0100011000110111", -- t[17975] = 2
      "000010" when "0100011000111000", -- t[17976] = 2
      "000010" when "0100011000111001", -- t[17977] = 2
      "000010" when "0100011000111010", -- t[17978] = 2
      "000010" when "0100011000111011", -- t[17979] = 2
      "000010" when "0100011000111100", -- t[17980] = 2
      "000010" when "0100011000111101", -- t[17981] = 2
      "000010" when "0100011000111110", -- t[17982] = 2
      "000010" when "0100011000111111", -- t[17983] = 2
      "000010" when "0100011001000000", -- t[17984] = 2
      "000010" when "0100011001000001", -- t[17985] = 2
      "000010" when "0100011001000010", -- t[17986] = 2
      "000010" when "0100011001000011", -- t[17987] = 2
      "000010" when "0100011001000100", -- t[17988] = 2
      "000010" when "0100011001000101", -- t[17989] = 2
      "000010" when "0100011001000110", -- t[17990] = 2
      "000010" when "0100011001000111", -- t[17991] = 2
      "000010" when "0100011001001000", -- t[17992] = 2
      "000010" when "0100011001001001", -- t[17993] = 2
      "000010" when "0100011001001010", -- t[17994] = 2
      "000010" when "0100011001001011", -- t[17995] = 2
      "000010" when "0100011001001100", -- t[17996] = 2
      "000010" when "0100011001001101", -- t[17997] = 2
      "000010" when "0100011001001110", -- t[17998] = 2
      "000010" when "0100011001001111", -- t[17999] = 2
      "000010" when "0100011001010000", -- t[18000] = 2
      "000010" when "0100011001010001", -- t[18001] = 2
      "000010" when "0100011001010010", -- t[18002] = 2
      "000010" when "0100011001010011", -- t[18003] = 2
      "000010" when "0100011001010100", -- t[18004] = 2
      "000010" when "0100011001010101", -- t[18005] = 2
      "000010" when "0100011001010110", -- t[18006] = 2
      "000010" when "0100011001010111", -- t[18007] = 2
      "000010" when "0100011001011000", -- t[18008] = 2
      "000010" when "0100011001011001", -- t[18009] = 2
      "000010" when "0100011001011010", -- t[18010] = 2
      "000010" when "0100011001011011", -- t[18011] = 2
      "000010" when "0100011001011100", -- t[18012] = 2
      "000010" when "0100011001011101", -- t[18013] = 2
      "000010" when "0100011001011110", -- t[18014] = 2
      "000010" when "0100011001011111", -- t[18015] = 2
      "000010" when "0100011001100000", -- t[18016] = 2
      "000010" when "0100011001100001", -- t[18017] = 2
      "000010" when "0100011001100010", -- t[18018] = 2
      "000010" when "0100011001100011", -- t[18019] = 2
      "000010" when "0100011001100100", -- t[18020] = 2
      "000010" when "0100011001100101", -- t[18021] = 2
      "000010" when "0100011001100110", -- t[18022] = 2
      "000010" when "0100011001100111", -- t[18023] = 2
      "000010" when "0100011001101000", -- t[18024] = 2
      "000010" when "0100011001101001", -- t[18025] = 2
      "000010" when "0100011001101010", -- t[18026] = 2
      "000010" when "0100011001101011", -- t[18027] = 2
      "000010" when "0100011001101100", -- t[18028] = 2
      "000010" when "0100011001101101", -- t[18029] = 2
      "000010" when "0100011001101110", -- t[18030] = 2
      "000010" when "0100011001101111", -- t[18031] = 2
      "000010" when "0100011001110000", -- t[18032] = 2
      "000010" when "0100011001110001", -- t[18033] = 2
      "000010" when "0100011001110010", -- t[18034] = 2
      "000010" when "0100011001110011", -- t[18035] = 2
      "000010" when "0100011001110100", -- t[18036] = 2
      "000010" when "0100011001110101", -- t[18037] = 2
      "000010" when "0100011001110110", -- t[18038] = 2
      "000010" when "0100011001110111", -- t[18039] = 2
      "000010" when "0100011001111000", -- t[18040] = 2
      "000010" when "0100011001111001", -- t[18041] = 2
      "000010" when "0100011001111010", -- t[18042] = 2
      "000010" when "0100011001111011", -- t[18043] = 2
      "000010" when "0100011001111100", -- t[18044] = 2
      "000010" when "0100011001111101", -- t[18045] = 2
      "000010" when "0100011001111110", -- t[18046] = 2
      "000010" when "0100011001111111", -- t[18047] = 2
      "000010" when "0100011010000000", -- t[18048] = 2
      "000010" when "0100011010000001", -- t[18049] = 2
      "000010" when "0100011010000010", -- t[18050] = 2
      "000010" when "0100011010000011", -- t[18051] = 2
      "000010" when "0100011010000100", -- t[18052] = 2
      "000010" when "0100011010000101", -- t[18053] = 2
      "000010" when "0100011010000110", -- t[18054] = 2
      "000010" when "0100011010000111", -- t[18055] = 2
      "000010" when "0100011010001000", -- t[18056] = 2
      "000010" when "0100011010001001", -- t[18057] = 2
      "000010" when "0100011010001010", -- t[18058] = 2
      "000010" when "0100011010001011", -- t[18059] = 2
      "000010" when "0100011010001100", -- t[18060] = 2
      "000010" when "0100011010001101", -- t[18061] = 2
      "000010" when "0100011010001110", -- t[18062] = 2
      "000010" when "0100011010001111", -- t[18063] = 2
      "000010" when "0100011010010000", -- t[18064] = 2
      "000010" when "0100011010010001", -- t[18065] = 2
      "000010" when "0100011010010010", -- t[18066] = 2
      "000010" when "0100011010010011", -- t[18067] = 2
      "000010" when "0100011010010100", -- t[18068] = 2
      "000010" when "0100011010010101", -- t[18069] = 2
      "000010" when "0100011010010110", -- t[18070] = 2
      "000010" when "0100011010010111", -- t[18071] = 2
      "000010" when "0100011010011000", -- t[18072] = 2
      "000010" when "0100011010011001", -- t[18073] = 2
      "000010" when "0100011010011010", -- t[18074] = 2
      "000010" when "0100011010011011", -- t[18075] = 2
      "000010" when "0100011010011100", -- t[18076] = 2
      "000010" when "0100011010011101", -- t[18077] = 2
      "000010" when "0100011010011110", -- t[18078] = 2
      "000010" when "0100011010011111", -- t[18079] = 2
      "000010" when "0100011010100000", -- t[18080] = 2
      "000010" when "0100011010100001", -- t[18081] = 2
      "000010" when "0100011010100010", -- t[18082] = 2
      "000010" when "0100011010100011", -- t[18083] = 2
      "000010" when "0100011010100100", -- t[18084] = 2
      "000010" when "0100011010100101", -- t[18085] = 2
      "000010" when "0100011010100110", -- t[18086] = 2
      "000010" when "0100011010100111", -- t[18087] = 2
      "000010" when "0100011010101000", -- t[18088] = 2
      "000010" when "0100011010101001", -- t[18089] = 2
      "000010" when "0100011010101010", -- t[18090] = 2
      "000010" when "0100011010101011", -- t[18091] = 2
      "000010" when "0100011010101100", -- t[18092] = 2
      "000010" when "0100011010101101", -- t[18093] = 2
      "000010" when "0100011010101110", -- t[18094] = 2
      "000010" when "0100011010101111", -- t[18095] = 2
      "000010" when "0100011010110000", -- t[18096] = 2
      "000010" when "0100011010110001", -- t[18097] = 2
      "000010" when "0100011010110010", -- t[18098] = 2
      "000010" when "0100011010110011", -- t[18099] = 2
      "000010" when "0100011010110100", -- t[18100] = 2
      "000010" when "0100011010110101", -- t[18101] = 2
      "000010" when "0100011010110110", -- t[18102] = 2
      "000010" when "0100011010110111", -- t[18103] = 2
      "000010" when "0100011010111000", -- t[18104] = 2
      "000010" when "0100011010111001", -- t[18105] = 2
      "000010" when "0100011010111010", -- t[18106] = 2
      "000010" when "0100011010111011", -- t[18107] = 2
      "000010" when "0100011010111100", -- t[18108] = 2
      "000010" when "0100011010111101", -- t[18109] = 2
      "000010" when "0100011010111110", -- t[18110] = 2
      "000010" when "0100011010111111", -- t[18111] = 2
      "000010" when "0100011011000000", -- t[18112] = 2
      "000010" when "0100011011000001", -- t[18113] = 2
      "000010" when "0100011011000010", -- t[18114] = 2
      "000010" when "0100011011000011", -- t[18115] = 2
      "000010" when "0100011011000100", -- t[18116] = 2
      "000010" when "0100011011000101", -- t[18117] = 2
      "000010" when "0100011011000110", -- t[18118] = 2
      "000010" when "0100011011000111", -- t[18119] = 2
      "000010" when "0100011011001000", -- t[18120] = 2
      "000010" when "0100011011001001", -- t[18121] = 2
      "000010" when "0100011011001010", -- t[18122] = 2
      "000010" when "0100011011001011", -- t[18123] = 2
      "000010" when "0100011011001100", -- t[18124] = 2
      "000010" when "0100011011001101", -- t[18125] = 2
      "000010" when "0100011011001110", -- t[18126] = 2
      "000010" when "0100011011001111", -- t[18127] = 2
      "000010" when "0100011011010000", -- t[18128] = 2
      "000010" when "0100011011010001", -- t[18129] = 2
      "000010" when "0100011011010010", -- t[18130] = 2
      "000010" when "0100011011010011", -- t[18131] = 2
      "000010" when "0100011011010100", -- t[18132] = 2
      "000010" when "0100011011010101", -- t[18133] = 2
      "000010" when "0100011011010110", -- t[18134] = 2
      "000010" when "0100011011010111", -- t[18135] = 2
      "000010" when "0100011011011000", -- t[18136] = 2
      "000010" when "0100011011011001", -- t[18137] = 2
      "000010" when "0100011011011010", -- t[18138] = 2
      "000010" when "0100011011011011", -- t[18139] = 2
      "000010" when "0100011011011100", -- t[18140] = 2
      "000010" when "0100011011011101", -- t[18141] = 2
      "000010" when "0100011011011110", -- t[18142] = 2
      "000010" when "0100011011011111", -- t[18143] = 2
      "000010" when "0100011011100000", -- t[18144] = 2
      "000010" when "0100011011100001", -- t[18145] = 2
      "000010" when "0100011011100010", -- t[18146] = 2
      "000010" when "0100011011100011", -- t[18147] = 2
      "000010" when "0100011011100100", -- t[18148] = 2
      "000010" when "0100011011100101", -- t[18149] = 2
      "000010" when "0100011011100110", -- t[18150] = 2
      "000010" when "0100011011100111", -- t[18151] = 2
      "000010" when "0100011011101000", -- t[18152] = 2
      "000010" when "0100011011101001", -- t[18153] = 2
      "000010" when "0100011011101010", -- t[18154] = 2
      "000010" when "0100011011101011", -- t[18155] = 2
      "000010" when "0100011011101100", -- t[18156] = 2
      "000010" when "0100011011101101", -- t[18157] = 2
      "000010" when "0100011011101110", -- t[18158] = 2
      "000010" when "0100011011101111", -- t[18159] = 2
      "000010" when "0100011011110000", -- t[18160] = 2
      "000010" when "0100011011110001", -- t[18161] = 2
      "000010" when "0100011011110010", -- t[18162] = 2
      "000010" when "0100011011110011", -- t[18163] = 2
      "000010" when "0100011011110100", -- t[18164] = 2
      "000010" when "0100011011110101", -- t[18165] = 2
      "000010" when "0100011011110110", -- t[18166] = 2
      "000010" when "0100011011110111", -- t[18167] = 2
      "000010" when "0100011011111000", -- t[18168] = 2
      "000010" when "0100011011111001", -- t[18169] = 2
      "000010" when "0100011011111010", -- t[18170] = 2
      "000010" when "0100011011111011", -- t[18171] = 2
      "000010" when "0100011011111100", -- t[18172] = 2
      "000010" when "0100011011111101", -- t[18173] = 2
      "000010" when "0100011011111110", -- t[18174] = 2
      "000010" when "0100011011111111", -- t[18175] = 2
      "000010" when "0100011100000000", -- t[18176] = 2
      "000010" when "0100011100000001", -- t[18177] = 2
      "000010" when "0100011100000010", -- t[18178] = 2
      "000010" when "0100011100000011", -- t[18179] = 2
      "000010" when "0100011100000100", -- t[18180] = 2
      "000010" when "0100011100000101", -- t[18181] = 2
      "000010" when "0100011100000110", -- t[18182] = 2
      "000010" when "0100011100000111", -- t[18183] = 2
      "000010" when "0100011100001000", -- t[18184] = 2
      "000010" when "0100011100001001", -- t[18185] = 2
      "000010" when "0100011100001010", -- t[18186] = 2
      "000010" when "0100011100001011", -- t[18187] = 2
      "000010" when "0100011100001100", -- t[18188] = 2
      "000010" when "0100011100001101", -- t[18189] = 2
      "000010" when "0100011100001110", -- t[18190] = 2
      "000010" when "0100011100001111", -- t[18191] = 2
      "000010" when "0100011100010000", -- t[18192] = 2
      "000010" when "0100011100010001", -- t[18193] = 2
      "000010" when "0100011100010010", -- t[18194] = 2
      "000010" when "0100011100010011", -- t[18195] = 2
      "000010" when "0100011100010100", -- t[18196] = 2
      "000010" when "0100011100010101", -- t[18197] = 2
      "000010" when "0100011100010110", -- t[18198] = 2
      "000010" when "0100011100010111", -- t[18199] = 2
      "000010" when "0100011100011000", -- t[18200] = 2
      "000010" when "0100011100011001", -- t[18201] = 2
      "000010" when "0100011100011010", -- t[18202] = 2
      "000010" when "0100011100011011", -- t[18203] = 2
      "000010" when "0100011100011100", -- t[18204] = 2
      "000010" when "0100011100011101", -- t[18205] = 2
      "000010" when "0100011100011110", -- t[18206] = 2
      "000010" when "0100011100011111", -- t[18207] = 2
      "000010" when "0100011100100000", -- t[18208] = 2
      "000010" when "0100011100100001", -- t[18209] = 2
      "000010" when "0100011100100010", -- t[18210] = 2
      "000010" when "0100011100100011", -- t[18211] = 2
      "000010" when "0100011100100100", -- t[18212] = 2
      "000010" when "0100011100100101", -- t[18213] = 2
      "000010" when "0100011100100110", -- t[18214] = 2
      "000010" when "0100011100100111", -- t[18215] = 2
      "000010" when "0100011100101000", -- t[18216] = 2
      "000010" when "0100011100101001", -- t[18217] = 2
      "000010" when "0100011100101010", -- t[18218] = 2
      "000010" when "0100011100101011", -- t[18219] = 2
      "000010" when "0100011100101100", -- t[18220] = 2
      "000010" when "0100011100101101", -- t[18221] = 2
      "000010" when "0100011100101110", -- t[18222] = 2
      "000010" when "0100011100101111", -- t[18223] = 2
      "000010" when "0100011100110000", -- t[18224] = 2
      "000010" when "0100011100110001", -- t[18225] = 2
      "000010" when "0100011100110010", -- t[18226] = 2
      "000010" when "0100011100110011", -- t[18227] = 2
      "000010" when "0100011100110100", -- t[18228] = 2
      "000010" when "0100011100110101", -- t[18229] = 2
      "000010" when "0100011100110110", -- t[18230] = 2
      "000010" when "0100011100110111", -- t[18231] = 2
      "000010" when "0100011100111000", -- t[18232] = 2
      "000010" when "0100011100111001", -- t[18233] = 2
      "000010" when "0100011100111010", -- t[18234] = 2
      "000010" when "0100011100111011", -- t[18235] = 2
      "000010" when "0100011100111100", -- t[18236] = 2
      "000010" when "0100011100111101", -- t[18237] = 2
      "000010" when "0100011100111110", -- t[18238] = 2
      "000010" when "0100011100111111", -- t[18239] = 2
      "000010" when "0100011101000000", -- t[18240] = 2
      "000010" when "0100011101000001", -- t[18241] = 2
      "000010" when "0100011101000010", -- t[18242] = 2
      "000010" when "0100011101000011", -- t[18243] = 2
      "000010" when "0100011101000100", -- t[18244] = 2
      "000010" when "0100011101000101", -- t[18245] = 2
      "000010" when "0100011101000110", -- t[18246] = 2
      "000010" when "0100011101000111", -- t[18247] = 2
      "000010" when "0100011101001000", -- t[18248] = 2
      "000010" when "0100011101001001", -- t[18249] = 2
      "000010" when "0100011101001010", -- t[18250] = 2
      "000010" when "0100011101001011", -- t[18251] = 2
      "000010" when "0100011101001100", -- t[18252] = 2
      "000010" when "0100011101001101", -- t[18253] = 2
      "000010" when "0100011101001110", -- t[18254] = 2
      "000010" when "0100011101001111", -- t[18255] = 2
      "000010" when "0100011101010000", -- t[18256] = 2
      "000010" when "0100011101010001", -- t[18257] = 2
      "000010" when "0100011101010010", -- t[18258] = 2
      "000010" when "0100011101010011", -- t[18259] = 2
      "000010" when "0100011101010100", -- t[18260] = 2
      "000010" when "0100011101010101", -- t[18261] = 2
      "000010" when "0100011101010110", -- t[18262] = 2
      "000010" when "0100011101010111", -- t[18263] = 2
      "000010" when "0100011101011000", -- t[18264] = 2
      "000010" when "0100011101011001", -- t[18265] = 2
      "000010" when "0100011101011010", -- t[18266] = 2
      "000010" when "0100011101011011", -- t[18267] = 2
      "000010" when "0100011101011100", -- t[18268] = 2
      "000010" when "0100011101011101", -- t[18269] = 2
      "000010" when "0100011101011110", -- t[18270] = 2
      "000010" when "0100011101011111", -- t[18271] = 2
      "000010" when "0100011101100000", -- t[18272] = 2
      "000010" when "0100011101100001", -- t[18273] = 2
      "000010" when "0100011101100010", -- t[18274] = 2
      "000010" when "0100011101100011", -- t[18275] = 2
      "000010" when "0100011101100100", -- t[18276] = 2
      "000010" when "0100011101100101", -- t[18277] = 2
      "000010" when "0100011101100110", -- t[18278] = 2
      "000010" when "0100011101100111", -- t[18279] = 2
      "000010" when "0100011101101000", -- t[18280] = 2
      "000010" when "0100011101101001", -- t[18281] = 2
      "000010" when "0100011101101010", -- t[18282] = 2
      "000010" when "0100011101101011", -- t[18283] = 2
      "000010" when "0100011101101100", -- t[18284] = 2
      "000010" when "0100011101101101", -- t[18285] = 2
      "000010" when "0100011101101110", -- t[18286] = 2
      "000010" when "0100011101101111", -- t[18287] = 2
      "000010" when "0100011101110000", -- t[18288] = 2
      "000010" when "0100011101110001", -- t[18289] = 2
      "000010" when "0100011101110010", -- t[18290] = 2
      "000010" when "0100011101110011", -- t[18291] = 2
      "000010" when "0100011101110100", -- t[18292] = 2
      "000010" when "0100011101110101", -- t[18293] = 2
      "000010" when "0100011101110110", -- t[18294] = 2
      "000010" when "0100011101110111", -- t[18295] = 2
      "000010" when "0100011101111000", -- t[18296] = 2
      "000010" when "0100011101111001", -- t[18297] = 2
      "000010" when "0100011101111010", -- t[18298] = 2
      "000010" when "0100011101111011", -- t[18299] = 2
      "000010" when "0100011101111100", -- t[18300] = 2
      "000010" when "0100011101111101", -- t[18301] = 2
      "000010" when "0100011101111110", -- t[18302] = 2
      "000010" when "0100011101111111", -- t[18303] = 2
      "000010" when "0100011110000000", -- t[18304] = 2
      "000010" when "0100011110000001", -- t[18305] = 2
      "000010" when "0100011110000010", -- t[18306] = 2
      "000010" when "0100011110000011", -- t[18307] = 2
      "000010" when "0100011110000100", -- t[18308] = 2
      "000010" when "0100011110000101", -- t[18309] = 2
      "000010" when "0100011110000110", -- t[18310] = 2
      "000010" when "0100011110000111", -- t[18311] = 2
      "000010" when "0100011110001000", -- t[18312] = 2
      "000010" when "0100011110001001", -- t[18313] = 2
      "000010" when "0100011110001010", -- t[18314] = 2
      "000010" when "0100011110001011", -- t[18315] = 2
      "000010" when "0100011110001100", -- t[18316] = 2
      "000010" when "0100011110001101", -- t[18317] = 2
      "000010" when "0100011110001110", -- t[18318] = 2
      "000010" when "0100011110001111", -- t[18319] = 2
      "000010" when "0100011110010000", -- t[18320] = 2
      "000010" when "0100011110010001", -- t[18321] = 2
      "000010" when "0100011110010010", -- t[18322] = 2
      "000010" when "0100011110010011", -- t[18323] = 2
      "000010" when "0100011110010100", -- t[18324] = 2
      "000010" when "0100011110010101", -- t[18325] = 2
      "000010" when "0100011110010110", -- t[18326] = 2
      "000010" when "0100011110010111", -- t[18327] = 2
      "000010" when "0100011110011000", -- t[18328] = 2
      "000010" when "0100011110011001", -- t[18329] = 2
      "000010" when "0100011110011010", -- t[18330] = 2
      "000010" when "0100011110011011", -- t[18331] = 2
      "000010" when "0100011110011100", -- t[18332] = 2
      "000010" when "0100011110011101", -- t[18333] = 2
      "000010" when "0100011110011110", -- t[18334] = 2
      "000010" when "0100011110011111", -- t[18335] = 2
      "000010" when "0100011110100000", -- t[18336] = 2
      "000010" when "0100011110100001", -- t[18337] = 2
      "000010" when "0100011110100010", -- t[18338] = 2
      "000010" when "0100011110100011", -- t[18339] = 2
      "000010" when "0100011110100100", -- t[18340] = 2
      "000010" when "0100011110100101", -- t[18341] = 2
      "000010" when "0100011110100110", -- t[18342] = 2
      "000010" when "0100011110100111", -- t[18343] = 2
      "000010" when "0100011110101000", -- t[18344] = 2
      "000010" when "0100011110101001", -- t[18345] = 2
      "000010" when "0100011110101010", -- t[18346] = 2
      "000010" when "0100011110101011", -- t[18347] = 2
      "000010" when "0100011110101100", -- t[18348] = 2
      "000010" when "0100011110101101", -- t[18349] = 2
      "000010" when "0100011110101110", -- t[18350] = 2
      "000010" when "0100011110101111", -- t[18351] = 2
      "000010" when "0100011110110000", -- t[18352] = 2
      "000010" when "0100011110110001", -- t[18353] = 2
      "000010" when "0100011110110010", -- t[18354] = 2
      "000010" when "0100011110110011", -- t[18355] = 2
      "000010" when "0100011110110100", -- t[18356] = 2
      "000010" when "0100011110110101", -- t[18357] = 2
      "000010" when "0100011110110110", -- t[18358] = 2
      "000010" when "0100011110110111", -- t[18359] = 2
      "000010" when "0100011110111000", -- t[18360] = 2
      "000010" when "0100011110111001", -- t[18361] = 2
      "000010" when "0100011110111010", -- t[18362] = 2
      "000010" when "0100011110111011", -- t[18363] = 2
      "000010" when "0100011110111100", -- t[18364] = 2
      "000010" when "0100011110111101", -- t[18365] = 2
      "000010" when "0100011110111110", -- t[18366] = 2
      "000010" when "0100011110111111", -- t[18367] = 2
      "000010" when "0100011111000000", -- t[18368] = 2
      "000010" when "0100011111000001", -- t[18369] = 2
      "000010" when "0100011111000010", -- t[18370] = 2
      "000010" when "0100011111000011", -- t[18371] = 2
      "000010" when "0100011111000100", -- t[18372] = 2
      "000010" when "0100011111000101", -- t[18373] = 2
      "000010" when "0100011111000110", -- t[18374] = 2
      "000010" when "0100011111000111", -- t[18375] = 2
      "000010" when "0100011111001000", -- t[18376] = 2
      "000010" when "0100011111001001", -- t[18377] = 2
      "000010" when "0100011111001010", -- t[18378] = 2
      "000010" when "0100011111001011", -- t[18379] = 2
      "000010" when "0100011111001100", -- t[18380] = 2
      "000010" when "0100011111001101", -- t[18381] = 2
      "000010" when "0100011111001110", -- t[18382] = 2
      "000010" when "0100011111001111", -- t[18383] = 2
      "000010" when "0100011111010000", -- t[18384] = 2
      "000010" when "0100011111010001", -- t[18385] = 2
      "000010" when "0100011111010010", -- t[18386] = 2
      "000010" when "0100011111010011", -- t[18387] = 2
      "000010" when "0100011111010100", -- t[18388] = 2
      "000010" when "0100011111010101", -- t[18389] = 2
      "000010" when "0100011111010110", -- t[18390] = 2
      "000010" when "0100011111010111", -- t[18391] = 2
      "000010" when "0100011111011000", -- t[18392] = 2
      "000010" when "0100011111011001", -- t[18393] = 2
      "000010" when "0100011111011010", -- t[18394] = 2
      "000010" when "0100011111011011", -- t[18395] = 2
      "000010" when "0100011111011100", -- t[18396] = 2
      "000010" when "0100011111011101", -- t[18397] = 2
      "000010" when "0100011111011110", -- t[18398] = 2
      "000010" when "0100011111011111", -- t[18399] = 2
      "000010" when "0100011111100000", -- t[18400] = 2
      "000010" when "0100011111100001", -- t[18401] = 2
      "000010" when "0100011111100010", -- t[18402] = 2
      "000010" when "0100011111100011", -- t[18403] = 2
      "000010" when "0100011111100100", -- t[18404] = 2
      "000010" when "0100011111100101", -- t[18405] = 2
      "000010" when "0100011111100110", -- t[18406] = 2
      "000010" when "0100011111100111", -- t[18407] = 2
      "000010" when "0100011111101000", -- t[18408] = 2
      "000010" when "0100011111101001", -- t[18409] = 2
      "000010" when "0100011111101010", -- t[18410] = 2
      "000010" when "0100011111101011", -- t[18411] = 2
      "000010" when "0100011111101100", -- t[18412] = 2
      "000010" when "0100011111101101", -- t[18413] = 2
      "000010" when "0100011111101110", -- t[18414] = 2
      "000010" when "0100011111101111", -- t[18415] = 2
      "000010" when "0100011111110000", -- t[18416] = 2
      "000010" when "0100011111110001", -- t[18417] = 2
      "000010" when "0100011111110010", -- t[18418] = 2
      "000010" when "0100011111110011", -- t[18419] = 2
      "000010" when "0100011111110100", -- t[18420] = 2
      "000010" when "0100011111110101", -- t[18421] = 2
      "000010" when "0100011111110110", -- t[18422] = 2
      "000010" when "0100011111110111", -- t[18423] = 2
      "000010" when "0100011111111000", -- t[18424] = 2
      "000010" when "0100011111111001", -- t[18425] = 2
      "000010" when "0100011111111010", -- t[18426] = 2
      "000010" when "0100011111111011", -- t[18427] = 2
      "000010" when "0100011111111100", -- t[18428] = 2
      "000010" when "0100011111111101", -- t[18429] = 2
      "000010" when "0100011111111110", -- t[18430] = 2
      "000010" when "0100011111111111", -- t[18431] = 2
      "000010" when "0100100000000000", -- t[18432] = 2
      "000010" when "0100100000000001", -- t[18433] = 2
      "000010" when "0100100000000010", -- t[18434] = 2
      "000010" when "0100100000000011", -- t[18435] = 2
      "000010" when "0100100000000100", -- t[18436] = 2
      "000010" when "0100100000000101", -- t[18437] = 2
      "000010" when "0100100000000110", -- t[18438] = 2
      "000010" when "0100100000000111", -- t[18439] = 2
      "000010" when "0100100000001000", -- t[18440] = 2
      "000010" when "0100100000001001", -- t[18441] = 2
      "000010" when "0100100000001010", -- t[18442] = 2
      "000010" when "0100100000001011", -- t[18443] = 2
      "000010" when "0100100000001100", -- t[18444] = 2
      "000010" when "0100100000001101", -- t[18445] = 2
      "000010" when "0100100000001110", -- t[18446] = 2
      "000010" when "0100100000001111", -- t[18447] = 2
      "000010" when "0100100000010000", -- t[18448] = 2
      "000010" when "0100100000010001", -- t[18449] = 2
      "000010" when "0100100000010010", -- t[18450] = 2
      "000010" when "0100100000010011", -- t[18451] = 2
      "000010" when "0100100000010100", -- t[18452] = 2
      "000010" when "0100100000010101", -- t[18453] = 2
      "000010" when "0100100000010110", -- t[18454] = 2
      "000010" when "0100100000010111", -- t[18455] = 2
      "000010" when "0100100000011000", -- t[18456] = 2
      "000010" when "0100100000011001", -- t[18457] = 2
      "000010" when "0100100000011010", -- t[18458] = 2
      "000010" when "0100100000011011", -- t[18459] = 2
      "000010" when "0100100000011100", -- t[18460] = 2
      "000010" when "0100100000011101", -- t[18461] = 2
      "000010" when "0100100000011110", -- t[18462] = 2
      "000010" when "0100100000011111", -- t[18463] = 2
      "000010" when "0100100000100000", -- t[18464] = 2
      "000010" when "0100100000100001", -- t[18465] = 2
      "000010" when "0100100000100010", -- t[18466] = 2
      "000010" when "0100100000100011", -- t[18467] = 2
      "000010" when "0100100000100100", -- t[18468] = 2
      "000010" when "0100100000100101", -- t[18469] = 2
      "000010" when "0100100000100110", -- t[18470] = 2
      "000010" when "0100100000100111", -- t[18471] = 2
      "000010" when "0100100000101000", -- t[18472] = 2
      "000010" when "0100100000101001", -- t[18473] = 2
      "000010" when "0100100000101010", -- t[18474] = 2
      "000010" when "0100100000101011", -- t[18475] = 2
      "000010" when "0100100000101100", -- t[18476] = 2
      "000010" when "0100100000101101", -- t[18477] = 2
      "000010" when "0100100000101110", -- t[18478] = 2
      "000010" when "0100100000101111", -- t[18479] = 2
      "000010" when "0100100000110000", -- t[18480] = 2
      "000010" when "0100100000110001", -- t[18481] = 2
      "000010" when "0100100000110010", -- t[18482] = 2
      "000010" when "0100100000110011", -- t[18483] = 2
      "000010" when "0100100000110100", -- t[18484] = 2
      "000010" when "0100100000110101", -- t[18485] = 2
      "000010" when "0100100000110110", -- t[18486] = 2
      "000010" when "0100100000110111", -- t[18487] = 2
      "000010" when "0100100000111000", -- t[18488] = 2
      "000010" when "0100100000111001", -- t[18489] = 2
      "000010" when "0100100000111010", -- t[18490] = 2
      "000010" when "0100100000111011", -- t[18491] = 2
      "000010" when "0100100000111100", -- t[18492] = 2
      "000010" when "0100100000111101", -- t[18493] = 2
      "000010" when "0100100000111110", -- t[18494] = 2
      "000010" when "0100100000111111", -- t[18495] = 2
      "000010" when "0100100001000000", -- t[18496] = 2
      "000010" when "0100100001000001", -- t[18497] = 2
      "000010" when "0100100001000010", -- t[18498] = 2
      "000010" when "0100100001000011", -- t[18499] = 2
      "000010" when "0100100001000100", -- t[18500] = 2
      "000010" when "0100100001000101", -- t[18501] = 2
      "000010" when "0100100001000110", -- t[18502] = 2
      "000010" when "0100100001000111", -- t[18503] = 2
      "000010" when "0100100001001000", -- t[18504] = 2
      "000010" when "0100100001001001", -- t[18505] = 2
      "000010" when "0100100001001010", -- t[18506] = 2
      "000010" when "0100100001001011", -- t[18507] = 2
      "000010" when "0100100001001100", -- t[18508] = 2
      "000010" when "0100100001001101", -- t[18509] = 2
      "000010" when "0100100001001110", -- t[18510] = 2
      "000010" when "0100100001001111", -- t[18511] = 2
      "000010" when "0100100001010000", -- t[18512] = 2
      "000010" when "0100100001010001", -- t[18513] = 2
      "000010" when "0100100001010010", -- t[18514] = 2
      "000010" when "0100100001010011", -- t[18515] = 2
      "000010" when "0100100001010100", -- t[18516] = 2
      "000010" when "0100100001010101", -- t[18517] = 2
      "000010" when "0100100001010110", -- t[18518] = 2
      "000010" when "0100100001010111", -- t[18519] = 2
      "000010" when "0100100001011000", -- t[18520] = 2
      "000010" when "0100100001011001", -- t[18521] = 2
      "000010" when "0100100001011010", -- t[18522] = 2
      "000010" when "0100100001011011", -- t[18523] = 2
      "000010" when "0100100001011100", -- t[18524] = 2
      "000010" when "0100100001011101", -- t[18525] = 2
      "000010" when "0100100001011110", -- t[18526] = 2
      "000010" when "0100100001011111", -- t[18527] = 2
      "000010" when "0100100001100000", -- t[18528] = 2
      "000010" when "0100100001100001", -- t[18529] = 2
      "000010" when "0100100001100010", -- t[18530] = 2
      "000010" when "0100100001100011", -- t[18531] = 2
      "000010" when "0100100001100100", -- t[18532] = 2
      "000010" when "0100100001100101", -- t[18533] = 2
      "000010" when "0100100001100110", -- t[18534] = 2
      "000010" when "0100100001100111", -- t[18535] = 2
      "000010" when "0100100001101000", -- t[18536] = 2
      "000010" when "0100100001101001", -- t[18537] = 2
      "000010" when "0100100001101010", -- t[18538] = 2
      "000010" when "0100100001101011", -- t[18539] = 2
      "000010" when "0100100001101100", -- t[18540] = 2
      "000010" when "0100100001101101", -- t[18541] = 2
      "000010" when "0100100001101110", -- t[18542] = 2
      "000010" when "0100100001101111", -- t[18543] = 2
      "000010" when "0100100001110000", -- t[18544] = 2
      "000010" when "0100100001110001", -- t[18545] = 2
      "000010" when "0100100001110010", -- t[18546] = 2
      "000010" when "0100100001110011", -- t[18547] = 2
      "000010" when "0100100001110100", -- t[18548] = 2
      "000010" when "0100100001110101", -- t[18549] = 2
      "000010" when "0100100001110110", -- t[18550] = 2
      "000010" when "0100100001110111", -- t[18551] = 2
      "000010" when "0100100001111000", -- t[18552] = 2
      "000010" when "0100100001111001", -- t[18553] = 2
      "000010" when "0100100001111010", -- t[18554] = 2
      "000010" when "0100100001111011", -- t[18555] = 2
      "000010" when "0100100001111100", -- t[18556] = 2
      "000010" when "0100100001111101", -- t[18557] = 2
      "000010" when "0100100001111110", -- t[18558] = 2
      "000010" when "0100100001111111", -- t[18559] = 2
      "000010" when "0100100010000000", -- t[18560] = 2
      "000010" when "0100100010000001", -- t[18561] = 2
      "000010" when "0100100010000010", -- t[18562] = 2
      "000010" when "0100100010000011", -- t[18563] = 2
      "000010" when "0100100010000100", -- t[18564] = 2
      "000010" when "0100100010000101", -- t[18565] = 2
      "000010" when "0100100010000110", -- t[18566] = 2
      "000010" when "0100100010000111", -- t[18567] = 2
      "000010" when "0100100010001000", -- t[18568] = 2
      "000010" when "0100100010001001", -- t[18569] = 2
      "000010" when "0100100010001010", -- t[18570] = 2
      "000010" when "0100100010001011", -- t[18571] = 2
      "000010" when "0100100010001100", -- t[18572] = 2
      "000010" when "0100100010001101", -- t[18573] = 2
      "000010" when "0100100010001110", -- t[18574] = 2
      "000010" when "0100100010001111", -- t[18575] = 2
      "000010" when "0100100010010000", -- t[18576] = 2
      "000010" when "0100100010010001", -- t[18577] = 2
      "000010" when "0100100010010010", -- t[18578] = 2
      "000010" when "0100100010010011", -- t[18579] = 2
      "000010" when "0100100010010100", -- t[18580] = 2
      "000010" when "0100100010010101", -- t[18581] = 2
      "000010" when "0100100010010110", -- t[18582] = 2
      "000010" when "0100100010010111", -- t[18583] = 2
      "000010" when "0100100010011000", -- t[18584] = 2
      "000010" when "0100100010011001", -- t[18585] = 2
      "000010" when "0100100010011010", -- t[18586] = 2
      "000010" when "0100100010011011", -- t[18587] = 2
      "000010" when "0100100010011100", -- t[18588] = 2
      "000010" when "0100100010011101", -- t[18589] = 2
      "000010" when "0100100010011110", -- t[18590] = 2
      "000010" when "0100100010011111", -- t[18591] = 2
      "000010" when "0100100010100000", -- t[18592] = 2
      "000010" when "0100100010100001", -- t[18593] = 2
      "000010" when "0100100010100010", -- t[18594] = 2
      "000010" when "0100100010100011", -- t[18595] = 2
      "000010" when "0100100010100100", -- t[18596] = 2
      "000010" when "0100100010100101", -- t[18597] = 2
      "000010" when "0100100010100110", -- t[18598] = 2
      "000010" when "0100100010100111", -- t[18599] = 2
      "000010" when "0100100010101000", -- t[18600] = 2
      "000010" when "0100100010101001", -- t[18601] = 2
      "000010" when "0100100010101010", -- t[18602] = 2
      "000010" when "0100100010101011", -- t[18603] = 2
      "000010" when "0100100010101100", -- t[18604] = 2
      "000010" when "0100100010101101", -- t[18605] = 2
      "000010" when "0100100010101110", -- t[18606] = 2
      "000010" when "0100100010101111", -- t[18607] = 2
      "000010" when "0100100010110000", -- t[18608] = 2
      "000010" when "0100100010110001", -- t[18609] = 2
      "000010" when "0100100010110010", -- t[18610] = 2
      "000010" when "0100100010110011", -- t[18611] = 2
      "000010" when "0100100010110100", -- t[18612] = 2
      "000010" when "0100100010110101", -- t[18613] = 2
      "000010" when "0100100010110110", -- t[18614] = 2
      "000010" when "0100100010110111", -- t[18615] = 2
      "000010" when "0100100010111000", -- t[18616] = 2
      "000010" when "0100100010111001", -- t[18617] = 2
      "000010" when "0100100010111010", -- t[18618] = 2
      "000010" when "0100100010111011", -- t[18619] = 2
      "000010" when "0100100010111100", -- t[18620] = 2
      "000010" when "0100100010111101", -- t[18621] = 2
      "000010" when "0100100010111110", -- t[18622] = 2
      "000010" when "0100100010111111", -- t[18623] = 2
      "000010" when "0100100011000000", -- t[18624] = 2
      "000010" when "0100100011000001", -- t[18625] = 2
      "000010" when "0100100011000010", -- t[18626] = 2
      "000010" when "0100100011000011", -- t[18627] = 2
      "000010" when "0100100011000100", -- t[18628] = 2
      "000010" when "0100100011000101", -- t[18629] = 2
      "000010" when "0100100011000110", -- t[18630] = 2
      "000010" when "0100100011000111", -- t[18631] = 2
      "000010" when "0100100011001000", -- t[18632] = 2
      "000010" when "0100100011001001", -- t[18633] = 2
      "000010" when "0100100011001010", -- t[18634] = 2
      "000010" when "0100100011001011", -- t[18635] = 2
      "000010" when "0100100011001100", -- t[18636] = 2
      "000010" when "0100100011001101", -- t[18637] = 2
      "000010" when "0100100011001110", -- t[18638] = 2
      "000010" when "0100100011001111", -- t[18639] = 2
      "000010" when "0100100011010000", -- t[18640] = 2
      "000010" when "0100100011010001", -- t[18641] = 2
      "000010" when "0100100011010010", -- t[18642] = 2
      "000010" when "0100100011010011", -- t[18643] = 2
      "000010" when "0100100011010100", -- t[18644] = 2
      "000010" when "0100100011010101", -- t[18645] = 2
      "000010" when "0100100011010110", -- t[18646] = 2
      "000010" when "0100100011010111", -- t[18647] = 2
      "000010" when "0100100011011000", -- t[18648] = 2
      "000010" when "0100100011011001", -- t[18649] = 2
      "000010" when "0100100011011010", -- t[18650] = 2
      "000010" when "0100100011011011", -- t[18651] = 2
      "000010" when "0100100011011100", -- t[18652] = 2
      "000010" when "0100100011011101", -- t[18653] = 2
      "000010" when "0100100011011110", -- t[18654] = 2
      "000010" when "0100100011011111", -- t[18655] = 2
      "000010" when "0100100011100000", -- t[18656] = 2
      "000010" when "0100100011100001", -- t[18657] = 2
      "000010" when "0100100011100010", -- t[18658] = 2
      "000010" when "0100100011100011", -- t[18659] = 2
      "000010" when "0100100011100100", -- t[18660] = 2
      "000010" when "0100100011100101", -- t[18661] = 2
      "000010" when "0100100011100110", -- t[18662] = 2
      "000010" when "0100100011100111", -- t[18663] = 2
      "000010" when "0100100011101000", -- t[18664] = 2
      "000010" when "0100100011101001", -- t[18665] = 2
      "000010" when "0100100011101010", -- t[18666] = 2
      "000010" when "0100100011101011", -- t[18667] = 2
      "000010" when "0100100011101100", -- t[18668] = 2
      "000010" when "0100100011101101", -- t[18669] = 2
      "000010" when "0100100011101110", -- t[18670] = 2
      "000010" when "0100100011101111", -- t[18671] = 2
      "000010" when "0100100011110000", -- t[18672] = 2
      "000010" when "0100100011110001", -- t[18673] = 2
      "000010" when "0100100011110010", -- t[18674] = 2
      "000010" when "0100100011110011", -- t[18675] = 2
      "000010" when "0100100011110100", -- t[18676] = 2
      "000010" when "0100100011110101", -- t[18677] = 2
      "000010" when "0100100011110110", -- t[18678] = 2
      "000010" when "0100100011110111", -- t[18679] = 2
      "000010" when "0100100011111000", -- t[18680] = 2
      "000010" when "0100100011111001", -- t[18681] = 2
      "000010" when "0100100011111010", -- t[18682] = 2
      "000010" when "0100100011111011", -- t[18683] = 2
      "000010" when "0100100011111100", -- t[18684] = 2
      "000010" when "0100100011111101", -- t[18685] = 2
      "000010" when "0100100011111110", -- t[18686] = 2
      "000010" when "0100100011111111", -- t[18687] = 2
      "000010" when "0100100100000000", -- t[18688] = 2
      "000010" when "0100100100000001", -- t[18689] = 2
      "000010" when "0100100100000010", -- t[18690] = 2
      "000010" when "0100100100000011", -- t[18691] = 2
      "000010" when "0100100100000100", -- t[18692] = 2
      "000010" when "0100100100000101", -- t[18693] = 2
      "000010" when "0100100100000110", -- t[18694] = 2
      "000010" when "0100100100000111", -- t[18695] = 2
      "000010" when "0100100100001000", -- t[18696] = 2
      "000010" when "0100100100001001", -- t[18697] = 2
      "000010" when "0100100100001010", -- t[18698] = 2
      "000010" when "0100100100001011", -- t[18699] = 2
      "000010" when "0100100100001100", -- t[18700] = 2
      "000010" when "0100100100001101", -- t[18701] = 2
      "000010" when "0100100100001110", -- t[18702] = 2
      "000010" when "0100100100001111", -- t[18703] = 2
      "000010" when "0100100100010000", -- t[18704] = 2
      "000010" when "0100100100010001", -- t[18705] = 2
      "000010" when "0100100100010010", -- t[18706] = 2
      "000010" when "0100100100010011", -- t[18707] = 2
      "000010" when "0100100100010100", -- t[18708] = 2
      "000010" when "0100100100010101", -- t[18709] = 2
      "000010" when "0100100100010110", -- t[18710] = 2
      "000010" when "0100100100010111", -- t[18711] = 2
      "000010" when "0100100100011000", -- t[18712] = 2
      "000010" when "0100100100011001", -- t[18713] = 2
      "000010" when "0100100100011010", -- t[18714] = 2
      "000010" when "0100100100011011", -- t[18715] = 2
      "000010" when "0100100100011100", -- t[18716] = 2
      "000010" when "0100100100011101", -- t[18717] = 2
      "000010" when "0100100100011110", -- t[18718] = 2
      "000010" when "0100100100011111", -- t[18719] = 2
      "000010" when "0100100100100000", -- t[18720] = 2
      "000010" when "0100100100100001", -- t[18721] = 2
      "000010" when "0100100100100010", -- t[18722] = 2
      "000010" when "0100100100100011", -- t[18723] = 2
      "000010" when "0100100100100100", -- t[18724] = 2
      "000010" when "0100100100100101", -- t[18725] = 2
      "000010" when "0100100100100110", -- t[18726] = 2
      "000010" when "0100100100100111", -- t[18727] = 2
      "000010" when "0100100100101000", -- t[18728] = 2
      "000010" when "0100100100101001", -- t[18729] = 2
      "000010" when "0100100100101010", -- t[18730] = 2
      "000010" when "0100100100101011", -- t[18731] = 2
      "000010" when "0100100100101100", -- t[18732] = 2
      "000010" when "0100100100101101", -- t[18733] = 2
      "000010" when "0100100100101110", -- t[18734] = 2
      "000010" when "0100100100101111", -- t[18735] = 2
      "000010" when "0100100100110000", -- t[18736] = 2
      "000010" when "0100100100110001", -- t[18737] = 2
      "000010" when "0100100100110010", -- t[18738] = 2
      "000010" when "0100100100110011", -- t[18739] = 2
      "000010" when "0100100100110100", -- t[18740] = 2
      "000010" when "0100100100110101", -- t[18741] = 2
      "000010" when "0100100100110110", -- t[18742] = 2
      "000010" when "0100100100110111", -- t[18743] = 2
      "000010" when "0100100100111000", -- t[18744] = 2
      "000010" when "0100100100111001", -- t[18745] = 2
      "000010" when "0100100100111010", -- t[18746] = 2
      "000010" when "0100100100111011", -- t[18747] = 2
      "000010" when "0100100100111100", -- t[18748] = 2
      "000010" when "0100100100111101", -- t[18749] = 2
      "000010" when "0100100100111110", -- t[18750] = 2
      "000010" when "0100100100111111", -- t[18751] = 2
      "000010" when "0100100101000000", -- t[18752] = 2
      "000010" when "0100100101000001", -- t[18753] = 2
      "000010" when "0100100101000010", -- t[18754] = 2
      "000010" when "0100100101000011", -- t[18755] = 2
      "000010" when "0100100101000100", -- t[18756] = 2
      "000010" when "0100100101000101", -- t[18757] = 2
      "000010" when "0100100101000110", -- t[18758] = 2
      "000010" when "0100100101000111", -- t[18759] = 2
      "000010" when "0100100101001000", -- t[18760] = 2
      "000010" when "0100100101001001", -- t[18761] = 2
      "000010" when "0100100101001010", -- t[18762] = 2
      "000010" when "0100100101001011", -- t[18763] = 2
      "000010" when "0100100101001100", -- t[18764] = 2
      "000010" when "0100100101001101", -- t[18765] = 2
      "000010" when "0100100101001110", -- t[18766] = 2
      "000010" when "0100100101001111", -- t[18767] = 2
      "000010" when "0100100101010000", -- t[18768] = 2
      "000010" when "0100100101010001", -- t[18769] = 2
      "000010" when "0100100101010010", -- t[18770] = 2
      "000010" when "0100100101010011", -- t[18771] = 2
      "000010" when "0100100101010100", -- t[18772] = 2
      "000010" when "0100100101010101", -- t[18773] = 2
      "000010" when "0100100101010110", -- t[18774] = 2
      "000010" when "0100100101010111", -- t[18775] = 2
      "000010" when "0100100101011000", -- t[18776] = 2
      "000010" when "0100100101011001", -- t[18777] = 2
      "000010" when "0100100101011010", -- t[18778] = 2
      "000010" when "0100100101011011", -- t[18779] = 2
      "000010" when "0100100101011100", -- t[18780] = 2
      "000010" when "0100100101011101", -- t[18781] = 2
      "000010" when "0100100101011110", -- t[18782] = 2
      "000010" when "0100100101011111", -- t[18783] = 2
      "000010" when "0100100101100000", -- t[18784] = 2
      "000010" when "0100100101100001", -- t[18785] = 2
      "000010" when "0100100101100010", -- t[18786] = 2
      "000010" when "0100100101100011", -- t[18787] = 2
      "000010" when "0100100101100100", -- t[18788] = 2
      "000010" when "0100100101100101", -- t[18789] = 2
      "000010" when "0100100101100110", -- t[18790] = 2
      "000010" when "0100100101100111", -- t[18791] = 2
      "000010" when "0100100101101000", -- t[18792] = 2
      "000010" when "0100100101101001", -- t[18793] = 2
      "000010" when "0100100101101010", -- t[18794] = 2
      "000010" when "0100100101101011", -- t[18795] = 2
      "000010" when "0100100101101100", -- t[18796] = 2
      "000010" when "0100100101101101", -- t[18797] = 2
      "000010" when "0100100101101110", -- t[18798] = 2
      "000010" when "0100100101101111", -- t[18799] = 2
      "000010" when "0100100101110000", -- t[18800] = 2
      "000010" when "0100100101110001", -- t[18801] = 2
      "000010" when "0100100101110010", -- t[18802] = 2
      "000010" when "0100100101110011", -- t[18803] = 2
      "000010" when "0100100101110100", -- t[18804] = 2
      "000010" when "0100100101110101", -- t[18805] = 2
      "000010" when "0100100101110110", -- t[18806] = 2
      "000010" when "0100100101110111", -- t[18807] = 2
      "000010" when "0100100101111000", -- t[18808] = 2
      "000010" when "0100100101111001", -- t[18809] = 2
      "000010" when "0100100101111010", -- t[18810] = 2
      "000010" when "0100100101111011", -- t[18811] = 2
      "000010" when "0100100101111100", -- t[18812] = 2
      "000010" when "0100100101111101", -- t[18813] = 2
      "000010" when "0100100101111110", -- t[18814] = 2
      "000010" when "0100100101111111", -- t[18815] = 2
      "000010" when "0100100110000000", -- t[18816] = 2
      "000010" when "0100100110000001", -- t[18817] = 2
      "000010" when "0100100110000010", -- t[18818] = 2
      "000010" when "0100100110000011", -- t[18819] = 2
      "000010" when "0100100110000100", -- t[18820] = 2
      "000010" when "0100100110000101", -- t[18821] = 2
      "000010" when "0100100110000110", -- t[18822] = 2
      "000010" when "0100100110000111", -- t[18823] = 2
      "000010" when "0100100110001000", -- t[18824] = 2
      "000010" when "0100100110001001", -- t[18825] = 2
      "000010" when "0100100110001010", -- t[18826] = 2
      "000010" when "0100100110001011", -- t[18827] = 2
      "000010" when "0100100110001100", -- t[18828] = 2
      "000010" when "0100100110001101", -- t[18829] = 2
      "000010" when "0100100110001110", -- t[18830] = 2
      "000010" when "0100100110001111", -- t[18831] = 2
      "000010" when "0100100110010000", -- t[18832] = 2
      "000010" when "0100100110010001", -- t[18833] = 2
      "000010" when "0100100110010010", -- t[18834] = 2
      "000010" when "0100100110010011", -- t[18835] = 2
      "000010" when "0100100110010100", -- t[18836] = 2
      "000010" when "0100100110010101", -- t[18837] = 2
      "000010" when "0100100110010110", -- t[18838] = 2
      "000010" when "0100100110010111", -- t[18839] = 2
      "000010" when "0100100110011000", -- t[18840] = 2
      "000010" when "0100100110011001", -- t[18841] = 2
      "000010" when "0100100110011010", -- t[18842] = 2
      "000010" when "0100100110011011", -- t[18843] = 2
      "000010" when "0100100110011100", -- t[18844] = 2
      "000010" when "0100100110011101", -- t[18845] = 2
      "000010" when "0100100110011110", -- t[18846] = 2
      "000010" when "0100100110011111", -- t[18847] = 2
      "000010" when "0100100110100000", -- t[18848] = 2
      "000010" when "0100100110100001", -- t[18849] = 2
      "000010" when "0100100110100010", -- t[18850] = 2
      "000010" when "0100100110100011", -- t[18851] = 2
      "000010" when "0100100110100100", -- t[18852] = 2
      "000010" when "0100100110100101", -- t[18853] = 2
      "000010" when "0100100110100110", -- t[18854] = 2
      "000010" when "0100100110100111", -- t[18855] = 2
      "000010" when "0100100110101000", -- t[18856] = 2
      "000010" when "0100100110101001", -- t[18857] = 2
      "000010" when "0100100110101010", -- t[18858] = 2
      "000010" when "0100100110101011", -- t[18859] = 2
      "000010" when "0100100110101100", -- t[18860] = 2
      "000010" when "0100100110101101", -- t[18861] = 2
      "000010" when "0100100110101110", -- t[18862] = 2
      "000010" when "0100100110101111", -- t[18863] = 2
      "000010" when "0100100110110000", -- t[18864] = 2
      "000010" when "0100100110110001", -- t[18865] = 2
      "000010" when "0100100110110010", -- t[18866] = 2
      "000010" when "0100100110110011", -- t[18867] = 2
      "000010" when "0100100110110100", -- t[18868] = 2
      "000010" when "0100100110110101", -- t[18869] = 2
      "000010" when "0100100110110110", -- t[18870] = 2
      "000010" when "0100100110110111", -- t[18871] = 2
      "000010" when "0100100110111000", -- t[18872] = 2
      "000010" when "0100100110111001", -- t[18873] = 2
      "000010" when "0100100110111010", -- t[18874] = 2
      "000010" when "0100100110111011", -- t[18875] = 2
      "000010" when "0100100110111100", -- t[18876] = 2
      "000010" when "0100100110111101", -- t[18877] = 2
      "000010" when "0100100110111110", -- t[18878] = 2
      "000010" when "0100100110111111", -- t[18879] = 2
      "000010" when "0100100111000000", -- t[18880] = 2
      "000010" when "0100100111000001", -- t[18881] = 2
      "000010" when "0100100111000010", -- t[18882] = 2
      "000010" when "0100100111000011", -- t[18883] = 2
      "000010" when "0100100111000100", -- t[18884] = 2
      "000010" when "0100100111000101", -- t[18885] = 2
      "000010" when "0100100111000110", -- t[18886] = 2
      "000010" when "0100100111000111", -- t[18887] = 2
      "000010" when "0100100111001000", -- t[18888] = 2
      "000010" when "0100100111001001", -- t[18889] = 2
      "000010" when "0100100111001010", -- t[18890] = 2
      "000010" when "0100100111001011", -- t[18891] = 2
      "000010" when "0100100111001100", -- t[18892] = 2
      "000010" when "0100100111001101", -- t[18893] = 2
      "000010" when "0100100111001110", -- t[18894] = 2
      "000010" when "0100100111001111", -- t[18895] = 2
      "000010" when "0100100111010000", -- t[18896] = 2
      "000010" when "0100100111010001", -- t[18897] = 2
      "000010" when "0100100111010010", -- t[18898] = 2
      "000010" when "0100100111010011", -- t[18899] = 2
      "000010" when "0100100111010100", -- t[18900] = 2
      "000010" when "0100100111010101", -- t[18901] = 2
      "000010" when "0100100111010110", -- t[18902] = 2
      "000010" when "0100100111010111", -- t[18903] = 2
      "000010" when "0100100111011000", -- t[18904] = 2
      "000010" when "0100100111011001", -- t[18905] = 2
      "000010" when "0100100111011010", -- t[18906] = 2
      "000010" when "0100100111011011", -- t[18907] = 2
      "000010" when "0100100111011100", -- t[18908] = 2
      "000010" when "0100100111011101", -- t[18909] = 2
      "000010" when "0100100111011110", -- t[18910] = 2
      "000010" when "0100100111011111", -- t[18911] = 2
      "000010" when "0100100111100000", -- t[18912] = 2
      "000010" when "0100100111100001", -- t[18913] = 2
      "000010" when "0100100111100010", -- t[18914] = 2
      "000010" when "0100100111100011", -- t[18915] = 2
      "000010" when "0100100111100100", -- t[18916] = 2
      "000010" when "0100100111100101", -- t[18917] = 2
      "000010" when "0100100111100110", -- t[18918] = 2
      "000010" when "0100100111100111", -- t[18919] = 2
      "000010" when "0100100111101000", -- t[18920] = 2
      "000010" when "0100100111101001", -- t[18921] = 2
      "000010" when "0100100111101010", -- t[18922] = 2
      "000010" when "0100100111101011", -- t[18923] = 2
      "000010" when "0100100111101100", -- t[18924] = 2
      "000010" when "0100100111101101", -- t[18925] = 2
      "000010" when "0100100111101110", -- t[18926] = 2
      "000010" when "0100100111101111", -- t[18927] = 2
      "000010" when "0100100111110000", -- t[18928] = 2
      "000010" when "0100100111110001", -- t[18929] = 2
      "000010" when "0100100111110010", -- t[18930] = 2
      "000010" when "0100100111110011", -- t[18931] = 2
      "000010" when "0100100111110100", -- t[18932] = 2
      "000010" when "0100100111110101", -- t[18933] = 2
      "000010" when "0100100111110110", -- t[18934] = 2
      "000010" when "0100100111110111", -- t[18935] = 2
      "000010" when "0100100111111000", -- t[18936] = 2
      "000010" when "0100100111111001", -- t[18937] = 2
      "000010" when "0100100111111010", -- t[18938] = 2
      "000010" when "0100100111111011", -- t[18939] = 2
      "000010" when "0100100111111100", -- t[18940] = 2
      "000010" when "0100100111111101", -- t[18941] = 2
      "000010" when "0100100111111110", -- t[18942] = 2
      "000010" when "0100100111111111", -- t[18943] = 2
      "000010" when "0100101000000000", -- t[18944] = 2
      "000010" when "0100101000000001", -- t[18945] = 2
      "000010" when "0100101000000010", -- t[18946] = 2
      "000010" when "0100101000000011", -- t[18947] = 2
      "000010" when "0100101000000100", -- t[18948] = 2
      "000010" when "0100101000000101", -- t[18949] = 2
      "000010" when "0100101000000110", -- t[18950] = 2
      "000010" when "0100101000000111", -- t[18951] = 2
      "000010" when "0100101000001000", -- t[18952] = 2
      "000010" when "0100101000001001", -- t[18953] = 2
      "000010" when "0100101000001010", -- t[18954] = 2
      "000010" when "0100101000001011", -- t[18955] = 2
      "000010" when "0100101000001100", -- t[18956] = 2
      "000010" when "0100101000001101", -- t[18957] = 2
      "000010" when "0100101000001110", -- t[18958] = 2
      "000010" when "0100101000001111", -- t[18959] = 2
      "000010" when "0100101000010000", -- t[18960] = 2
      "000010" when "0100101000010001", -- t[18961] = 2
      "000010" when "0100101000010010", -- t[18962] = 2
      "000010" when "0100101000010011", -- t[18963] = 2
      "000010" when "0100101000010100", -- t[18964] = 2
      "000010" when "0100101000010101", -- t[18965] = 2
      "000010" when "0100101000010110", -- t[18966] = 2
      "000010" when "0100101000010111", -- t[18967] = 2
      "000010" when "0100101000011000", -- t[18968] = 2
      "000010" when "0100101000011001", -- t[18969] = 2
      "000010" when "0100101000011010", -- t[18970] = 2
      "000010" when "0100101000011011", -- t[18971] = 2
      "000010" when "0100101000011100", -- t[18972] = 2
      "000010" when "0100101000011101", -- t[18973] = 2
      "000010" when "0100101000011110", -- t[18974] = 2
      "000010" when "0100101000011111", -- t[18975] = 2
      "000010" when "0100101000100000", -- t[18976] = 2
      "000010" when "0100101000100001", -- t[18977] = 2
      "000010" when "0100101000100010", -- t[18978] = 2
      "000010" when "0100101000100011", -- t[18979] = 2
      "000010" when "0100101000100100", -- t[18980] = 2
      "000010" when "0100101000100101", -- t[18981] = 2
      "000010" when "0100101000100110", -- t[18982] = 2
      "000010" when "0100101000100111", -- t[18983] = 2
      "000010" when "0100101000101000", -- t[18984] = 2
      "000010" when "0100101000101001", -- t[18985] = 2
      "000010" when "0100101000101010", -- t[18986] = 2
      "000010" when "0100101000101011", -- t[18987] = 2
      "000010" when "0100101000101100", -- t[18988] = 2
      "000010" when "0100101000101101", -- t[18989] = 2
      "000010" when "0100101000101110", -- t[18990] = 2
      "000010" when "0100101000101111", -- t[18991] = 2
      "000010" when "0100101000110000", -- t[18992] = 2
      "000010" when "0100101000110001", -- t[18993] = 2
      "000010" when "0100101000110010", -- t[18994] = 2
      "000010" when "0100101000110011", -- t[18995] = 2
      "000010" when "0100101000110100", -- t[18996] = 2
      "000010" when "0100101000110101", -- t[18997] = 2
      "000010" when "0100101000110110", -- t[18998] = 2
      "000010" when "0100101000110111", -- t[18999] = 2
      "000010" when "0100101000111000", -- t[19000] = 2
      "000010" when "0100101000111001", -- t[19001] = 2
      "000010" when "0100101000111010", -- t[19002] = 2
      "000010" when "0100101000111011", -- t[19003] = 2
      "000010" when "0100101000111100", -- t[19004] = 2
      "000010" when "0100101000111101", -- t[19005] = 2
      "000010" when "0100101000111110", -- t[19006] = 2
      "000010" when "0100101000111111", -- t[19007] = 2
      "000010" when "0100101001000000", -- t[19008] = 2
      "000010" when "0100101001000001", -- t[19009] = 2
      "000010" when "0100101001000010", -- t[19010] = 2
      "000010" when "0100101001000011", -- t[19011] = 2
      "000010" when "0100101001000100", -- t[19012] = 2
      "000010" when "0100101001000101", -- t[19013] = 2
      "000010" when "0100101001000110", -- t[19014] = 2
      "000010" when "0100101001000111", -- t[19015] = 2
      "000010" when "0100101001001000", -- t[19016] = 2
      "000010" when "0100101001001001", -- t[19017] = 2
      "000010" when "0100101001001010", -- t[19018] = 2
      "000010" when "0100101001001011", -- t[19019] = 2
      "000010" when "0100101001001100", -- t[19020] = 2
      "000010" when "0100101001001101", -- t[19021] = 2
      "000010" when "0100101001001110", -- t[19022] = 2
      "000010" when "0100101001001111", -- t[19023] = 2
      "000010" when "0100101001010000", -- t[19024] = 2
      "000010" when "0100101001010001", -- t[19025] = 2
      "000010" when "0100101001010010", -- t[19026] = 2
      "000010" when "0100101001010011", -- t[19027] = 2
      "000010" when "0100101001010100", -- t[19028] = 2
      "000010" when "0100101001010101", -- t[19029] = 2
      "000010" when "0100101001010110", -- t[19030] = 2
      "000010" when "0100101001010111", -- t[19031] = 2
      "000010" when "0100101001011000", -- t[19032] = 2
      "000010" when "0100101001011001", -- t[19033] = 2
      "000010" when "0100101001011010", -- t[19034] = 2
      "000010" when "0100101001011011", -- t[19035] = 2
      "000010" when "0100101001011100", -- t[19036] = 2
      "000010" when "0100101001011101", -- t[19037] = 2
      "000010" when "0100101001011110", -- t[19038] = 2
      "000010" when "0100101001011111", -- t[19039] = 2
      "000010" when "0100101001100000", -- t[19040] = 2
      "000010" when "0100101001100001", -- t[19041] = 2
      "000010" when "0100101001100010", -- t[19042] = 2
      "000010" when "0100101001100011", -- t[19043] = 2
      "000010" when "0100101001100100", -- t[19044] = 2
      "000010" when "0100101001100101", -- t[19045] = 2
      "000010" when "0100101001100110", -- t[19046] = 2
      "000010" when "0100101001100111", -- t[19047] = 2
      "000010" when "0100101001101000", -- t[19048] = 2
      "000010" when "0100101001101001", -- t[19049] = 2
      "000010" when "0100101001101010", -- t[19050] = 2
      "000010" when "0100101001101011", -- t[19051] = 2
      "000010" when "0100101001101100", -- t[19052] = 2
      "000010" when "0100101001101101", -- t[19053] = 2
      "000010" when "0100101001101110", -- t[19054] = 2
      "000010" when "0100101001101111", -- t[19055] = 2
      "000010" when "0100101001110000", -- t[19056] = 2
      "000010" when "0100101001110001", -- t[19057] = 2
      "000010" when "0100101001110010", -- t[19058] = 2
      "000010" when "0100101001110011", -- t[19059] = 2
      "000010" when "0100101001110100", -- t[19060] = 2
      "000010" when "0100101001110101", -- t[19061] = 2
      "000010" when "0100101001110110", -- t[19062] = 2
      "000010" when "0100101001110111", -- t[19063] = 2
      "000010" when "0100101001111000", -- t[19064] = 2
      "000010" when "0100101001111001", -- t[19065] = 2
      "000010" when "0100101001111010", -- t[19066] = 2
      "000010" when "0100101001111011", -- t[19067] = 2
      "000010" when "0100101001111100", -- t[19068] = 2
      "000010" when "0100101001111101", -- t[19069] = 2
      "000010" when "0100101001111110", -- t[19070] = 2
      "000010" when "0100101001111111", -- t[19071] = 2
      "000010" when "0100101010000000", -- t[19072] = 2
      "000010" when "0100101010000001", -- t[19073] = 2
      "000010" when "0100101010000010", -- t[19074] = 2
      "000010" when "0100101010000011", -- t[19075] = 2
      "000010" when "0100101010000100", -- t[19076] = 2
      "000010" when "0100101010000101", -- t[19077] = 2
      "000010" when "0100101010000110", -- t[19078] = 2
      "000010" when "0100101010000111", -- t[19079] = 2
      "000010" when "0100101010001000", -- t[19080] = 2
      "000010" when "0100101010001001", -- t[19081] = 2
      "000010" when "0100101010001010", -- t[19082] = 2
      "000010" when "0100101010001011", -- t[19083] = 2
      "000010" when "0100101010001100", -- t[19084] = 2
      "000010" when "0100101010001101", -- t[19085] = 2
      "000010" when "0100101010001110", -- t[19086] = 2
      "000010" when "0100101010001111", -- t[19087] = 2
      "000010" when "0100101010010000", -- t[19088] = 2
      "000010" when "0100101010010001", -- t[19089] = 2
      "000010" when "0100101010010010", -- t[19090] = 2
      "000010" when "0100101010010011", -- t[19091] = 2
      "000010" when "0100101010010100", -- t[19092] = 2
      "000010" when "0100101010010101", -- t[19093] = 2
      "000010" when "0100101010010110", -- t[19094] = 2
      "000010" when "0100101010010111", -- t[19095] = 2
      "000010" when "0100101010011000", -- t[19096] = 2
      "000010" when "0100101010011001", -- t[19097] = 2
      "000010" when "0100101010011010", -- t[19098] = 2
      "000010" when "0100101010011011", -- t[19099] = 2
      "000010" when "0100101010011100", -- t[19100] = 2
      "000010" when "0100101010011101", -- t[19101] = 2
      "000010" when "0100101010011110", -- t[19102] = 2
      "000010" when "0100101010011111", -- t[19103] = 2
      "000010" when "0100101010100000", -- t[19104] = 2
      "000010" when "0100101010100001", -- t[19105] = 2
      "000010" when "0100101010100010", -- t[19106] = 2
      "000010" when "0100101010100011", -- t[19107] = 2
      "000010" when "0100101010100100", -- t[19108] = 2
      "000010" when "0100101010100101", -- t[19109] = 2
      "000010" when "0100101010100110", -- t[19110] = 2
      "000010" when "0100101010100111", -- t[19111] = 2
      "000010" when "0100101010101000", -- t[19112] = 2
      "000010" when "0100101010101001", -- t[19113] = 2
      "000010" when "0100101010101010", -- t[19114] = 2
      "000010" when "0100101010101011", -- t[19115] = 2
      "000010" when "0100101010101100", -- t[19116] = 2
      "000010" when "0100101010101101", -- t[19117] = 2
      "000010" when "0100101010101110", -- t[19118] = 2
      "000010" when "0100101010101111", -- t[19119] = 2
      "000010" when "0100101010110000", -- t[19120] = 2
      "000010" when "0100101010110001", -- t[19121] = 2
      "000010" when "0100101010110010", -- t[19122] = 2
      "000010" when "0100101010110011", -- t[19123] = 2
      "000010" when "0100101010110100", -- t[19124] = 2
      "000010" when "0100101010110101", -- t[19125] = 2
      "000010" when "0100101010110110", -- t[19126] = 2
      "000010" when "0100101010110111", -- t[19127] = 2
      "000010" when "0100101010111000", -- t[19128] = 2
      "000010" when "0100101010111001", -- t[19129] = 2
      "000010" when "0100101010111010", -- t[19130] = 2
      "000010" when "0100101010111011", -- t[19131] = 2
      "000010" when "0100101010111100", -- t[19132] = 2
      "000010" when "0100101010111101", -- t[19133] = 2
      "000010" when "0100101010111110", -- t[19134] = 2
      "000010" when "0100101010111111", -- t[19135] = 2
      "000010" when "0100101011000000", -- t[19136] = 2
      "000010" when "0100101011000001", -- t[19137] = 2
      "000010" when "0100101011000010", -- t[19138] = 2
      "000010" when "0100101011000011", -- t[19139] = 2
      "000010" when "0100101011000100", -- t[19140] = 2
      "000010" when "0100101011000101", -- t[19141] = 2
      "000010" when "0100101011000110", -- t[19142] = 2
      "000010" when "0100101011000111", -- t[19143] = 2
      "000010" when "0100101011001000", -- t[19144] = 2
      "000010" when "0100101011001001", -- t[19145] = 2
      "000010" when "0100101011001010", -- t[19146] = 2
      "000010" when "0100101011001011", -- t[19147] = 2
      "000010" when "0100101011001100", -- t[19148] = 2
      "000010" when "0100101011001101", -- t[19149] = 2
      "000010" when "0100101011001110", -- t[19150] = 2
      "000010" when "0100101011001111", -- t[19151] = 2
      "000010" when "0100101011010000", -- t[19152] = 2
      "000010" when "0100101011010001", -- t[19153] = 2
      "000010" when "0100101011010010", -- t[19154] = 2
      "000010" when "0100101011010011", -- t[19155] = 2
      "000010" when "0100101011010100", -- t[19156] = 2
      "000010" when "0100101011010101", -- t[19157] = 2
      "000010" when "0100101011010110", -- t[19158] = 2
      "000010" when "0100101011010111", -- t[19159] = 2
      "000010" when "0100101011011000", -- t[19160] = 2
      "000010" when "0100101011011001", -- t[19161] = 2
      "000010" when "0100101011011010", -- t[19162] = 2
      "000010" when "0100101011011011", -- t[19163] = 2
      "000010" when "0100101011011100", -- t[19164] = 2
      "000010" when "0100101011011101", -- t[19165] = 2
      "000010" when "0100101011011110", -- t[19166] = 2
      "000010" when "0100101011011111", -- t[19167] = 2
      "000010" when "0100101011100000", -- t[19168] = 2
      "000010" when "0100101011100001", -- t[19169] = 2
      "000010" when "0100101011100010", -- t[19170] = 2
      "000010" when "0100101011100011", -- t[19171] = 2
      "000010" when "0100101011100100", -- t[19172] = 2
      "000010" when "0100101011100101", -- t[19173] = 2
      "000010" when "0100101011100110", -- t[19174] = 2
      "000010" when "0100101011100111", -- t[19175] = 2
      "000010" when "0100101011101000", -- t[19176] = 2
      "000010" when "0100101011101001", -- t[19177] = 2
      "000010" when "0100101011101010", -- t[19178] = 2
      "000010" when "0100101011101011", -- t[19179] = 2
      "000010" when "0100101011101100", -- t[19180] = 2
      "000010" when "0100101011101101", -- t[19181] = 2
      "000010" when "0100101011101110", -- t[19182] = 2
      "000010" when "0100101011101111", -- t[19183] = 2
      "000010" when "0100101011110000", -- t[19184] = 2
      "000010" when "0100101011110001", -- t[19185] = 2
      "000010" when "0100101011110010", -- t[19186] = 2
      "000010" when "0100101011110011", -- t[19187] = 2
      "000010" when "0100101011110100", -- t[19188] = 2
      "000010" when "0100101011110101", -- t[19189] = 2
      "000010" when "0100101011110110", -- t[19190] = 2
      "000010" when "0100101011110111", -- t[19191] = 2
      "000010" when "0100101011111000", -- t[19192] = 2
      "000010" when "0100101011111001", -- t[19193] = 2
      "000010" when "0100101011111010", -- t[19194] = 2
      "000010" when "0100101011111011", -- t[19195] = 2
      "000010" when "0100101011111100", -- t[19196] = 2
      "000010" when "0100101011111101", -- t[19197] = 2
      "000010" when "0100101011111110", -- t[19198] = 2
      "000010" when "0100101011111111", -- t[19199] = 2
      "000010" when "0100101100000000", -- t[19200] = 2
      "000010" when "0100101100000001", -- t[19201] = 2
      "000010" when "0100101100000010", -- t[19202] = 2
      "000010" when "0100101100000011", -- t[19203] = 2
      "000010" when "0100101100000100", -- t[19204] = 2
      "000010" when "0100101100000101", -- t[19205] = 2
      "000010" when "0100101100000110", -- t[19206] = 2
      "000010" when "0100101100000111", -- t[19207] = 2
      "000010" when "0100101100001000", -- t[19208] = 2
      "000010" when "0100101100001001", -- t[19209] = 2
      "000010" when "0100101100001010", -- t[19210] = 2
      "000010" when "0100101100001011", -- t[19211] = 2
      "000010" when "0100101100001100", -- t[19212] = 2
      "000010" when "0100101100001101", -- t[19213] = 2
      "000010" when "0100101100001110", -- t[19214] = 2
      "000010" when "0100101100001111", -- t[19215] = 2
      "000010" when "0100101100010000", -- t[19216] = 2
      "000010" when "0100101100010001", -- t[19217] = 2
      "000010" when "0100101100010010", -- t[19218] = 2
      "000010" when "0100101100010011", -- t[19219] = 2
      "000010" when "0100101100010100", -- t[19220] = 2
      "000010" when "0100101100010101", -- t[19221] = 2
      "000010" when "0100101100010110", -- t[19222] = 2
      "000010" when "0100101100010111", -- t[19223] = 2
      "000010" when "0100101100011000", -- t[19224] = 2
      "000010" when "0100101100011001", -- t[19225] = 2
      "000010" when "0100101100011010", -- t[19226] = 2
      "000010" when "0100101100011011", -- t[19227] = 2
      "000010" when "0100101100011100", -- t[19228] = 2
      "000010" when "0100101100011101", -- t[19229] = 2
      "000010" when "0100101100011110", -- t[19230] = 2
      "000010" when "0100101100011111", -- t[19231] = 2
      "000010" when "0100101100100000", -- t[19232] = 2
      "000010" when "0100101100100001", -- t[19233] = 2
      "000010" when "0100101100100010", -- t[19234] = 2
      "000010" when "0100101100100011", -- t[19235] = 2
      "000010" when "0100101100100100", -- t[19236] = 2
      "000010" when "0100101100100101", -- t[19237] = 2
      "000010" when "0100101100100110", -- t[19238] = 2
      "000010" when "0100101100100111", -- t[19239] = 2
      "000010" when "0100101100101000", -- t[19240] = 2
      "000010" when "0100101100101001", -- t[19241] = 2
      "000010" when "0100101100101010", -- t[19242] = 2
      "000010" when "0100101100101011", -- t[19243] = 2
      "000010" when "0100101100101100", -- t[19244] = 2
      "000010" when "0100101100101101", -- t[19245] = 2
      "000010" when "0100101100101110", -- t[19246] = 2
      "000010" when "0100101100101111", -- t[19247] = 2
      "000010" when "0100101100110000", -- t[19248] = 2
      "000010" when "0100101100110001", -- t[19249] = 2
      "000010" when "0100101100110010", -- t[19250] = 2
      "000010" when "0100101100110011", -- t[19251] = 2
      "000010" when "0100101100110100", -- t[19252] = 2
      "000010" when "0100101100110101", -- t[19253] = 2
      "000010" when "0100101100110110", -- t[19254] = 2
      "000010" when "0100101100110111", -- t[19255] = 2
      "000010" when "0100101100111000", -- t[19256] = 2
      "000010" when "0100101100111001", -- t[19257] = 2
      "000010" when "0100101100111010", -- t[19258] = 2
      "000010" when "0100101100111011", -- t[19259] = 2
      "000010" when "0100101100111100", -- t[19260] = 2
      "000010" when "0100101100111101", -- t[19261] = 2
      "000010" when "0100101100111110", -- t[19262] = 2
      "000010" when "0100101100111111", -- t[19263] = 2
      "000010" when "0100101101000000", -- t[19264] = 2
      "000010" when "0100101101000001", -- t[19265] = 2
      "000010" when "0100101101000010", -- t[19266] = 2
      "000010" when "0100101101000011", -- t[19267] = 2
      "000010" when "0100101101000100", -- t[19268] = 2
      "000010" when "0100101101000101", -- t[19269] = 2
      "000010" when "0100101101000110", -- t[19270] = 2
      "000010" when "0100101101000111", -- t[19271] = 2
      "000010" when "0100101101001000", -- t[19272] = 2
      "000010" when "0100101101001001", -- t[19273] = 2
      "000010" when "0100101101001010", -- t[19274] = 2
      "000010" when "0100101101001011", -- t[19275] = 2
      "000010" when "0100101101001100", -- t[19276] = 2
      "000010" when "0100101101001101", -- t[19277] = 2
      "000010" when "0100101101001110", -- t[19278] = 2
      "000010" when "0100101101001111", -- t[19279] = 2
      "000010" when "0100101101010000", -- t[19280] = 2
      "000010" when "0100101101010001", -- t[19281] = 2
      "000010" when "0100101101010010", -- t[19282] = 2
      "000010" when "0100101101010011", -- t[19283] = 2
      "000010" when "0100101101010100", -- t[19284] = 2
      "000010" when "0100101101010101", -- t[19285] = 2
      "000010" when "0100101101010110", -- t[19286] = 2
      "000010" when "0100101101010111", -- t[19287] = 2
      "000010" when "0100101101011000", -- t[19288] = 2
      "000010" when "0100101101011001", -- t[19289] = 2
      "000010" when "0100101101011010", -- t[19290] = 2
      "000010" when "0100101101011011", -- t[19291] = 2
      "000010" when "0100101101011100", -- t[19292] = 2
      "000010" when "0100101101011101", -- t[19293] = 2
      "000010" when "0100101101011110", -- t[19294] = 2
      "000010" when "0100101101011111", -- t[19295] = 2
      "000010" when "0100101101100000", -- t[19296] = 2
      "000010" when "0100101101100001", -- t[19297] = 2
      "000010" when "0100101101100010", -- t[19298] = 2
      "000010" when "0100101101100011", -- t[19299] = 2
      "000010" when "0100101101100100", -- t[19300] = 2
      "000010" when "0100101101100101", -- t[19301] = 2
      "000010" when "0100101101100110", -- t[19302] = 2
      "000010" when "0100101101100111", -- t[19303] = 2
      "000010" when "0100101101101000", -- t[19304] = 2
      "000010" when "0100101101101001", -- t[19305] = 2
      "000010" when "0100101101101010", -- t[19306] = 2
      "000010" when "0100101101101011", -- t[19307] = 2
      "000010" when "0100101101101100", -- t[19308] = 2
      "000010" when "0100101101101101", -- t[19309] = 2
      "000010" when "0100101101101110", -- t[19310] = 2
      "000010" when "0100101101101111", -- t[19311] = 2
      "000010" when "0100101101110000", -- t[19312] = 2
      "000010" when "0100101101110001", -- t[19313] = 2
      "000010" when "0100101101110010", -- t[19314] = 2
      "000010" when "0100101101110011", -- t[19315] = 2
      "000010" when "0100101101110100", -- t[19316] = 2
      "000010" when "0100101101110101", -- t[19317] = 2
      "000010" when "0100101101110110", -- t[19318] = 2
      "000010" when "0100101101110111", -- t[19319] = 2
      "000010" when "0100101101111000", -- t[19320] = 2
      "000010" when "0100101101111001", -- t[19321] = 2
      "000010" when "0100101101111010", -- t[19322] = 2
      "000010" when "0100101101111011", -- t[19323] = 2
      "000010" when "0100101101111100", -- t[19324] = 2
      "000010" when "0100101101111101", -- t[19325] = 2
      "000010" when "0100101101111110", -- t[19326] = 2
      "000010" when "0100101101111111", -- t[19327] = 2
      "000010" when "0100101110000000", -- t[19328] = 2
      "000010" when "0100101110000001", -- t[19329] = 2
      "000010" when "0100101110000010", -- t[19330] = 2
      "000010" when "0100101110000011", -- t[19331] = 2
      "000010" when "0100101110000100", -- t[19332] = 2
      "000010" when "0100101110000101", -- t[19333] = 2
      "000010" when "0100101110000110", -- t[19334] = 2
      "000010" when "0100101110000111", -- t[19335] = 2
      "000010" when "0100101110001000", -- t[19336] = 2
      "000010" when "0100101110001001", -- t[19337] = 2
      "000010" when "0100101110001010", -- t[19338] = 2
      "000010" when "0100101110001011", -- t[19339] = 2
      "000010" when "0100101110001100", -- t[19340] = 2
      "000010" when "0100101110001101", -- t[19341] = 2
      "000010" when "0100101110001110", -- t[19342] = 2
      "000010" when "0100101110001111", -- t[19343] = 2
      "000010" when "0100101110010000", -- t[19344] = 2
      "000010" when "0100101110010001", -- t[19345] = 2
      "000010" when "0100101110010010", -- t[19346] = 2
      "000010" when "0100101110010011", -- t[19347] = 2
      "000010" when "0100101110010100", -- t[19348] = 2
      "000010" when "0100101110010101", -- t[19349] = 2
      "000010" when "0100101110010110", -- t[19350] = 2
      "000010" when "0100101110010111", -- t[19351] = 2
      "000010" when "0100101110011000", -- t[19352] = 2
      "000010" when "0100101110011001", -- t[19353] = 2
      "000010" when "0100101110011010", -- t[19354] = 2
      "000010" when "0100101110011011", -- t[19355] = 2
      "000010" when "0100101110011100", -- t[19356] = 2
      "000010" when "0100101110011101", -- t[19357] = 2
      "000010" when "0100101110011110", -- t[19358] = 2
      "000010" when "0100101110011111", -- t[19359] = 2
      "000010" when "0100101110100000", -- t[19360] = 2
      "000010" when "0100101110100001", -- t[19361] = 2
      "000010" when "0100101110100010", -- t[19362] = 2
      "000010" when "0100101110100011", -- t[19363] = 2
      "000010" when "0100101110100100", -- t[19364] = 2
      "000010" when "0100101110100101", -- t[19365] = 2
      "000010" when "0100101110100110", -- t[19366] = 2
      "000010" when "0100101110100111", -- t[19367] = 2
      "000010" when "0100101110101000", -- t[19368] = 2
      "000010" when "0100101110101001", -- t[19369] = 2
      "000010" when "0100101110101010", -- t[19370] = 2
      "000010" when "0100101110101011", -- t[19371] = 2
      "000010" when "0100101110101100", -- t[19372] = 2
      "000010" when "0100101110101101", -- t[19373] = 2
      "000010" when "0100101110101110", -- t[19374] = 2
      "000010" when "0100101110101111", -- t[19375] = 2
      "000010" when "0100101110110000", -- t[19376] = 2
      "000010" when "0100101110110001", -- t[19377] = 2
      "000010" when "0100101110110010", -- t[19378] = 2
      "000010" when "0100101110110011", -- t[19379] = 2
      "000010" when "0100101110110100", -- t[19380] = 2
      "000010" when "0100101110110101", -- t[19381] = 2
      "000010" when "0100101110110110", -- t[19382] = 2
      "000010" when "0100101110110111", -- t[19383] = 2
      "000010" when "0100101110111000", -- t[19384] = 2
      "000010" when "0100101110111001", -- t[19385] = 2
      "000010" when "0100101110111010", -- t[19386] = 2
      "000010" when "0100101110111011", -- t[19387] = 2
      "000010" when "0100101110111100", -- t[19388] = 2
      "000010" when "0100101110111101", -- t[19389] = 2
      "000010" when "0100101110111110", -- t[19390] = 2
      "000010" when "0100101110111111", -- t[19391] = 2
      "000010" when "0100101111000000", -- t[19392] = 2
      "000010" when "0100101111000001", -- t[19393] = 2
      "000010" when "0100101111000010", -- t[19394] = 2
      "000010" when "0100101111000011", -- t[19395] = 2
      "000010" when "0100101111000100", -- t[19396] = 2
      "000010" when "0100101111000101", -- t[19397] = 2
      "000010" when "0100101111000110", -- t[19398] = 2
      "000010" when "0100101111000111", -- t[19399] = 2
      "000010" when "0100101111001000", -- t[19400] = 2
      "000010" when "0100101111001001", -- t[19401] = 2
      "000010" when "0100101111001010", -- t[19402] = 2
      "000010" when "0100101111001011", -- t[19403] = 2
      "000010" when "0100101111001100", -- t[19404] = 2
      "000010" when "0100101111001101", -- t[19405] = 2
      "000010" when "0100101111001110", -- t[19406] = 2
      "000010" when "0100101111001111", -- t[19407] = 2
      "000010" when "0100101111010000", -- t[19408] = 2
      "000010" when "0100101111010001", -- t[19409] = 2
      "000010" when "0100101111010010", -- t[19410] = 2
      "000010" when "0100101111010011", -- t[19411] = 2
      "000010" when "0100101111010100", -- t[19412] = 2
      "000010" when "0100101111010101", -- t[19413] = 2
      "000010" when "0100101111010110", -- t[19414] = 2
      "000010" when "0100101111010111", -- t[19415] = 2
      "000010" when "0100101111011000", -- t[19416] = 2
      "000010" when "0100101111011001", -- t[19417] = 2
      "000010" when "0100101111011010", -- t[19418] = 2
      "000010" when "0100101111011011", -- t[19419] = 2
      "000010" when "0100101111011100", -- t[19420] = 2
      "000010" when "0100101111011101", -- t[19421] = 2
      "000010" when "0100101111011110", -- t[19422] = 2
      "000010" when "0100101111011111", -- t[19423] = 2
      "000010" when "0100101111100000", -- t[19424] = 2
      "000010" when "0100101111100001", -- t[19425] = 2
      "000010" when "0100101111100010", -- t[19426] = 2
      "000010" when "0100101111100011", -- t[19427] = 2
      "000010" when "0100101111100100", -- t[19428] = 2
      "000010" when "0100101111100101", -- t[19429] = 2
      "000010" when "0100101111100110", -- t[19430] = 2
      "000010" when "0100101111100111", -- t[19431] = 2
      "000010" when "0100101111101000", -- t[19432] = 2
      "000010" when "0100101111101001", -- t[19433] = 2
      "000010" when "0100101111101010", -- t[19434] = 2
      "000010" when "0100101111101011", -- t[19435] = 2
      "000010" when "0100101111101100", -- t[19436] = 2
      "000010" when "0100101111101101", -- t[19437] = 2
      "000010" when "0100101111101110", -- t[19438] = 2
      "000010" when "0100101111101111", -- t[19439] = 2
      "000010" when "0100101111110000", -- t[19440] = 2
      "000010" when "0100101111110001", -- t[19441] = 2
      "000010" when "0100101111110010", -- t[19442] = 2
      "000010" when "0100101111110011", -- t[19443] = 2
      "000010" when "0100101111110100", -- t[19444] = 2
      "000010" when "0100101111110101", -- t[19445] = 2
      "000010" when "0100101111110110", -- t[19446] = 2
      "000010" when "0100101111110111", -- t[19447] = 2
      "000010" when "0100101111111000", -- t[19448] = 2
      "000010" when "0100101111111001", -- t[19449] = 2
      "000010" when "0100101111111010", -- t[19450] = 2
      "000010" when "0100101111111011", -- t[19451] = 2
      "000010" when "0100101111111100", -- t[19452] = 2
      "000010" when "0100101111111101", -- t[19453] = 2
      "000010" when "0100101111111110", -- t[19454] = 2
      "000010" when "0100101111111111", -- t[19455] = 2
      "000010" when "0100110000000000", -- t[19456] = 2
      "000010" when "0100110000000001", -- t[19457] = 2
      "000010" when "0100110000000010", -- t[19458] = 2
      "000010" when "0100110000000011", -- t[19459] = 2
      "000010" when "0100110000000100", -- t[19460] = 2
      "000010" when "0100110000000101", -- t[19461] = 2
      "000010" when "0100110000000110", -- t[19462] = 2
      "000010" when "0100110000000111", -- t[19463] = 2
      "000010" when "0100110000001000", -- t[19464] = 2
      "000010" when "0100110000001001", -- t[19465] = 2
      "000010" when "0100110000001010", -- t[19466] = 2
      "000010" when "0100110000001011", -- t[19467] = 2
      "000010" when "0100110000001100", -- t[19468] = 2
      "000010" when "0100110000001101", -- t[19469] = 2
      "000010" when "0100110000001110", -- t[19470] = 2
      "000010" when "0100110000001111", -- t[19471] = 2
      "000010" when "0100110000010000", -- t[19472] = 2
      "000010" when "0100110000010001", -- t[19473] = 2
      "000010" when "0100110000010010", -- t[19474] = 2
      "000010" when "0100110000010011", -- t[19475] = 2
      "000010" when "0100110000010100", -- t[19476] = 2
      "000010" when "0100110000010101", -- t[19477] = 2
      "000010" when "0100110000010110", -- t[19478] = 2
      "000010" when "0100110000010111", -- t[19479] = 2
      "000010" when "0100110000011000", -- t[19480] = 2
      "000010" when "0100110000011001", -- t[19481] = 2
      "000010" when "0100110000011010", -- t[19482] = 2
      "000010" when "0100110000011011", -- t[19483] = 2
      "000010" when "0100110000011100", -- t[19484] = 2
      "000010" when "0100110000011101", -- t[19485] = 2
      "000010" when "0100110000011110", -- t[19486] = 2
      "000010" when "0100110000011111", -- t[19487] = 2
      "000010" when "0100110000100000", -- t[19488] = 2
      "000010" when "0100110000100001", -- t[19489] = 2
      "000010" when "0100110000100010", -- t[19490] = 2
      "000010" when "0100110000100011", -- t[19491] = 2
      "000010" when "0100110000100100", -- t[19492] = 2
      "000010" when "0100110000100101", -- t[19493] = 2
      "000010" when "0100110000100110", -- t[19494] = 2
      "000010" when "0100110000100111", -- t[19495] = 2
      "000010" when "0100110000101000", -- t[19496] = 2
      "000010" when "0100110000101001", -- t[19497] = 2
      "000010" when "0100110000101010", -- t[19498] = 2
      "000010" when "0100110000101011", -- t[19499] = 2
      "000010" when "0100110000101100", -- t[19500] = 2
      "000010" when "0100110000101101", -- t[19501] = 2
      "000010" when "0100110000101110", -- t[19502] = 2
      "000010" when "0100110000101111", -- t[19503] = 2
      "000010" when "0100110000110000", -- t[19504] = 2
      "000010" when "0100110000110001", -- t[19505] = 2
      "000010" when "0100110000110010", -- t[19506] = 2
      "000010" when "0100110000110011", -- t[19507] = 2
      "000010" when "0100110000110100", -- t[19508] = 2
      "000010" when "0100110000110101", -- t[19509] = 2
      "000010" when "0100110000110110", -- t[19510] = 2
      "000010" when "0100110000110111", -- t[19511] = 2
      "000010" when "0100110000111000", -- t[19512] = 2
      "000010" when "0100110000111001", -- t[19513] = 2
      "000010" when "0100110000111010", -- t[19514] = 2
      "000010" when "0100110000111011", -- t[19515] = 2
      "000010" when "0100110000111100", -- t[19516] = 2
      "000010" when "0100110000111101", -- t[19517] = 2
      "000010" when "0100110000111110", -- t[19518] = 2
      "000010" when "0100110000111111", -- t[19519] = 2
      "000010" when "0100110001000000", -- t[19520] = 2
      "000010" when "0100110001000001", -- t[19521] = 2
      "000010" when "0100110001000010", -- t[19522] = 2
      "000010" when "0100110001000011", -- t[19523] = 2
      "000010" when "0100110001000100", -- t[19524] = 2
      "000010" when "0100110001000101", -- t[19525] = 2
      "000010" when "0100110001000110", -- t[19526] = 2
      "000010" when "0100110001000111", -- t[19527] = 2
      "000010" when "0100110001001000", -- t[19528] = 2
      "000010" when "0100110001001001", -- t[19529] = 2
      "000010" when "0100110001001010", -- t[19530] = 2
      "000010" when "0100110001001011", -- t[19531] = 2
      "000010" when "0100110001001100", -- t[19532] = 2
      "000010" when "0100110001001101", -- t[19533] = 2
      "000010" when "0100110001001110", -- t[19534] = 2
      "000010" when "0100110001001111", -- t[19535] = 2
      "000010" when "0100110001010000", -- t[19536] = 2
      "000010" when "0100110001010001", -- t[19537] = 2
      "000010" when "0100110001010010", -- t[19538] = 2
      "000010" when "0100110001010011", -- t[19539] = 2
      "000010" when "0100110001010100", -- t[19540] = 2
      "000010" when "0100110001010101", -- t[19541] = 2
      "000010" when "0100110001010110", -- t[19542] = 2
      "000010" when "0100110001010111", -- t[19543] = 2
      "000010" when "0100110001011000", -- t[19544] = 2
      "000010" when "0100110001011001", -- t[19545] = 2
      "000010" when "0100110001011010", -- t[19546] = 2
      "000010" when "0100110001011011", -- t[19547] = 2
      "000010" when "0100110001011100", -- t[19548] = 2
      "000010" when "0100110001011101", -- t[19549] = 2
      "000010" when "0100110001011110", -- t[19550] = 2
      "000010" when "0100110001011111", -- t[19551] = 2
      "000010" when "0100110001100000", -- t[19552] = 2
      "000010" when "0100110001100001", -- t[19553] = 2
      "000010" when "0100110001100010", -- t[19554] = 2
      "000010" when "0100110001100011", -- t[19555] = 2
      "000010" when "0100110001100100", -- t[19556] = 2
      "000010" when "0100110001100101", -- t[19557] = 2
      "000010" when "0100110001100110", -- t[19558] = 2
      "000010" when "0100110001100111", -- t[19559] = 2
      "000010" when "0100110001101000", -- t[19560] = 2
      "000010" when "0100110001101001", -- t[19561] = 2
      "000010" when "0100110001101010", -- t[19562] = 2
      "000010" when "0100110001101011", -- t[19563] = 2
      "000010" when "0100110001101100", -- t[19564] = 2
      "000010" when "0100110001101101", -- t[19565] = 2
      "000010" when "0100110001101110", -- t[19566] = 2
      "000010" when "0100110001101111", -- t[19567] = 2
      "000010" when "0100110001110000", -- t[19568] = 2
      "000010" when "0100110001110001", -- t[19569] = 2
      "000010" when "0100110001110010", -- t[19570] = 2
      "000010" when "0100110001110011", -- t[19571] = 2
      "000010" when "0100110001110100", -- t[19572] = 2
      "000010" when "0100110001110101", -- t[19573] = 2
      "000010" when "0100110001110110", -- t[19574] = 2
      "000010" when "0100110001110111", -- t[19575] = 2
      "000010" when "0100110001111000", -- t[19576] = 2
      "000010" when "0100110001111001", -- t[19577] = 2
      "000010" when "0100110001111010", -- t[19578] = 2
      "000010" when "0100110001111011", -- t[19579] = 2
      "000010" when "0100110001111100", -- t[19580] = 2
      "000010" when "0100110001111101", -- t[19581] = 2
      "000010" when "0100110001111110", -- t[19582] = 2
      "000010" when "0100110001111111", -- t[19583] = 2
      "000010" when "0100110010000000", -- t[19584] = 2
      "000010" when "0100110010000001", -- t[19585] = 2
      "000010" when "0100110010000010", -- t[19586] = 2
      "000010" when "0100110010000011", -- t[19587] = 2
      "000010" when "0100110010000100", -- t[19588] = 2
      "000010" when "0100110010000101", -- t[19589] = 2
      "000010" when "0100110010000110", -- t[19590] = 2
      "000010" when "0100110010000111", -- t[19591] = 2
      "000010" when "0100110010001000", -- t[19592] = 2
      "000010" when "0100110010001001", -- t[19593] = 2
      "000010" when "0100110010001010", -- t[19594] = 2
      "000010" when "0100110010001011", -- t[19595] = 2
      "000010" when "0100110010001100", -- t[19596] = 2
      "000010" when "0100110010001101", -- t[19597] = 2
      "000010" when "0100110010001110", -- t[19598] = 2
      "000010" when "0100110010001111", -- t[19599] = 2
      "000010" when "0100110010010000", -- t[19600] = 2
      "000010" when "0100110010010001", -- t[19601] = 2
      "000010" when "0100110010010010", -- t[19602] = 2
      "000010" when "0100110010010011", -- t[19603] = 2
      "000010" when "0100110010010100", -- t[19604] = 2
      "000010" when "0100110010010101", -- t[19605] = 2
      "000010" when "0100110010010110", -- t[19606] = 2
      "000010" when "0100110010010111", -- t[19607] = 2
      "000010" when "0100110010011000", -- t[19608] = 2
      "000010" when "0100110010011001", -- t[19609] = 2
      "000010" when "0100110010011010", -- t[19610] = 2
      "000010" when "0100110010011011", -- t[19611] = 2
      "000010" when "0100110010011100", -- t[19612] = 2
      "000010" when "0100110010011101", -- t[19613] = 2
      "000010" when "0100110010011110", -- t[19614] = 2
      "000010" when "0100110010011111", -- t[19615] = 2
      "000010" when "0100110010100000", -- t[19616] = 2
      "000010" when "0100110010100001", -- t[19617] = 2
      "000010" when "0100110010100010", -- t[19618] = 2
      "000010" when "0100110010100011", -- t[19619] = 2
      "000010" when "0100110010100100", -- t[19620] = 2
      "000010" when "0100110010100101", -- t[19621] = 2
      "000010" when "0100110010100110", -- t[19622] = 2
      "000010" when "0100110010100111", -- t[19623] = 2
      "000010" when "0100110010101000", -- t[19624] = 2
      "000010" when "0100110010101001", -- t[19625] = 2
      "000010" when "0100110010101010", -- t[19626] = 2
      "000010" when "0100110010101011", -- t[19627] = 2
      "000010" when "0100110010101100", -- t[19628] = 2
      "000010" when "0100110010101101", -- t[19629] = 2
      "000010" when "0100110010101110", -- t[19630] = 2
      "000010" when "0100110010101111", -- t[19631] = 2
      "000011" when "0100110010110000", -- t[19632] = 3
      "000011" when "0100110010110001", -- t[19633] = 3
      "000011" when "0100110010110010", -- t[19634] = 3
      "000011" when "0100110010110011", -- t[19635] = 3
      "000011" when "0100110010110100", -- t[19636] = 3
      "000011" when "0100110010110101", -- t[19637] = 3
      "000011" when "0100110010110110", -- t[19638] = 3
      "000011" when "0100110010110111", -- t[19639] = 3
      "000011" when "0100110010111000", -- t[19640] = 3
      "000011" when "0100110010111001", -- t[19641] = 3
      "000011" when "0100110010111010", -- t[19642] = 3
      "000011" when "0100110010111011", -- t[19643] = 3
      "000011" when "0100110010111100", -- t[19644] = 3
      "000011" when "0100110010111101", -- t[19645] = 3
      "000011" when "0100110010111110", -- t[19646] = 3
      "000011" when "0100110010111111", -- t[19647] = 3
      "000011" when "0100110011000000", -- t[19648] = 3
      "000011" when "0100110011000001", -- t[19649] = 3
      "000011" when "0100110011000010", -- t[19650] = 3
      "000011" when "0100110011000011", -- t[19651] = 3
      "000011" when "0100110011000100", -- t[19652] = 3
      "000011" when "0100110011000101", -- t[19653] = 3
      "000011" when "0100110011000110", -- t[19654] = 3
      "000011" when "0100110011000111", -- t[19655] = 3
      "000011" when "0100110011001000", -- t[19656] = 3
      "000011" when "0100110011001001", -- t[19657] = 3
      "000011" when "0100110011001010", -- t[19658] = 3
      "000011" when "0100110011001011", -- t[19659] = 3
      "000011" when "0100110011001100", -- t[19660] = 3
      "000011" when "0100110011001101", -- t[19661] = 3
      "000011" when "0100110011001110", -- t[19662] = 3
      "000011" when "0100110011001111", -- t[19663] = 3
      "000011" when "0100110011010000", -- t[19664] = 3
      "000011" when "0100110011010001", -- t[19665] = 3
      "000011" when "0100110011010010", -- t[19666] = 3
      "000011" when "0100110011010011", -- t[19667] = 3
      "000011" when "0100110011010100", -- t[19668] = 3
      "000011" when "0100110011010101", -- t[19669] = 3
      "000011" when "0100110011010110", -- t[19670] = 3
      "000011" when "0100110011010111", -- t[19671] = 3
      "000011" when "0100110011011000", -- t[19672] = 3
      "000011" when "0100110011011001", -- t[19673] = 3
      "000011" when "0100110011011010", -- t[19674] = 3
      "000011" when "0100110011011011", -- t[19675] = 3
      "000011" when "0100110011011100", -- t[19676] = 3
      "000011" when "0100110011011101", -- t[19677] = 3
      "000011" when "0100110011011110", -- t[19678] = 3
      "000011" when "0100110011011111", -- t[19679] = 3
      "000011" when "0100110011100000", -- t[19680] = 3
      "000011" when "0100110011100001", -- t[19681] = 3
      "000011" when "0100110011100010", -- t[19682] = 3
      "000011" when "0100110011100011", -- t[19683] = 3
      "000011" when "0100110011100100", -- t[19684] = 3
      "000011" when "0100110011100101", -- t[19685] = 3
      "000011" when "0100110011100110", -- t[19686] = 3
      "000011" when "0100110011100111", -- t[19687] = 3
      "000011" when "0100110011101000", -- t[19688] = 3
      "000011" when "0100110011101001", -- t[19689] = 3
      "000011" when "0100110011101010", -- t[19690] = 3
      "000011" when "0100110011101011", -- t[19691] = 3
      "000011" when "0100110011101100", -- t[19692] = 3
      "000011" when "0100110011101101", -- t[19693] = 3
      "000011" when "0100110011101110", -- t[19694] = 3
      "000011" when "0100110011101111", -- t[19695] = 3
      "000011" when "0100110011110000", -- t[19696] = 3
      "000011" when "0100110011110001", -- t[19697] = 3
      "000011" when "0100110011110010", -- t[19698] = 3
      "000011" when "0100110011110011", -- t[19699] = 3
      "000011" when "0100110011110100", -- t[19700] = 3
      "000011" when "0100110011110101", -- t[19701] = 3
      "000011" when "0100110011110110", -- t[19702] = 3
      "000011" when "0100110011110111", -- t[19703] = 3
      "000011" when "0100110011111000", -- t[19704] = 3
      "000011" when "0100110011111001", -- t[19705] = 3
      "000011" when "0100110011111010", -- t[19706] = 3
      "000011" when "0100110011111011", -- t[19707] = 3
      "000011" when "0100110011111100", -- t[19708] = 3
      "000011" when "0100110011111101", -- t[19709] = 3
      "000011" when "0100110011111110", -- t[19710] = 3
      "000011" when "0100110011111111", -- t[19711] = 3
      "000011" when "0100110100000000", -- t[19712] = 3
      "000011" when "0100110100000001", -- t[19713] = 3
      "000011" when "0100110100000010", -- t[19714] = 3
      "000011" when "0100110100000011", -- t[19715] = 3
      "000011" when "0100110100000100", -- t[19716] = 3
      "000011" when "0100110100000101", -- t[19717] = 3
      "000011" when "0100110100000110", -- t[19718] = 3
      "000011" when "0100110100000111", -- t[19719] = 3
      "000011" when "0100110100001000", -- t[19720] = 3
      "000011" when "0100110100001001", -- t[19721] = 3
      "000011" when "0100110100001010", -- t[19722] = 3
      "000011" when "0100110100001011", -- t[19723] = 3
      "000011" when "0100110100001100", -- t[19724] = 3
      "000011" when "0100110100001101", -- t[19725] = 3
      "000011" when "0100110100001110", -- t[19726] = 3
      "000011" when "0100110100001111", -- t[19727] = 3
      "000011" when "0100110100010000", -- t[19728] = 3
      "000011" when "0100110100010001", -- t[19729] = 3
      "000011" when "0100110100010010", -- t[19730] = 3
      "000011" when "0100110100010011", -- t[19731] = 3
      "000011" when "0100110100010100", -- t[19732] = 3
      "000011" when "0100110100010101", -- t[19733] = 3
      "000011" when "0100110100010110", -- t[19734] = 3
      "000011" when "0100110100010111", -- t[19735] = 3
      "000011" when "0100110100011000", -- t[19736] = 3
      "000011" when "0100110100011001", -- t[19737] = 3
      "000011" when "0100110100011010", -- t[19738] = 3
      "000011" when "0100110100011011", -- t[19739] = 3
      "000011" when "0100110100011100", -- t[19740] = 3
      "000011" when "0100110100011101", -- t[19741] = 3
      "000011" when "0100110100011110", -- t[19742] = 3
      "000011" when "0100110100011111", -- t[19743] = 3
      "000011" when "0100110100100000", -- t[19744] = 3
      "000011" when "0100110100100001", -- t[19745] = 3
      "000011" when "0100110100100010", -- t[19746] = 3
      "000011" when "0100110100100011", -- t[19747] = 3
      "000011" when "0100110100100100", -- t[19748] = 3
      "000011" when "0100110100100101", -- t[19749] = 3
      "000011" when "0100110100100110", -- t[19750] = 3
      "000011" when "0100110100100111", -- t[19751] = 3
      "000011" when "0100110100101000", -- t[19752] = 3
      "000011" when "0100110100101001", -- t[19753] = 3
      "000011" when "0100110100101010", -- t[19754] = 3
      "000011" when "0100110100101011", -- t[19755] = 3
      "000011" when "0100110100101100", -- t[19756] = 3
      "000011" when "0100110100101101", -- t[19757] = 3
      "000011" when "0100110100101110", -- t[19758] = 3
      "000011" when "0100110100101111", -- t[19759] = 3
      "000011" when "0100110100110000", -- t[19760] = 3
      "000011" when "0100110100110001", -- t[19761] = 3
      "000011" when "0100110100110010", -- t[19762] = 3
      "000011" when "0100110100110011", -- t[19763] = 3
      "000011" when "0100110100110100", -- t[19764] = 3
      "000011" when "0100110100110101", -- t[19765] = 3
      "000011" when "0100110100110110", -- t[19766] = 3
      "000011" when "0100110100110111", -- t[19767] = 3
      "000011" when "0100110100111000", -- t[19768] = 3
      "000011" when "0100110100111001", -- t[19769] = 3
      "000011" when "0100110100111010", -- t[19770] = 3
      "000011" when "0100110100111011", -- t[19771] = 3
      "000011" when "0100110100111100", -- t[19772] = 3
      "000011" when "0100110100111101", -- t[19773] = 3
      "000011" when "0100110100111110", -- t[19774] = 3
      "000011" when "0100110100111111", -- t[19775] = 3
      "000011" when "0100110101000000", -- t[19776] = 3
      "000011" when "0100110101000001", -- t[19777] = 3
      "000011" when "0100110101000010", -- t[19778] = 3
      "000011" when "0100110101000011", -- t[19779] = 3
      "000011" when "0100110101000100", -- t[19780] = 3
      "000011" when "0100110101000101", -- t[19781] = 3
      "000011" when "0100110101000110", -- t[19782] = 3
      "000011" when "0100110101000111", -- t[19783] = 3
      "000011" when "0100110101001000", -- t[19784] = 3
      "000011" when "0100110101001001", -- t[19785] = 3
      "000011" when "0100110101001010", -- t[19786] = 3
      "000011" when "0100110101001011", -- t[19787] = 3
      "000011" when "0100110101001100", -- t[19788] = 3
      "000011" when "0100110101001101", -- t[19789] = 3
      "000011" when "0100110101001110", -- t[19790] = 3
      "000011" when "0100110101001111", -- t[19791] = 3
      "000011" when "0100110101010000", -- t[19792] = 3
      "000011" when "0100110101010001", -- t[19793] = 3
      "000011" when "0100110101010010", -- t[19794] = 3
      "000011" when "0100110101010011", -- t[19795] = 3
      "000011" when "0100110101010100", -- t[19796] = 3
      "000011" when "0100110101010101", -- t[19797] = 3
      "000011" when "0100110101010110", -- t[19798] = 3
      "000011" when "0100110101010111", -- t[19799] = 3
      "000011" when "0100110101011000", -- t[19800] = 3
      "000011" when "0100110101011001", -- t[19801] = 3
      "000011" when "0100110101011010", -- t[19802] = 3
      "000011" when "0100110101011011", -- t[19803] = 3
      "000011" when "0100110101011100", -- t[19804] = 3
      "000011" when "0100110101011101", -- t[19805] = 3
      "000011" when "0100110101011110", -- t[19806] = 3
      "000011" when "0100110101011111", -- t[19807] = 3
      "000011" when "0100110101100000", -- t[19808] = 3
      "000011" when "0100110101100001", -- t[19809] = 3
      "000011" when "0100110101100010", -- t[19810] = 3
      "000011" when "0100110101100011", -- t[19811] = 3
      "000011" when "0100110101100100", -- t[19812] = 3
      "000011" when "0100110101100101", -- t[19813] = 3
      "000011" when "0100110101100110", -- t[19814] = 3
      "000011" when "0100110101100111", -- t[19815] = 3
      "000011" when "0100110101101000", -- t[19816] = 3
      "000011" when "0100110101101001", -- t[19817] = 3
      "000011" when "0100110101101010", -- t[19818] = 3
      "000011" when "0100110101101011", -- t[19819] = 3
      "000011" when "0100110101101100", -- t[19820] = 3
      "000011" when "0100110101101101", -- t[19821] = 3
      "000011" when "0100110101101110", -- t[19822] = 3
      "000011" when "0100110101101111", -- t[19823] = 3
      "000011" when "0100110101110000", -- t[19824] = 3
      "000011" when "0100110101110001", -- t[19825] = 3
      "000011" when "0100110101110010", -- t[19826] = 3
      "000011" when "0100110101110011", -- t[19827] = 3
      "000011" when "0100110101110100", -- t[19828] = 3
      "000011" when "0100110101110101", -- t[19829] = 3
      "000011" when "0100110101110110", -- t[19830] = 3
      "000011" when "0100110101110111", -- t[19831] = 3
      "000011" when "0100110101111000", -- t[19832] = 3
      "000011" when "0100110101111001", -- t[19833] = 3
      "000011" when "0100110101111010", -- t[19834] = 3
      "000011" when "0100110101111011", -- t[19835] = 3
      "000011" when "0100110101111100", -- t[19836] = 3
      "000011" when "0100110101111101", -- t[19837] = 3
      "000011" when "0100110101111110", -- t[19838] = 3
      "000011" when "0100110101111111", -- t[19839] = 3
      "000011" when "0100110110000000", -- t[19840] = 3
      "000011" when "0100110110000001", -- t[19841] = 3
      "000011" when "0100110110000010", -- t[19842] = 3
      "000011" when "0100110110000011", -- t[19843] = 3
      "000011" when "0100110110000100", -- t[19844] = 3
      "000011" when "0100110110000101", -- t[19845] = 3
      "000011" when "0100110110000110", -- t[19846] = 3
      "000011" when "0100110110000111", -- t[19847] = 3
      "000011" when "0100110110001000", -- t[19848] = 3
      "000011" when "0100110110001001", -- t[19849] = 3
      "000011" when "0100110110001010", -- t[19850] = 3
      "000011" when "0100110110001011", -- t[19851] = 3
      "000011" when "0100110110001100", -- t[19852] = 3
      "000011" when "0100110110001101", -- t[19853] = 3
      "000011" when "0100110110001110", -- t[19854] = 3
      "000011" when "0100110110001111", -- t[19855] = 3
      "000011" when "0100110110010000", -- t[19856] = 3
      "000011" when "0100110110010001", -- t[19857] = 3
      "000011" when "0100110110010010", -- t[19858] = 3
      "000011" when "0100110110010011", -- t[19859] = 3
      "000011" when "0100110110010100", -- t[19860] = 3
      "000011" when "0100110110010101", -- t[19861] = 3
      "000011" when "0100110110010110", -- t[19862] = 3
      "000011" when "0100110110010111", -- t[19863] = 3
      "000011" when "0100110110011000", -- t[19864] = 3
      "000011" when "0100110110011001", -- t[19865] = 3
      "000011" when "0100110110011010", -- t[19866] = 3
      "000011" when "0100110110011011", -- t[19867] = 3
      "000011" when "0100110110011100", -- t[19868] = 3
      "000011" when "0100110110011101", -- t[19869] = 3
      "000011" when "0100110110011110", -- t[19870] = 3
      "000011" when "0100110110011111", -- t[19871] = 3
      "000011" when "0100110110100000", -- t[19872] = 3
      "000011" when "0100110110100001", -- t[19873] = 3
      "000011" when "0100110110100010", -- t[19874] = 3
      "000011" when "0100110110100011", -- t[19875] = 3
      "000011" when "0100110110100100", -- t[19876] = 3
      "000011" when "0100110110100101", -- t[19877] = 3
      "000011" when "0100110110100110", -- t[19878] = 3
      "000011" when "0100110110100111", -- t[19879] = 3
      "000011" when "0100110110101000", -- t[19880] = 3
      "000011" when "0100110110101001", -- t[19881] = 3
      "000011" when "0100110110101010", -- t[19882] = 3
      "000011" when "0100110110101011", -- t[19883] = 3
      "000011" when "0100110110101100", -- t[19884] = 3
      "000011" when "0100110110101101", -- t[19885] = 3
      "000011" when "0100110110101110", -- t[19886] = 3
      "000011" when "0100110110101111", -- t[19887] = 3
      "000011" when "0100110110110000", -- t[19888] = 3
      "000011" when "0100110110110001", -- t[19889] = 3
      "000011" when "0100110110110010", -- t[19890] = 3
      "000011" when "0100110110110011", -- t[19891] = 3
      "000011" when "0100110110110100", -- t[19892] = 3
      "000011" when "0100110110110101", -- t[19893] = 3
      "000011" when "0100110110110110", -- t[19894] = 3
      "000011" when "0100110110110111", -- t[19895] = 3
      "000011" when "0100110110111000", -- t[19896] = 3
      "000011" when "0100110110111001", -- t[19897] = 3
      "000011" when "0100110110111010", -- t[19898] = 3
      "000011" when "0100110110111011", -- t[19899] = 3
      "000011" when "0100110110111100", -- t[19900] = 3
      "000011" when "0100110110111101", -- t[19901] = 3
      "000011" when "0100110110111110", -- t[19902] = 3
      "000011" when "0100110110111111", -- t[19903] = 3
      "000011" when "0100110111000000", -- t[19904] = 3
      "000011" when "0100110111000001", -- t[19905] = 3
      "000011" when "0100110111000010", -- t[19906] = 3
      "000011" when "0100110111000011", -- t[19907] = 3
      "000011" when "0100110111000100", -- t[19908] = 3
      "000011" when "0100110111000101", -- t[19909] = 3
      "000011" when "0100110111000110", -- t[19910] = 3
      "000011" when "0100110111000111", -- t[19911] = 3
      "000011" when "0100110111001000", -- t[19912] = 3
      "000011" when "0100110111001001", -- t[19913] = 3
      "000011" when "0100110111001010", -- t[19914] = 3
      "000011" when "0100110111001011", -- t[19915] = 3
      "000011" when "0100110111001100", -- t[19916] = 3
      "000011" when "0100110111001101", -- t[19917] = 3
      "000011" when "0100110111001110", -- t[19918] = 3
      "000011" when "0100110111001111", -- t[19919] = 3
      "000011" when "0100110111010000", -- t[19920] = 3
      "000011" when "0100110111010001", -- t[19921] = 3
      "000011" when "0100110111010010", -- t[19922] = 3
      "000011" when "0100110111010011", -- t[19923] = 3
      "000011" when "0100110111010100", -- t[19924] = 3
      "000011" when "0100110111010101", -- t[19925] = 3
      "000011" when "0100110111010110", -- t[19926] = 3
      "000011" when "0100110111010111", -- t[19927] = 3
      "000011" when "0100110111011000", -- t[19928] = 3
      "000011" when "0100110111011001", -- t[19929] = 3
      "000011" when "0100110111011010", -- t[19930] = 3
      "000011" when "0100110111011011", -- t[19931] = 3
      "000011" when "0100110111011100", -- t[19932] = 3
      "000011" when "0100110111011101", -- t[19933] = 3
      "000011" when "0100110111011110", -- t[19934] = 3
      "000011" when "0100110111011111", -- t[19935] = 3
      "000011" when "0100110111100000", -- t[19936] = 3
      "000011" when "0100110111100001", -- t[19937] = 3
      "000011" when "0100110111100010", -- t[19938] = 3
      "000011" when "0100110111100011", -- t[19939] = 3
      "000011" when "0100110111100100", -- t[19940] = 3
      "000011" when "0100110111100101", -- t[19941] = 3
      "000011" when "0100110111100110", -- t[19942] = 3
      "000011" when "0100110111100111", -- t[19943] = 3
      "000011" when "0100110111101000", -- t[19944] = 3
      "000011" when "0100110111101001", -- t[19945] = 3
      "000011" when "0100110111101010", -- t[19946] = 3
      "000011" when "0100110111101011", -- t[19947] = 3
      "000011" when "0100110111101100", -- t[19948] = 3
      "000011" when "0100110111101101", -- t[19949] = 3
      "000011" when "0100110111101110", -- t[19950] = 3
      "000011" when "0100110111101111", -- t[19951] = 3
      "000011" when "0100110111110000", -- t[19952] = 3
      "000011" when "0100110111110001", -- t[19953] = 3
      "000011" when "0100110111110010", -- t[19954] = 3
      "000011" when "0100110111110011", -- t[19955] = 3
      "000011" when "0100110111110100", -- t[19956] = 3
      "000011" when "0100110111110101", -- t[19957] = 3
      "000011" when "0100110111110110", -- t[19958] = 3
      "000011" when "0100110111110111", -- t[19959] = 3
      "000011" when "0100110111111000", -- t[19960] = 3
      "000011" when "0100110111111001", -- t[19961] = 3
      "000011" when "0100110111111010", -- t[19962] = 3
      "000011" when "0100110111111011", -- t[19963] = 3
      "000011" when "0100110111111100", -- t[19964] = 3
      "000011" when "0100110111111101", -- t[19965] = 3
      "000011" when "0100110111111110", -- t[19966] = 3
      "000011" when "0100110111111111", -- t[19967] = 3
      "000011" when "0100111000000000", -- t[19968] = 3
      "000011" when "0100111000000001", -- t[19969] = 3
      "000011" when "0100111000000010", -- t[19970] = 3
      "000011" when "0100111000000011", -- t[19971] = 3
      "000011" when "0100111000000100", -- t[19972] = 3
      "000011" when "0100111000000101", -- t[19973] = 3
      "000011" when "0100111000000110", -- t[19974] = 3
      "000011" when "0100111000000111", -- t[19975] = 3
      "000011" when "0100111000001000", -- t[19976] = 3
      "000011" when "0100111000001001", -- t[19977] = 3
      "000011" when "0100111000001010", -- t[19978] = 3
      "000011" when "0100111000001011", -- t[19979] = 3
      "000011" when "0100111000001100", -- t[19980] = 3
      "000011" when "0100111000001101", -- t[19981] = 3
      "000011" when "0100111000001110", -- t[19982] = 3
      "000011" when "0100111000001111", -- t[19983] = 3
      "000011" when "0100111000010000", -- t[19984] = 3
      "000011" when "0100111000010001", -- t[19985] = 3
      "000011" when "0100111000010010", -- t[19986] = 3
      "000011" when "0100111000010011", -- t[19987] = 3
      "000011" when "0100111000010100", -- t[19988] = 3
      "000011" when "0100111000010101", -- t[19989] = 3
      "000011" when "0100111000010110", -- t[19990] = 3
      "000011" when "0100111000010111", -- t[19991] = 3
      "000011" when "0100111000011000", -- t[19992] = 3
      "000011" when "0100111000011001", -- t[19993] = 3
      "000011" when "0100111000011010", -- t[19994] = 3
      "000011" when "0100111000011011", -- t[19995] = 3
      "000011" when "0100111000011100", -- t[19996] = 3
      "000011" when "0100111000011101", -- t[19997] = 3
      "000011" when "0100111000011110", -- t[19998] = 3
      "000011" when "0100111000011111", -- t[19999] = 3
      "000011" when "0100111000100000", -- t[20000] = 3
      "000011" when "0100111000100001", -- t[20001] = 3
      "000011" when "0100111000100010", -- t[20002] = 3
      "000011" when "0100111000100011", -- t[20003] = 3
      "000011" when "0100111000100100", -- t[20004] = 3
      "000011" when "0100111000100101", -- t[20005] = 3
      "000011" when "0100111000100110", -- t[20006] = 3
      "000011" when "0100111000100111", -- t[20007] = 3
      "000011" when "0100111000101000", -- t[20008] = 3
      "000011" when "0100111000101001", -- t[20009] = 3
      "000011" when "0100111000101010", -- t[20010] = 3
      "000011" when "0100111000101011", -- t[20011] = 3
      "000011" when "0100111000101100", -- t[20012] = 3
      "000011" when "0100111000101101", -- t[20013] = 3
      "000011" when "0100111000101110", -- t[20014] = 3
      "000011" when "0100111000101111", -- t[20015] = 3
      "000011" when "0100111000110000", -- t[20016] = 3
      "000011" when "0100111000110001", -- t[20017] = 3
      "000011" when "0100111000110010", -- t[20018] = 3
      "000011" when "0100111000110011", -- t[20019] = 3
      "000011" when "0100111000110100", -- t[20020] = 3
      "000011" when "0100111000110101", -- t[20021] = 3
      "000011" when "0100111000110110", -- t[20022] = 3
      "000011" when "0100111000110111", -- t[20023] = 3
      "000011" when "0100111000111000", -- t[20024] = 3
      "000011" when "0100111000111001", -- t[20025] = 3
      "000011" when "0100111000111010", -- t[20026] = 3
      "000011" when "0100111000111011", -- t[20027] = 3
      "000011" when "0100111000111100", -- t[20028] = 3
      "000011" when "0100111000111101", -- t[20029] = 3
      "000011" when "0100111000111110", -- t[20030] = 3
      "000011" when "0100111000111111", -- t[20031] = 3
      "000011" when "0100111001000000", -- t[20032] = 3
      "000011" when "0100111001000001", -- t[20033] = 3
      "000011" when "0100111001000010", -- t[20034] = 3
      "000011" when "0100111001000011", -- t[20035] = 3
      "000011" when "0100111001000100", -- t[20036] = 3
      "000011" when "0100111001000101", -- t[20037] = 3
      "000011" when "0100111001000110", -- t[20038] = 3
      "000011" when "0100111001000111", -- t[20039] = 3
      "000011" when "0100111001001000", -- t[20040] = 3
      "000011" when "0100111001001001", -- t[20041] = 3
      "000011" when "0100111001001010", -- t[20042] = 3
      "000011" when "0100111001001011", -- t[20043] = 3
      "000011" when "0100111001001100", -- t[20044] = 3
      "000011" when "0100111001001101", -- t[20045] = 3
      "000011" when "0100111001001110", -- t[20046] = 3
      "000011" when "0100111001001111", -- t[20047] = 3
      "000011" when "0100111001010000", -- t[20048] = 3
      "000011" when "0100111001010001", -- t[20049] = 3
      "000011" when "0100111001010010", -- t[20050] = 3
      "000011" when "0100111001010011", -- t[20051] = 3
      "000011" when "0100111001010100", -- t[20052] = 3
      "000011" when "0100111001010101", -- t[20053] = 3
      "000011" when "0100111001010110", -- t[20054] = 3
      "000011" when "0100111001010111", -- t[20055] = 3
      "000011" when "0100111001011000", -- t[20056] = 3
      "000011" when "0100111001011001", -- t[20057] = 3
      "000011" when "0100111001011010", -- t[20058] = 3
      "000011" when "0100111001011011", -- t[20059] = 3
      "000011" when "0100111001011100", -- t[20060] = 3
      "000011" when "0100111001011101", -- t[20061] = 3
      "000011" when "0100111001011110", -- t[20062] = 3
      "000011" when "0100111001011111", -- t[20063] = 3
      "000011" when "0100111001100000", -- t[20064] = 3
      "000011" when "0100111001100001", -- t[20065] = 3
      "000011" when "0100111001100010", -- t[20066] = 3
      "000011" when "0100111001100011", -- t[20067] = 3
      "000011" when "0100111001100100", -- t[20068] = 3
      "000011" when "0100111001100101", -- t[20069] = 3
      "000011" when "0100111001100110", -- t[20070] = 3
      "000011" when "0100111001100111", -- t[20071] = 3
      "000011" when "0100111001101000", -- t[20072] = 3
      "000011" when "0100111001101001", -- t[20073] = 3
      "000011" when "0100111001101010", -- t[20074] = 3
      "000011" when "0100111001101011", -- t[20075] = 3
      "000011" when "0100111001101100", -- t[20076] = 3
      "000011" when "0100111001101101", -- t[20077] = 3
      "000011" when "0100111001101110", -- t[20078] = 3
      "000011" when "0100111001101111", -- t[20079] = 3
      "000011" when "0100111001110000", -- t[20080] = 3
      "000011" when "0100111001110001", -- t[20081] = 3
      "000011" when "0100111001110010", -- t[20082] = 3
      "000011" when "0100111001110011", -- t[20083] = 3
      "000011" when "0100111001110100", -- t[20084] = 3
      "000011" when "0100111001110101", -- t[20085] = 3
      "000011" when "0100111001110110", -- t[20086] = 3
      "000011" when "0100111001110111", -- t[20087] = 3
      "000011" when "0100111001111000", -- t[20088] = 3
      "000011" when "0100111001111001", -- t[20089] = 3
      "000011" when "0100111001111010", -- t[20090] = 3
      "000011" when "0100111001111011", -- t[20091] = 3
      "000011" when "0100111001111100", -- t[20092] = 3
      "000011" when "0100111001111101", -- t[20093] = 3
      "000011" when "0100111001111110", -- t[20094] = 3
      "000011" when "0100111001111111", -- t[20095] = 3
      "000011" when "0100111010000000", -- t[20096] = 3
      "000011" when "0100111010000001", -- t[20097] = 3
      "000011" when "0100111010000010", -- t[20098] = 3
      "000011" when "0100111010000011", -- t[20099] = 3
      "000011" when "0100111010000100", -- t[20100] = 3
      "000011" when "0100111010000101", -- t[20101] = 3
      "000011" when "0100111010000110", -- t[20102] = 3
      "000011" when "0100111010000111", -- t[20103] = 3
      "000011" when "0100111010001000", -- t[20104] = 3
      "000011" when "0100111010001001", -- t[20105] = 3
      "000011" when "0100111010001010", -- t[20106] = 3
      "000011" when "0100111010001011", -- t[20107] = 3
      "000011" when "0100111010001100", -- t[20108] = 3
      "000011" when "0100111010001101", -- t[20109] = 3
      "000011" when "0100111010001110", -- t[20110] = 3
      "000011" when "0100111010001111", -- t[20111] = 3
      "000011" when "0100111010010000", -- t[20112] = 3
      "000011" when "0100111010010001", -- t[20113] = 3
      "000011" when "0100111010010010", -- t[20114] = 3
      "000011" when "0100111010010011", -- t[20115] = 3
      "000011" when "0100111010010100", -- t[20116] = 3
      "000011" when "0100111010010101", -- t[20117] = 3
      "000011" when "0100111010010110", -- t[20118] = 3
      "000011" when "0100111010010111", -- t[20119] = 3
      "000011" when "0100111010011000", -- t[20120] = 3
      "000011" when "0100111010011001", -- t[20121] = 3
      "000011" when "0100111010011010", -- t[20122] = 3
      "000011" when "0100111010011011", -- t[20123] = 3
      "000011" when "0100111010011100", -- t[20124] = 3
      "000011" when "0100111010011101", -- t[20125] = 3
      "000011" when "0100111010011110", -- t[20126] = 3
      "000011" when "0100111010011111", -- t[20127] = 3
      "000011" when "0100111010100000", -- t[20128] = 3
      "000011" when "0100111010100001", -- t[20129] = 3
      "000011" when "0100111010100010", -- t[20130] = 3
      "000011" when "0100111010100011", -- t[20131] = 3
      "000011" when "0100111010100100", -- t[20132] = 3
      "000011" when "0100111010100101", -- t[20133] = 3
      "000011" when "0100111010100110", -- t[20134] = 3
      "000011" when "0100111010100111", -- t[20135] = 3
      "000011" when "0100111010101000", -- t[20136] = 3
      "000011" when "0100111010101001", -- t[20137] = 3
      "000011" when "0100111010101010", -- t[20138] = 3
      "000011" when "0100111010101011", -- t[20139] = 3
      "000011" when "0100111010101100", -- t[20140] = 3
      "000011" when "0100111010101101", -- t[20141] = 3
      "000011" when "0100111010101110", -- t[20142] = 3
      "000011" when "0100111010101111", -- t[20143] = 3
      "000011" when "0100111010110000", -- t[20144] = 3
      "000011" when "0100111010110001", -- t[20145] = 3
      "000011" when "0100111010110010", -- t[20146] = 3
      "000011" when "0100111010110011", -- t[20147] = 3
      "000011" when "0100111010110100", -- t[20148] = 3
      "000011" when "0100111010110101", -- t[20149] = 3
      "000011" when "0100111010110110", -- t[20150] = 3
      "000011" when "0100111010110111", -- t[20151] = 3
      "000011" when "0100111010111000", -- t[20152] = 3
      "000011" when "0100111010111001", -- t[20153] = 3
      "000011" when "0100111010111010", -- t[20154] = 3
      "000011" when "0100111010111011", -- t[20155] = 3
      "000011" when "0100111010111100", -- t[20156] = 3
      "000011" when "0100111010111101", -- t[20157] = 3
      "000011" when "0100111010111110", -- t[20158] = 3
      "000011" when "0100111010111111", -- t[20159] = 3
      "000011" when "0100111011000000", -- t[20160] = 3
      "000011" when "0100111011000001", -- t[20161] = 3
      "000011" when "0100111011000010", -- t[20162] = 3
      "000011" when "0100111011000011", -- t[20163] = 3
      "000011" when "0100111011000100", -- t[20164] = 3
      "000011" when "0100111011000101", -- t[20165] = 3
      "000011" when "0100111011000110", -- t[20166] = 3
      "000011" when "0100111011000111", -- t[20167] = 3
      "000011" when "0100111011001000", -- t[20168] = 3
      "000011" when "0100111011001001", -- t[20169] = 3
      "000011" when "0100111011001010", -- t[20170] = 3
      "000011" when "0100111011001011", -- t[20171] = 3
      "000011" when "0100111011001100", -- t[20172] = 3
      "000011" when "0100111011001101", -- t[20173] = 3
      "000011" when "0100111011001110", -- t[20174] = 3
      "000011" when "0100111011001111", -- t[20175] = 3
      "000011" when "0100111011010000", -- t[20176] = 3
      "000011" when "0100111011010001", -- t[20177] = 3
      "000011" when "0100111011010010", -- t[20178] = 3
      "000011" when "0100111011010011", -- t[20179] = 3
      "000011" when "0100111011010100", -- t[20180] = 3
      "000011" when "0100111011010101", -- t[20181] = 3
      "000011" when "0100111011010110", -- t[20182] = 3
      "000011" when "0100111011010111", -- t[20183] = 3
      "000011" when "0100111011011000", -- t[20184] = 3
      "000011" when "0100111011011001", -- t[20185] = 3
      "000011" when "0100111011011010", -- t[20186] = 3
      "000011" when "0100111011011011", -- t[20187] = 3
      "000011" when "0100111011011100", -- t[20188] = 3
      "000011" when "0100111011011101", -- t[20189] = 3
      "000011" when "0100111011011110", -- t[20190] = 3
      "000011" when "0100111011011111", -- t[20191] = 3
      "000011" when "0100111011100000", -- t[20192] = 3
      "000011" when "0100111011100001", -- t[20193] = 3
      "000011" when "0100111011100010", -- t[20194] = 3
      "000011" when "0100111011100011", -- t[20195] = 3
      "000011" when "0100111011100100", -- t[20196] = 3
      "000011" when "0100111011100101", -- t[20197] = 3
      "000011" when "0100111011100110", -- t[20198] = 3
      "000011" when "0100111011100111", -- t[20199] = 3
      "000011" when "0100111011101000", -- t[20200] = 3
      "000011" when "0100111011101001", -- t[20201] = 3
      "000011" when "0100111011101010", -- t[20202] = 3
      "000011" when "0100111011101011", -- t[20203] = 3
      "000011" when "0100111011101100", -- t[20204] = 3
      "000011" when "0100111011101101", -- t[20205] = 3
      "000011" when "0100111011101110", -- t[20206] = 3
      "000011" when "0100111011101111", -- t[20207] = 3
      "000011" when "0100111011110000", -- t[20208] = 3
      "000011" when "0100111011110001", -- t[20209] = 3
      "000011" when "0100111011110010", -- t[20210] = 3
      "000011" when "0100111011110011", -- t[20211] = 3
      "000011" when "0100111011110100", -- t[20212] = 3
      "000011" when "0100111011110101", -- t[20213] = 3
      "000011" when "0100111011110110", -- t[20214] = 3
      "000011" when "0100111011110111", -- t[20215] = 3
      "000011" when "0100111011111000", -- t[20216] = 3
      "000011" when "0100111011111001", -- t[20217] = 3
      "000011" when "0100111011111010", -- t[20218] = 3
      "000011" when "0100111011111011", -- t[20219] = 3
      "000011" when "0100111011111100", -- t[20220] = 3
      "000011" when "0100111011111101", -- t[20221] = 3
      "000011" when "0100111011111110", -- t[20222] = 3
      "000011" when "0100111011111111", -- t[20223] = 3
      "000011" when "0100111100000000", -- t[20224] = 3
      "000011" when "0100111100000001", -- t[20225] = 3
      "000011" when "0100111100000010", -- t[20226] = 3
      "000011" when "0100111100000011", -- t[20227] = 3
      "000011" when "0100111100000100", -- t[20228] = 3
      "000011" when "0100111100000101", -- t[20229] = 3
      "000011" when "0100111100000110", -- t[20230] = 3
      "000011" when "0100111100000111", -- t[20231] = 3
      "000011" when "0100111100001000", -- t[20232] = 3
      "000011" when "0100111100001001", -- t[20233] = 3
      "000011" when "0100111100001010", -- t[20234] = 3
      "000011" when "0100111100001011", -- t[20235] = 3
      "000011" when "0100111100001100", -- t[20236] = 3
      "000011" when "0100111100001101", -- t[20237] = 3
      "000011" when "0100111100001110", -- t[20238] = 3
      "000011" when "0100111100001111", -- t[20239] = 3
      "000011" when "0100111100010000", -- t[20240] = 3
      "000011" when "0100111100010001", -- t[20241] = 3
      "000011" when "0100111100010010", -- t[20242] = 3
      "000011" when "0100111100010011", -- t[20243] = 3
      "000011" when "0100111100010100", -- t[20244] = 3
      "000011" when "0100111100010101", -- t[20245] = 3
      "000011" when "0100111100010110", -- t[20246] = 3
      "000011" when "0100111100010111", -- t[20247] = 3
      "000011" when "0100111100011000", -- t[20248] = 3
      "000011" when "0100111100011001", -- t[20249] = 3
      "000011" when "0100111100011010", -- t[20250] = 3
      "000011" when "0100111100011011", -- t[20251] = 3
      "000011" when "0100111100011100", -- t[20252] = 3
      "000011" when "0100111100011101", -- t[20253] = 3
      "000011" when "0100111100011110", -- t[20254] = 3
      "000011" when "0100111100011111", -- t[20255] = 3
      "000011" when "0100111100100000", -- t[20256] = 3
      "000011" when "0100111100100001", -- t[20257] = 3
      "000011" when "0100111100100010", -- t[20258] = 3
      "000011" when "0100111100100011", -- t[20259] = 3
      "000011" when "0100111100100100", -- t[20260] = 3
      "000011" when "0100111100100101", -- t[20261] = 3
      "000011" when "0100111100100110", -- t[20262] = 3
      "000011" when "0100111100100111", -- t[20263] = 3
      "000011" when "0100111100101000", -- t[20264] = 3
      "000011" when "0100111100101001", -- t[20265] = 3
      "000011" when "0100111100101010", -- t[20266] = 3
      "000011" when "0100111100101011", -- t[20267] = 3
      "000011" when "0100111100101100", -- t[20268] = 3
      "000011" when "0100111100101101", -- t[20269] = 3
      "000011" when "0100111100101110", -- t[20270] = 3
      "000011" when "0100111100101111", -- t[20271] = 3
      "000011" when "0100111100110000", -- t[20272] = 3
      "000011" when "0100111100110001", -- t[20273] = 3
      "000011" when "0100111100110010", -- t[20274] = 3
      "000011" when "0100111100110011", -- t[20275] = 3
      "000011" when "0100111100110100", -- t[20276] = 3
      "000011" when "0100111100110101", -- t[20277] = 3
      "000011" when "0100111100110110", -- t[20278] = 3
      "000011" when "0100111100110111", -- t[20279] = 3
      "000011" when "0100111100111000", -- t[20280] = 3
      "000011" when "0100111100111001", -- t[20281] = 3
      "000011" when "0100111100111010", -- t[20282] = 3
      "000011" when "0100111100111011", -- t[20283] = 3
      "000011" when "0100111100111100", -- t[20284] = 3
      "000011" when "0100111100111101", -- t[20285] = 3
      "000011" when "0100111100111110", -- t[20286] = 3
      "000011" when "0100111100111111", -- t[20287] = 3
      "000011" when "0100111101000000", -- t[20288] = 3
      "000011" when "0100111101000001", -- t[20289] = 3
      "000011" when "0100111101000010", -- t[20290] = 3
      "000011" when "0100111101000011", -- t[20291] = 3
      "000011" when "0100111101000100", -- t[20292] = 3
      "000011" when "0100111101000101", -- t[20293] = 3
      "000011" when "0100111101000110", -- t[20294] = 3
      "000011" when "0100111101000111", -- t[20295] = 3
      "000011" when "0100111101001000", -- t[20296] = 3
      "000011" when "0100111101001001", -- t[20297] = 3
      "000011" when "0100111101001010", -- t[20298] = 3
      "000011" when "0100111101001011", -- t[20299] = 3
      "000011" when "0100111101001100", -- t[20300] = 3
      "000011" when "0100111101001101", -- t[20301] = 3
      "000011" when "0100111101001110", -- t[20302] = 3
      "000011" when "0100111101001111", -- t[20303] = 3
      "000011" when "0100111101010000", -- t[20304] = 3
      "000011" when "0100111101010001", -- t[20305] = 3
      "000011" when "0100111101010010", -- t[20306] = 3
      "000011" when "0100111101010011", -- t[20307] = 3
      "000011" when "0100111101010100", -- t[20308] = 3
      "000011" when "0100111101010101", -- t[20309] = 3
      "000011" when "0100111101010110", -- t[20310] = 3
      "000011" when "0100111101010111", -- t[20311] = 3
      "000011" when "0100111101011000", -- t[20312] = 3
      "000011" when "0100111101011001", -- t[20313] = 3
      "000011" when "0100111101011010", -- t[20314] = 3
      "000011" when "0100111101011011", -- t[20315] = 3
      "000011" when "0100111101011100", -- t[20316] = 3
      "000011" when "0100111101011101", -- t[20317] = 3
      "000011" when "0100111101011110", -- t[20318] = 3
      "000011" when "0100111101011111", -- t[20319] = 3
      "000011" when "0100111101100000", -- t[20320] = 3
      "000011" when "0100111101100001", -- t[20321] = 3
      "000011" when "0100111101100010", -- t[20322] = 3
      "000011" when "0100111101100011", -- t[20323] = 3
      "000011" when "0100111101100100", -- t[20324] = 3
      "000011" when "0100111101100101", -- t[20325] = 3
      "000011" when "0100111101100110", -- t[20326] = 3
      "000011" when "0100111101100111", -- t[20327] = 3
      "000011" when "0100111101101000", -- t[20328] = 3
      "000011" when "0100111101101001", -- t[20329] = 3
      "000011" when "0100111101101010", -- t[20330] = 3
      "000011" when "0100111101101011", -- t[20331] = 3
      "000011" when "0100111101101100", -- t[20332] = 3
      "000011" when "0100111101101101", -- t[20333] = 3
      "000011" when "0100111101101110", -- t[20334] = 3
      "000011" when "0100111101101111", -- t[20335] = 3
      "000011" when "0100111101110000", -- t[20336] = 3
      "000011" when "0100111101110001", -- t[20337] = 3
      "000011" when "0100111101110010", -- t[20338] = 3
      "000011" when "0100111101110011", -- t[20339] = 3
      "000011" when "0100111101110100", -- t[20340] = 3
      "000011" when "0100111101110101", -- t[20341] = 3
      "000011" when "0100111101110110", -- t[20342] = 3
      "000011" when "0100111101110111", -- t[20343] = 3
      "000011" when "0100111101111000", -- t[20344] = 3
      "000011" when "0100111101111001", -- t[20345] = 3
      "000011" when "0100111101111010", -- t[20346] = 3
      "000011" when "0100111101111011", -- t[20347] = 3
      "000011" when "0100111101111100", -- t[20348] = 3
      "000011" when "0100111101111101", -- t[20349] = 3
      "000011" when "0100111101111110", -- t[20350] = 3
      "000011" when "0100111101111111", -- t[20351] = 3
      "000011" when "0100111110000000", -- t[20352] = 3
      "000011" when "0100111110000001", -- t[20353] = 3
      "000011" when "0100111110000010", -- t[20354] = 3
      "000011" when "0100111110000011", -- t[20355] = 3
      "000011" when "0100111110000100", -- t[20356] = 3
      "000011" when "0100111110000101", -- t[20357] = 3
      "000011" when "0100111110000110", -- t[20358] = 3
      "000011" when "0100111110000111", -- t[20359] = 3
      "000011" when "0100111110001000", -- t[20360] = 3
      "000011" when "0100111110001001", -- t[20361] = 3
      "000011" when "0100111110001010", -- t[20362] = 3
      "000011" when "0100111110001011", -- t[20363] = 3
      "000011" when "0100111110001100", -- t[20364] = 3
      "000011" when "0100111110001101", -- t[20365] = 3
      "000011" when "0100111110001110", -- t[20366] = 3
      "000011" when "0100111110001111", -- t[20367] = 3
      "000011" when "0100111110010000", -- t[20368] = 3
      "000011" when "0100111110010001", -- t[20369] = 3
      "000011" when "0100111110010010", -- t[20370] = 3
      "000011" when "0100111110010011", -- t[20371] = 3
      "000011" when "0100111110010100", -- t[20372] = 3
      "000011" when "0100111110010101", -- t[20373] = 3
      "000011" when "0100111110010110", -- t[20374] = 3
      "000011" when "0100111110010111", -- t[20375] = 3
      "000011" when "0100111110011000", -- t[20376] = 3
      "000011" when "0100111110011001", -- t[20377] = 3
      "000011" when "0100111110011010", -- t[20378] = 3
      "000011" when "0100111110011011", -- t[20379] = 3
      "000011" when "0100111110011100", -- t[20380] = 3
      "000011" when "0100111110011101", -- t[20381] = 3
      "000011" when "0100111110011110", -- t[20382] = 3
      "000011" when "0100111110011111", -- t[20383] = 3
      "000011" when "0100111110100000", -- t[20384] = 3
      "000011" when "0100111110100001", -- t[20385] = 3
      "000011" when "0100111110100010", -- t[20386] = 3
      "000011" when "0100111110100011", -- t[20387] = 3
      "000011" when "0100111110100100", -- t[20388] = 3
      "000011" when "0100111110100101", -- t[20389] = 3
      "000011" when "0100111110100110", -- t[20390] = 3
      "000011" when "0100111110100111", -- t[20391] = 3
      "000011" when "0100111110101000", -- t[20392] = 3
      "000011" when "0100111110101001", -- t[20393] = 3
      "000011" when "0100111110101010", -- t[20394] = 3
      "000011" when "0100111110101011", -- t[20395] = 3
      "000011" when "0100111110101100", -- t[20396] = 3
      "000011" when "0100111110101101", -- t[20397] = 3
      "000011" when "0100111110101110", -- t[20398] = 3
      "000011" when "0100111110101111", -- t[20399] = 3
      "000011" when "0100111110110000", -- t[20400] = 3
      "000011" when "0100111110110001", -- t[20401] = 3
      "000011" when "0100111110110010", -- t[20402] = 3
      "000011" when "0100111110110011", -- t[20403] = 3
      "000011" when "0100111110110100", -- t[20404] = 3
      "000011" when "0100111110110101", -- t[20405] = 3
      "000011" when "0100111110110110", -- t[20406] = 3
      "000011" when "0100111110110111", -- t[20407] = 3
      "000011" when "0100111110111000", -- t[20408] = 3
      "000011" when "0100111110111001", -- t[20409] = 3
      "000011" when "0100111110111010", -- t[20410] = 3
      "000011" when "0100111110111011", -- t[20411] = 3
      "000011" when "0100111110111100", -- t[20412] = 3
      "000011" when "0100111110111101", -- t[20413] = 3
      "000011" when "0100111110111110", -- t[20414] = 3
      "000011" when "0100111110111111", -- t[20415] = 3
      "000011" when "0100111111000000", -- t[20416] = 3
      "000011" when "0100111111000001", -- t[20417] = 3
      "000011" when "0100111111000010", -- t[20418] = 3
      "000011" when "0100111111000011", -- t[20419] = 3
      "000011" when "0100111111000100", -- t[20420] = 3
      "000011" when "0100111111000101", -- t[20421] = 3
      "000011" when "0100111111000110", -- t[20422] = 3
      "000011" when "0100111111000111", -- t[20423] = 3
      "000011" when "0100111111001000", -- t[20424] = 3
      "000011" when "0100111111001001", -- t[20425] = 3
      "000011" when "0100111111001010", -- t[20426] = 3
      "000011" when "0100111111001011", -- t[20427] = 3
      "000011" when "0100111111001100", -- t[20428] = 3
      "000011" when "0100111111001101", -- t[20429] = 3
      "000011" when "0100111111001110", -- t[20430] = 3
      "000011" when "0100111111001111", -- t[20431] = 3
      "000011" when "0100111111010000", -- t[20432] = 3
      "000011" when "0100111111010001", -- t[20433] = 3
      "000011" when "0100111111010010", -- t[20434] = 3
      "000011" when "0100111111010011", -- t[20435] = 3
      "000011" when "0100111111010100", -- t[20436] = 3
      "000011" when "0100111111010101", -- t[20437] = 3
      "000011" when "0100111111010110", -- t[20438] = 3
      "000011" when "0100111111010111", -- t[20439] = 3
      "000011" when "0100111111011000", -- t[20440] = 3
      "000011" when "0100111111011001", -- t[20441] = 3
      "000011" when "0100111111011010", -- t[20442] = 3
      "000011" when "0100111111011011", -- t[20443] = 3
      "000011" when "0100111111011100", -- t[20444] = 3
      "000011" when "0100111111011101", -- t[20445] = 3
      "000011" when "0100111111011110", -- t[20446] = 3
      "000011" when "0100111111011111", -- t[20447] = 3
      "000011" when "0100111111100000", -- t[20448] = 3
      "000011" when "0100111111100001", -- t[20449] = 3
      "000011" when "0100111111100010", -- t[20450] = 3
      "000011" when "0100111111100011", -- t[20451] = 3
      "000011" when "0100111111100100", -- t[20452] = 3
      "000011" when "0100111111100101", -- t[20453] = 3
      "000011" when "0100111111100110", -- t[20454] = 3
      "000011" when "0100111111100111", -- t[20455] = 3
      "000011" when "0100111111101000", -- t[20456] = 3
      "000011" when "0100111111101001", -- t[20457] = 3
      "000011" when "0100111111101010", -- t[20458] = 3
      "000011" when "0100111111101011", -- t[20459] = 3
      "000011" when "0100111111101100", -- t[20460] = 3
      "000011" when "0100111111101101", -- t[20461] = 3
      "000011" when "0100111111101110", -- t[20462] = 3
      "000011" when "0100111111101111", -- t[20463] = 3
      "000011" when "0100111111110000", -- t[20464] = 3
      "000011" when "0100111111110001", -- t[20465] = 3
      "000011" when "0100111111110010", -- t[20466] = 3
      "000011" when "0100111111110011", -- t[20467] = 3
      "000011" when "0100111111110100", -- t[20468] = 3
      "000011" when "0100111111110101", -- t[20469] = 3
      "000011" when "0100111111110110", -- t[20470] = 3
      "000011" when "0100111111110111", -- t[20471] = 3
      "000011" when "0100111111111000", -- t[20472] = 3
      "000011" when "0100111111111001", -- t[20473] = 3
      "000011" when "0100111111111010", -- t[20474] = 3
      "000011" when "0100111111111011", -- t[20475] = 3
      "000011" when "0100111111111100", -- t[20476] = 3
      "000011" when "0100111111111101", -- t[20477] = 3
      "000011" when "0100111111111110", -- t[20478] = 3
      "000011" when "0100111111111111", -- t[20479] = 3
      "000011" when "0101000000000000", -- t[20480] = 3
      "000011" when "0101000000000001", -- t[20481] = 3
      "000011" when "0101000000000010", -- t[20482] = 3
      "000011" when "0101000000000011", -- t[20483] = 3
      "000011" when "0101000000000100", -- t[20484] = 3
      "000011" when "0101000000000101", -- t[20485] = 3
      "000011" when "0101000000000110", -- t[20486] = 3
      "000011" when "0101000000000111", -- t[20487] = 3
      "000011" when "0101000000001000", -- t[20488] = 3
      "000011" when "0101000000001001", -- t[20489] = 3
      "000011" when "0101000000001010", -- t[20490] = 3
      "000011" when "0101000000001011", -- t[20491] = 3
      "000011" when "0101000000001100", -- t[20492] = 3
      "000011" when "0101000000001101", -- t[20493] = 3
      "000011" when "0101000000001110", -- t[20494] = 3
      "000011" when "0101000000001111", -- t[20495] = 3
      "000011" when "0101000000010000", -- t[20496] = 3
      "000011" when "0101000000010001", -- t[20497] = 3
      "000011" when "0101000000010010", -- t[20498] = 3
      "000011" when "0101000000010011", -- t[20499] = 3
      "000011" when "0101000000010100", -- t[20500] = 3
      "000011" when "0101000000010101", -- t[20501] = 3
      "000011" when "0101000000010110", -- t[20502] = 3
      "000011" when "0101000000010111", -- t[20503] = 3
      "000011" when "0101000000011000", -- t[20504] = 3
      "000011" when "0101000000011001", -- t[20505] = 3
      "000011" when "0101000000011010", -- t[20506] = 3
      "000011" when "0101000000011011", -- t[20507] = 3
      "000011" when "0101000000011100", -- t[20508] = 3
      "000011" when "0101000000011101", -- t[20509] = 3
      "000011" when "0101000000011110", -- t[20510] = 3
      "000011" when "0101000000011111", -- t[20511] = 3
      "000011" when "0101000000100000", -- t[20512] = 3
      "000011" when "0101000000100001", -- t[20513] = 3
      "000011" when "0101000000100010", -- t[20514] = 3
      "000011" when "0101000000100011", -- t[20515] = 3
      "000011" when "0101000000100100", -- t[20516] = 3
      "000011" when "0101000000100101", -- t[20517] = 3
      "000011" when "0101000000100110", -- t[20518] = 3
      "000011" when "0101000000100111", -- t[20519] = 3
      "000011" when "0101000000101000", -- t[20520] = 3
      "000011" when "0101000000101001", -- t[20521] = 3
      "000011" when "0101000000101010", -- t[20522] = 3
      "000011" when "0101000000101011", -- t[20523] = 3
      "000011" when "0101000000101100", -- t[20524] = 3
      "000011" when "0101000000101101", -- t[20525] = 3
      "000011" when "0101000000101110", -- t[20526] = 3
      "000011" when "0101000000101111", -- t[20527] = 3
      "000011" when "0101000000110000", -- t[20528] = 3
      "000011" when "0101000000110001", -- t[20529] = 3
      "000011" when "0101000000110010", -- t[20530] = 3
      "000011" when "0101000000110011", -- t[20531] = 3
      "000011" when "0101000000110100", -- t[20532] = 3
      "000011" when "0101000000110101", -- t[20533] = 3
      "000011" when "0101000000110110", -- t[20534] = 3
      "000011" when "0101000000110111", -- t[20535] = 3
      "000011" when "0101000000111000", -- t[20536] = 3
      "000011" when "0101000000111001", -- t[20537] = 3
      "000011" when "0101000000111010", -- t[20538] = 3
      "000011" when "0101000000111011", -- t[20539] = 3
      "000011" when "0101000000111100", -- t[20540] = 3
      "000011" when "0101000000111101", -- t[20541] = 3
      "000011" when "0101000000111110", -- t[20542] = 3
      "000011" when "0101000000111111", -- t[20543] = 3
      "000011" when "0101000001000000", -- t[20544] = 3
      "000011" when "0101000001000001", -- t[20545] = 3
      "000011" when "0101000001000010", -- t[20546] = 3
      "000011" when "0101000001000011", -- t[20547] = 3
      "000011" when "0101000001000100", -- t[20548] = 3
      "000011" when "0101000001000101", -- t[20549] = 3
      "000011" when "0101000001000110", -- t[20550] = 3
      "000011" when "0101000001000111", -- t[20551] = 3
      "000011" when "0101000001001000", -- t[20552] = 3
      "000011" when "0101000001001001", -- t[20553] = 3
      "000011" when "0101000001001010", -- t[20554] = 3
      "000011" when "0101000001001011", -- t[20555] = 3
      "000011" when "0101000001001100", -- t[20556] = 3
      "000011" when "0101000001001101", -- t[20557] = 3
      "000011" when "0101000001001110", -- t[20558] = 3
      "000011" when "0101000001001111", -- t[20559] = 3
      "000011" when "0101000001010000", -- t[20560] = 3
      "000011" when "0101000001010001", -- t[20561] = 3
      "000011" when "0101000001010010", -- t[20562] = 3
      "000011" when "0101000001010011", -- t[20563] = 3
      "000011" when "0101000001010100", -- t[20564] = 3
      "000011" when "0101000001010101", -- t[20565] = 3
      "000011" when "0101000001010110", -- t[20566] = 3
      "000011" when "0101000001010111", -- t[20567] = 3
      "000011" when "0101000001011000", -- t[20568] = 3
      "000011" when "0101000001011001", -- t[20569] = 3
      "000011" when "0101000001011010", -- t[20570] = 3
      "000011" when "0101000001011011", -- t[20571] = 3
      "000011" when "0101000001011100", -- t[20572] = 3
      "000011" when "0101000001011101", -- t[20573] = 3
      "000011" when "0101000001011110", -- t[20574] = 3
      "000011" when "0101000001011111", -- t[20575] = 3
      "000011" when "0101000001100000", -- t[20576] = 3
      "000011" when "0101000001100001", -- t[20577] = 3
      "000011" when "0101000001100010", -- t[20578] = 3
      "000011" when "0101000001100011", -- t[20579] = 3
      "000011" when "0101000001100100", -- t[20580] = 3
      "000011" when "0101000001100101", -- t[20581] = 3
      "000011" when "0101000001100110", -- t[20582] = 3
      "000011" when "0101000001100111", -- t[20583] = 3
      "000011" when "0101000001101000", -- t[20584] = 3
      "000011" when "0101000001101001", -- t[20585] = 3
      "000011" when "0101000001101010", -- t[20586] = 3
      "000011" when "0101000001101011", -- t[20587] = 3
      "000011" when "0101000001101100", -- t[20588] = 3
      "000011" when "0101000001101101", -- t[20589] = 3
      "000011" when "0101000001101110", -- t[20590] = 3
      "000011" when "0101000001101111", -- t[20591] = 3
      "000011" when "0101000001110000", -- t[20592] = 3
      "000011" when "0101000001110001", -- t[20593] = 3
      "000011" when "0101000001110010", -- t[20594] = 3
      "000011" when "0101000001110011", -- t[20595] = 3
      "000011" when "0101000001110100", -- t[20596] = 3
      "000011" when "0101000001110101", -- t[20597] = 3
      "000011" when "0101000001110110", -- t[20598] = 3
      "000011" when "0101000001110111", -- t[20599] = 3
      "000011" when "0101000001111000", -- t[20600] = 3
      "000011" when "0101000001111001", -- t[20601] = 3
      "000011" when "0101000001111010", -- t[20602] = 3
      "000011" when "0101000001111011", -- t[20603] = 3
      "000011" when "0101000001111100", -- t[20604] = 3
      "000011" when "0101000001111101", -- t[20605] = 3
      "000011" when "0101000001111110", -- t[20606] = 3
      "000011" when "0101000001111111", -- t[20607] = 3
      "000011" when "0101000010000000", -- t[20608] = 3
      "000011" when "0101000010000001", -- t[20609] = 3
      "000011" when "0101000010000010", -- t[20610] = 3
      "000011" when "0101000010000011", -- t[20611] = 3
      "000011" when "0101000010000100", -- t[20612] = 3
      "000011" when "0101000010000101", -- t[20613] = 3
      "000011" when "0101000010000110", -- t[20614] = 3
      "000011" when "0101000010000111", -- t[20615] = 3
      "000011" when "0101000010001000", -- t[20616] = 3
      "000011" when "0101000010001001", -- t[20617] = 3
      "000011" when "0101000010001010", -- t[20618] = 3
      "000011" when "0101000010001011", -- t[20619] = 3
      "000011" when "0101000010001100", -- t[20620] = 3
      "000011" when "0101000010001101", -- t[20621] = 3
      "000011" when "0101000010001110", -- t[20622] = 3
      "000011" when "0101000010001111", -- t[20623] = 3
      "000011" when "0101000010010000", -- t[20624] = 3
      "000011" when "0101000010010001", -- t[20625] = 3
      "000011" when "0101000010010010", -- t[20626] = 3
      "000011" when "0101000010010011", -- t[20627] = 3
      "000011" when "0101000010010100", -- t[20628] = 3
      "000011" when "0101000010010101", -- t[20629] = 3
      "000011" when "0101000010010110", -- t[20630] = 3
      "000011" when "0101000010010111", -- t[20631] = 3
      "000011" when "0101000010011000", -- t[20632] = 3
      "000011" when "0101000010011001", -- t[20633] = 3
      "000011" when "0101000010011010", -- t[20634] = 3
      "000011" when "0101000010011011", -- t[20635] = 3
      "000011" when "0101000010011100", -- t[20636] = 3
      "000011" when "0101000010011101", -- t[20637] = 3
      "000011" when "0101000010011110", -- t[20638] = 3
      "000011" when "0101000010011111", -- t[20639] = 3
      "000011" when "0101000010100000", -- t[20640] = 3
      "000011" when "0101000010100001", -- t[20641] = 3
      "000011" when "0101000010100010", -- t[20642] = 3
      "000011" when "0101000010100011", -- t[20643] = 3
      "000011" when "0101000010100100", -- t[20644] = 3
      "000011" when "0101000010100101", -- t[20645] = 3
      "000011" when "0101000010100110", -- t[20646] = 3
      "000011" when "0101000010100111", -- t[20647] = 3
      "000011" when "0101000010101000", -- t[20648] = 3
      "000011" when "0101000010101001", -- t[20649] = 3
      "000011" when "0101000010101010", -- t[20650] = 3
      "000011" when "0101000010101011", -- t[20651] = 3
      "000011" when "0101000010101100", -- t[20652] = 3
      "000011" when "0101000010101101", -- t[20653] = 3
      "000011" when "0101000010101110", -- t[20654] = 3
      "000011" when "0101000010101111", -- t[20655] = 3
      "000011" when "0101000010110000", -- t[20656] = 3
      "000011" when "0101000010110001", -- t[20657] = 3
      "000011" when "0101000010110010", -- t[20658] = 3
      "000011" when "0101000010110011", -- t[20659] = 3
      "000011" when "0101000010110100", -- t[20660] = 3
      "000011" when "0101000010110101", -- t[20661] = 3
      "000011" when "0101000010110110", -- t[20662] = 3
      "000011" when "0101000010110111", -- t[20663] = 3
      "000011" when "0101000010111000", -- t[20664] = 3
      "000011" when "0101000010111001", -- t[20665] = 3
      "000011" when "0101000010111010", -- t[20666] = 3
      "000011" when "0101000010111011", -- t[20667] = 3
      "000011" when "0101000010111100", -- t[20668] = 3
      "000011" when "0101000010111101", -- t[20669] = 3
      "000011" when "0101000010111110", -- t[20670] = 3
      "000011" when "0101000010111111", -- t[20671] = 3
      "000011" when "0101000011000000", -- t[20672] = 3
      "000011" when "0101000011000001", -- t[20673] = 3
      "000011" when "0101000011000010", -- t[20674] = 3
      "000011" when "0101000011000011", -- t[20675] = 3
      "000011" when "0101000011000100", -- t[20676] = 3
      "000011" when "0101000011000101", -- t[20677] = 3
      "000011" when "0101000011000110", -- t[20678] = 3
      "000011" when "0101000011000111", -- t[20679] = 3
      "000011" when "0101000011001000", -- t[20680] = 3
      "000011" when "0101000011001001", -- t[20681] = 3
      "000011" when "0101000011001010", -- t[20682] = 3
      "000011" when "0101000011001011", -- t[20683] = 3
      "000011" when "0101000011001100", -- t[20684] = 3
      "000011" when "0101000011001101", -- t[20685] = 3
      "000011" when "0101000011001110", -- t[20686] = 3
      "000011" when "0101000011001111", -- t[20687] = 3
      "000011" when "0101000011010000", -- t[20688] = 3
      "000011" when "0101000011010001", -- t[20689] = 3
      "000011" when "0101000011010010", -- t[20690] = 3
      "000011" when "0101000011010011", -- t[20691] = 3
      "000011" when "0101000011010100", -- t[20692] = 3
      "000011" when "0101000011010101", -- t[20693] = 3
      "000011" when "0101000011010110", -- t[20694] = 3
      "000011" when "0101000011010111", -- t[20695] = 3
      "000011" when "0101000011011000", -- t[20696] = 3
      "000011" when "0101000011011001", -- t[20697] = 3
      "000011" when "0101000011011010", -- t[20698] = 3
      "000011" when "0101000011011011", -- t[20699] = 3
      "000011" when "0101000011011100", -- t[20700] = 3
      "000011" when "0101000011011101", -- t[20701] = 3
      "000011" when "0101000011011110", -- t[20702] = 3
      "000011" when "0101000011011111", -- t[20703] = 3
      "000011" when "0101000011100000", -- t[20704] = 3
      "000011" when "0101000011100001", -- t[20705] = 3
      "000011" when "0101000011100010", -- t[20706] = 3
      "000011" when "0101000011100011", -- t[20707] = 3
      "000011" when "0101000011100100", -- t[20708] = 3
      "000011" when "0101000011100101", -- t[20709] = 3
      "000011" when "0101000011100110", -- t[20710] = 3
      "000011" when "0101000011100111", -- t[20711] = 3
      "000011" when "0101000011101000", -- t[20712] = 3
      "000011" when "0101000011101001", -- t[20713] = 3
      "000011" when "0101000011101010", -- t[20714] = 3
      "000011" when "0101000011101011", -- t[20715] = 3
      "000011" when "0101000011101100", -- t[20716] = 3
      "000011" when "0101000011101101", -- t[20717] = 3
      "000011" when "0101000011101110", -- t[20718] = 3
      "000011" when "0101000011101111", -- t[20719] = 3
      "000011" when "0101000011110000", -- t[20720] = 3
      "000011" when "0101000011110001", -- t[20721] = 3
      "000011" when "0101000011110010", -- t[20722] = 3
      "000011" when "0101000011110011", -- t[20723] = 3
      "000011" when "0101000011110100", -- t[20724] = 3
      "000011" when "0101000011110101", -- t[20725] = 3
      "000011" when "0101000011110110", -- t[20726] = 3
      "000011" when "0101000011110111", -- t[20727] = 3
      "000011" when "0101000011111000", -- t[20728] = 3
      "000011" when "0101000011111001", -- t[20729] = 3
      "000011" when "0101000011111010", -- t[20730] = 3
      "000011" when "0101000011111011", -- t[20731] = 3
      "000011" when "0101000011111100", -- t[20732] = 3
      "000011" when "0101000011111101", -- t[20733] = 3
      "000011" when "0101000011111110", -- t[20734] = 3
      "000011" when "0101000011111111", -- t[20735] = 3
      "000011" when "0101000100000000", -- t[20736] = 3
      "000011" when "0101000100000001", -- t[20737] = 3
      "000011" when "0101000100000010", -- t[20738] = 3
      "000011" when "0101000100000011", -- t[20739] = 3
      "000011" when "0101000100000100", -- t[20740] = 3
      "000011" when "0101000100000101", -- t[20741] = 3
      "000011" when "0101000100000110", -- t[20742] = 3
      "000011" when "0101000100000111", -- t[20743] = 3
      "000011" when "0101000100001000", -- t[20744] = 3
      "000011" when "0101000100001001", -- t[20745] = 3
      "000011" when "0101000100001010", -- t[20746] = 3
      "000011" when "0101000100001011", -- t[20747] = 3
      "000011" when "0101000100001100", -- t[20748] = 3
      "000011" when "0101000100001101", -- t[20749] = 3
      "000011" when "0101000100001110", -- t[20750] = 3
      "000011" when "0101000100001111", -- t[20751] = 3
      "000011" when "0101000100010000", -- t[20752] = 3
      "000011" when "0101000100010001", -- t[20753] = 3
      "000011" when "0101000100010010", -- t[20754] = 3
      "000011" when "0101000100010011", -- t[20755] = 3
      "000011" when "0101000100010100", -- t[20756] = 3
      "000011" when "0101000100010101", -- t[20757] = 3
      "000011" when "0101000100010110", -- t[20758] = 3
      "000011" when "0101000100010111", -- t[20759] = 3
      "000011" when "0101000100011000", -- t[20760] = 3
      "000011" when "0101000100011001", -- t[20761] = 3
      "000011" when "0101000100011010", -- t[20762] = 3
      "000011" when "0101000100011011", -- t[20763] = 3
      "000011" when "0101000100011100", -- t[20764] = 3
      "000011" when "0101000100011101", -- t[20765] = 3
      "000011" when "0101000100011110", -- t[20766] = 3
      "000011" when "0101000100011111", -- t[20767] = 3
      "000011" when "0101000100100000", -- t[20768] = 3
      "000011" when "0101000100100001", -- t[20769] = 3
      "000011" when "0101000100100010", -- t[20770] = 3
      "000011" when "0101000100100011", -- t[20771] = 3
      "000011" when "0101000100100100", -- t[20772] = 3
      "000011" when "0101000100100101", -- t[20773] = 3
      "000011" when "0101000100100110", -- t[20774] = 3
      "000011" when "0101000100100111", -- t[20775] = 3
      "000011" when "0101000100101000", -- t[20776] = 3
      "000011" when "0101000100101001", -- t[20777] = 3
      "000011" when "0101000100101010", -- t[20778] = 3
      "000011" when "0101000100101011", -- t[20779] = 3
      "000011" when "0101000100101100", -- t[20780] = 3
      "000011" when "0101000100101101", -- t[20781] = 3
      "000011" when "0101000100101110", -- t[20782] = 3
      "000011" when "0101000100101111", -- t[20783] = 3
      "000011" when "0101000100110000", -- t[20784] = 3
      "000011" when "0101000100110001", -- t[20785] = 3
      "000011" when "0101000100110010", -- t[20786] = 3
      "000011" when "0101000100110011", -- t[20787] = 3
      "000011" when "0101000100110100", -- t[20788] = 3
      "000011" when "0101000100110101", -- t[20789] = 3
      "000011" when "0101000100110110", -- t[20790] = 3
      "000011" when "0101000100110111", -- t[20791] = 3
      "000011" when "0101000100111000", -- t[20792] = 3
      "000011" when "0101000100111001", -- t[20793] = 3
      "000011" when "0101000100111010", -- t[20794] = 3
      "000011" when "0101000100111011", -- t[20795] = 3
      "000011" when "0101000100111100", -- t[20796] = 3
      "000011" when "0101000100111101", -- t[20797] = 3
      "000011" when "0101000100111110", -- t[20798] = 3
      "000011" when "0101000100111111", -- t[20799] = 3
      "000011" when "0101000101000000", -- t[20800] = 3
      "000011" when "0101000101000001", -- t[20801] = 3
      "000011" when "0101000101000010", -- t[20802] = 3
      "000011" when "0101000101000011", -- t[20803] = 3
      "000011" when "0101000101000100", -- t[20804] = 3
      "000011" when "0101000101000101", -- t[20805] = 3
      "000011" when "0101000101000110", -- t[20806] = 3
      "000011" when "0101000101000111", -- t[20807] = 3
      "000011" when "0101000101001000", -- t[20808] = 3
      "000011" when "0101000101001001", -- t[20809] = 3
      "000011" when "0101000101001010", -- t[20810] = 3
      "000011" when "0101000101001011", -- t[20811] = 3
      "000011" when "0101000101001100", -- t[20812] = 3
      "000011" when "0101000101001101", -- t[20813] = 3
      "000011" when "0101000101001110", -- t[20814] = 3
      "000011" when "0101000101001111", -- t[20815] = 3
      "000011" when "0101000101010000", -- t[20816] = 3
      "000011" when "0101000101010001", -- t[20817] = 3
      "000011" when "0101000101010010", -- t[20818] = 3
      "000011" when "0101000101010011", -- t[20819] = 3
      "000011" when "0101000101010100", -- t[20820] = 3
      "000011" when "0101000101010101", -- t[20821] = 3
      "000011" when "0101000101010110", -- t[20822] = 3
      "000011" when "0101000101010111", -- t[20823] = 3
      "000011" when "0101000101011000", -- t[20824] = 3
      "000011" when "0101000101011001", -- t[20825] = 3
      "000011" when "0101000101011010", -- t[20826] = 3
      "000011" when "0101000101011011", -- t[20827] = 3
      "000011" when "0101000101011100", -- t[20828] = 3
      "000011" when "0101000101011101", -- t[20829] = 3
      "000011" when "0101000101011110", -- t[20830] = 3
      "000011" when "0101000101011111", -- t[20831] = 3
      "000011" when "0101000101100000", -- t[20832] = 3
      "000011" when "0101000101100001", -- t[20833] = 3
      "000011" when "0101000101100010", -- t[20834] = 3
      "000011" when "0101000101100011", -- t[20835] = 3
      "000011" when "0101000101100100", -- t[20836] = 3
      "000011" when "0101000101100101", -- t[20837] = 3
      "000011" when "0101000101100110", -- t[20838] = 3
      "000011" when "0101000101100111", -- t[20839] = 3
      "000011" when "0101000101101000", -- t[20840] = 3
      "000011" when "0101000101101001", -- t[20841] = 3
      "000011" when "0101000101101010", -- t[20842] = 3
      "000011" when "0101000101101011", -- t[20843] = 3
      "000011" when "0101000101101100", -- t[20844] = 3
      "000011" when "0101000101101101", -- t[20845] = 3
      "000011" when "0101000101101110", -- t[20846] = 3
      "000011" when "0101000101101111", -- t[20847] = 3
      "000011" when "0101000101110000", -- t[20848] = 3
      "000011" when "0101000101110001", -- t[20849] = 3
      "000011" when "0101000101110010", -- t[20850] = 3
      "000011" when "0101000101110011", -- t[20851] = 3
      "000011" when "0101000101110100", -- t[20852] = 3
      "000011" when "0101000101110101", -- t[20853] = 3
      "000011" when "0101000101110110", -- t[20854] = 3
      "000011" when "0101000101110111", -- t[20855] = 3
      "000011" when "0101000101111000", -- t[20856] = 3
      "000011" when "0101000101111001", -- t[20857] = 3
      "000011" when "0101000101111010", -- t[20858] = 3
      "000011" when "0101000101111011", -- t[20859] = 3
      "000011" when "0101000101111100", -- t[20860] = 3
      "000011" when "0101000101111101", -- t[20861] = 3
      "000011" when "0101000101111110", -- t[20862] = 3
      "000011" when "0101000101111111", -- t[20863] = 3
      "000011" when "0101000110000000", -- t[20864] = 3
      "000011" when "0101000110000001", -- t[20865] = 3
      "000011" when "0101000110000010", -- t[20866] = 3
      "000011" when "0101000110000011", -- t[20867] = 3
      "000011" when "0101000110000100", -- t[20868] = 3
      "000011" when "0101000110000101", -- t[20869] = 3
      "000011" when "0101000110000110", -- t[20870] = 3
      "000011" when "0101000110000111", -- t[20871] = 3
      "000011" when "0101000110001000", -- t[20872] = 3
      "000011" when "0101000110001001", -- t[20873] = 3
      "000011" when "0101000110001010", -- t[20874] = 3
      "000011" when "0101000110001011", -- t[20875] = 3
      "000011" when "0101000110001100", -- t[20876] = 3
      "000011" when "0101000110001101", -- t[20877] = 3
      "000011" when "0101000110001110", -- t[20878] = 3
      "000011" when "0101000110001111", -- t[20879] = 3
      "000011" when "0101000110010000", -- t[20880] = 3
      "000011" when "0101000110010001", -- t[20881] = 3
      "000011" when "0101000110010010", -- t[20882] = 3
      "000011" when "0101000110010011", -- t[20883] = 3
      "000011" when "0101000110010100", -- t[20884] = 3
      "000011" when "0101000110010101", -- t[20885] = 3
      "000011" when "0101000110010110", -- t[20886] = 3
      "000011" when "0101000110010111", -- t[20887] = 3
      "000011" when "0101000110011000", -- t[20888] = 3
      "000011" when "0101000110011001", -- t[20889] = 3
      "000011" when "0101000110011010", -- t[20890] = 3
      "000011" when "0101000110011011", -- t[20891] = 3
      "000011" when "0101000110011100", -- t[20892] = 3
      "000011" when "0101000110011101", -- t[20893] = 3
      "000011" when "0101000110011110", -- t[20894] = 3
      "000011" when "0101000110011111", -- t[20895] = 3
      "000011" when "0101000110100000", -- t[20896] = 3
      "000011" when "0101000110100001", -- t[20897] = 3
      "000011" when "0101000110100010", -- t[20898] = 3
      "000011" when "0101000110100011", -- t[20899] = 3
      "000011" when "0101000110100100", -- t[20900] = 3
      "000011" when "0101000110100101", -- t[20901] = 3
      "000011" when "0101000110100110", -- t[20902] = 3
      "000011" when "0101000110100111", -- t[20903] = 3
      "000011" when "0101000110101000", -- t[20904] = 3
      "000011" when "0101000110101001", -- t[20905] = 3
      "000011" when "0101000110101010", -- t[20906] = 3
      "000011" when "0101000110101011", -- t[20907] = 3
      "000011" when "0101000110101100", -- t[20908] = 3
      "000011" when "0101000110101101", -- t[20909] = 3
      "000011" when "0101000110101110", -- t[20910] = 3
      "000011" when "0101000110101111", -- t[20911] = 3
      "000011" when "0101000110110000", -- t[20912] = 3
      "000011" when "0101000110110001", -- t[20913] = 3
      "000011" when "0101000110110010", -- t[20914] = 3
      "000011" when "0101000110110011", -- t[20915] = 3
      "000011" when "0101000110110100", -- t[20916] = 3
      "000011" when "0101000110110101", -- t[20917] = 3
      "000011" when "0101000110110110", -- t[20918] = 3
      "000011" when "0101000110110111", -- t[20919] = 3
      "000011" when "0101000110111000", -- t[20920] = 3
      "000011" when "0101000110111001", -- t[20921] = 3
      "000011" when "0101000110111010", -- t[20922] = 3
      "000011" when "0101000110111011", -- t[20923] = 3
      "000011" when "0101000110111100", -- t[20924] = 3
      "000011" when "0101000110111101", -- t[20925] = 3
      "000011" when "0101000110111110", -- t[20926] = 3
      "000011" when "0101000110111111", -- t[20927] = 3
      "000011" when "0101000111000000", -- t[20928] = 3
      "000011" when "0101000111000001", -- t[20929] = 3
      "000011" when "0101000111000010", -- t[20930] = 3
      "000011" when "0101000111000011", -- t[20931] = 3
      "000011" when "0101000111000100", -- t[20932] = 3
      "000011" when "0101000111000101", -- t[20933] = 3
      "000011" when "0101000111000110", -- t[20934] = 3
      "000011" when "0101000111000111", -- t[20935] = 3
      "000011" when "0101000111001000", -- t[20936] = 3
      "000011" when "0101000111001001", -- t[20937] = 3
      "000011" when "0101000111001010", -- t[20938] = 3
      "000011" when "0101000111001011", -- t[20939] = 3
      "000011" when "0101000111001100", -- t[20940] = 3
      "000011" when "0101000111001101", -- t[20941] = 3
      "000011" when "0101000111001110", -- t[20942] = 3
      "000011" when "0101000111001111", -- t[20943] = 3
      "000011" when "0101000111010000", -- t[20944] = 3
      "000011" when "0101000111010001", -- t[20945] = 3
      "000011" when "0101000111010010", -- t[20946] = 3
      "000011" when "0101000111010011", -- t[20947] = 3
      "000011" when "0101000111010100", -- t[20948] = 3
      "000011" when "0101000111010101", -- t[20949] = 3
      "000011" when "0101000111010110", -- t[20950] = 3
      "000011" when "0101000111010111", -- t[20951] = 3
      "000011" when "0101000111011000", -- t[20952] = 3
      "000011" when "0101000111011001", -- t[20953] = 3
      "000011" when "0101000111011010", -- t[20954] = 3
      "000011" when "0101000111011011", -- t[20955] = 3
      "000011" when "0101000111011100", -- t[20956] = 3
      "000011" when "0101000111011101", -- t[20957] = 3
      "000011" when "0101000111011110", -- t[20958] = 3
      "000011" when "0101000111011111", -- t[20959] = 3
      "000011" when "0101000111100000", -- t[20960] = 3
      "000011" when "0101000111100001", -- t[20961] = 3
      "000011" when "0101000111100010", -- t[20962] = 3
      "000011" when "0101000111100011", -- t[20963] = 3
      "000011" when "0101000111100100", -- t[20964] = 3
      "000011" when "0101000111100101", -- t[20965] = 3
      "000011" when "0101000111100110", -- t[20966] = 3
      "000011" when "0101000111100111", -- t[20967] = 3
      "000011" when "0101000111101000", -- t[20968] = 3
      "000011" when "0101000111101001", -- t[20969] = 3
      "000011" when "0101000111101010", -- t[20970] = 3
      "000011" when "0101000111101011", -- t[20971] = 3
      "000011" when "0101000111101100", -- t[20972] = 3
      "000011" when "0101000111101101", -- t[20973] = 3
      "000011" when "0101000111101110", -- t[20974] = 3
      "000011" when "0101000111101111", -- t[20975] = 3
      "000011" when "0101000111110000", -- t[20976] = 3
      "000011" when "0101000111110001", -- t[20977] = 3
      "000011" when "0101000111110010", -- t[20978] = 3
      "000011" when "0101000111110011", -- t[20979] = 3
      "000011" when "0101000111110100", -- t[20980] = 3
      "000011" when "0101000111110101", -- t[20981] = 3
      "000011" when "0101000111110110", -- t[20982] = 3
      "000011" when "0101000111110111", -- t[20983] = 3
      "000011" when "0101000111111000", -- t[20984] = 3
      "000011" when "0101000111111001", -- t[20985] = 3
      "000011" when "0101000111111010", -- t[20986] = 3
      "000011" when "0101000111111011", -- t[20987] = 3
      "000011" when "0101000111111100", -- t[20988] = 3
      "000011" when "0101000111111101", -- t[20989] = 3
      "000011" when "0101000111111110", -- t[20990] = 3
      "000011" when "0101000111111111", -- t[20991] = 3
      "000011" when "0101001000000000", -- t[20992] = 3
      "000011" when "0101001000000001", -- t[20993] = 3
      "000011" when "0101001000000010", -- t[20994] = 3
      "000011" when "0101001000000011", -- t[20995] = 3
      "000011" when "0101001000000100", -- t[20996] = 3
      "000011" when "0101001000000101", -- t[20997] = 3
      "000011" when "0101001000000110", -- t[20998] = 3
      "000011" when "0101001000000111", -- t[20999] = 3
      "000011" when "0101001000001000", -- t[21000] = 3
      "000011" when "0101001000001001", -- t[21001] = 3
      "000011" when "0101001000001010", -- t[21002] = 3
      "000011" when "0101001000001011", -- t[21003] = 3
      "000011" when "0101001000001100", -- t[21004] = 3
      "000011" when "0101001000001101", -- t[21005] = 3
      "000011" when "0101001000001110", -- t[21006] = 3
      "000011" when "0101001000001111", -- t[21007] = 3
      "000011" when "0101001000010000", -- t[21008] = 3
      "000011" when "0101001000010001", -- t[21009] = 3
      "000011" when "0101001000010010", -- t[21010] = 3
      "000011" when "0101001000010011", -- t[21011] = 3
      "000011" when "0101001000010100", -- t[21012] = 3
      "000011" when "0101001000010101", -- t[21013] = 3
      "000011" when "0101001000010110", -- t[21014] = 3
      "000011" when "0101001000010111", -- t[21015] = 3
      "000011" when "0101001000011000", -- t[21016] = 3
      "000011" when "0101001000011001", -- t[21017] = 3
      "000011" when "0101001000011010", -- t[21018] = 3
      "000011" when "0101001000011011", -- t[21019] = 3
      "000011" when "0101001000011100", -- t[21020] = 3
      "000011" when "0101001000011101", -- t[21021] = 3
      "000011" when "0101001000011110", -- t[21022] = 3
      "000011" when "0101001000011111", -- t[21023] = 3
      "000011" when "0101001000100000", -- t[21024] = 3
      "000011" when "0101001000100001", -- t[21025] = 3
      "000011" when "0101001000100010", -- t[21026] = 3
      "000011" when "0101001000100011", -- t[21027] = 3
      "000011" when "0101001000100100", -- t[21028] = 3
      "000011" when "0101001000100101", -- t[21029] = 3
      "000011" when "0101001000100110", -- t[21030] = 3
      "000011" when "0101001000100111", -- t[21031] = 3
      "000011" when "0101001000101000", -- t[21032] = 3
      "000011" when "0101001000101001", -- t[21033] = 3
      "000011" when "0101001000101010", -- t[21034] = 3
      "000011" when "0101001000101011", -- t[21035] = 3
      "000011" when "0101001000101100", -- t[21036] = 3
      "000011" when "0101001000101101", -- t[21037] = 3
      "000011" when "0101001000101110", -- t[21038] = 3
      "000011" when "0101001000101111", -- t[21039] = 3
      "000011" when "0101001000110000", -- t[21040] = 3
      "000011" when "0101001000110001", -- t[21041] = 3
      "000011" when "0101001000110010", -- t[21042] = 3
      "000011" when "0101001000110011", -- t[21043] = 3
      "000011" when "0101001000110100", -- t[21044] = 3
      "000011" when "0101001000110101", -- t[21045] = 3
      "000011" when "0101001000110110", -- t[21046] = 3
      "000011" when "0101001000110111", -- t[21047] = 3
      "000011" when "0101001000111000", -- t[21048] = 3
      "000011" when "0101001000111001", -- t[21049] = 3
      "000011" when "0101001000111010", -- t[21050] = 3
      "000011" when "0101001000111011", -- t[21051] = 3
      "000011" when "0101001000111100", -- t[21052] = 3
      "000011" when "0101001000111101", -- t[21053] = 3
      "000011" when "0101001000111110", -- t[21054] = 3
      "000011" when "0101001000111111", -- t[21055] = 3
      "000011" when "0101001001000000", -- t[21056] = 3
      "000011" when "0101001001000001", -- t[21057] = 3
      "000011" when "0101001001000010", -- t[21058] = 3
      "000011" when "0101001001000011", -- t[21059] = 3
      "000011" when "0101001001000100", -- t[21060] = 3
      "000011" when "0101001001000101", -- t[21061] = 3
      "000011" when "0101001001000110", -- t[21062] = 3
      "000011" when "0101001001000111", -- t[21063] = 3
      "000011" when "0101001001001000", -- t[21064] = 3
      "000011" when "0101001001001001", -- t[21065] = 3
      "000011" when "0101001001001010", -- t[21066] = 3
      "000011" when "0101001001001011", -- t[21067] = 3
      "000011" when "0101001001001100", -- t[21068] = 3
      "000011" when "0101001001001101", -- t[21069] = 3
      "000011" when "0101001001001110", -- t[21070] = 3
      "000011" when "0101001001001111", -- t[21071] = 3
      "000011" when "0101001001010000", -- t[21072] = 3
      "000011" when "0101001001010001", -- t[21073] = 3
      "000011" when "0101001001010010", -- t[21074] = 3
      "000011" when "0101001001010011", -- t[21075] = 3
      "000011" when "0101001001010100", -- t[21076] = 3
      "000011" when "0101001001010101", -- t[21077] = 3
      "000011" when "0101001001010110", -- t[21078] = 3
      "000011" when "0101001001010111", -- t[21079] = 3
      "000011" when "0101001001011000", -- t[21080] = 3
      "000011" when "0101001001011001", -- t[21081] = 3
      "000011" when "0101001001011010", -- t[21082] = 3
      "000011" when "0101001001011011", -- t[21083] = 3
      "000011" when "0101001001011100", -- t[21084] = 3
      "000011" when "0101001001011101", -- t[21085] = 3
      "000011" when "0101001001011110", -- t[21086] = 3
      "000011" when "0101001001011111", -- t[21087] = 3
      "000011" when "0101001001100000", -- t[21088] = 3
      "000011" when "0101001001100001", -- t[21089] = 3
      "000011" when "0101001001100010", -- t[21090] = 3
      "000011" when "0101001001100011", -- t[21091] = 3
      "000011" when "0101001001100100", -- t[21092] = 3
      "000011" when "0101001001100101", -- t[21093] = 3
      "000011" when "0101001001100110", -- t[21094] = 3
      "000011" when "0101001001100111", -- t[21095] = 3
      "000011" when "0101001001101000", -- t[21096] = 3
      "000011" when "0101001001101001", -- t[21097] = 3
      "000011" when "0101001001101010", -- t[21098] = 3
      "000011" when "0101001001101011", -- t[21099] = 3
      "000011" when "0101001001101100", -- t[21100] = 3
      "000011" when "0101001001101101", -- t[21101] = 3
      "000011" when "0101001001101110", -- t[21102] = 3
      "000011" when "0101001001101111", -- t[21103] = 3
      "000011" when "0101001001110000", -- t[21104] = 3
      "000011" when "0101001001110001", -- t[21105] = 3
      "000011" when "0101001001110010", -- t[21106] = 3
      "000011" when "0101001001110011", -- t[21107] = 3
      "000011" when "0101001001110100", -- t[21108] = 3
      "000011" when "0101001001110101", -- t[21109] = 3
      "000011" when "0101001001110110", -- t[21110] = 3
      "000011" when "0101001001110111", -- t[21111] = 3
      "000011" when "0101001001111000", -- t[21112] = 3
      "000011" when "0101001001111001", -- t[21113] = 3
      "000011" when "0101001001111010", -- t[21114] = 3
      "000011" when "0101001001111011", -- t[21115] = 3
      "000011" when "0101001001111100", -- t[21116] = 3
      "000011" when "0101001001111101", -- t[21117] = 3
      "000011" when "0101001001111110", -- t[21118] = 3
      "000011" when "0101001001111111", -- t[21119] = 3
      "000011" when "0101001010000000", -- t[21120] = 3
      "000011" when "0101001010000001", -- t[21121] = 3
      "000011" when "0101001010000010", -- t[21122] = 3
      "000011" when "0101001010000011", -- t[21123] = 3
      "000011" when "0101001010000100", -- t[21124] = 3
      "000011" when "0101001010000101", -- t[21125] = 3
      "000011" when "0101001010000110", -- t[21126] = 3
      "000011" when "0101001010000111", -- t[21127] = 3
      "000011" when "0101001010001000", -- t[21128] = 3
      "000011" when "0101001010001001", -- t[21129] = 3
      "000011" when "0101001010001010", -- t[21130] = 3
      "000011" when "0101001010001011", -- t[21131] = 3
      "000011" when "0101001010001100", -- t[21132] = 3
      "000011" when "0101001010001101", -- t[21133] = 3
      "000011" when "0101001010001110", -- t[21134] = 3
      "000011" when "0101001010001111", -- t[21135] = 3
      "000011" when "0101001010010000", -- t[21136] = 3
      "000011" when "0101001010010001", -- t[21137] = 3
      "000011" when "0101001010010010", -- t[21138] = 3
      "000011" when "0101001010010011", -- t[21139] = 3
      "000011" when "0101001010010100", -- t[21140] = 3
      "000011" when "0101001010010101", -- t[21141] = 3
      "000011" when "0101001010010110", -- t[21142] = 3
      "000011" when "0101001010010111", -- t[21143] = 3
      "000011" when "0101001010011000", -- t[21144] = 3
      "000011" when "0101001010011001", -- t[21145] = 3
      "000011" when "0101001010011010", -- t[21146] = 3
      "000011" when "0101001010011011", -- t[21147] = 3
      "000011" when "0101001010011100", -- t[21148] = 3
      "000011" when "0101001010011101", -- t[21149] = 3
      "000011" when "0101001010011110", -- t[21150] = 3
      "000011" when "0101001010011111", -- t[21151] = 3
      "000011" when "0101001010100000", -- t[21152] = 3
      "000011" when "0101001010100001", -- t[21153] = 3
      "000011" when "0101001010100010", -- t[21154] = 3
      "000011" when "0101001010100011", -- t[21155] = 3
      "000011" when "0101001010100100", -- t[21156] = 3
      "000011" when "0101001010100101", -- t[21157] = 3
      "000011" when "0101001010100110", -- t[21158] = 3
      "000011" when "0101001010100111", -- t[21159] = 3
      "000011" when "0101001010101000", -- t[21160] = 3
      "000011" when "0101001010101001", -- t[21161] = 3
      "000011" when "0101001010101010", -- t[21162] = 3
      "000011" when "0101001010101011", -- t[21163] = 3
      "000011" when "0101001010101100", -- t[21164] = 3
      "000011" when "0101001010101101", -- t[21165] = 3
      "000011" when "0101001010101110", -- t[21166] = 3
      "000011" when "0101001010101111", -- t[21167] = 3
      "000011" when "0101001010110000", -- t[21168] = 3
      "000011" when "0101001010110001", -- t[21169] = 3
      "000011" when "0101001010110010", -- t[21170] = 3
      "000011" when "0101001010110011", -- t[21171] = 3
      "000011" when "0101001010110100", -- t[21172] = 3
      "000011" when "0101001010110101", -- t[21173] = 3
      "000011" when "0101001010110110", -- t[21174] = 3
      "000011" when "0101001010110111", -- t[21175] = 3
      "000011" when "0101001010111000", -- t[21176] = 3
      "000011" when "0101001010111001", -- t[21177] = 3
      "000011" when "0101001010111010", -- t[21178] = 3
      "000011" when "0101001010111011", -- t[21179] = 3
      "000011" when "0101001010111100", -- t[21180] = 3
      "000011" when "0101001010111101", -- t[21181] = 3
      "000011" when "0101001010111110", -- t[21182] = 3
      "000011" when "0101001010111111", -- t[21183] = 3
      "000011" when "0101001011000000", -- t[21184] = 3
      "000011" when "0101001011000001", -- t[21185] = 3
      "000011" when "0101001011000010", -- t[21186] = 3
      "000011" when "0101001011000011", -- t[21187] = 3
      "000011" when "0101001011000100", -- t[21188] = 3
      "000011" when "0101001011000101", -- t[21189] = 3
      "000011" when "0101001011000110", -- t[21190] = 3
      "000011" when "0101001011000111", -- t[21191] = 3
      "000011" when "0101001011001000", -- t[21192] = 3
      "000011" when "0101001011001001", -- t[21193] = 3
      "000011" when "0101001011001010", -- t[21194] = 3
      "000011" when "0101001011001011", -- t[21195] = 3
      "000011" when "0101001011001100", -- t[21196] = 3
      "000011" when "0101001011001101", -- t[21197] = 3
      "000011" when "0101001011001110", -- t[21198] = 3
      "000011" when "0101001011001111", -- t[21199] = 3
      "000011" when "0101001011010000", -- t[21200] = 3
      "000011" when "0101001011010001", -- t[21201] = 3
      "000011" when "0101001011010010", -- t[21202] = 3
      "000011" when "0101001011010011", -- t[21203] = 3
      "000011" when "0101001011010100", -- t[21204] = 3
      "000011" when "0101001011010101", -- t[21205] = 3
      "000011" when "0101001011010110", -- t[21206] = 3
      "000011" when "0101001011010111", -- t[21207] = 3
      "000011" when "0101001011011000", -- t[21208] = 3
      "000011" when "0101001011011001", -- t[21209] = 3
      "000011" when "0101001011011010", -- t[21210] = 3
      "000011" when "0101001011011011", -- t[21211] = 3
      "000011" when "0101001011011100", -- t[21212] = 3
      "000011" when "0101001011011101", -- t[21213] = 3
      "000011" when "0101001011011110", -- t[21214] = 3
      "000011" when "0101001011011111", -- t[21215] = 3
      "000011" when "0101001011100000", -- t[21216] = 3
      "000011" when "0101001011100001", -- t[21217] = 3
      "000011" when "0101001011100010", -- t[21218] = 3
      "000011" when "0101001011100011", -- t[21219] = 3
      "000011" when "0101001011100100", -- t[21220] = 3
      "000011" when "0101001011100101", -- t[21221] = 3
      "000011" when "0101001011100110", -- t[21222] = 3
      "000011" when "0101001011100111", -- t[21223] = 3
      "000011" when "0101001011101000", -- t[21224] = 3
      "000011" when "0101001011101001", -- t[21225] = 3
      "000011" when "0101001011101010", -- t[21226] = 3
      "000011" when "0101001011101011", -- t[21227] = 3
      "000011" when "0101001011101100", -- t[21228] = 3
      "000011" when "0101001011101101", -- t[21229] = 3
      "000011" when "0101001011101110", -- t[21230] = 3
      "000011" when "0101001011101111", -- t[21231] = 3
      "000011" when "0101001011110000", -- t[21232] = 3
      "000011" when "0101001011110001", -- t[21233] = 3
      "000011" when "0101001011110010", -- t[21234] = 3
      "000011" when "0101001011110011", -- t[21235] = 3
      "000011" when "0101001011110100", -- t[21236] = 3
      "000011" when "0101001011110101", -- t[21237] = 3
      "000011" when "0101001011110110", -- t[21238] = 3
      "000011" when "0101001011110111", -- t[21239] = 3
      "000011" when "0101001011111000", -- t[21240] = 3
      "000011" when "0101001011111001", -- t[21241] = 3
      "000011" when "0101001011111010", -- t[21242] = 3
      "000011" when "0101001011111011", -- t[21243] = 3
      "000011" when "0101001011111100", -- t[21244] = 3
      "000011" when "0101001011111101", -- t[21245] = 3
      "000011" when "0101001011111110", -- t[21246] = 3
      "000011" when "0101001011111111", -- t[21247] = 3
      "000011" when "0101001100000000", -- t[21248] = 3
      "000011" when "0101001100000001", -- t[21249] = 3
      "000011" when "0101001100000010", -- t[21250] = 3
      "000011" when "0101001100000011", -- t[21251] = 3
      "000011" when "0101001100000100", -- t[21252] = 3
      "000011" when "0101001100000101", -- t[21253] = 3
      "000011" when "0101001100000110", -- t[21254] = 3
      "000011" when "0101001100000111", -- t[21255] = 3
      "000011" when "0101001100001000", -- t[21256] = 3
      "000011" when "0101001100001001", -- t[21257] = 3
      "000011" when "0101001100001010", -- t[21258] = 3
      "000011" when "0101001100001011", -- t[21259] = 3
      "000011" when "0101001100001100", -- t[21260] = 3
      "000011" when "0101001100001101", -- t[21261] = 3
      "000011" when "0101001100001110", -- t[21262] = 3
      "000011" when "0101001100001111", -- t[21263] = 3
      "000011" when "0101001100010000", -- t[21264] = 3
      "000011" when "0101001100010001", -- t[21265] = 3
      "000011" when "0101001100010010", -- t[21266] = 3
      "000011" when "0101001100010011", -- t[21267] = 3
      "000011" when "0101001100010100", -- t[21268] = 3
      "000011" when "0101001100010101", -- t[21269] = 3
      "000011" when "0101001100010110", -- t[21270] = 3
      "000011" when "0101001100010111", -- t[21271] = 3
      "000011" when "0101001100011000", -- t[21272] = 3
      "000011" when "0101001100011001", -- t[21273] = 3
      "000011" when "0101001100011010", -- t[21274] = 3
      "000011" when "0101001100011011", -- t[21275] = 3
      "000011" when "0101001100011100", -- t[21276] = 3
      "000011" when "0101001100011101", -- t[21277] = 3
      "000011" when "0101001100011110", -- t[21278] = 3
      "000011" when "0101001100011111", -- t[21279] = 3
      "000011" when "0101001100100000", -- t[21280] = 3
      "000011" when "0101001100100001", -- t[21281] = 3
      "000011" when "0101001100100010", -- t[21282] = 3
      "000011" when "0101001100100011", -- t[21283] = 3
      "000011" when "0101001100100100", -- t[21284] = 3
      "000011" when "0101001100100101", -- t[21285] = 3
      "000011" when "0101001100100110", -- t[21286] = 3
      "000011" when "0101001100100111", -- t[21287] = 3
      "000011" when "0101001100101000", -- t[21288] = 3
      "000011" when "0101001100101001", -- t[21289] = 3
      "000011" when "0101001100101010", -- t[21290] = 3
      "000011" when "0101001100101011", -- t[21291] = 3
      "000011" when "0101001100101100", -- t[21292] = 3
      "000011" when "0101001100101101", -- t[21293] = 3
      "000011" when "0101001100101110", -- t[21294] = 3
      "000011" when "0101001100101111", -- t[21295] = 3
      "000011" when "0101001100110000", -- t[21296] = 3
      "000011" when "0101001100110001", -- t[21297] = 3
      "000011" when "0101001100110010", -- t[21298] = 3
      "000011" when "0101001100110011", -- t[21299] = 3
      "000011" when "0101001100110100", -- t[21300] = 3
      "000011" when "0101001100110101", -- t[21301] = 3
      "000011" when "0101001100110110", -- t[21302] = 3
      "000011" when "0101001100110111", -- t[21303] = 3
      "000011" when "0101001100111000", -- t[21304] = 3
      "000011" when "0101001100111001", -- t[21305] = 3
      "000011" when "0101001100111010", -- t[21306] = 3
      "000011" when "0101001100111011", -- t[21307] = 3
      "000011" when "0101001100111100", -- t[21308] = 3
      "000011" when "0101001100111101", -- t[21309] = 3
      "000011" when "0101001100111110", -- t[21310] = 3
      "000011" when "0101001100111111", -- t[21311] = 3
      "000011" when "0101001101000000", -- t[21312] = 3
      "000011" when "0101001101000001", -- t[21313] = 3
      "000011" when "0101001101000010", -- t[21314] = 3
      "000011" when "0101001101000011", -- t[21315] = 3
      "000011" when "0101001101000100", -- t[21316] = 3
      "000011" when "0101001101000101", -- t[21317] = 3
      "000011" when "0101001101000110", -- t[21318] = 3
      "000011" when "0101001101000111", -- t[21319] = 3
      "000011" when "0101001101001000", -- t[21320] = 3
      "000011" when "0101001101001001", -- t[21321] = 3
      "000011" when "0101001101001010", -- t[21322] = 3
      "000011" when "0101001101001011", -- t[21323] = 3
      "000011" when "0101001101001100", -- t[21324] = 3
      "000011" when "0101001101001101", -- t[21325] = 3
      "000011" when "0101001101001110", -- t[21326] = 3
      "000011" when "0101001101001111", -- t[21327] = 3
      "000011" when "0101001101010000", -- t[21328] = 3
      "000011" when "0101001101010001", -- t[21329] = 3
      "000011" when "0101001101010010", -- t[21330] = 3
      "000011" when "0101001101010011", -- t[21331] = 3
      "000011" when "0101001101010100", -- t[21332] = 3
      "000011" when "0101001101010101", -- t[21333] = 3
      "000011" when "0101001101010110", -- t[21334] = 3
      "000011" when "0101001101010111", -- t[21335] = 3
      "000011" when "0101001101011000", -- t[21336] = 3
      "000011" when "0101001101011001", -- t[21337] = 3
      "000011" when "0101001101011010", -- t[21338] = 3
      "000011" when "0101001101011011", -- t[21339] = 3
      "000011" when "0101001101011100", -- t[21340] = 3
      "000011" when "0101001101011101", -- t[21341] = 3
      "000011" when "0101001101011110", -- t[21342] = 3
      "000011" when "0101001101011111", -- t[21343] = 3
      "000011" when "0101001101100000", -- t[21344] = 3
      "000011" when "0101001101100001", -- t[21345] = 3
      "000011" when "0101001101100010", -- t[21346] = 3
      "000011" when "0101001101100011", -- t[21347] = 3
      "000011" when "0101001101100100", -- t[21348] = 3
      "000011" when "0101001101100101", -- t[21349] = 3
      "000011" when "0101001101100110", -- t[21350] = 3
      "000011" when "0101001101100111", -- t[21351] = 3
      "000011" when "0101001101101000", -- t[21352] = 3
      "000011" when "0101001101101001", -- t[21353] = 3
      "000011" when "0101001101101010", -- t[21354] = 3
      "000011" when "0101001101101011", -- t[21355] = 3
      "000011" when "0101001101101100", -- t[21356] = 3
      "000011" when "0101001101101101", -- t[21357] = 3
      "000011" when "0101001101101110", -- t[21358] = 3
      "000011" when "0101001101101111", -- t[21359] = 3
      "000011" when "0101001101110000", -- t[21360] = 3
      "000011" when "0101001101110001", -- t[21361] = 3
      "000011" when "0101001101110010", -- t[21362] = 3
      "000011" when "0101001101110011", -- t[21363] = 3
      "000011" when "0101001101110100", -- t[21364] = 3
      "000011" when "0101001101110101", -- t[21365] = 3
      "000011" when "0101001101110110", -- t[21366] = 3
      "000011" when "0101001101110111", -- t[21367] = 3
      "000011" when "0101001101111000", -- t[21368] = 3
      "000011" when "0101001101111001", -- t[21369] = 3
      "000011" when "0101001101111010", -- t[21370] = 3
      "000011" when "0101001101111011", -- t[21371] = 3
      "000011" when "0101001101111100", -- t[21372] = 3
      "000011" when "0101001101111101", -- t[21373] = 3
      "000011" when "0101001101111110", -- t[21374] = 3
      "000011" when "0101001101111111", -- t[21375] = 3
      "000011" when "0101001110000000", -- t[21376] = 3
      "000011" when "0101001110000001", -- t[21377] = 3
      "000011" when "0101001110000010", -- t[21378] = 3
      "000011" when "0101001110000011", -- t[21379] = 3
      "000011" when "0101001110000100", -- t[21380] = 3
      "000011" when "0101001110000101", -- t[21381] = 3
      "000011" when "0101001110000110", -- t[21382] = 3
      "000011" when "0101001110000111", -- t[21383] = 3
      "000011" when "0101001110001000", -- t[21384] = 3
      "000011" when "0101001110001001", -- t[21385] = 3
      "000011" when "0101001110001010", -- t[21386] = 3
      "000011" when "0101001110001011", -- t[21387] = 3
      "000011" when "0101001110001100", -- t[21388] = 3
      "000011" when "0101001110001101", -- t[21389] = 3
      "000011" when "0101001110001110", -- t[21390] = 3
      "000011" when "0101001110001111", -- t[21391] = 3
      "000011" when "0101001110010000", -- t[21392] = 3
      "000011" when "0101001110010001", -- t[21393] = 3
      "000011" when "0101001110010010", -- t[21394] = 3
      "000011" when "0101001110010011", -- t[21395] = 3
      "000011" when "0101001110010100", -- t[21396] = 3
      "000011" when "0101001110010101", -- t[21397] = 3
      "000011" when "0101001110010110", -- t[21398] = 3
      "000011" when "0101001110010111", -- t[21399] = 3
      "000011" when "0101001110011000", -- t[21400] = 3
      "000011" when "0101001110011001", -- t[21401] = 3
      "000011" when "0101001110011010", -- t[21402] = 3
      "000011" when "0101001110011011", -- t[21403] = 3
      "000011" when "0101001110011100", -- t[21404] = 3
      "000011" when "0101001110011101", -- t[21405] = 3
      "000011" when "0101001110011110", -- t[21406] = 3
      "000011" when "0101001110011111", -- t[21407] = 3
      "000011" when "0101001110100000", -- t[21408] = 3
      "000011" when "0101001110100001", -- t[21409] = 3
      "000011" when "0101001110100010", -- t[21410] = 3
      "000011" when "0101001110100011", -- t[21411] = 3
      "000011" when "0101001110100100", -- t[21412] = 3
      "000011" when "0101001110100101", -- t[21413] = 3
      "000011" when "0101001110100110", -- t[21414] = 3
      "000011" when "0101001110100111", -- t[21415] = 3
      "000011" when "0101001110101000", -- t[21416] = 3
      "000011" when "0101001110101001", -- t[21417] = 3
      "000011" when "0101001110101010", -- t[21418] = 3
      "000011" when "0101001110101011", -- t[21419] = 3
      "000011" when "0101001110101100", -- t[21420] = 3
      "000011" when "0101001110101101", -- t[21421] = 3
      "000011" when "0101001110101110", -- t[21422] = 3
      "000011" when "0101001110101111", -- t[21423] = 3
      "000011" when "0101001110110000", -- t[21424] = 3
      "000011" when "0101001110110001", -- t[21425] = 3
      "000011" when "0101001110110010", -- t[21426] = 3
      "000011" when "0101001110110011", -- t[21427] = 3
      "000011" when "0101001110110100", -- t[21428] = 3
      "000011" when "0101001110110101", -- t[21429] = 3
      "000011" when "0101001110110110", -- t[21430] = 3
      "000011" when "0101001110110111", -- t[21431] = 3
      "000011" when "0101001110111000", -- t[21432] = 3
      "000011" when "0101001110111001", -- t[21433] = 3
      "000011" when "0101001110111010", -- t[21434] = 3
      "000011" when "0101001110111011", -- t[21435] = 3
      "000011" when "0101001110111100", -- t[21436] = 3
      "000011" when "0101001110111101", -- t[21437] = 3
      "000011" when "0101001110111110", -- t[21438] = 3
      "000011" when "0101001110111111", -- t[21439] = 3
      "000011" when "0101001111000000", -- t[21440] = 3
      "000011" when "0101001111000001", -- t[21441] = 3
      "000011" when "0101001111000010", -- t[21442] = 3
      "000011" when "0101001111000011", -- t[21443] = 3
      "000011" when "0101001111000100", -- t[21444] = 3
      "000011" when "0101001111000101", -- t[21445] = 3
      "000011" when "0101001111000110", -- t[21446] = 3
      "000011" when "0101001111000111", -- t[21447] = 3
      "000011" when "0101001111001000", -- t[21448] = 3
      "000011" when "0101001111001001", -- t[21449] = 3
      "000011" when "0101001111001010", -- t[21450] = 3
      "000011" when "0101001111001011", -- t[21451] = 3
      "000011" when "0101001111001100", -- t[21452] = 3
      "000011" when "0101001111001101", -- t[21453] = 3
      "000011" when "0101001111001110", -- t[21454] = 3
      "000011" when "0101001111001111", -- t[21455] = 3
      "000011" when "0101001111010000", -- t[21456] = 3
      "000011" when "0101001111010001", -- t[21457] = 3
      "000011" when "0101001111010010", -- t[21458] = 3
      "000011" when "0101001111010011", -- t[21459] = 3
      "000011" when "0101001111010100", -- t[21460] = 3
      "000011" when "0101001111010101", -- t[21461] = 3
      "000011" when "0101001111010110", -- t[21462] = 3
      "000011" when "0101001111010111", -- t[21463] = 3
      "000011" when "0101001111011000", -- t[21464] = 3
      "000011" when "0101001111011001", -- t[21465] = 3
      "000011" when "0101001111011010", -- t[21466] = 3
      "000011" when "0101001111011011", -- t[21467] = 3
      "000011" when "0101001111011100", -- t[21468] = 3
      "000011" when "0101001111011101", -- t[21469] = 3
      "000011" when "0101001111011110", -- t[21470] = 3
      "000011" when "0101001111011111", -- t[21471] = 3
      "000011" when "0101001111100000", -- t[21472] = 3
      "000011" when "0101001111100001", -- t[21473] = 3
      "000011" when "0101001111100010", -- t[21474] = 3
      "000011" when "0101001111100011", -- t[21475] = 3
      "000011" when "0101001111100100", -- t[21476] = 3
      "000011" when "0101001111100101", -- t[21477] = 3
      "000011" when "0101001111100110", -- t[21478] = 3
      "000011" when "0101001111100111", -- t[21479] = 3
      "000011" when "0101001111101000", -- t[21480] = 3
      "000011" when "0101001111101001", -- t[21481] = 3
      "000011" when "0101001111101010", -- t[21482] = 3
      "000011" when "0101001111101011", -- t[21483] = 3
      "000011" when "0101001111101100", -- t[21484] = 3
      "000011" when "0101001111101101", -- t[21485] = 3
      "000011" when "0101001111101110", -- t[21486] = 3
      "000011" when "0101001111101111", -- t[21487] = 3
      "000011" when "0101001111110000", -- t[21488] = 3
      "000011" when "0101001111110001", -- t[21489] = 3
      "000011" when "0101001111110010", -- t[21490] = 3
      "000011" when "0101001111110011", -- t[21491] = 3
      "000011" when "0101001111110100", -- t[21492] = 3
      "000011" when "0101001111110101", -- t[21493] = 3
      "000011" when "0101001111110110", -- t[21494] = 3
      "000011" when "0101001111110111", -- t[21495] = 3
      "000011" when "0101001111111000", -- t[21496] = 3
      "000011" when "0101001111111001", -- t[21497] = 3
      "000011" when "0101001111111010", -- t[21498] = 3
      "000011" when "0101001111111011", -- t[21499] = 3
      "000011" when "0101001111111100", -- t[21500] = 3
      "000011" when "0101001111111101", -- t[21501] = 3
      "000011" when "0101001111111110", -- t[21502] = 3
      "000011" when "0101001111111111", -- t[21503] = 3
      "000011" when "0101010000000000", -- t[21504] = 3
      "000011" when "0101010000000001", -- t[21505] = 3
      "000011" when "0101010000000010", -- t[21506] = 3
      "000011" when "0101010000000011", -- t[21507] = 3
      "000011" when "0101010000000100", -- t[21508] = 3
      "000011" when "0101010000000101", -- t[21509] = 3
      "000011" when "0101010000000110", -- t[21510] = 3
      "000011" when "0101010000000111", -- t[21511] = 3
      "000011" when "0101010000001000", -- t[21512] = 3
      "000011" when "0101010000001001", -- t[21513] = 3
      "000011" when "0101010000001010", -- t[21514] = 3
      "000011" when "0101010000001011", -- t[21515] = 3
      "000011" when "0101010000001100", -- t[21516] = 3
      "000011" when "0101010000001101", -- t[21517] = 3
      "000011" when "0101010000001110", -- t[21518] = 3
      "000011" when "0101010000001111", -- t[21519] = 3
      "000011" when "0101010000010000", -- t[21520] = 3
      "000011" when "0101010000010001", -- t[21521] = 3
      "000011" when "0101010000010010", -- t[21522] = 3
      "000011" when "0101010000010011", -- t[21523] = 3
      "000011" when "0101010000010100", -- t[21524] = 3
      "000011" when "0101010000010101", -- t[21525] = 3
      "000011" when "0101010000010110", -- t[21526] = 3
      "000011" when "0101010000010111", -- t[21527] = 3
      "000011" when "0101010000011000", -- t[21528] = 3
      "000011" when "0101010000011001", -- t[21529] = 3
      "000011" when "0101010000011010", -- t[21530] = 3
      "000011" when "0101010000011011", -- t[21531] = 3
      "000011" when "0101010000011100", -- t[21532] = 3
      "000011" when "0101010000011101", -- t[21533] = 3
      "000011" when "0101010000011110", -- t[21534] = 3
      "000011" when "0101010000011111", -- t[21535] = 3
      "000011" when "0101010000100000", -- t[21536] = 3
      "000011" when "0101010000100001", -- t[21537] = 3
      "000011" when "0101010000100010", -- t[21538] = 3
      "000011" when "0101010000100011", -- t[21539] = 3
      "000011" when "0101010000100100", -- t[21540] = 3
      "000011" when "0101010000100101", -- t[21541] = 3
      "000011" when "0101010000100110", -- t[21542] = 3
      "000011" when "0101010000100111", -- t[21543] = 3
      "000011" when "0101010000101000", -- t[21544] = 3
      "000011" when "0101010000101001", -- t[21545] = 3
      "000011" when "0101010000101010", -- t[21546] = 3
      "000011" when "0101010000101011", -- t[21547] = 3
      "000011" when "0101010000101100", -- t[21548] = 3
      "000011" when "0101010000101101", -- t[21549] = 3
      "000011" when "0101010000101110", -- t[21550] = 3
      "000011" when "0101010000101111", -- t[21551] = 3
      "000011" when "0101010000110000", -- t[21552] = 3
      "000011" when "0101010000110001", -- t[21553] = 3
      "000011" when "0101010000110010", -- t[21554] = 3
      "000011" when "0101010000110011", -- t[21555] = 3
      "000011" when "0101010000110100", -- t[21556] = 3
      "000011" when "0101010000110101", -- t[21557] = 3
      "000011" when "0101010000110110", -- t[21558] = 3
      "000011" when "0101010000110111", -- t[21559] = 3
      "000011" when "0101010000111000", -- t[21560] = 3
      "000011" when "0101010000111001", -- t[21561] = 3
      "000011" when "0101010000111010", -- t[21562] = 3
      "000011" when "0101010000111011", -- t[21563] = 3
      "000011" when "0101010000111100", -- t[21564] = 3
      "000011" when "0101010000111101", -- t[21565] = 3
      "000011" when "0101010000111110", -- t[21566] = 3
      "000011" when "0101010000111111", -- t[21567] = 3
      "000011" when "0101010001000000", -- t[21568] = 3
      "000011" when "0101010001000001", -- t[21569] = 3
      "000011" when "0101010001000010", -- t[21570] = 3
      "000011" when "0101010001000011", -- t[21571] = 3
      "000011" when "0101010001000100", -- t[21572] = 3
      "000011" when "0101010001000101", -- t[21573] = 3
      "000011" when "0101010001000110", -- t[21574] = 3
      "000011" when "0101010001000111", -- t[21575] = 3
      "000011" when "0101010001001000", -- t[21576] = 3
      "000011" when "0101010001001001", -- t[21577] = 3
      "000011" when "0101010001001010", -- t[21578] = 3
      "000011" when "0101010001001011", -- t[21579] = 3
      "000011" when "0101010001001100", -- t[21580] = 3
      "000011" when "0101010001001101", -- t[21581] = 3
      "000011" when "0101010001001110", -- t[21582] = 3
      "000011" when "0101010001001111", -- t[21583] = 3
      "000011" when "0101010001010000", -- t[21584] = 3
      "000011" when "0101010001010001", -- t[21585] = 3
      "000011" when "0101010001010010", -- t[21586] = 3
      "000011" when "0101010001010011", -- t[21587] = 3
      "000011" when "0101010001010100", -- t[21588] = 3
      "000011" when "0101010001010101", -- t[21589] = 3
      "000011" when "0101010001010110", -- t[21590] = 3
      "000011" when "0101010001010111", -- t[21591] = 3
      "000011" when "0101010001011000", -- t[21592] = 3
      "000011" when "0101010001011001", -- t[21593] = 3
      "000011" when "0101010001011010", -- t[21594] = 3
      "000011" when "0101010001011011", -- t[21595] = 3
      "000011" when "0101010001011100", -- t[21596] = 3
      "000011" when "0101010001011101", -- t[21597] = 3
      "000011" when "0101010001011110", -- t[21598] = 3
      "000011" when "0101010001011111", -- t[21599] = 3
      "000011" when "0101010001100000", -- t[21600] = 3
      "000011" when "0101010001100001", -- t[21601] = 3
      "000011" when "0101010001100010", -- t[21602] = 3
      "000011" when "0101010001100011", -- t[21603] = 3
      "000011" when "0101010001100100", -- t[21604] = 3
      "000011" when "0101010001100101", -- t[21605] = 3
      "000011" when "0101010001100110", -- t[21606] = 3
      "000011" when "0101010001100111", -- t[21607] = 3
      "000011" when "0101010001101000", -- t[21608] = 3
      "000011" when "0101010001101001", -- t[21609] = 3
      "000011" when "0101010001101010", -- t[21610] = 3
      "000011" when "0101010001101011", -- t[21611] = 3
      "000011" when "0101010001101100", -- t[21612] = 3
      "000011" when "0101010001101101", -- t[21613] = 3
      "000011" when "0101010001101110", -- t[21614] = 3
      "000011" when "0101010001101111", -- t[21615] = 3
      "000011" when "0101010001110000", -- t[21616] = 3
      "000011" when "0101010001110001", -- t[21617] = 3
      "000011" when "0101010001110010", -- t[21618] = 3
      "000011" when "0101010001110011", -- t[21619] = 3
      "000100" when "0101010001110100", -- t[21620] = 4
      "000100" when "0101010001110101", -- t[21621] = 4
      "000100" when "0101010001110110", -- t[21622] = 4
      "000100" when "0101010001110111", -- t[21623] = 4
      "000100" when "0101010001111000", -- t[21624] = 4
      "000100" when "0101010001111001", -- t[21625] = 4
      "000100" when "0101010001111010", -- t[21626] = 4
      "000100" when "0101010001111011", -- t[21627] = 4
      "000100" when "0101010001111100", -- t[21628] = 4
      "000100" when "0101010001111101", -- t[21629] = 4
      "000100" when "0101010001111110", -- t[21630] = 4
      "000100" when "0101010001111111", -- t[21631] = 4
      "000100" when "0101010010000000", -- t[21632] = 4
      "000100" when "0101010010000001", -- t[21633] = 4
      "000100" when "0101010010000010", -- t[21634] = 4
      "000100" when "0101010010000011", -- t[21635] = 4
      "000100" when "0101010010000100", -- t[21636] = 4
      "000100" when "0101010010000101", -- t[21637] = 4
      "000100" when "0101010010000110", -- t[21638] = 4
      "000100" when "0101010010000111", -- t[21639] = 4
      "000100" when "0101010010001000", -- t[21640] = 4
      "000100" when "0101010010001001", -- t[21641] = 4
      "000100" when "0101010010001010", -- t[21642] = 4
      "000100" when "0101010010001011", -- t[21643] = 4
      "000100" when "0101010010001100", -- t[21644] = 4
      "000100" when "0101010010001101", -- t[21645] = 4
      "000100" when "0101010010001110", -- t[21646] = 4
      "000100" when "0101010010001111", -- t[21647] = 4
      "000100" when "0101010010010000", -- t[21648] = 4
      "000100" when "0101010010010001", -- t[21649] = 4
      "000100" when "0101010010010010", -- t[21650] = 4
      "000100" when "0101010010010011", -- t[21651] = 4
      "000100" when "0101010010010100", -- t[21652] = 4
      "000100" when "0101010010010101", -- t[21653] = 4
      "000100" when "0101010010010110", -- t[21654] = 4
      "000100" when "0101010010010111", -- t[21655] = 4
      "000100" when "0101010010011000", -- t[21656] = 4
      "000100" when "0101010010011001", -- t[21657] = 4
      "000100" when "0101010010011010", -- t[21658] = 4
      "000100" when "0101010010011011", -- t[21659] = 4
      "000100" when "0101010010011100", -- t[21660] = 4
      "000100" when "0101010010011101", -- t[21661] = 4
      "000100" when "0101010010011110", -- t[21662] = 4
      "000100" when "0101010010011111", -- t[21663] = 4
      "000100" when "0101010010100000", -- t[21664] = 4
      "000100" when "0101010010100001", -- t[21665] = 4
      "000100" when "0101010010100010", -- t[21666] = 4
      "000100" when "0101010010100011", -- t[21667] = 4
      "000100" when "0101010010100100", -- t[21668] = 4
      "000100" when "0101010010100101", -- t[21669] = 4
      "000100" when "0101010010100110", -- t[21670] = 4
      "000100" when "0101010010100111", -- t[21671] = 4
      "000100" when "0101010010101000", -- t[21672] = 4
      "000100" when "0101010010101001", -- t[21673] = 4
      "000100" when "0101010010101010", -- t[21674] = 4
      "000100" when "0101010010101011", -- t[21675] = 4
      "000100" when "0101010010101100", -- t[21676] = 4
      "000100" when "0101010010101101", -- t[21677] = 4
      "000100" when "0101010010101110", -- t[21678] = 4
      "000100" when "0101010010101111", -- t[21679] = 4
      "000100" when "0101010010110000", -- t[21680] = 4
      "000100" when "0101010010110001", -- t[21681] = 4
      "000100" when "0101010010110010", -- t[21682] = 4
      "000100" when "0101010010110011", -- t[21683] = 4
      "000100" when "0101010010110100", -- t[21684] = 4
      "000100" when "0101010010110101", -- t[21685] = 4
      "000100" when "0101010010110110", -- t[21686] = 4
      "000100" when "0101010010110111", -- t[21687] = 4
      "000100" when "0101010010111000", -- t[21688] = 4
      "000100" when "0101010010111001", -- t[21689] = 4
      "000100" when "0101010010111010", -- t[21690] = 4
      "000100" when "0101010010111011", -- t[21691] = 4
      "000100" when "0101010010111100", -- t[21692] = 4
      "000100" when "0101010010111101", -- t[21693] = 4
      "000100" when "0101010010111110", -- t[21694] = 4
      "000100" when "0101010010111111", -- t[21695] = 4
      "000100" when "0101010011000000", -- t[21696] = 4
      "000100" when "0101010011000001", -- t[21697] = 4
      "000100" when "0101010011000010", -- t[21698] = 4
      "000100" when "0101010011000011", -- t[21699] = 4
      "000100" when "0101010011000100", -- t[21700] = 4
      "000100" when "0101010011000101", -- t[21701] = 4
      "000100" when "0101010011000110", -- t[21702] = 4
      "000100" when "0101010011000111", -- t[21703] = 4
      "000100" when "0101010011001000", -- t[21704] = 4
      "000100" when "0101010011001001", -- t[21705] = 4
      "000100" when "0101010011001010", -- t[21706] = 4
      "000100" when "0101010011001011", -- t[21707] = 4
      "000100" when "0101010011001100", -- t[21708] = 4
      "000100" when "0101010011001101", -- t[21709] = 4
      "000100" when "0101010011001110", -- t[21710] = 4
      "000100" when "0101010011001111", -- t[21711] = 4
      "000100" when "0101010011010000", -- t[21712] = 4
      "000100" when "0101010011010001", -- t[21713] = 4
      "000100" when "0101010011010010", -- t[21714] = 4
      "000100" when "0101010011010011", -- t[21715] = 4
      "000100" when "0101010011010100", -- t[21716] = 4
      "000100" when "0101010011010101", -- t[21717] = 4
      "000100" when "0101010011010110", -- t[21718] = 4
      "000100" when "0101010011010111", -- t[21719] = 4
      "000100" when "0101010011011000", -- t[21720] = 4
      "000100" when "0101010011011001", -- t[21721] = 4
      "000100" when "0101010011011010", -- t[21722] = 4
      "000100" when "0101010011011011", -- t[21723] = 4
      "000100" when "0101010011011100", -- t[21724] = 4
      "000100" when "0101010011011101", -- t[21725] = 4
      "000100" when "0101010011011110", -- t[21726] = 4
      "000100" when "0101010011011111", -- t[21727] = 4
      "000100" when "0101010011100000", -- t[21728] = 4
      "000100" when "0101010011100001", -- t[21729] = 4
      "000100" when "0101010011100010", -- t[21730] = 4
      "000100" when "0101010011100011", -- t[21731] = 4
      "000100" when "0101010011100100", -- t[21732] = 4
      "000100" when "0101010011100101", -- t[21733] = 4
      "000100" when "0101010011100110", -- t[21734] = 4
      "000100" when "0101010011100111", -- t[21735] = 4
      "000100" when "0101010011101000", -- t[21736] = 4
      "000100" when "0101010011101001", -- t[21737] = 4
      "000100" when "0101010011101010", -- t[21738] = 4
      "000100" when "0101010011101011", -- t[21739] = 4
      "000100" when "0101010011101100", -- t[21740] = 4
      "000100" when "0101010011101101", -- t[21741] = 4
      "000100" when "0101010011101110", -- t[21742] = 4
      "000100" when "0101010011101111", -- t[21743] = 4
      "000100" when "0101010011110000", -- t[21744] = 4
      "000100" when "0101010011110001", -- t[21745] = 4
      "000100" when "0101010011110010", -- t[21746] = 4
      "000100" when "0101010011110011", -- t[21747] = 4
      "000100" when "0101010011110100", -- t[21748] = 4
      "000100" when "0101010011110101", -- t[21749] = 4
      "000100" when "0101010011110110", -- t[21750] = 4
      "000100" when "0101010011110111", -- t[21751] = 4
      "000100" when "0101010011111000", -- t[21752] = 4
      "000100" when "0101010011111001", -- t[21753] = 4
      "000100" when "0101010011111010", -- t[21754] = 4
      "000100" when "0101010011111011", -- t[21755] = 4
      "000100" when "0101010011111100", -- t[21756] = 4
      "000100" when "0101010011111101", -- t[21757] = 4
      "000100" when "0101010011111110", -- t[21758] = 4
      "000100" when "0101010011111111", -- t[21759] = 4
      "000100" when "0101010100000000", -- t[21760] = 4
      "000100" when "0101010100000001", -- t[21761] = 4
      "000100" when "0101010100000010", -- t[21762] = 4
      "000100" when "0101010100000011", -- t[21763] = 4
      "000100" when "0101010100000100", -- t[21764] = 4
      "000100" when "0101010100000101", -- t[21765] = 4
      "000100" when "0101010100000110", -- t[21766] = 4
      "000100" when "0101010100000111", -- t[21767] = 4
      "000100" when "0101010100001000", -- t[21768] = 4
      "000100" when "0101010100001001", -- t[21769] = 4
      "000100" when "0101010100001010", -- t[21770] = 4
      "000100" when "0101010100001011", -- t[21771] = 4
      "000100" when "0101010100001100", -- t[21772] = 4
      "000100" when "0101010100001101", -- t[21773] = 4
      "000100" when "0101010100001110", -- t[21774] = 4
      "000100" when "0101010100001111", -- t[21775] = 4
      "000100" when "0101010100010000", -- t[21776] = 4
      "000100" when "0101010100010001", -- t[21777] = 4
      "000100" when "0101010100010010", -- t[21778] = 4
      "000100" when "0101010100010011", -- t[21779] = 4
      "000100" when "0101010100010100", -- t[21780] = 4
      "000100" when "0101010100010101", -- t[21781] = 4
      "000100" when "0101010100010110", -- t[21782] = 4
      "000100" when "0101010100010111", -- t[21783] = 4
      "000100" when "0101010100011000", -- t[21784] = 4
      "000100" when "0101010100011001", -- t[21785] = 4
      "000100" when "0101010100011010", -- t[21786] = 4
      "000100" when "0101010100011011", -- t[21787] = 4
      "000100" when "0101010100011100", -- t[21788] = 4
      "000100" when "0101010100011101", -- t[21789] = 4
      "000100" when "0101010100011110", -- t[21790] = 4
      "000100" when "0101010100011111", -- t[21791] = 4
      "000100" when "0101010100100000", -- t[21792] = 4
      "000100" when "0101010100100001", -- t[21793] = 4
      "000100" when "0101010100100010", -- t[21794] = 4
      "000100" when "0101010100100011", -- t[21795] = 4
      "000100" when "0101010100100100", -- t[21796] = 4
      "000100" when "0101010100100101", -- t[21797] = 4
      "000100" when "0101010100100110", -- t[21798] = 4
      "000100" when "0101010100100111", -- t[21799] = 4
      "000100" when "0101010100101000", -- t[21800] = 4
      "000100" when "0101010100101001", -- t[21801] = 4
      "000100" when "0101010100101010", -- t[21802] = 4
      "000100" when "0101010100101011", -- t[21803] = 4
      "000100" when "0101010100101100", -- t[21804] = 4
      "000100" when "0101010100101101", -- t[21805] = 4
      "000100" when "0101010100101110", -- t[21806] = 4
      "000100" when "0101010100101111", -- t[21807] = 4
      "000100" when "0101010100110000", -- t[21808] = 4
      "000100" when "0101010100110001", -- t[21809] = 4
      "000100" when "0101010100110010", -- t[21810] = 4
      "000100" when "0101010100110011", -- t[21811] = 4
      "000100" when "0101010100110100", -- t[21812] = 4
      "000100" when "0101010100110101", -- t[21813] = 4
      "000100" when "0101010100110110", -- t[21814] = 4
      "000100" when "0101010100110111", -- t[21815] = 4
      "000100" when "0101010100111000", -- t[21816] = 4
      "000100" when "0101010100111001", -- t[21817] = 4
      "000100" when "0101010100111010", -- t[21818] = 4
      "000100" when "0101010100111011", -- t[21819] = 4
      "000100" when "0101010100111100", -- t[21820] = 4
      "000100" when "0101010100111101", -- t[21821] = 4
      "000100" when "0101010100111110", -- t[21822] = 4
      "000100" when "0101010100111111", -- t[21823] = 4
      "000100" when "0101010101000000", -- t[21824] = 4
      "000100" when "0101010101000001", -- t[21825] = 4
      "000100" when "0101010101000010", -- t[21826] = 4
      "000100" when "0101010101000011", -- t[21827] = 4
      "000100" when "0101010101000100", -- t[21828] = 4
      "000100" when "0101010101000101", -- t[21829] = 4
      "000100" when "0101010101000110", -- t[21830] = 4
      "000100" when "0101010101000111", -- t[21831] = 4
      "000100" when "0101010101001000", -- t[21832] = 4
      "000100" when "0101010101001001", -- t[21833] = 4
      "000100" when "0101010101001010", -- t[21834] = 4
      "000100" when "0101010101001011", -- t[21835] = 4
      "000100" when "0101010101001100", -- t[21836] = 4
      "000100" when "0101010101001101", -- t[21837] = 4
      "000100" when "0101010101001110", -- t[21838] = 4
      "000100" when "0101010101001111", -- t[21839] = 4
      "000100" when "0101010101010000", -- t[21840] = 4
      "000100" when "0101010101010001", -- t[21841] = 4
      "000100" when "0101010101010010", -- t[21842] = 4
      "000100" when "0101010101010011", -- t[21843] = 4
      "000100" when "0101010101010100", -- t[21844] = 4
      "000100" when "0101010101010101", -- t[21845] = 4
      "000100" when "0101010101010110", -- t[21846] = 4
      "000100" when "0101010101010111", -- t[21847] = 4
      "000100" when "0101010101011000", -- t[21848] = 4
      "000100" when "0101010101011001", -- t[21849] = 4
      "000100" when "0101010101011010", -- t[21850] = 4
      "000100" when "0101010101011011", -- t[21851] = 4
      "000100" when "0101010101011100", -- t[21852] = 4
      "000100" when "0101010101011101", -- t[21853] = 4
      "000100" when "0101010101011110", -- t[21854] = 4
      "000100" when "0101010101011111", -- t[21855] = 4
      "000100" when "0101010101100000", -- t[21856] = 4
      "000100" when "0101010101100001", -- t[21857] = 4
      "000100" when "0101010101100010", -- t[21858] = 4
      "000100" when "0101010101100011", -- t[21859] = 4
      "000100" when "0101010101100100", -- t[21860] = 4
      "000100" when "0101010101100101", -- t[21861] = 4
      "000100" when "0101010101100110", -- t[21862] = 4
      "000100" when "0101010101100111", -- t[21863] = 4
      "000100" when "0101010101101000", -- t[21864] = 4
      "000100" when "0101010101101001", -- t[21865] = 4
      "000100" when "0101010101101010", -- t[21866] = 4
      "000100" when "0101010101101011", -- t[21867] = 4
      "000100" when "0101010101101100", -- t[21868] = 4
      "000100" when "0101010101101101", -- t[21869] = 4
      "000100" when "0101010101101110", -- t[21870] = 4
      "000100" when "0101010101101111", -- t[21871] = 4
      "000100" when "0101010101110000", -- t[21872] = 4
      "000100" when "0101010101110001", -- t[21873] = 4
      "000100" when "0101010101110010", -- t[21874] = 4
      "000100" when "0101010101110011", -- t[21875] = 4
      "000100" when "0101010101110100", -- t[21876] = 4
      "000100" when "0101010101110101", -- t[21877] = 4
      "000100" when "0101010101110110", -- t[21878] = 4
      "000100" when "0101010101110111", -- t[21879] = 4
      "000100" when "0101010101111000", -- t[21880] = 4
      "000100" when "0101010101111001", -- t[21881] = 4
      "000100" when "0101010101111010", -- t[21882] = 4
      "000100" when "0101010101111011", -- t[21883] = 4
      "000100" when "0101010101111100", -- t[21884] = 4
      "000100" when "0101010101111101", -- t[21885] = 4
      "000100" when "0101010101111110", -- t[21886] = 4
      "000100" when "0101010101111111", -- t[21887] = 4
      "000100" when "0101010110000000", -- t[21888] = 4
      "000100" when "0101010110000001", -- t[21889] = 4
      "000100" when "0101010110000010", -- t[21890] = 4
      "000100" when "0101010110000011", -- t[21891] = 4
      "000100" when "0101010110000100", -- t[21892] = 4
      "000100" when "0101010110000101", -- t[21893] = 4
      "000100" when "0101010110000110", -- t[21894] = 4
      "000100" when "0101010110000111", -- t[21895] = 4
      "000100" when "0101010110001000", -- t[21896] = 4
      "000100" when "0101010110001001", -- t[21897] = 4
      "000100" when "0101010110001010", -- t[21898] = 4
      "000100" when "0101010110001011", -- t[21899] = 4
      "000100" when "0101010110001100", -- t[21900] = 4
      "000100" when "0101010110001101", -- t[21901] = 4
      "000100" when "0101010110001110", -- t[21902] = 4
      "000100" when "0101010110001111", -- t[21903] = 4
      "000100" when "0101010110010000", -- t[21904] = 4
      "000100" when "0101010110010001", -- t[21905] = 4
      "000100" when "0101010110010010", -- t[21906] = 4
      "000100" when "0101010110010011", -- t[21907] = 4
      "000100" when "0101010110010100", -- t[21908] = 4
      "000100" when "0101010110010101", -- t[21909] = 4
      "000100" when "0101010110010110", -- t[21910] = 4
      "000100" when "0101010110010111", -- t[21911] = 4
      "000100" when "0101010110011000", -- t[21912] = 4
      "000100" when "0101010110011001", -- t[21913] = 4
      "000100" when "0101010110011010", -- t[21914] = 4
      "000100" when "0101010110011011", -- t[21915] = 4
      "000100" when "0101010110011100", -- t[21916] = 4
      "000100" when "0101010110011101", -- t[21917] = 4
      "000100" when "0101010110011110", -- t[21918] = 4
      "000100" when "0101010110011111", -- t[21919] = 4
      "000100" when "0101010110100000", -- t[21920] = 4
      "000100" when "0101010110100001", -- t[21921] = 4
      "000100" when "0101010110100010", -- t[21922] = 4
      "000100" when "0101010110100011", -- t[21923] = 4
      "000100" when "0101010110100100", -- t[21924] = 4
      "000100" when "0101010110100101", -- t[21925] = 4
      "000100" when "0101010110100110", -- t[21926] = 4
      "000100" when "0101010110100111", -- t[21927] = 4
      "000100" when "0101010110101000", -- t[21928] = 4
      "000100" when "0101010110101001", -- t[21929] = 4
      "000100" when "0101010110101010", -- t[21930] = 4
      "000100" when "0101010110101011", -- t[21931] = 4
      "000100" when "0101010110101100", -- t[21932] = 4
      "000100" when "0101010110101101", -- t[21933] = 4
      "000100" when "0101010110101110", -- t[21934] = 4
      "000100" when "0101010110101111", -- t[21935] = 4
      "000100" when "0101010110110000", -- t[21936] = 4
      "000100" when "0101010110110001", -- t[21937] = 4
      "000100" when "0101010110110010", -- t[21938] = 4
      "000100" when "0101010110110011", -- t[21939] = 4
      "000100" when "0101010110110100", -- t[21940] = 4
      "000100" when "0101010110110101", -- t[21941] = 4
      "000100" when "0101010110110110", -- t[21942] = 4
      "000100" when "0101010110110111", -- t[21943] = 4
      "000100" when "0101010110111000", -- t[21944] = 4
      "000100" when "0101010110111001", -- t[21945] = 4
      "000100" when "0101010110111010", -- t[21946] = 4
      "000100" when "0101010110111011", -- t[21947] = 4
      "000100" when "0101010110111100", -- t[21948] = 4
      "000100" when "0101010110111101", -- t[21949] = 4
      "000100" when "0101010110111110", -- t[21950] = 4
      "000100" when "0101010110111111", -- t[21951] = 4
      "000100" when "0101010111000000", -- t[21952] = 4
      "000100" when "0101010111000001", -- t[21953] = 4
      "000100" when "0101010111000010", -- t[21954] = 4
      "000100" when "0101010111000011", -- t[21955] = 4
      "000100" when "0101010111000100", -- t[21956] = 4
      "000100" when "0101010111000101", -- t[21957] = 4
      "000100" when "0101010111000110", -- t[21958] = 4
      "000100" when "0101010111000111", -- t[21959] = 4
      "000100" when "0101010111001000", -- t[21960] = 4
      "000100" when "0101010111001001", -- t[21961] = 4
      "000100" when "0101010111001010", -- t[21962] = 4
      "000100" when "0101010111001011", -- t[21963] = 4
      "000100" when "0101010111001100", -- t[21964] = 4
      "000100" when "0101010111001101", -- t[21965] = 4
      "000100" when "0101010111001110", -- t[21966] = 4
      "000100" when "0101010111001111", -- t[21967] = 4
      "000100" when "0101010111010000", -- t[21968] = 4
      "000100" when "0101010111010001", -- t[21969] = 4
      "000100" when "0101010111010010", -- t[21970] = 4
      "000100" when "0101010111010011", -- t[21971] = 4
      "000100" when "0101010111010100", -- t[21972] = 4
      "000100" when "0101010111010101", -- t[21973] = 4
      "000100" when "0101010111010110", -- t[21974] = 4
      "000100" when "0101010111010111", -- t[21975] = 4
      "000100" when "0101010111011000", -- t[21976] = 4
      "000100" when "0101010111011001", -- t[21977] = 4
      "000100" when "0101010111011010", -- t[21978] = 4
      "000100" when "0101010111011011", -- t[21979] = 4
      "000100" when "0101010111011100", -- t[21980] = 4
      "000100" when "0101010111011101", -- t[21981] = 4
      "000100" when "0101010111011110", -- t[21982] = 4
      "000100" when "0101010111011111", -- t[21983] = 4
      "000100" when "0101010111100000", -- t[21984] = 4
      "000100" when "0101010111100001", -- t[21985] = 4
      "000100" when "0101010111100010", -- t[21986] = 4
      "000100" when "0101010111100011", -- t[21987] = 4
      "000100" when "0101010111100100", -- t[21988] = 4
      "000100" when "0101010111100101", -- t[21989] = 4
      "000100" when "0101010111100110", -- t[21990] = 4
      "000100" when "0101010111100111", -- t[21991] = 4
      "000100" when "0101010111101000", -- t[21992] = 4
      "000100" when "0101010111101001", -- t[21993] = 4
      "000100" when "0101010111101010", -- t[21994] = 4
      "000100" when "0101010111101011", -- t[21995] = 4
      "000100" when "0101010111101100", -- t[21996] = 4
      "000100" when "0101010111101101", -- t[21997] = 4
      "000100" when "0101010111101110", -- t[21998] = 4
      "000100" when "0101010111101111", -- t[21999] = 4
      "000100" when "0101010111110000", -- t[22000] = 4
      "000100" when "0101010111110001", -- t[22001] = 4
      "000100" when "0101010111110010", -- t[22002] = 4
      "000100" when "0101010111110011", -- t[22003] = 4
      "000100" when "0101010111110100", -- t[22004] = 4
      "000100" when "0101010111110101", -- t[22005] = 4
      "000100" when "0101010111110110", -- t[22006] = 4
      "000100" when "0101010111110111", -- t[22007] = 4
      "000100" when "0101010111111000", -- t[22008] = 4
      "000100" when "0101010111111001", -- t[22009] = 4
      "000100" when "0101010111111010", -- t[22010] = 4
      "000100" when "0101010111111011", -- t[22011] = 4
      "000100" when "0101010111111100", -- t[22012] = 4
      "000100" when "0101010111111101", -- t[22013] = 4
      "000100" when "0101010111111110", -- t[22014] = 4
      "000100" when "0101010111111111", -- t[22015] = 4
      "000100" when "0101011000000000", -- t[22016] = 4
      "000100" when "0101011000000001", -- t[22017] = 4
      "000100" when "0101011000000010", -- t[22018] = 4
      "000100" when "0101011000000011", -- t[22019] = 4
      "000100" when "0101011000000100", -- t[22020] = 4
      "000100" when "0101011000000101", -- t[22021] = 4
      "000100" when "0101011000000110", -- t[22022] = 4
      "000100" when "0101011000000111", -- t[22023] = 4
      "000100" when "0101011000001000", -- t[22024] = 4
      "000100" when "0101011000001001", -- t[22025] = 4
      "000100" when "0101011000001010", -- t[22026] = 4
      "000100" when "0101011000001011", -- t[22027] = 4
      "000100" when "0101011000001100", -- t[22028] = 4
      "000100" when "0101011000001101", -- t[22029] = 4
      "000100" when "0101011000001110", -- t[22030] = 4
      "000100" when "0101011000001111", -- t[22031] = 4
      "000100" when "0101011000010000", -- t[22032] = 4
      "000100" when "0101011000010001", -- t[22033] = 4
      "000100" when "0101011000010010", -- t[22034] = 4
      "000100" when "0101011000010011", -- t[22035] = 4
      "000100" when "0101011000010100", -- t[22036] = 4
      "000100" when "0101011000010101", -- t[22037] = 4
      "000100" when "0101011000010110", -- t[22038] = 4
      "000100" when "0101011000010111", -- t[22039] = 4
      "000100" when "0101011000011000", -- t[22040] = 4
      "000100" when "0101011000011001", -- t[22041] = 4
      "000100" when "0101011000011010", -- t[22042] = 4
      "000100" when "0101011000011011", -- t[22043] = 4
      "000100" when "0101011000011100", -- t[22044] = 4
      "000100" when "0101011000011101", -- t[22045] = 4
      "000100" when "0101011000011110", -- t[22046] = 4
      "000100" when "0101011000011111", -- t[22047] = 4
      "000100" when "0101011000100000", -- t[22048] = 4
      "000100" when "0101011000100001", -- t[22049] = 4
      "000100" when "0101011000100010", -- t[22050] = 4
      "000100" when "0101011000100011", -- t[22051] = 4
      "000100" when "0101011000100100", -- t[22052] = 4
      "000100" when "0101011000100101", -- t[22053] = 4
      "000100" when "0101011000100110", -- t[22054] = 4
      "000100" when "0101011000100111", -- t[22055] = 4
      "000100" when "0101011000101000", -- t[22056] = 4
      "000100" when "0101011000101001", -- t[22057] = 4
      "000100" when "0101011000101010", -- t[22058] = 4
      "000100" when "0101011000101011", -- t[22059] = 4
      "000100" when "0101011000101100", -- t[22060] = 4
      "000100" when "0101011000101101", -- t[22061] = 4
      "000100" when "0101011000101110", -- t[22062] = 4
      "000100" when "0101011000101111", -- t[22063] = 4
      "000100" when "0101011000110000", -- t[22064] = 4
      "000100" when "0101011000110001", -- t[22065] = 4
      "000100" when "0101011000110010", -- t[22066] = 4
      "000100" when "0101011000110011", -- t[22067] = 4
      "000100" when "0101011000110100", -- t[22068] = 4
      "000100" when "0101011000110101", -- t[22069] = 4
      "000100" when "0101011000110110", -- t[22070] = 4
      "000100" when "0101011000110111", -- t[22071] = 4
      "000100" when "0101011000111000", -- t[22072] = 4
      "000100" when "0101011000111001", -- t[22073] = 4
      "000100" when "0101011000111010", -- t[22074] = 4
      "000100" when "0101011000111011", -- t[22075] = 4
      "000100" when "0101011000111100", -- t[22076] = 4
      "000100" when "0101011000111101", -- t[22077] = 4
      "000100" when "0101011000111110", -- t[22078] = 4
      "000100" when "0101011000111111", -- t[22079] = 4
      "000100" when "0101011001000000", -- t[22080] = 4
      "000100" when "0101011001000001", -- t[22081] = 4
      "000100" when "0101011001000010", -- t[22082] = 4
      "000100" when "0101011001000011", -- t[22083] = 4
      "000100" when "0101011001000100", -- t[22084] = 4
      "000100" when "0101011001000101", -- t[22085] = 4
      "000100" when "0101011001000110", -- t[22086] = 4
      "000100" when "0101011001000111", -- t[22087] = 4
      "000100" when "0101011001001000", -- t[22088] = 4
      "000100" when "0101011001001001", -- t[22089] = 4
      "000100" when "0101011001001010", -- t[22090] = 4
      "000100" when "0101011001001011", -- t[22091] = 4
      "000100" when "0101011001001100", -- t[22092] = 4
      "000100" when "0101011001001101", -- t[22093] = 4
      "000100" when "0101011001001110", -- t[22094] = 4
      "000100" when "0101011001001111", -- t[22095] = 4
      "000100" when "0101011001010000", -- t[22096] = 4
      "000100" when "0101011001010001", -- t[22097] = 4
      "000100" when "0101011001010010", -- t[22098] = 4
      "000100" when "0101011001010011", -- t[22099] = 4
      "000100" when "0101011001010100", -- t[22100] = 4
      "000100" when "0101011001010101", -- t[22101] = 4
      "000100" when "0101011001010110", -- t[22102] = 4
      "000100" when "0101011001010111", -- t[22103] = 4
      "000100" when "0101011001011000", -- t[22104] = 4
      "000100" when "0101011001011001", -- t[22105] = 4
      "000100" when "0101011001011010", -- t[22106] = 4
      "000100" when "0101011001011011", -- t[22107] = 4
      "000100" when "0101011001011100", -- t[22108] = 4
      "000100" when "0101011001011101", -- t[22109] = 4
      "000100" when "0101011001011110", -- t[22110] = 4
      "000100" when "0101011001011111", -- t[22111] = 4
      "000100" when "0101011001100000", -- t[22112] = 4
      "000100" when "0101011001100001", -- t[22113] = 4
      "000100" when "0101011001100010", -- t[22114] = 4
      "000100" when "0101011001100011", -- t[22115] = 4
      "000100" when "0101011001100100", -- t[22116] = 4
      "000100" when "0101011001100101", -- t[22117] = 4
      "000100" when "0101011001100110", -- t[22118] = 4
      "000100" when "0101011001100111", -- t[22119] = 4
      "000100" when "0101011001101000", -- t[22120] = 4
      "000100" when "0101011001101001", -- t[22121] = 4
      "000100" when "0101011001101010", -- t[22122] = 4
      "000100" when "0101011001101011", -- t[22123] = 4
      "000100" when "0101011001101100", -- t[22124] = 4
      "000100" when "0101011001101101", -- t[22125] = 4
      "000100" when "0101011001101110", -- t[22126] = 4
      "000100" when "0101011001101111", -- t[22127] = 4
      "000100" when "0101011001110000", -- t[22128] = 4
      "000100" when "0101011001110001", -- t[22129] = 4
      "000100" when "0101011001110010", -- t[22130] = 4
      "000100" when "0101011001110011", -- t[22131] = 4
      "000100" when "0101011001110100", -- t[22132] = 4
      "000100" when "0101011001110101", -- t[22133] = 4
      "000100" when "0101011001110110", -- t[22134] = 4
      "000100" when "0101011001110111", -- t[22135] = 4
      "000100" when "0101011001111000", -- t[22136] = 4
      "000100" when "0101011001111001", -- t[22137] = 4
      "000100" when "0101011001111010", -- t[22138] = 4
      "000100" when "0101011001111011", -- t[22139] = 4
      "000100" when "0101011001111100", -- t[22140] = 4
      "000100" when "0101011001111101", -- t[22141] = 4
      "000100" when "0101011001111110", -- t[22142] = 4
      "000100" when "0101011001111111", -- t[22143] = 4
      "000100" when "0101011010000000", -- t[22144] = 4
      "000100" when "0101011010000001", -- t[22145] = 4
      "000100" when "0101011010000010", -- t[22146] = 4
      "000100" when "0101011010000011", -- t[22147] = 4
      "000100" when "0101011010000100", -- t[22148] = 4
      "000100" when "0101011010000101", -- t[22149] = 4
      "000100" when "0101011010000110", -- t[22150] = 4
      "000100" when "0101011010000111", -- t[22151] = 4
      "000100" when "0101011010001000", -- t[22152] = 4
      "000100" when "0101011010001001", -- t[22153] = 4
      "000100" when "0101011010001010", -- t[22154] = 4
      "000100" when "0101011010001011", -- t[22155] = 4
      "000100" when "0101011010001100", -- t[22156] = 4
      "000100" when "0101011010001101", -- t[22157] = 4
      "000100" when "0101011010001110", -- t[22158] = 4
      "000100" when "0101011010001111", -- t[22159] = 4
      "000100" when "0101011010010000", -- t[22160] = 4
      "000100" when "0101011010010001", -- t[22161] = 4
      "000100" when "0101011010010010", -- t[22162] = 4
      "000100" when "0101011010010011", -- t[22163] = 4
      "000100" when "0101011010010100", -- t[22164] = 4
      "000100" when "0101011010010101", -- t[22165] = 4
      "000100" when "0101011010010110", -- t[22166] = 4
      "000100" when "0101011010010111", -- t[22167] = 4
      "000100" when "0101011010011000", -- t[22168] = 4
      "000100" when "0101011010011001", -- t[22169] = 4
      "000100" when "0101011010011010", -- t[22170] = 4
      "000100" when "0101011010011011", -- t[22171] = 4
      "000100" when "0101011010011100", -- t[22172] = 4
      "000100" when "0101011010011101", -- t[22173] = 4
      "000100" when "0101011010011110", -- t[22174] = 4
      "000100" when "0101011010011111", -- t[22175] = 4
      "000100" when "0101011010100000", -- t[22176] = 4
      "000100" when "0101011010100001", -- t[22177] = 4
      "000100" when "0101011010100010", -- t[22178] = 4
      "000100" when "0101011010100011", -- t[22179] = 4
      "000100" when "0101011010100100", -- t[22180] = 4
      "000100" when "0101011010100101", -- t[22181] = 4
      "000100" when "0101011010100110", -- t[22182] = 4
      "000100" when "0101011010100111", -- t[22183] = 4
      "000100" when "0101011010101000", -- t[22184] = 4
      "000100" when "0101011010101001", -- t[22185] = 4
      "000100" when "0101011010101010", -- t[22186] = 4
      "000100" when "0101011010101011", -- t[22187] = 4
      "000100" when "0101011010101100", -- t[22188] = 4
      "000100" when "0101011010101101", -- t[22189] = 4
      "000100" when "0101011010101110", -- t[22190] = 4
      "000100" when "0101011010101111", -- t[22191] = 4
      "000100" when "0101011010110000", -- t[22192] = 4
      "000100" when "0101011010110001", -- t[22193] = 4
      "000100" when "0101011010110010", -- t[22194] = 4
      "000100" when "0101011010110011", -- t[22195] = 4
      "000100" when "0101011010110100", -- t[22196] = 4
      "000100" when "0101011010110101", -- t[22197] = 4
      "000100" when "0101011010110110", -- t[22198] = 4
      "000100" when "0101011010110111", -- t[22199] = 4
      "000100" when "0101011010111000", -- t[22200] = 4
      "000100" when "0101011010111001", -- t[22201] = 4
      "000100" when "0101011010111010", -- t[22202] = 4
      "000100" when "0101011010111011", -- t[22203] = 4
      "000100" when "0101011010111100", -- t[22204] = 4
      "000100" when "0101011010111101", -- t[22205] = 4
      "000100" when "0101011010111110", -- t[22206] = 4
      "000100" when "0101011010111111", -- t[22207] = 4
      "000100" when "0101011011000000", -- t[22208] = 4
      "000100" when "0101011011000001", -- t[22209] = 4
      "000100" when "0101011011000010", -- t[22210] = 4
      "000100" when "0101011011000011", -- t[22211] = 4
      "000100" when "0101011011000100", -- t[22212] = 4
      "000100" when "0101011011000101", -- t[22213] = 4
      "000100" when "0101011011000110", -- t[22214] = 4
      "000100" when "0101011011000111", -- t[22215] = 4
      "000100" when "0101011011001000", -- t[22216] = 4
      "000100" when "0101011011001001", -- t[22217] = 4
      "000100" when "0101011011001010", -- t[22218] = 4
      "000100" when "0101011011001011", -- t[22219] = 4
      "000100" when "0101011011001100", -- t[22220] = 4
      "000100" when "0101011011001101", -- t[22221] = 4
      "000100" when "0101011011001110", -- t[22222] = 4
      "000100" when "0101011011001111", -- t[22223] = 4
      "000100" when "0101011011010000", -- t[22224] = 4
      "000100" when "0101011011010001", -- t[22225] = 4
      "000100" when "0101011011010010", -- t[22226] = 4
      "000100" when "0101011011010011", -- t[22227] = 4
      "000100" when "0101011011010100", -- t[22228] = 4
      "000100" when "0101011011010101", -- t[22229] = 4
      "000100" when "0101011011010110", -- t[22230] = 4
      "000100" when "0101011011010111", -- t[22231] = 4
      "000100" when "0101011011011000", -- t[22232] = 4
      "000100" when "0101011011011001", -- t[22233] = 4
      "000100" when "0101011011011010", -- t[22234] = 4
      "000100" when "0101011011011011", -- t[22235] = 4
      "000100" when "0101011011011100", -- t[22236] = 4
      "000100" when "0101011011011101", -- t[22237] = 4
      "000100" when "0101011011011110", -- t[22238] = 4
      "000100" when "0101011011011111", -- t[22239] = 4
      "000100" when "0101011011100000", -- t[22240] = 4
      "000100" when "0101011011100001", -- t[22241] = 4
      "000100" when "0101011011100010", -- t[22242] = 4
      "000100" when "0101011011100011", -- t[22243] = 4
      "000100" when "0101011011100100", -- t[22244] = 4
      "000100" when "0101011011100101", -- t[22245] = 4
      "000100" when "0101011011100110", -- t[22246] = 4
      "000100" when "0101011011100111", -- t[22247] = 4
      "000100" when "0101011011101000", -- t[22248] = 4
      "000100" when "0101011011101001", -- t[22249] = 4
      "000100" when "0101011011101010", -- t[22250] = 4
      "000100" when "0101011011101011", -- t[22251] = 4
      "000100" when "0101011011101100", -- t[22252] = 4
      "000100" when "0101011011101101", -- t[22253] = 4
      "000100" when "0101011011101110", -- t[22254] = 4
      "000100" when "0101011011101111", -- t[22255] = 4
      "000100" when "0101011011110000", -- t[22256] = 4
      "000100" when "0101011011110001", -- t[22257] = 4
      "000100" when "0101011011110010", -- t[22258] = 4
      "000100" when "0101011011110011", -- t[22259] = 4
      "000100" when "0101011011110100", -- t[22260] = 4
      "000100" when "0101011011110101", -- t[22261] = 4
      "000100" when "0101011011110110", -- t[22262] = 4
      "000100" when "0101011011110111", -- t[22263] = 4
      "000100" when "0101011011111000", -- t[22264] = 4
      "000100" when "0101011011111001", -- t[22265] = 4
      "000100" when "0101011011111010", -- t[22266] = 4
      "000100" when "0101011011111011", -- t[22267] = 4
      "000100" when "0101011011111100", -- t[22268] = 4
      "000100" when "0101011011111101", -- t[22269] = 4
      "000100" when "0101011011111110", -- t[22270] = 4
      "000100" when "0101011011111111", -- t[22271] = 4
      "000100" when "0101011100000000", -- t[22272] = 4
      "000100" when "0101011100000001", -- t[22273] = 4
      "000100" when "0101011100000010", -- t[22274] = 4
      "000100" when "0101011100000011", -- t[22275] = 4
      "000100" when "0101011100000100", -- t[22276] = 4
      "000100" when "0101011100000101", -- t[22277] = 4
      "000100" when "0101011100000110", -- t[22278] = 4
      "000100" when "0101011100000111", -- t[22279] = 4
      "000100" when "0101011100001000", -- t[22280] = 4
      "000100" when "0101011100001001", -- t[22281] = 4
      "000100" when "0101011100001010", -- t[22282] = 4
      "000100" when "0101011100001011", -- t[22283] = 4
      "000100" when "0101011100001100", -- t[22284] = 4
      "000100" when "0101011100001101", -- t[22285] = 4
      "000100" when "0101011100001110", -- t[22286] = 4
      "000100" when "0101011100001111", -- t[22287] = 4
      "000100" when "0101011100010000", -- t[22288] = 4
      "000100" when "0101011100010001", -- t[22289] = 4
      "000100" when "0101011100010010", -- t[22290] = 4
      "000100" when "0101011100010011", -- t[22291] = 4
      "000100" when "0101011100010100", -- t[22292] = 4
      "000100" when "0101011100010101", -- t[22293] = 4
      "000100" when "0101011100010110", -- t[22294] = 4
      "000100" when "0101011100010111", -- t[22295] = 4
      "000100" when "0101011100011000", -- t[22296] = 4
      "000100" when "0101011100011001", -- t[22297] = 4
      "000100" when "0101011100011010", -- t[22298] = 4
      "000100" when "0101011100011011", -- t[22299] = 4
      "000100" when "0101011100011100", -- t[22300] = 4
      "000100" when "0101011100011101", -- t[22301] = 4
      "000100" when "0101011100011110", -- t[22302] = 4
      "000100" when "0101011100011111", -- t[22303] = 4
      "000100" when "0101011100100000", -- t[22304] = 4
      "000100" when "0101011100100001", -- t[22305] = 4
      "000100" when "0101011100100010", -- t[22306] = 4
      "000100" when "0101011100100011", -- t[22307] = 4
      "000100" when "0101011100100100", -- t[22308] = 4
      "000100" when "0101011100100101", -- t[22309] = 4
      "000100" when "0101011100100110", -- t[22310] = 4
      "000100" when "0101011100100111", -- t[22311] = 4
      "000100" when "0101011100101000", -- t[22312] = 4
      "000100" when "0101011100101001", -- t[22313] = 4
      "000100" when "0101011100101010", -- t[22314] = 4
      "000100" when "0101011100101011", -- t[22315] = 4
      "000100" when "0101011100101100", -- t[22316] = 4
      "000100" when "0101011100101101", -- t[22317] = 4
      "000100" when "0101011100101110", -- t[22318] = 4
      "000100" when "0101011100101111", -- t[22319] = 4
      "000100" when "0101011100110000", -- t[22320] = 4
      "000100" when "0101011100110001", -- t[22321] = 4
      "000100" when "0101011100110010", -- t[22322] = 4
      "000100" when "0101011100110011", -- t[22323] = 4
      "000100" when "0101011100110100", -- t[22324] = 4
      "000100" when "0101011100110101", -- t[22325] = 4
      "000100" when "0101011100110110", -- t[22326] = 4
      "000100" when "0101011100110111", -- t[22327] = 4
      "000100" when "0101011100111000", -- t[22328] = 4
      "000100" when "0101011100111001", -- t[22329] = 4
      "000100" when "0101011100111010", -- t[22330] = 4
      "000100" when "0101011100111011", -- t[22331] = 4
      "000100" when "0101011100111100", -- t[22332] = 4
      "000100" when "0101011100111101", -- t[22333] = 4
      "000100" when "0101011100111110", -- t[22334] = 4
      "000100" when "0101011100111111", -- t[22335] = 4
      "000100" when "0101011101000000", -- t[22336] = 4
      "000100" when "0101011101000001", -- t[22337] = 4
      "000100" when "0101011101000010", -- t[22338] = 4
      "000100" when "0101011101000011", -- t[22339] = 4
      "000100" when "0101011101000100", -- t[22340] = 4
      "000100" when "0101011101000101", -- t[22341] = 4
      "000100" when "0101011101000110", -- t[22342] = 4
      "000100" when "0101011101000111", -- t[22343] = 4
      "000100" when "0101011101001000", -- t[22344] = 4
      "000100" when "0101011101001001", -- t[22345] = 4
      "000100" when "0101011101001010", -- t[22346] = 4
      "000100" when "0101011101001011", -- t[22347] = 4
      "000100" when "0101011101001100", -- t[22348] = 4
      "000100" when "0101011101001101", -- t[22349] = 4
      "000100" when "0101011101001110", -- t[22350] = 4
      "000100" when "0101011101001111", -- t[22351] = 4
      "000100" when "0101011101010000", -- t[22352] = 4
      "000100" when "0101011101010001", -- t[22353] = 4
      "000100" when "0101011101010010", -- t[22354] = 4
      "000100" when "0101011101010011", -- t[22355] = 4
      "000100" when "0101011101010100", -- t[22356] = 4
      "000100" when "0101011101010101", -- t[22357] = 4
      "000100" when "0101011101010110", -- t[22358] = 4
      "000100" when "0101011101010111", -- t[22359] = 4
      "000100" when "0101011101011000", -- t[22360] = 4
      "000100" when "0101011101011001", -- t[22361] = 4
      "000100" when "0101011101011010", -- t[22362] = 4
      "000100" when "0101011101011011", -- t[22363] = 4
      "000100" when "0101011101011100", -- t[22364] = 4
      "000100" when "0101011101011101", -- t[22365] = 4
      "000100" when "0101011101011110", -- t[22366] = 4
      "000100" when "0101011101011111", -- t[22367] = 4
      "000100" when "0101011101100000", -- t[22368] = 4
      "000100" when "0101011101100001", -- t[22369] = 4
      "000100" when "0101011101100010", -- t[22370] = 4
      "000100" when "0101011101100011", -- t[22371] = 4
      "000100" when "0101011101100100", -- t[22372] = 4
      "000100" when "0101011101100101", -- t[22373] = 4
      "000100" when "0101011101100110", -- t[22374] = 4
      "000100" when "0101011101100111", -- t[22375] = 4
      "000100" when "0101011101101000", -- t[22376] = 4
      "000100" when "0101011101101001", -- t[22377] = 4
      "000100" when "0101011101101010", -- t[22378] = 4
      "000100" when "0101011101101011", -- t[22379] = 4
      "000100" when "0101011101101100", -- t[22380] = 4
      "000100" when "0101011101101101", -- t[22381] = 4
      "000100" when "0101011101101110", -- t[22382] = 4
      "000100" when "0101011101101111", -- t[22383] = 4
      "000100" when "0101011101110000", -- t[22384] = 4
      "000100" when "0101011101110001", -- t[22385] = 4
      "000100" when "0101011101110010", -- t[22386] = 4
      "000100" when "0101011101110011", -- t[22387] = 4
      "000100" when "0101011101110100", -- t[22388] = 4
      "000100" when "0101011101110101", -- t[22389] = 4
      "000100" when "0101011101110110", -- t[22390] = 4
      "000100" when "0101011101110111", -- t[22391] = 4
      "000100" when "0101011101111000", -- t[22392] = 4
      "000100" when "0101011101111001", -- t[22393] = 4
      "000100" when "0101011101111010", -- t[22394] = 4
      "000100" when "0101011101111011", -- t[22395] = 4
      "000100" when "0101011101111100", -- t[22396] = 4
      "000100" when "0101011101111101", -- t[22397] = 4
      "000100" when "0101011101111110", -- t[22398] = 4
      "000100" when "0101011101111111", -- t[22399] = 4
      "000100" when "0101011110000000", -- t[22400] = 4
      "000100" when "0101011110000001", -- t[22401] = 4
      "000100" when "0101011110000010", -- t[22402] = 4
      "000100" when "0101011110000011", -- t[22403] = 4
      "000100" when "0101011110000100", -- t[22404] = 4
      "000100" when "0101011110000101", -- t[22405] = 4
      "000100" when "0101011110000110", -- t[22406] = 4
      "000100" when "0101011110000111", -- t[22407] = 4
      "000100" when "0101011110001000", -- t[22408] = 4
      "000100" when "0101011110001001", -- t[22409] = 4
      "000100" when "0101011110001010", -- t[22410] = 4
      "000100" when "0101011110001011", -- t[22411] = 4
      "000100" when "0101011110001100", -- t[22412] = 4
      "000100" when "0101011110001101", -- t[22413] = 4
      "000100" when "0101011110001110", -- t[22414] = 4
      "000100" when "0101011110001111", -- t[22415] = 4
      "000100" when "0101011110010000", -- t[22416] = 4
      "000100" when "0101011110010001", -- t[22417] = 4
      "000100" when "0101011110010010", -- t[22418] = 4
      "000100" when "0101011110010011", -- t[22419] = 4
      "000100" when "0101011110010100", -- t[22420] = 4
      "000100" when "0101011110010101", -- t[22421] = 4
      "000100" when "0101011110010110", -- t[22422] = 4
      "000100" when "0101011110010111", -- t[22423] = 4
      "000100" when "0101011110011000", -- t[22424] = 4
      "000100" when "0101011110011001", -- t[22425] = 4
      "000100" when "0101011110011010", -- t[22426] = 4
      "000100" when "0101011110011011", -- t[22427] = 4
      "000100" when "0101011110011100", -- t[22428] = 4
      "000100" when "0101011110011101", -- t[22429] = 4
      "000100" when "0101011110011110", -- t[22430] = 4
      "000100" when "0101011110011111", -- t[22431] = 4
      "000100" when "0101011110100000", -- t[22432] = 4
      "000100" when "0101011110100001", -- t[22433] = 4
      "000100" when "0101011110100010", -- t[22434] = 4
      "000100" when "0101011110100011", -- t[22435] = 4
      "000100" when "0101011110100100", -- t[22436] = 4
      "000100" when "0101011110100101", -- t[22437] = 4
      "000100" when "0101011110100110", -- t[22438] = 4
      "000100" when "0101011110100111", -- t[22439] = 4
      "000100" when "0101011110101000", -- t[22440] = 4
      "000100" when "0101011110101001", -- t[22441] = 4
      "000100" when "0101011110101010", -- t[22442] = 4
      "000100" when "0101011110101011", -- t[22443] = 4
      "000100" when "0101011110101100", -- t[22444] = 4
      "000100" when "0101011110101101", -- t[22445] = 4
      "000100" when "0101011110101110", -- t[22446] = 4
      "000100" when "0101011110101111", -- t[22447] = 4
      "000100" when "0101011110110000", -- t[22448] = 4
      "000100" when "0101011110110001", -- t[22449] = 4
      "000100" when "0101011110110010", -- t[22450] = 4
      "000100" when "0101011110110011", -- t[22451] = 4
      "000100" when "0101011110110100", -- t[22452] = 4
      "000100" when "0101011110110101", -- t[22453] = 4
      "000100" when "0101011110110110", -- t[22454] = 4
      "000100" when "0101011110110111", -- t[22455] = 4
      "000100" when "0101011110111000", -- t[22456] = 4
      "000100" when "0101011110111001", -- t[22457] = 4
      "000100" when "0101011110111010", -- t[22458] = 4
      "000100" when "0101011110111011", -- t[22459] = 4
      "000100" when "0101011110111100", -- t[22460] = 4
      "000100" when "0101011110111101", -- t[22461] = 4
      "000100" when "0101011110111110", -- t[22462] = 4
      "000100" when "0101011110111111", -- t[22463] = 4
      "000100" when "0101011111000000", -- t[22464] = 4
      "000100" when "0101011111000001", -- t[22465] = 4
      "000100" when "0101011111000010", -- t[22466] = 4
      "000100" when "0101011111000011", -- t[22467] = 4
      "000100" when "0101011111000100", -- t[22468] = 4
      "000100" when "0101011111000101", -- t[22469] = 4
      "000100" when "0101011111000110", -- t[22470] = 4
      "000100" when "0101011111000111", -- t[22471] = 4
      "000100" when "0101011111001000", -- t[22472] = 4
      "000100" when "0101011111001001", -- t[22473] = 4
      "000100" when "0101011111001010", -- t[22474] = 4
      "000100" when "0101011111001011", -- t[22475] = 4
      "000100" when "0101011111001100", -- t[22476] = 4
      "000100" when "0101011111001101", -- t[22477] = 4
      "000100" when "0101011111001110", -- t[22478] = 4
      "000100" when "0101011111001111", -- t[22479] = 4
      "000100" when "0101011111010000", -- t[22480] = 4
      "000100" when "0101011111010001", -- t[22481] = 4
      "000100" when "0101011111010010", -- t[22482] = 4
      "000100" when "0101011111010011", -- t[22483] = 4
      "000100" when "0101011111010100", -- t[22484] = 4
      "000100" when "0101011111010101", -- t[22485] = 4
      "000100" when "0101011111010110", -- t[22486] = 4
      "000100" when "0101011111010111", -- t[22487] = 4
      "000100" when "0101011111011000", -- t[22488] = 4
      "000100" when "0101011111011001", -- t[22489] = 4
      "000100" when "0101011111011010", -- t[22490] = 4
      "000100" when "0101011111011011", -- t[22491] = 4
      "000100" when "0101011111011100", -- t[22492] = 4
      "000100" when "0101011111011101", -- t[22493] = 4
      "000100" when "0101011111011110", -- t[22494] = 4
      "000100" when "0101011111011111", -- t[22495] = 4
      "000100" when "0101011111100000", -- t[22496] = 4
      "000100" when "0101011111100001", -- t[22497] = 4
      "000100" when "0101011111100010", -- t[22498] = 4
      "000100" when "0101011111100011", -- t[22499] = 4
      "000100" when "0101011111100100", -- t[22500] = 4
      "000100" when "0101011111100101", -- t[22501] = 4
      "000100" when "0101011111100110", -- t[22502] = 4
      "000100" when "0101011111100111", -- t[22503] = 4
      "000100" when "0101011111101000", -- t[22504] = 4
      "000100" when "0101011111101001", -- t[22505] = 4
      "000100" when "0101011111101010", -- t[22506] = 4
      "000100" when "0101011111101011", -- t[22507] = 4
      "000100" when "0101011111101100", -- t[22508] = 4
      "000100" when "0101011111101101", -- t[22509] = 4
      "000100" when "0101011111101110", -- t[22510] = 4
      "000100" when "0101011111101111", -- t[22511] = 4
      "000100" when "0101011111110000", -- t[22512] = 4
      "000100" when "0101011111110001", -- t[22513] = 4
      "000100" when "0101011111110010", -- t[22514] = 4
      "000100" when "0101011111110011", -- t[22515] = 4
      "000100" when "0101011111110100", -- t[22516] = 4
      "000100" when "0101011111110101", -- t[22517] = 4
      "000100" when "0101011111110110", -- t[22518] = 4
      "000100" when "0101011111110111", -- t[22519] = 4
      "000100" when "0101011111111000", -- t[22520] = 4
      "000100" when "0101011111111001", -- t[22521] = 4
      "000100" when "0101011111111010", -- t[22522] = 4
      "000100" when "0101011111111011", -- t[22523] = 4
      "000100" when "0101011111111100", -- t[22524] = 4
      "000100" when "0101011111111101", -- t[22525] = 4
      "000100" when "0101011111111110", -- t[22526] = 4
      "000100" when "0101011111111111", -- t[22527] = 4
      "000100" when "0101100000000000", -- t[22528] = 4
      "000100" when "0101100000000001", -- t[22529] = 4
      "000100" when "0101100000000010", -- t[22530] = 4
      "000100" when "0101100000000011", -- t[22531] = 4
      "000100" when "0101100000000100", -- t[22532] = 4
      "000100" when "0101100000000101", -- t[22533] = 4
      "000100" when "0101100000000110", -- t[22534] = 4
      "000100" when "0101100000000111", -- t[22535] = 4
      "000100" when "0101100000001000", -- t[22536] = 4
      "000100" when "0101100000001001", -- t[22537] = 4
      "000100" when "0101100000001010", -- t[22538] = 4
      "000100" when "0101100000001011", -- t[22539] = 4
      "000100" when "0101100000001100", -- t[22540] = 4
      "000100" when "0101100000001101", -- t[22541] = 4
      "000100" when "0101100000001110", -- t[22542] = 4
      "000100" when "0101100000001111", -- t[22543] = 4
      "000100" when "0101100000010000", -- t[22544] = 4
      "000100" when "0101100000010001", -- t[22545] = 4
      "000100" when "0101100000010010", -- t[22546] = 4
      "000100" when "0101100000010011", -- t[22547] = 4
      "000100" when "0101100000010100", -- t[22548] = 4
      "000100" when "0101100000010101", -- t[22549] = 4
      "000100" when "0101100000010110", -- t[22550] = 4
      "000100" when "0101100000010111", -- t[22551] = 4
      "000100" when "0101100000011000", -- t[22552] = 4
      "000100" when "0101100000011001", -- t[22553] = 4
      "000100" when "0101100000011010", -- t[22554] = 4
      "000100" when "0101100000011011", -- t[22555] = 4
      "000100" when "0101100000011100", -- t[22556] = 4
      "000100" when "0101100000011101", -- t[22557] = 4
      "000100" when "0101100000011110", -- t[22558] = 4
      "000100" when "0101100000011111", -- t[22559] = 4
      "000100" when "0101100000100000", -- t[22560] = 4
      "000100" when "0101100000100001", -- t[22561] = 4
      "000100" when "0101100000100010", -- t[22562] = 4
      "000100" when "0101100000100011", -- t[22563] = 4
      "000100" when "0101100000100100", -- t[22564] = 4
      "000100" when "0101100000100101", -- t[22565] = 4
      "000100" when "0101100000100110", -- t[22566] = 4
      "000100" when "0101100000100111", -- t[22567] = 4
      "000100" when "0101100000101000", -- t[22568] = 4
      "000100" when "0101100000101001", -- t[22569] = 4
      "000100" when "0101100000101010", -- t[22570] = 4
      "000100" when "0101100000101011", -- t[22571] = 4
      "000100" when "0101100000101100", -- t[22572] = 4
      "000100" when "0101100000101101", -- t[22573] = 4
      "000100" when "0101100000101110", -- t[22574] = 4
      "000100" when "0101100000101111", -- t[22575] = 4
      "000100" when "0101100000110000", -- t[22576] = 4
      "000100" when "0101100000110001", -- t[22577] = 4
      "000100" when "0101100000110010", -- t[22578] = 4
      "000100" when "0101100000110011", -- t[22579] = 4
      "000100" when "0101100000110100", -- t[22580] = 4
      "000100" when "0101100000110101", -- t[22581] = 4
      "000100" when "0101100000110110", -- t[22582] = 4
      "000100" when "0101100000110111", -- t[22583] = 4
      "000100" when "0101100000111000", -- t[22584] = 4
      "000100" when "0101100000111001", -- t[22585] = 4
      "000100" when "0101100000111010", -- t[22586] = 4
      "000100" when "0101100000111011", -- t[22587] = 4
      "000100" when "0101100000111100", -- t[22588] = 4
      "000100" when "0101100000111101", -- t[22589] = 4
      "000100" when "0101100000111110", -- t[22590] = 4
      "000100" when "0101100000111111", -- t[22591] = 4
      "000100" when "0101100001000000", -- t[22592] = 4
      "000100" when "0101100001000001", -- t[22593] = 4
      "000100" when "0101100001000010", -- t[22594] = 4
      "000100" when "0101100001000011", -- t[22595] = 4
      "000100" when "0101100001000100", -- t[22596] = 4
      "000100" when "0101100001000101", -- t[22597] = 4
      "000100" when "0101100001000110", -- t[22598] = 4
      "000100" when "0101100001000111", -- t[22599] = 4
      "000100" when "0101100001001000", -- t[22600] = 4
      "000100" when "0101100001001001", -- t[22601] = 4
      "000100" when "0101100001001010", -- t[22602] = 4
      "000100" when "0101100001001011", -- t[22603] = 4
      "000100" when "0101100001001100", -- t[22604] = 4
      "000100" when "0101100001001101", -- t[22605] = 4
      "000100" when "0101100001001110", -- t[22606] = 4
      "000100" when "0101100001001111", -- t[22607] = 4
      "000100" when "0101100001010000", -- t[22608] = 4
      "000100" when "0101100001010001", -- t[22609] = 4
      "000100" when "0101100001010010", -- t[22610] = 4
      "000100" when "0101100001010011", -- t[22611] = 4
      "000100" when "0101100001010100", -- t[22612] = 4
      "000100" when "0101100001010101", -- t[22613] = 4
      "000100" when "0101100001010110", -- t[22614] = 4
      "000100" when "0101100001010111", -- t[22615] = 4
      "000100" when "0101100001011000", -- t[22616] = 4
      "000100" when "0101100001011001", -- t[22617] = 4
      "000100" when "0101100001011010", -- t[22618] = 4
      "000100" when "0101100001011011", -- t[22619] = 4
      "000100" when "0101100001011100", -- t[22620] = 4
      "000100" when "0101100001011101", -- t[22621] = 4
      "000100" when "0101100001011110", -- t[22622] = 4
      "000100" when "0101100001011111", -- t[22623] = 4
      "000100" when "0101100001100000", -- t[22624] = 4
      "000100" when "0101100001100001", -- t[22625] = 4
      "000100" when "0101100001100010", -- t[22626] = 4
      "000100" when "0101100001100011", -- t[22627] = 4
      "000100" when "0101100001100100", -- t[22628] = 4
      "000100" when "0101100001100101", -- t[22629] = 4
      "000100" when "0101100001100110", -- t[22630] = 4
      "000100" when "0101100001100111", -- t[22631] = 4
      "000100" when "0101100001101000", -- t[22632] = 4
      "000100" when "0101100001101001", -- t[22633] = 4
      "000100" when "0101100001101010", -- t[22634] = 4
      "000100" when "0101100001101011", -- t[22635] = 4
      "000100" when "0101100001101100", -- t[22636] = 4
      "000100" when "0101100001101101", -- t[22637] = 4
      "000100" when "0101100001101110", -- t[22638] = 4
      "000100" when "0101100001101111", -- t[22639] = 4
      "000100" when "0101100001110000", -- t[22640] = 4
      "000100" when "0101100001110001", -- t[22641] = 4
      "000100" when "0101100001110010", -- t[22642] = 4
      "000100" when "0101100001110011", -- t[22643] = 4
      "000100" when "0101100001110100", -- t[22644] = 4
      "000100" when "0101100001110101", -- t[22645] = 4
      "000100" when "0101100001110110", -- t[22646] = 4
      "000100" when "0101100001110111", -- t[22647] = 4
      "000100" when "0101100001111000", -- t[22648] = 4
      "000100" when "0101100001111001", -- t[22649] = 4
      "000100" when "0101100001111010", -- t[22650] = 4
      "000100" when "0101100001111011", -- t[22651] = 4
      "000100" when "0101100001111100", -- t[22652] = 4
      "000100" when "0101100001111101", -- t[22653] = 4
      "000100" when "0101100001111110", -- t[22654] = 4
      "000100" when "0101100001111111", -- t[22655] = 4
      "000100" when "0101100010000000", -- t[22656] = 4
      "000100" when "0101100010000001", -- t[22657] = 4
      "000100" when "0101100010000010", -- t[22658] = 4
      "000100" when "0101100010000011", -- t[22659] = 4
      "000100" when "0101100010000100", -- t[22660] = 4
      "000100" when "0101100010000101", -- t[22661] = 4
      "000100" when "0101100010000110", -- t[22662] = 4
      "000100" when "0101100010000111", -- t[22663] = 4
      "000100" when "0101100010001000", -- t[22664] = 4
      "000100" when "0101100010001001", -- t[22665] = 4
      "000100" when "0101100010001010", -- t[22666] = 4
      "000100" when "0101100010001011", -- t[22667] = 4
      "000100" when "0101100010001100", -- t[22668] = 4
      "000100" when "0101100010001101", -- t[22669] = 4
      "000100" when "0101100010001110", -- t[22670] = 4
      "000100" when "0101100010001111", -- t[22671] = 4
      "000100" when "0101100010010000", -- t[22672] = 4
      "000100" when "0101100010010001", -- t[22673] = 4
      "000100" when "0101100010010010", -- t[22674] = 4
      "000100" when "0101100010010011", -- t[22675] = 4
      "000100" when "0101100010010100", -- t[22676] = 4
      "000100" when "0101100010010101", -- t[22677] = 4
      "000100" when "0101100010010110", -- t[22678] = 4
      "000100" when "0101100010010111", -- t[22679] = 4
      "000100" when "0101100010011000", -- t[22680] = 4
      "000100" when "0101100010011001", -- t[22681] = 4
      "000100" when "0101100010011010", -- t[22682] = 4
      "000100" when "0101100010011011", -- t[22683] = 4
      "000100" when "0101100010011100", -- t[22684] = 4
      "000100" when "0101100010011101", -- t[22685] = 4
      "000100" when "0101100010011110", -- t[22686] = 4
      "000100" when "0101100010011111", -- t[22687] = 4
      "000100" when "0101100010100000", -- t[22688] = 4
      "000100" when "0101100010100001", -- t[22689] = 4
      "000100" when "0101100010100010", -- t[22690] = 4
      "000100" when "0101100010100011", -- t[22691] = 4
      "000100" when "0101100010100100", -- t[22692] = 4
      "000100" when "0101100010100101", -- t[22693] = 4
      "000100" when "0101100010100110", -- t[22694] = 4
      "000100" when "0101100010100111", -- t[22695] = 4
      "000100" when "0101100010101000", -- t[22696] = 4
      "000100" when "0101100010101001", -- t[22697] = 4
      "000100" when "0101100010101010", -- t[22698] = 4
      "000100" when "0101100010101011", -- t[22699] = 4
      "000100" when "0101100010101100", -- t[22700] = 4
      "000100" when "0101100010101101", -- t[22701] = 4
      "000100" when "0101100010101110", -- t[22702] = 4
      "000100" when "0101100010101111", -- t[22703] = 4
      "000100" when "0101100010110000", -- t[22704] = 4
      "000100" when "0101100010110001", -- t[22705] = 4
      "000100" when "0101100010110010", -- t[22706] = 4
      "000100" when "0101100010110011", -- t[22707] = 4
      "000100" when "0101100010110100", -- t[22708] = 4
      "000100" when "0101100010110101", -- t[22709] = 4
      "000100" when "0101100010110110", -- t[22710] = 4
      "000100" when "0101100010110111", -- t[22711] = 4
      "000100" when "0101100010111000", -- t[22712] = 4
      "000100" when "0101100010111001", -- t[22713] = 4
      "000100" when "0101100010111010", -- t[22714] = 4
      "000100" when "0101100010111011", -- t[22715] = 4
      "000100" when "0101100010111100", -- t[22716] = 4
      "000100" when "0101100010111101", -- t[22717] = 4
      "000100" when "0101100010111110", -- t[22718] = 4
      "000100" when "0101100010111111", -- t[22719] = 4
      "000100" when "0101100011000000", -- t[22720] = 4
      "000100" when "0101100011000001", -- t[22721] = 4
      "000100" when "0101100011000010", -- t[22722] = 4
      "000100" when "0101100011000011", -- t[22723] = 4
      "000100" when "0101100011000100", -- t[22724] = 4
      "000100" when "0101100011000101", -- t[22725] = 4
      "000100" when "0101100011000110", -- t[22726] = 4
      "000100" when "0101100011000111", -- t[22727] = 4
      "000100" when "0101100011001000", -- t[22728] = 4
      "000100" when "0101100011001001", -- t[22729] = 4
      "000100" when "0101100011001010", -- t[22730] = 4
      "000100" when "0101100011001011", -- t[22731] = 4
      "000100" when "0101100011001100", -- t[22732] = 4
      "000100" when "0101100011001101", -- t[22733] = 4
      "000100" when "0101100011001110", -- t[22734] = 4
      "000100" when "0101100011001111", -- t[22735] = 4
      "000100" when "0101100011010000", -- t[22736] = 4
      "000100" when "0101100011010001", -- t[22737] = 4
      "000100" when "0101100011010010", -- t[22738] = 4
      "000100" when "0101100011010011", -- t[22739] = 4
      "000100" when "0101100011010100", -- t[22740] = 4
      "000100" when "0101100011010101", -- t[22741] = 4
      "000100" when "0101100011010110", -- t[22742] = 4
      "000100" when "0101100011010111", -- t[22743] = 4
      "000100" when "0101100011011000", -- t[22744] = 4
      "000100" when "0101100011011001", -- t[22745] = 4
      "000100" when "0101100011011010", -- t[22746] = 4
      "000100" when "0101100011011011", -- t[22747] = 4
      "000100" when "0101100011011100", -- t[22748] = 4
      "000100" when "0101100011011101", -- t[22749] = 4
      "000100" when "0101100011011110", -- t[22750] = 4
      "000100" when "0101100011011111", -- t[22751] = 4
      "000100" when "0101100011100000", -- t[22752] = 4
      "000100" when "0101100011100001", -- t[22753] = 4
      "000100" when "0101100011100010", -- t[22754] = 4
      "000100" when "0101100011100011", -- t[22755] = 4
      "000100" when "0101100011100100", -- t[22756] = 4
      "000100" when "0101100011100101", -- t[22757] = 4
      "000100" when "0101100011100110", -- t[22758] = 4
      "000100" when "0101100011100111", -- t[22759] = 4
      "000100" when "0101100011101000", -- t[22760] = 4
      "000100" when "0101100011101001", -- t[22761] = 4
      "000100" when "0101100011101010", -- t[22762] = 4
      "000100" when "0101100011101011", -- t[22763] = 4
      "000100" when "0101100011101100", -- t[22764] = 4
      "000100" when "0101100011101101", -- t[22765] = 4
      "000100" when "0101100011101110", -- t[22766] = 4
      "000100" when "0101100011101111", -- t[22767] = 4
      "000100" when "0101100011110000", -- t[22768] = 4
      "000100" when "0101100011110001", -- t[22769] = 4
      "000100" when "0101100011110010", -- t[22770] = 4
      "000100" when "0101100011110011", -- t[22771] = 4
      "000100" when "0101100011110100", -- t[22772] = 4
      "000100" when "0101100011110101", -- t[22773] = 4
      "000100" when "0101100011110110", -- t[22774] = 4
      "000100" when "0101100011110111", -- t[22775] = 4
      "000100" when "0101100011111000", -- t[22776] = 4
      "000100" when "0101100011111001", -- t[22777] = 4
      "000100" when "0101100011111010", -- t[22778] = 4
      "000100" when "0101100011111011", -- t[22779] = 4
      "000100" when "0101100011111100", -- t[22780] = 4
      "000100" when "0101100011111101", -- t[22781] = 4
      "000100" when "0101100011111110", -- t[22782] = 4
      "000100" when "0101100011111111", -- t[22783] = 4
      "000100" when "0101100100000000", -- t[22784] = 4
      "000100" when "0101100100000001", -- t[22785] = 4
      "000100" when "0101100100000010", -- t[22786] = 4
      "000100" when "0101100100000011", -- t[22787] = 4
      "000100" when "0101100100000100", -- t[22788] = 4
      "000100" when "0101100100000101", -- t[22789] = 4
      "000100" when "0101100100000110", -- t[22790] = 4
      "000100" when "0101100100000111", -- t[22791] = 4
      "000100" when "0101100100001000", -- t[22792] = 4
      "000100" when "0101100100001001", -- t[22793] = 4
      "000100" when "0101100100001010", -- t[22794] = 4
      "000100" when "0101100100001011", -- t[22795] = 4
      "000100" when "0101100100001100", -- t[22796] = 4
      "000100" when "0101100100001101", -- t[22797] = 4
      "000100" when "0101100100001110", -- t[22798] = 4
      "000100" when "0101100100001111", -- t[22799] = 4
      "000100" when "0101100100010000", -- t[22800] = 4
      "000100" when "0101100100010001", -- t[22801] = 4
      "000100" when "0101100100010010", -- t[22802] = 4
      "000100" when "0101100100010011", -- t[22803] = 4
      "000100" when "0101100100010100", -- t[22804] = 4
      "000100" when "0101100100010101", -- t[22805] = 4
      "000100" when "0101100100010110", -- t[22806] = 4
      "000100" when "0101100100010111", -- t[22807] = 4
      "000100" when "0101100100011000", -- t[22808] = 4
      "000100" when "0101100100011001", -- t[22809] = 4
      "000100" when "0101100100011010", -- t[22810] = 4
      "000100" when "0101100100011011", -- t[22811] = 4
      "000100" when "0101100100011100", -- t[22812] = 4
      "000100" when "0101100100011101", -- t[22813] = 4
      "000100" when "0101100100011110", -- t[22814] = 4
      "000100" when "0101100100011111", -- t[22815] = 4
      "000100" when "0101100100100000", -- t[22816] = 4
      "000100" when "0101100100100001", -- t[22817] = 4
      "000100" when "0101100100100010", -- t[22818] = 4
      "000100" when "0101100100100011", -- t[22819] = 4
      "000100" when "0101100100100100", -- t[22820] = 4
      "000100" when "0101100100100101", -- t[22821] = 4
      "000100" when "0101100100100110", -- t[22822] = 4
      "000100" when "0101100100100111", -- t[22823] = 4
      "000100" when "0101100100101000", -- t[22824] = 4
      "000100" when "0101100100101001", -- t[22825] = 4
      "000100" when "0101100100101010", -- t[22826] = 4
      "000100" when "0101100100101011", -- t[22827] = 4
      "000100" when "0101100100101100", -- t[22828] = 4
      "000100" when "0101100100101101", -- t[22829] = 4
      "000100" when "0101100100101110", -- t[22830] = 4
      "000100" when "0101100100101111", -- t[22831] = 4
      "000100" when "0101100100110000", -- t[22832] = 4
      "000100" when "0101100100110001", -- t[22833] = 4
      "000100" when "0101100100110010", -- t[22834] = 4
      "000100" when "0101100100110011", -- t[22835] = 4
      "000100" when "0101100100110100", -- t[22836] = 4
      "000100" when "0101100100110101", -- t[22837] = 4
      "000100" when "0101100100110110", -- t[22838] = 4
      "000100" when "0101100100110111", -- t[22839] = 4
      "000100" when "0101100100111000", -- t[22840] = 4
      "000100" when "0101100100111001", -- t[22841] = 4
      "000100" when "0101100100111010", -- t[22842] = 4
      "000100" when "0101100100111011", -- t[22843] = 4
      "000100" when "0101100100111100", -- t[22844] = 4
      "000100" when "0101100100111101", -- t[22845] = 4
      "000100" when "0101100100111110", -- t[22846] = 4
      "000100" when "0101100100111111", -- t[22847] = 4
      "000100" when "0101100101000000", -- t[22848] = 4
      "000100" when "0101100101000001", -- t[22849] = 4
      "000100" when "0101100101000010", -- t[22850] = 4
      "000100" when "0101100101000011", -- t[22851] = 4
      "000100" when "0101100101000100", -- t[22852] = 4
      "000100" when "0101100101000101", -- t[22853] = 4
      "000100" when "0101100101000110", -- t[22854] = 4
      "000100" when "0101100101000111", -- t[22855] = 4
      "000100" when "0101100101001000", -- t[22856] = 4
      "000100" when "0101100101001001", -- t[22857] = 4
      "000100" when "0101100101001010", -- t[22858] = 4
      "000100" when "0101100101001011", -- t[22859] = 4
      "000100" when "0101100101001100", -- t[22860] = 4
      "000100" when "0101100101001101", -- t[22861] = 4
      "000100" when "0101100101001110", -- t[22862] = 4
      "000100" when "0101100101001111", -- t[22863] = 4
      "000100" when "0101100101010000", -- t[22864] = 4
      "000100" when "0101100101010001", -- t[22865] = 4
      "000100" when "0101100101010010", -- t[22866] = 4
      "000100" when "0101100101010011", -- t[22867] = 4
      "000100" when "0101100101010100", -- t[22868] = 4
      "000100" when "0101100101010101", -- t[22869] = 4
      "000100" when "0101100101010110", -- t[22870] = 4
      "000100" when "0101100101010111", -- t[22871] = 4
      "000100" when "0101100101011000", -- t[22872] = 4
      "000100" when "0101100101011001", -- t[22873] = 4
      "000100" when "0101100101011010", -- t[22874] = 4
      "000100" when "0101100101011011", -- t[22875] = 4
      "000100" when "0101100101011100", -- t[22876] = 4
      "000100" when "0101100101011101", -- t[22877] = 4
      "000100" when "0101100101011110", -- t[22878] = 4
      "000100" when "0101100101011111", -- t[22879] = 4
      "000100" when "0101100101100000", -- t[22880] = 4
      "000100" when "0101100101100001", -- t[22881] = 4
      "000100" when "0101100101100010", -- t[22882] = 4
      "000100" when "0101100101100011", -- t[22883] = 4
      "000100" when "0101100101100100", -- t[22884] = 4
      "000100" when "0101100101100101", -- t[22885] = 4
      "000100" when "0101100101100110", -- t[22886] = 4
      "000100" when "0101100101100111", -- t[22887] = 4
      "000100" when "0101100101101000", -- t[22888] = 4
      "000100" when "0101100101101001", -- t[22889] = 4
      "000100" when "0101100101101010", -- t[22890] = 4
      "000100" when "0101100101101011", -- t[22891] = 4
      "000100" when "0101100101101100", -- t[22892] = 4
      "000100" when "0101100101101101", -- t[22893] = 4
      "000100" when "0101100101101110", -- t[22894] = 4
      "000100" when "0101100101101111", -- t[22895] = 4
      "000100" when "0101100101110000", -- t[22896] = 4
      "000100" when "0101100101110001", -- t[22897] = 4
      "000100" when "0101100101110010", -- t[22898] = 4
      "000100" when "0101100101110011", -- t[22899] = 4
      "000100" when "0101100101110100", -- t[22900] = 4
      "000100" when "0101100101110101", -- t[22901] = 4
      "000100" when "0101100101110110", -- t[22902] = 4
      "000100" when "0101100101110111", -- t[22903] = 4
      "000100" when "0101100101111000", -- t[22904] = 4
      "000100" when "0101100101111001", -- t[22905] = 4
      "000100" when "0101100101111010", -- t[22906] = 4
      "000100" when "0101100101111011", -- t[22907] = 4
      "000100" when "0101100101111100", -- t[22908] = 4
      "000100" when "0101100101111101", -- t[22909] = 4
      "000100" when "0101100101111110", -- t[22910] = 4
      "000100" when "0101100101111111", -- t[22911] = 4
      "000100" when "0101100110000000", -- t[22912] = 4
      "000100" when "0101100110000001", -- t[22913] = 4
      "000100" when "0101100110000010", -- t[22914] = 4
      "000100" when "0101100110000011", -- t[22915] = 4
      "000100" when "0101100110000100", -- t[22916] = 4
      "000100" when "0101100110000101", -- t[22917] = 4
      "000100" when "0101100110000110", -- t[22918] = 4
      "000100" when "0101100110000111", -- t[22919] = 4
      "000100" when "0101100110001000", -- t[22920] = 4
      "000100" when "0101100110001001", -- t[22921] = 4
      "000100" when "0101100110001010", -- t[22922] = 4
      "000100" when "0101100110001011", -- t[22923] = 4
      "000100" when "0101100110001100", -- t[22924] = 4
      "000100" when "0101100110001101", -- t[22925] = 4
      "000100" when "0101100110001110", -- t[22926] = 4
      "000100" when "0101100110001111", -- t[22927] = 4
      "000100" when "0101100110010000", -- t[22928] = 4
      "000100" when "0101100110010001", -- t[22929] = 4
      "000100" when "0101100110010010", -- t[22930] = 4
      "000100" when "0101100110010011", -- t[22931] = 4
      "000100" when "0101100110010100", -- t[22932] = 4
      "000100" when "0101100110010101", -- t[22933] = 4
      "000100" when "0101100110010110", -- t[22934] = 4
      "000100" when "0101100110010111", -- t[22935] = 4
      "000100" when "0101100110011000", -- t[22936] = 4
      "000100" when "0101100110011001", -- t[22937] = 4
      "000100" when "0101100110011010", -- t[22938] = 4
      "000100" when "0101100110011011", -- t[22939] = 4
      "000100" when "0101100110011100", -- t[22940] = 4
      "000100" when "0101100110011101", -- t[22941] = 4
      "000100" when "0101100110011110", -- t[22942] = 4
      "000100" when "0101100110011111", -- t[22943] = 4
      "000100" when "0101100110100000", -- t[22944] = 4
      "000100" when "0101100110100001", -- t[22945] = 4
      "000100" when "0101100110100010", -- t[22946] = 4
      "000100" when "0101100110100011", -- t[22947] = 4
      "000100" when "0101100110100100", -- t[22948] = 4
      "000100" when "0101100110100101", -- t[22949] = 4
      "000100" when "0101100110100110", -- t[22950] = 4
      "000100" when "0101100110100111", -- t[22951] = 4
      "000100" when "0101100110101000", -- t[22952] = 4
      "000100" when "0101100110101001", -- t[22953] = 4
      "000100" when "0101100110101010", -- t[22954] = 4
      "000100" when "0101100110101011", -- t[22955] = 4
      "000100" when "0101100110101100", -- t[22956] = 4
      "000100" when "0101100110101101", -- t[22957] = 4
      "000100" when "0101100110101110", -- t[22958] = 4
      "000100" when "0101100110101111", -- t[22959] = 4
      "000100" when "0101100110110000", -- t[22960] = 4
      "000100" when "0101100110110001", -- t[22961] = 4
      "000100" when "0101100110110010", -- t[22962] = 4
      "000100" when "0101100110110011", -- t[22963] = 4
      "000100" when "0101100110110100", -- t[22964] = 4
      "000100" when "0101100110110101", -- t[22965] = 4
      "000100" when "0101100110110110", -- t[22966] = 4
      "000100" when "0101100110110111", -- t[22967] = 4
      "000100" when "0101100110111000", -- t[22968] = 4
      "000100" when "0101100110111001", -- t[22969] = 4
      "000100" when "0101100110111010", -- t[22970] = 4
      "000100" when "0101100110111011", -- t[22971] = 4
      "000100" when "0101100110111100", -- t[22972] = 4
      "000100" when "0101100110111101", -- t[22973] = 4
      "000100" when "0101100110111110", -- t[22974] = 4
      "000100" when "0101100110111111", -- t[22975] = 4
      "000100" when "0101100111000000", -- t[22976] = 4
      "000100" when "0101100111000001", -- t[22977] = 4
      "000100" when "0101100111000010", -- t[22978] = 4
      "000100" when "0101100111000011", -- t[22979] = 4
      "000100" when "0101100111000100", -- t[22980] = 4
      "000100" when "0101100111000101", -- t[22981] = 4
      "000100" when "0101100111000110", -- t[22982] = 4
      "000100" when "0101100111000111", -- t[22983] = 4
      "000100" when "0101100111001000", -- t[22984] = 4
      "000100" when "0101100111001001", -- t[22985] = 4
      "000100" when "0101100111001010", -- t[22986] = 4
      "000100" when "0101100111001011", -- t[22987] = 4
      "000100" when "0101100111001100", -- t[22988] = 4
      "000100" when "0101100111001101", -- t[22989] = 4
      "000100" when "0101100111001110", -- t[22990] = 4
      "000100" when "0101100111001111", -- t[22991] = 4
      "000100" when "0101100111010000", -- t[22992] = 4
      "000100" when "0101100111010001", -- t[22993] = 4
      "000100" when "0101100111010010", -- t[22994] = 4
      "000100" when "0101100111010011", -- t[22995] = 4
      "000100" when "0101100111010100", -- t[22996] = 4
      "000100" when "0101100111010101", -- t[22997] = 4
      "000100" when "0101100111010110", -- t[22998] = 4
      "000100" when "0101100111010111", -- t[22999] = 4
      "000100" when "0101100111011000", -- t[23000] = 4
      "000100" when "0101100111011001", -- t[23001] = 4
      "000100" when "0101100111011010", -- t[23002] = 4
      "000100" when "0101100111011011", -- t[23003] = 4
      "000100" when "0101100111011100", -- t[23004] = 4
      "000100" when "0101100111011101", -- t[23005] = 4
      "000100" when "0101100111011110", -- t[23006] = 4
      "000100" when "0101100111011111", -- t[23007] = 4
      "000100" when "0101100111100000", -- t[23008] = 4
      "000100" when "0101100111100001", -- t[23009] = 4
      "000100" when "0101100111100010", -- t[23010] = 4
      "000100" when "0101100111100011", -- t[23011] = 4
      "000100" when "0101100111100100", -- t[23012] = 4
      "000100" when "0101100111100101", -- t[23013] = 4
      "000100" when "0101100111100110", -- t[23014] = 4
      "000100" when "0101100111100111", -- t[23015] = 4
      "000100" when "0101100111101000", -- t[23016] = 4
      "000100" when "0101100111101001", -- t[23017] = 4
      "000100" when "0101100111101010", -- t[23018] = 4
      "000100" when "0101100111101011", -- t[23019] = 4
      "000100" when "0101100111101100", -- t[23020] = 4
      "000100" when "0101100111101101", -- t[23021] = 4
      "000100" when "0101100111101110", -- t[23022] = 4
      "000100" when "0101100111101111", -- t[23023] = 4
      "000100" when "0101100111110000", -- t[23024] = 4
      "000100" when "0101100111110001", -- t[23025] = 4
      "000100" when "0101100111110010", -- t[23026] = 4
      "000100" when "0101100111110011", -- t[23027] = 4
      "000100" when "0101100111110100", -- t[23028] = 4
      "000100" when "0101100111110101", -- t[23029] = 4
      "000100" when "0101100111110110", -- t[23030] = 4
      "000100" when "0101100111110111", -- t[23031] = 4
      "000100" when "0101100111111000", -- t[23032] = 4
      "000100" when "0101100111111001", -- t[23033] = 4
      "000100" when "0101100111111010", -- t[23034] = 4
      "000100" when "0101100111111011", -- t[23035] = 4
      "000100" when "0101100111111100", -- t[23036] = 4
      "000100" when "0101100111111101", -- t[23037] = 4
      "000100" when "0101100111111110", -- t[23038] = 4
      "000100" when "0101100111111111", -- t[23039] = 4
      "000100" when "0101101000000000", -- t[23040] = 4
      "000100" when "0101101000000001", -- t[23041] = 4
      "000100" when "0101101000000010", -- t[23042] = 4
      "000100" when "0101101000000011", -- t[23043] = 4
      "000100" when "0101101000000100", -- t[23044] = 4
      "000100" when "0101101000000101", -- t[23045] = 4
      "000100" when "0101101000000110", -- t[23046] = 4
      "000100" when "0101101000000111", -- t[23047] = 4
      "000100" when "0101101000001000", -- t[23048] = 4
      "000100" when "0101101000001001", -- t[23049] = 4
      "000100" when "0101101000001010", -- t[23050] = 4
      "000100" when "0101101000001011", -- t[23051] = 4
      "000100" when "0101101000001100", -- t[23052] = 4
      "000100" when "0101101000001101", -- t[23053] = 4
      "000100" when "0101101000001110", -- t[23054] = 4
      "000100" when "0101101000001111", -- t[23055] = 4
      "000100" when "0101101000010000", -- t[23056] = 4
      "000100" when "0101101000010001", -- t[23057] = 4
      "000100" when "0101101000010010", -- t[23058] = 4
      "000100" when "0101101000010011", -- t[23059] = 4
      "000100" when "0101101000010100", -- t[23060] = 4
      "000100" when "0101101000010101", -- t[23061] = 4
      "000100" when "0101101000010110", -- t[23062] = 4
      "000100" when "0101101000010111", -- t[23063] = 4
      "000100" when "0101101000011000", -- t[23064] = 4
      "000100" when "0101101000011001", -- t[23065] = 4
      "000100" when "0101101000011010", -- t[23066] = 4
      "000100" when "0101101000011011", -- t[23067] = 4
      "000100" when "0101101000011100", -- t[23068] = 4
      "000100" when "0101101000011101", -- t[23069] = 4
      "000100" when "0101101000011110", -- t[23070] = 4
      "000100" when "0101101000011111", -- t[23071] = 4
      "000100" when "0101101000100000", -- t[23072] = 4
      "000100" when "0101101000100001", -- t[23073] = 4
      "000100" when "0101101000100010", -- t[23074] = 4
      "000100" when "0101101000100011", -- t[23075] = 4
      "000100" when "0101101000100100", -- t[23076] = 4
      "000100" when "0101101000100101", -- t[23077] = 4
      "000100" when "0101101000100110", -- t[23078] = 4
      "000100" when "0101101000100111", -- t[23079] = 4
      "000100" when "0101101000101000", -- t[23080] = 4
      "000100" when "0101101000101001", -- t[23081] = 4
      "000100" when "0101101000101010", -- t[23082] = 4
      "000100" when "0101101000101011", -- t[23083] = 4
      "000100" when "0101101000101100", -- t[23084] = 4
      "000100" when "0101101000101101", -- t[23085] = 4
      "000100" when "0101101000101110", -- t[23086] = 4
      "000100" when "0101101000101111", -- t[23087] = 4
      "000100" when "0101101000110000", -- t[23088] = 4
      "000100" when "0101101000110001", -- t[23089] = 4
      "000100" when "0101101000110010", -- t[23090] = 4
      "000100" when "0101101000110011", -- t[23091] = 4
      "000100" when "0101101000110100", -- t[23092] = 4
      "000100" when "0101101000110101", -- t[23093] = 4
      "000100" when "0101101000110110", -- t[23094] = 4
      "000100" when "0101101000110111", -- t[23095] = 4
      "000100" when "0101101000111000", -- t[23096] = 4
      "000100" when "0101101000111001", -- t[23097] = 4
      "000100" when "0101101000111010", -- t[23098] = 4
      "000100" when "0101101000111011", -- t[23099] = 4
      "000100" when "0101101000111100", -- t[23100] = 4
      "000100" when "0101101000111101", -- t[23101] = 4
      "000100" when "0101101000111110", -- t[23102] = 4
      "000100" when "0101101000111111", -- t[23103] = 4
      "000101" when "0101101001000000", -- t[23104] = 5
      "000101" when "0101101001000001", -- t[23105] = 5
      "000101" when "0101101001000010", -- t[23106] = 5
      "000101" when "0101101001000011", -- t[23107] = 5
      "000101" when "0101101001000100", -- t[23108] = 5
      "000101" when "0101101001000101", -- t[23109] = 5
      "000101" when "0101101001000110", -- t[23110] = 5
      "000101" when "0101101001000111", -- t[23111] = 5
      "000101" when "0101101001001000", -- t[23112] = 5
      "000101" when "0101101001001001", -- t[23113] = 5
      "000101" when "0101101001001010", -- t[23114] = 5
      "000101" when "0101101001001011", -- t[23115] = 5
      "000101" when "0101101001001100", -- t[23116] = 5
      "000101" when "0101101001001101", -- t[23117] = 5
      "000101" when "0101101001001110", -- t[23118] = 5
      "000101" when "0101101001001111", -- t[23119] = 5
      "000101" when "0101101001010000", -- t[23120] = 5
      "000101" when "0101101001010001", -- t[23121] = 5
      "000101" when "0101101001010010", -- t[23122] = 5
      "000101" when "0101101001010011", -- t[23123] = 5
      "000101" when "0101101001010100", -- t[23124] = 5
      "000101" when "0101101001010101", -- t[23125] = 5
      "000101" when "0101101001010110", -- t[23126] = 5
      "000101" when "0101101001010111", -- t[23127] = 5
      "000101" when "0101101001011000", -- t[23128] = 5
      "000101" when "0101101001011001", -- t[23129] = 5
      "000101" when "0101101001011010", -- t[23130] = 5
      "000101" when "0101101001011011", -- t[23131] = 5
      "000101" when "0101101001011100", -- t[23132] = 5
      "000101" when "0101101001011101", -- t[23133] = 5
      "000101" when "0101101001011110", -- t[23134] = 5
      "000101" when "0101101001011111", -- t[23135] = 5
      "000101" when "0101101001100000", -- t[23136] = 5
      "000101" when "0101101001100001", -- t[23137] = 5
      "000101" when "0101101001100010", -- t[23138] = 5
      "000101" when "0101101001100011", -- t[23139] = 5
      "000101" when "0101101001100100", -- t[23140] = 5
      "000101" when "0101101001100101", -- t[23141] = 5
      "000101" when "0101101001100110", -- t[23142] = 5
      "000101" when "0101101001100111", -- t[23143] = 5
      "000101" when "0101101001101000", -- t[23144] = 5
      "000101" when "0101101001101001", -- t[23145] = 5
      "000101" when "0101101001101010", -- t[23146] = 5
      "000101" when "0101101001101011", -- t[23147] = 5
      "000101" when "0101101001101100", -- t[23148] = 5
      "000101" when "0101101001101101", -- t[23149] = 5
      "000101" when "0101101001101110", -- t[23150] = 5
      "000101" when "0101101001101111", -- t[23151] = 5
      "000101" when "0101101001110000", -- t[23152] = 5
      "000101" when "0101101001110001", -- t[23153] = 5
      "000101" when "0101101001110010", -- t[23154] = 5
      "000101" when "0101101001110011", -- t[23155] = 5
      "000101" when "0101101001110100", -- t[23156] = 5
      "000101" when "0101101001110101", -- t[23157] = 5
      "000101" when "0101101001110110", -- t[23158] = 5
      "000101" when "0101101001110111", -- t[23159] = 5
      "000101" when "0101101001111000", -- t[23160] = 5
      "000101" when "0101101001111001", -- t[23161] = 5
      "000101" when "0101101001111010", -- t[23162] = 5
      "000101" when "0101101001111011", -- t[23163] = 5
      "000101" when "0101101001111100", -- t[23164] = 5
      "000101" when "0101101001111101", -- t[23165] = 5
      "000101" when "0101101001111110", -- t[23166] = 5
      "000101" when "0101101001111111", -- t[23167] = 5
      "000101" when "0101101010000000", -- t[23168] = 5
      "000101" when "0101101010000001", -- t[23169] = 5
      "000101" when "0101101010000010", -- t[23170] = 5
      "000101" when "0101101010000011", -- t[23171] = 5
      "000101" when "0101101010000100", -- t[23172] = 5
      "000101" when "0101101010000101", -- t[23173] = 5
      "000101" when "0101101010000110", -- t[23174] = 5
      "000101" when "0101101010000111", -- t[23175] = 5
      "000101" when "0101101010001000", -- t[23176] = 5
      "000101" when "0101101010001001", -- t[23177] = 5
      "000101" when "0101101010001010", -- t[23178] = 5
      "000101" when "0101101010001011", -- t[23179] = 5
      "000101" when "0101101010001100", -- t[23180] = 5
      "000101" when "0101101010001101", -- t[23181] = 5
      "000101" when "0101101010001110", -- t[23182] = 5
      "000101" when "0101101010001111", -- t[23183] = 5
      "000101" when "0101101010010000", -- t[23184] = 5
      "000101" when "0101101010010001", -- t[23185] = 5
      "000101" when "0101101010010010", -- t[23186] = 5
      "000101" when "0101101010010011", -- t[23187] = 5
      "000101" when "0101101010010100", -- t[23188] = 5
      "000101" when "0101101010010101", -- t[23189] = 5
      "000101" when "0101101010010110", -- t[23190] = 5
      "000101" when "0101101010010111", -- t[23191] = 5
      "000101" when "0101101010011000", -- t[23192] = 5
      "000101" when "0101101010011001", -- t[23193] = 5
      "000101" when "0101101010011010", -- t[23194] = 5
      "000101" when "0101101010011011", -- t[23195] = 5
      "000101" when "0101101010011100", -- t[23196] = 5
      "000101" when "0101101010011101", -- t[23197] = 5
      "000101" when "0101101010011110", -- t[23198] = 5
      "000101" when "0101101010011111", -- t[23199] = 5
      "000101" when "0101101010100000", -- t[23200] = 5
      "000101" when "0101101010100001", -- t[23201] = 5
      "000101" when "0101101010100010", -- t[23202] = 5
      "000101" when "0101101010100011", -- t[23203] = 5
      "000101" when "0101101010100100", -- t[23204] = 5
      "000101" when "0101101010100101", -- t[23205] = 5
      "000101" when "0101101010100110", -- t[23206] = 5
      "000101" when "0101101010100111", -- t[23207] = 5
      "000101" when "0101101010101000", -- t[23208] = 5
      "000101" when "0101101010101001", -- t[23209] = 5
      "000101" when "0101101010101010", -- t[23210] = 5
      "000101" when "0101101010101011", -- t[23211] = 5
      "000101" when "0101101010101100", -- t[23212] = 5
      "000101" when "0101101010101101", -- t[23213] = 5
      "000101" when "0101101010101110", -- t[23214] = 5
      "000101" when "0101101010101111", -- t[23215] = 5
      "000101" when "0101101010110000", -- t[23216] = 5
      "000101" when "0101101010110001", -- t[23217] = 5
      "000101" when "0101101010110010", -- t[23218] = 5
      "000101" when "0101101010110011", -- t[23219] = 5
      "000101" when "0101101010110100", -- t[23220] = 5
      "000101" when "0101101010110101", -- t[23221] = 5
      "000101" when "0101101010110110", -- t[23222] = 5
      "000101" when "0101101010110111", -- t[23223] = 5
      "000101" when "0101101010111000", -- t[23224] = 5
      "000101" when "0101101010111001", -- t[23225] = 5
      "000101" when "0101101010111010", -- t[23226] = 5
      "000101" when "0101101010111011", -- t[23227] = 5
      "000101" when "0101101010111100", -- t[23228] = 5
      "000101" when "0101101010111101", -- t[23229] = 5
      "000101" when "0101101010111110", -- t[23230] = 5
      "000101" when "0101101010111111", -- t[23231] = 5
      "000101" when "0101101011000000", -- t[23232] = 5
      "000101" when "0101101011000001", -- t[23233] = 5
      "000101" when "0101101011000010", -- t[23234] = 5
      "000101" when "0101101011000011", -- t[23235] = 5
      "000101" when "0101101011000100", -- t[23236] = 5
      "000101" when "0101101011000101", -- t[23237] = 5
      "000101" when "0101101011000110", -- t[23238] = 5
      "000101" when "0101101011000111", -- t[23239] = 5
      "000101" when "0101101011001000", -- t[23240] = 5
      "000101" when "0101101011001001", -- t[23241] = 5
      "000101" when "0101101011001010", -- t[23242] = 5
      "000101" when "0101101011001011", -- t[23243] = 5
      "000101" when "0101101011001100", -- t[23244] = 5
      "000101" when "0101101011001101", -- t[23245] = 5
      "000101" when "0101101011001110", -- t[23246] = 5
      "000101" when "0101101011001111", -- t[23247] = 5
      "000101" when "0101101011010000", -- t[23248] = 5
      "000101" when "0101101011010001", -- t[23249] = 5
      "000101" when "0101101011010010", -- t[23250] = 5
      "000101" when "0101101011010011", -- t[23251] = 5
      "000101" when "0101101011010100", -- t[23252] = 5
      "000101" when "0101101011010101", -- t[23253] = 5
      "000101" when "0101101011010110", -- t[23254] = 5
      "000101" when "0101101011010111", -- t[23255] = 5
      "000101" when "0101101011011000", -- t[23256] = 5
      "000101" when "0101101011011001", -- t[23257] = 5
      "000101" when "0101101011011010", -- t[23258] = 5
      "000101" when "0101101011011011", -- t[23259] = 5
      "000101" when "0101101011011100", -- t[23260] = 5
      "000101" when "0101101011011101", -- t[23261] = 5
      "000101" when "0101101011011110", -- t[23262] = 5
      "000101" when "0101101011011111", -- t[23263] = 5
      "000101" when "0101101011100000", -- t[23264] = 5
      "000101" when "0101101011100001", -- t[23265] = 5
      "000101" when "0101101011100010", -- t[23266] = 5
      "000101" when "0101101011100011", -- t[23267] = 5
      "000101" when "0101101011100100", -- t[23268] = 5
      "000101" when "0101101011100101", -- t[23269] = 5
      "000101" when "0101101011100110", -- t[23270] = 5
      "000101" when "0101101011100111", -- t[23271] = 5
      "000101" when "0101101011101000", -- t[23272] = 5
      "000101" when "0101101011101001", -- t[23273] = 5
      "000101" when "0101101011101010", -- t[23274] = 5
      "000101" when "0101101011101011", -- t[23275] = 5
      "000101" when "0101101011101100", -- t[23276] = 5
      "000101" when "0101101011101101", -- t[23277] = 5
      "000101" when "0101101011101110", -- t[23278] = 5
      "000101" when "0101101011101111", -- t[23279] = 5
      "000101" when "0101101011110000", -- t[23280] = 5
      "000101" when "0101101011110001", -- t[23281] = 5
      "000101" when "0101101011110010", -- t[23282] = 5
      "000101" when "0101101011110011", -- t[23283] = 5
      "000101" when "0101101011110100", -- t[23284] = 5
      "000101" when "0101101011110101", -- t[23285] = 5
      "000101" when "0101101011110110", -- t[23286] = 5
      "000101" when "0101101011110111", -- t[23287] = 5
      "000101" when "0101101011111000", -- t[23288] = 5
      "000101" when "0101101011111001", -- t[23289] = 5
      "000101" when "0101101011111010", -- t[23290] = 5
      "000101" when "0101101011111011", -- t[23291] = 5
      "000101" when "0101101011111100", -- t[23292] = 5
      "000101" when "0101101011111101", -- t[23293] = 5
      "000101" when "0101101011111110", -- t[23294] = 5
      "000101" when "0101101011111111", -- t[23295] = 5
      "000101" when "0101101100000000", -- t[23296] = 5
      "000101" when "0101101100000001", -- t[23297] = 5
      "000101" when "0101101100000010", -- t[23298] = 5
      "000101" when "0101101100000011", -- t[23299] = 5
      "000101" when "0101101100000100", -- t[23300] = 5
      "000101" when "0101101100000101", -- t[23301] = 5
      "000101" when "0101101100000110", -- t[23302] = 5
      "000101" when "0101101100000111", -- t[23303] = 5
      "000101" when "0101101100001000", -- t[23304] = 5
      "000101" when "0101101100001001", -- t[23305] = 5
      "000101" when "0101101100001010", -- t[23306] = 5
      "000101" when "0101101100001011", -- t[23307] = 5
      "000101" when "0101101100001100", -- t[23308] = 5
      "000101" when "0101101100001101", -- t[23309] = 5
      "000101" when "0101101100001110", -- t[23310] = 5
      "000101" when "0101101100001111", -- t[23311] = 5
      "000101" when "0101101100010000", -- t[23312] = 5
      "000101" when "0101101100010001", -- t[23313] = 5
      "000101" when "0101101100010010", -- t[23314] = 5
      "000101" when "0101101100010011", -- t[23315] = 5
      "000101" when "0101101100010100", -- t[23316] = 5
      "000101" when "0101101100010101", -- t[23317] = 5
      "000101" when "0101101100010110", -- t[23318] = 5
      "000101" when "0101101100010111", -- t[23319] = 5
      "000101" when "0101101100011000", -- t[23320] = 5
      "000101" when "0101101100011001", -- t[23321] = 5
      "000101" when "0101101100011010", -- t[23322] = 5
      "000101" when "0101101100011011", -- t[23323] = 5
      "000101" when "0101101100011100", -- t[23324] = 5
      "000101" when "0101101100011101", -- t[23325] = 5
      "000101" when "0101101100011110", -- t[23326] = 5
      "000101" when "0101101100011111", -- t[23327] = 5
      "000101" when "0101101100100000", -- t[23328] = 5
      "000101" when "0101101100100001", -- t[23329] = 5
      "000101" when "0101101100100010", -- t[23330] = 5
      "000101" when "0101101100100011", -- t[23331] = 5
      "000101" when "0101101100100100", -- t[23332] = 5
      "000101" when "0101101100100101", -- t[23333] = 5
      "000101" when "0101101100100110", -- t[23334] = 5
      "000101" when "0101101100100111", -- t[23335] = 5
      "000101" when "0101101100101000", -- t[23336] = 5
      "000101" when "0101101100101001", -- t[23337] = 5
      "000101" when "0101101100101010", -- t[23338] = 5
      "000101" when "0101101100101011", -- t[23339] = 5
      "000101" when "0101101100101100", -- t[23340] = 5
      "000101" when "0101101100101101", -- t[23341] = 5
      "000101" when "0101101100101110", -- t[23342] = 5
      "000101" when "0101101100101111", -- t[23343] = 5
      "000101" when "0101101100110000", -- t[23344] = 5
      "000101" when "0101101100110001", -- t[23345] = 5
      "000101" when "0101101100110010", -- t[23346] = 5
      "000101" when "0101101100110011", -- t[23347] = 5
      "000101" when "0101101100110100", -- t[23348] = 5
      "000101" when "0101101100110101", -- t[23349] = 5
      "000101" when "0101101100110110", -- t[23350] = 5
      "000101" when "0101101100110111", -- t[23351] = 5
      "000101" when "0101101100111000", -- t[23352] = 5
      "000101" when "0101101100111001", -- t[23353] = 5
      "000101" when "0101101100111010", -- t[23354] = 5
      "000101" when "0101101100111011", -- t[23355] = 5
      "000101" when "0101101100111100", -- t[23356] = 5
      "000101" when "0101101100111101", -- t[23357] = 5
      "000101" when "0101101100111110", -- t[23358] = 5
      "000101" when "0101101100111111", -- t[23359] = 5
      "000101" when "0101101101000000", -- t[23360] = 5
      "000101" when "0101101101000001", -- t[23361] = 5
      "000101" when "0101101101000010", -- t[23362] = 5
      "000101" when "0101101101000011", -- t[23363] = 5
      "000101" when "0101101101000100", -- t[23364] = 5
      "000101" when "0101101101000101", -- t[23365] = 5
      "000101" when "0101101101000110", -- t[23366] = 5
      "000101" when "0101101101000111", -- t[23367] = 5
      "000101" when "0101101101001000", -- t[23368] = 5
      "000101" when "0101101101001001", -- t[23369] = 5
      "000101" when "0101101101001010", -- t[23370] = 5
      "000101" when "0101101101001011", -- t[23371] = 5
      "000101" when "0101101101001100", -- t[23372] = 5
      "000101" when "0101101101001101", -- t[23373] = 5
      "000101" when "0101101101001110", -- t[23374] = 5
      "000101" when "0101101101001111", -- t[23375] = 5
      "000101" when "0101101101010000", -- t[23376] = 5
      "000101" when "0101101101010001", -- t[23377] = 5
      "000101" when "0101101101010010", -- t[23378] = 5
      "000101" when "0101101101010011", -- t[23379] = 5
      "000101" when "0101101101010100", -- t[23380] = 5
      "000101" when "0101101101010101", -- t[23381] = 5
      "000101" when "0101101101010110", -- t[23382] = 5
      "000101" when "0101101101010111", -- t[23383] = 5
      "000101" when "0101101101011000", -- t[23384] = 5
      "000101" when "0101101101011001", -- t[23385] = 5
      "000101" when "0101101101011010", -- t[23386] = 5
      "000101" when "0101101101011011", -- t[23387] = 5
      "000101" when "0101101101011100", -- t[23388] = 5
      "000101" when "0101101101011101", -- t[23389] = 5
      "000101" when "0101101101011110", -- t[23390] = 5
      "000101" when "0101101101011111", -- t[23391] = 5
      "000101" when "0101101101100000", -- t[23392] = 5
      "000101" when "0101101101100001", -- t[23393] = 5
      "000101" when "0101101101100010", -- t[23394] = 5
      "000101" when "0101101101100011", -- t[23395] = 5
      "000101" when "0101101101100100", -- t[23396] = 5
      "000101" when "0101101101100101", -- t[23397] = 5
      "000101" when "0101101101100110", -- t[23398] = 5
      "000101" when "0101101101100111", -- t[23399] = 5
      "000101" when "0101101101101000", -- t[23400] = 5
      "000101" when "0101101101101001", -- t[23401] = 5
      "000101" when "0101101101101010", -- t[23402] = 5
      "000101" when "0101101101101011", -- t[23403] = 5
      "000101" when "0101101101101100", -- t[23404] = 5
      "000101" when "0101101101101101", -- t[23405] = 5
      "000101" when "0101101101101110", -- t[23406] = 5
      "000101" when "0101101101101111", -- t[23407] = 5
      "000101" when "0101101101110000", -- t[23408] = 5
      "000101" when "0101101101110001", -- t[23409] = 5
      "000101" when "0101101101110010", -- t[23410] = 5
      "000101" when "0101101101110011", -- t[23411] = 5
      "000101" when "0101101101110100", -- t[23412] = 5
      "000101" when "0101101101110101", -- t[23413] = 5
      "000101" when "0101101101110110", -- t[23414] = 5
      "000101" when "0101101101110111", -- t[23415] = 5
      "000101" when "0101101101111000", -- t[23416] = 5
      "000101" when "0101101101111001", -- t[23417] = 5
      "000101" when "0101101101111010", -- t[23418] = 5
      "000101" when "0101101101111011", -- t[23419] = 5
      "000101" when "0101101101111100", -- t[23420] = 5
      "000101" when "0101101101111101", -- t[23421] = 5
      "000101" when "0101101101111110", -- t[23422] = 5
      "000101" when "0101101101111111", -- t[23423] = 5
      "000101" when "0101101110000000", -- t[23424] = 5
      "000101" when "0101101110000001", -- t[23425] = 5
      "000101" when "0101101110000010", -- t[23426] = 5
      "000101" when "0101101110000011", -- t[23427] = 5
      "000101" when "0101101110000100", -- t[23428] = 5
      "000101" when "0101101110000101", -- t[23429] = 5
      "000101" when "0101101110000110", -- t[23430] = 5
      "000101" when "0101101110000111", -- t[23431] = 5
      "000101" when "0101101110001000", -- t[23432] = 5
      "000101" when "0101101110001001", -- t[23433] = 5
      "000101" when "0101101110001010", -- t[23434] = 5
      "000101" when "0101101110001011", -- t[23435] = 5
      "000101" when "0101101110001100", -- t[23436] = 5
      "000101" when "0101101110001101", -- t[23437] = 5
      "000101" when "0101101110001110", -- t[23438] = 5
      "000101" when "0101101110001111", -- t[23439] = 5
      "000101" when "0101101110010000", -- t[23440] = 5
      "000101" when "0101101110010001", -- t[23441] = 5
      "000101" when "0101101110010010", -- t[23442] = 5
      "000101" when "0101101110010011", -- t[23443] = 5
      "000101" when "0101101110010100", -- t[23444] = 5
      "000101" when "0101101110010101", -- t[23445] = 5
      "000101" when "0101101110010110", -- t[23446] = 5
      "000101" when "0101101110010111", -- t[23447] = 5
      "000101" when "0101101110011000", -- t[23448] = 5
      "000101" when "0101101110011001", -- t[23449] = 5
      "000101" when "0101101110011010", -- t[23450] = 5
      "000101" when "0101101110011011", -- t[23451] = 5
      "000101" when "0101101110011100", -- t[23452] = 5
      "000101" when "0101101110011101", -- t[23453] = 5
      "000101" when "0101101110011110", -- t[23454] = 5
      "000101" when "0101101110011111", -- t[23455] = 5
      "000101" when "0101101110100000", -- t[23456] = 5
      "000101" when "0101101110100001", -- t[23457] = 5
      "000101" when "0101101110100010", -- t[23458] = 5
      "000101" when "0101101110100011", -- t[23459] = 5
      "000101" when "0101101110100100", -- t[23460] = 5
      "000101" when "0101101110100101", -- t[23461] = 5
      "000101" when "0101101110100110", -- t[23462] = 5
      "000101" when "0101101110100111", -- t[23463] = 5
      "000101" when "0101101110101000", -- t[23464] = 5
      "000101" when "0101101110101001", -- t[23465] = 5
      "000101" when "0101101110101010", -- t[23466] = 5
      "000101" when "0101101110101011", -- t[23467] = 5
      "000101" when "0101101110101100", -- t[23468] = 5
      "000101" when "0101101110101101", -- t[23469] = 5
      "000101" when "0101101110101110", -- t[23470] = 5
      "000101" when "0101101110101111", -- t[23471] = 5
      "000101" when "0101101110110000", -- t[23472] = 5
      "000101" when "0101101110110001", -- t[23473] = 5
      "000101" when "0101101110110010", -- t[23474] = 5
      "000101" when "0101101110110011", -- t[23475] = 5
      "000101" when "0101101110110100", -- t[23476] = 5
      "000101" when "0101101110110101", -- t[23477] = 5
      "000101" when "0101101110110110", -- t[23478] = 5
      "000101" when "0101101110110111", -- t[23479] = 5
      "000101" when "0101101110111000", -- t[23480] = 5
      "000101" when "0101101110111001", -- t[23481] = 5
      "000101" when "0101101110111010", -- t[23482] = 5
      "000101" when "0101101110111011", -- t[23483] = 5
      "000101" when "0101101110111100", -- t[23484] = 5
      "000101" when "0101101110111101", -- t[23485] = 5
      "000101" when "0101101110111110", -- t[23486] = 5
      "000101" when "0101101110111111", -- t[23487] = 5
      "000101" when "0101101111000000", -- t[23488] = 5
      "000101" when "0101101111000001", -- t[23489] = 5
      "000101" when "0101101111000010", -- t[23490] = 5
      "000101" when "0101101111000011", -- t[23491] = 5
      "000101" when "0101101111000100", -- t[23492] = 5
      "000101" when "0101101111000101", -- t[23493] = 5
      "000101" when "0101101111000110", -- t[23494] = 5
      "000101" when "0101101111000111", -- t[23495] = 5
      "000101" when "0101101111001000", -- t[23496] = 5
      "000101" when "0101101111001001", -- t[23497] = 5
      "000101" when "0101101111001010", -- t[23498] = 5
      "000101" when "0101101111001011", -- t[23499] = 5
      "000101" when "0101101111001100", -- t[23500] = 5
      "000101" when "0101101111001101", -- t[23501] = 5
      "000101" when "0101101111001110", -- t[23502] = 5
      "000101" when "0101101111001111", -- t[23503] = 5
      "000101" when "0101101111010000", -- t[23504] = 5
      "000101" when "0101101111010001", -- t[23505] = 5
      "000101" when "0101101111010010", -- t[23506] = 5
      "000101" when "0101101111010011", -- t[23507] = 5
      "000101" when "0101101111010100", -- t[23508] = 5
      "000101" when "0101101111010101", -- t[23509] = 5
      "000101" when "0101101111010110", -- t[23510] = 5
      "000101" when "0101101111010111", -- t[23511] = 5
      "000101" when "0101101111011000", -- t[23512] = 5
      "000101" when "0101101111011001", -- t[23513] = 5
      "000101" when "0101101111011010", -- t[23514] = 5
      "000101" when "0101101111011011", -- t[23515] = 5
      "000101" when "0101101111011100", -- t[23516] = 5
      "000101" when "0101101111011101", -- t[23517] = 5
      "000101" when "0101101111011110", -- t[23518] = 5
      "000101" when "0101101111011111", -- t[23519] = 5
      "000101" when "0101101111100000", -- t[23520] = 5
      "000101" when "0101101111100001", -- t[23521] = 5
      "000101" when "0101101111100010", -- t[23522] = 5
      "000101" when "0101101111100011", -- t[23523] = 5
      "000101" when "0101101111100100", -- t[23524] = 5
      "000101" when "0101101111100101", -- t[23525] = 5
      "000101" when "0101101111100110", -- t[23526] = 5
      "000101" when "0101101111100111", -- t[23527] = 5
      "000101" when "0101101111101000", -- t[23528] = 5
      "000101" when "0101101111101001", -- t[23529] = 5
      "000101" when "0101101111101010", -- t[23530] = 5
      "000101" when "0101101111101011", -- t[23531] = 5
      "000101" when "0101101111101100", -- t[23532] = 5
      "000101" when "0101101111101101", -- t[23533] = 5
      "000101" when "0101101111101110", -- t[23534] = 5
      "000101" when "0101101111101111", -- t[23535] = 5
      "000101" when "0101101111110000", -- t[23536] = 5
      "000101" when "0101101111110001", -- t[23537] = 5
      "000101" when "0101101111110010", -- t[23538] = 5
      "000101" when "0101101111110011", -- t[23539] = 5
      "000101" when "0101101111110100", -- t[23540] = 5
      "000101" when "0101101111110101", -- t[23541] = 5
      "000101" when "0101101111110110", -- t[23542] = 5
      "000101" when "0101101111110111", -- t[23543] = 5
      "000101" when "0101101111111000", -- t[23544] = 5
      "000101" when "0101101111111001", -- t[23545] = 5
      "000101" when "0101101111111010", -- t[23546] = 5
      "000101" when "0101101111111011", -- t[23547] = 5
      "000101" when "0101101111111100", -- t[23548] = 5
      "000101" when "0101101111111101", -- t[23549] = 5
      "000101" when "0101101111111110", -- t[23550] = 5
      "000101" when "0101101111111111", -- t[23551] = 5
      "000101" when "0101110000000000", -- t[23552] = 5
      "000101" when "0101110000000001", -- t[23553] = 5
      "000101" when "0101110000000010", -- t[23554] = 5
      "000101" when "0101110000000011", -- t[23555] = 5
      "000101" when "0101110000000100", -- t[23556] = 5
      "000101" when "0101110000000101", -- t[23557] = 5
      "000101" when "0101110000000110", -- t[23558] = 5
      "000101" when "0101110000000111", -- t[23559] = 5
      "000101" when "0101110000001000", -- t[23560] = 5
      "000101" when "0101110000001001", -- t[23561] = 5
      "000101" when "0101110000001010", -- t[23562] = 5
      "000101" when "0101110000001011", -- t[23563] = 5
      "000101" when "0101110000001100", -- t[23564] = 5
      "000101" when "0101110000001101", -- t[23565] = 5
      "000101" when "0101110000001110", -- t[23566] = 5
      "000101" when "0101110000001111", -- t[23567] = 5
      "000101" when "0101110000010000", -- t[23568] = 5
      "000101" when "0101110000010001", -- t[23569] = 5
      "000101" when "0101110000010010", -- t[23570] = 5
      "000101" when "0101110000010011", -- t[23571] = 5
      "000101" when "0101110000010100", -- t[23572] = 5
      "000101" when "0101110000010101", -- t[23573] = 5
      "000101" when "0101110000010110", -- t[23574] = 5
      "000101" when "0101110000010111", -- t[23575] = 5
      "000101" when "0101110000011000", -- t[23576] = 5
      "000101" when "0101110000011001", -- t[23577] = 5
      "000101" when "0101110000011010", -- t[23578] = 5
      "000101" when "0101110000011011", -- t[23579] = 5
      "000101" when "0101110000011100", -- t[23580] = 5
      "000101" when "0101110000011101", -- t[23581] = 5
      "000101" when "0101110000011110", -- t[23582] = 5
      "000101" when "0101110000011111", -- t[23583] = 5
      "000101" when "0101110000100000", -- t[23584] = 5
      "000101" when "0101110000100001", -- t[23585] = 5
      "000101" when "0101110000100010", -- t[23586] = 5
      "000101" when "0101110000100011", -- t[23587] = 5
      "000101" when "0101110000100100", -- t[23588] = 5
      "000101" when "0101110000100101", -- t[23589] = 5
      "000101" when "0101110000100110", -- t[23590] = 5
      "000101" when "0101110000100111", -- t[23591] = 5
      "000101" when "0101110000101000", -- t[23592] = 5
      "000101" when "0101110000101001", -- t[23593] = 5
      "000101" when "0101110000101010", -- t[23594] = 5
      "000101" when "0101110000101011", -- t[23595] = 5
      "000101" when "0101110000101100", -- t[23596] = 5
      "000101" when "0101110000101101", -- t[23597] = 5
      "000101" when "0101110000101110", -- t[23598] = 5
      "000101" when "0101110000101111", -- t[23599] = 5
      "000101" when "0101110000110000", -- t[23600] = 5
      "000101" when "0101110000110001", -- t[23601] = 5
      "000101" when "0101110000110010", -- t[23602] = 5
      "000101" when "0101110000110011", -- t[23603] = 5
      "000101" when "0101110000110100", -- t[23604] = 5
      "000101" when "0101110000110101", -- t[23605] = 5
      "000101" when "0101110000110110", -- t[23606] = 5
      "000101" when "0101110000110111", -- t[23607] = 5
      "000101" when "0101110000111000", -- t[23608] = 5
      "000101" when "0101110000111001", -- t[23609] = 5
      "000101" when "0101110000111010", -- t[23610] = 5
      "000101" when "0101110000111011", -- t[23611] = 5
      "000101" when "0101110000111100", -- t[23612] = 5
      "000101" when "0101110000111101", -- t[23613] = 5
      "000101" when "0101110000111110", -- t[23614] = 5
      "000101" when "0101110000111111", -- t[23615] = 5
      "000101" when "0101110001000000", -- t[23616] = 5
      "000101" when "0101110001000001", -- t[23617] = 5
      "000101" when "0101110001000010", -- t[23618] = 5
      "000101" when "0101110001000011", -- t[23619] = 5
      "000101" when "0101110001000100", -- t[23620] = 5
      "000101" when "0101110001000101", -- t[23621] = 5
      "000101" when "0101110001000110", -- t[23622] = 5
      "000101" when "0101110001000111", -- t[23623] = 5
      "000101" when "0101110001001000", -- t[23624] = 5
      "000101" when "0101110001001001", -- t[23625] = 5
      "000101" when "0101110001001010", -- t[23626] = 5
      "000101" when "0101110001001011", -- t[23627] = 5
      "000101" when "0101110001001100", -- t[23628] = 5
      "000101" when "0101110001001101", -- t[23629] = 5
      "000101" when "0101110001001110", -- t[23630] = 5
      "000101" when "0101110001001111", -- t[23631] = 5
      "000101" when "0101110001010000", -- t[23632] = 5
      "000101" when "0101110001010001", -- t[23633] = 5
      "000101" when "0101110001010010", -- t[23634] = 5
      "000101" when "0101110001010011", -- t[23635] = 5
      "000101" when "0101110001010100", -- t[23636] = 5
      "000101" when "0101110001010101", -- t[23637] = 5
      "000101" when "0101110001010110", -- t[23638] = 5
      "000101" when "0101110001010111", -- t[23639] = 5
      "000101" when "0101110001011000", -- t[23640] = 5
      "000101" when "0101110001011001", -- t[23641] = 5
      "000101" when "0101110001011010", -- t[23642] = 5
      "000101" when "0101110001011011", -- t[23643] = 5
      "000101" when "0101110001011100", -- t[23644] = 5
      "000101" when "0101110001011101", -- t[23645] = 5
      "000101" when "0101110001011110", -- t[23646] = 5
      "000101" when "0101110001011111", -- t[23647] = 5
      "000101" when "0101110001100000", -- t[23648] = 5
      "000101" when "0101110001100001", -- t[23649] = 5
      "000101" when "0101110001100010", -- t[23650] = 5
      "000101" when "0101110001100011", -- t[23651] = 5
      "000101" when "0101110001100100", -- t[23652] = 5
      "000101" when "0101110001100101", -- t[23653] = 5
      "000101" when "0101110001100110", -- t[23654] = 5
      "000101" when "0101110001100111", -- t[23655] = 5
      "000101" when "0101110001101000", -- t[23656] = 5
      "000101" when "0101110001101001", -- t[23657] = 5
      "000101" when "0101110001101010", -- t[23658] = 5
      "000101" when "0101110001101011", -- t[23659] = 5
      "000101" when "0101110001101100", -- t[23660] = 5
      "000101" when "0101110001101101", -- t[23661] = 5
      "000101" when "0101110001101110", -- t[23662] = 5
      "000101" when "0101110001101111", -- t[23663] = 5
      "000101" when "0101110001110000", -- t[23664] = 5
      "000101" when "0101110001110001", -- t[23665] = 5
      "000101" when "0101110001110010", -- t[23666] = 5
      "000101" when "0101110001110011", -- t[23667] = 5
      "000101" when "0101110001110100", -- t[23668] = 5
      "000101" when "0101110001110101", -- t[23669] = 5
      "000101" when "0101110001110110", -- t[23670] = 5
      "000101" when "0101110001110111", -- t[23671] = 5
      "000101" when "0101110001111000", -- t[23672] = 5
      "000101" when "0101110001111001", -- t[23673] = 5
      "000101" when "0101110001111010", -- t[23674] = 5
      "000101" when "0101110001111011", -- t[23675] = 5
      "000101" when "0101110001111100", -- t[23676] = 5
      "000101" when "0101110001111101", -- t[23677] = 5
      "000101" when "0101110001111110", -- t[23678] = 5
      "000101" when "0101110001111111", -- t[23679] = 5
      "000101" when "0101110010000000", -- t[23680] = 5
      "000101" when "0101110010000001", -- t[23681] = 5
      "000101" when "0101110010000010", -- t[23682] = 5
      "000101" when "0101110010000011", -- t[23683] = 5
      "000101" when "0101110010000100", -- t[23684] = 5
      "000101" when "0101110010000101", -- t[23685] = 5
      "000101" when "0101110010000110", -- t[23686] = 5
      "000101" when "0101110010000111", -- t[23687] = 5
      "000101" when "0101110010001000", -- t[23688] = 5
      "000101" when "0101110010001001", -- t[23689] = 5
      "000101" when "0101110010001010", -- t[23690] = 5
      "000101" when "0101110010001011", -- t[23691] = 5
      "000101" when "0101110010001100", -- t[23692] = 5
      "000101" when "0101110010001101", -- t[23693] = 5
      "000101" when "0101110010001110", -- t[23694] = 5
      "000101" when "0101110010001111", -- t[23695] = 5
      "000101" when "0101110010010000", -- t[23696] = 5
      "000101" when "0101110010010001", -- t[23697] = 5
      "000101" when "0101110010010010", -- t[23698] = 5
      "000101" when "0101110010010011", -- t[23699] = 5
      "000101" when "0101110010010100", -- t[23700] = 5
      "000101" when "0101110010010101", -- t[23701] = 5
      "000101" when "0101110010010110", -- t[23702] = 5
      "000101" when "0101110010010111", -- t[23703] = 5
      "000101" when "0101110010011000", -- t[23704] = 5
      "000101" when "0101110010011001", -- t[23705] = 5
      "000101" when "0101110010011010", -- t[23706] = 5
      "000101" when "0101110010011011", -- t[23707] = 5
      "000101" when "0101110010011100", -- t[23708] = 5
      "000101" when "0101110010011101", -- t[23709] = 5
      "000101" when "0101110010011110", -- t[23710] = 5
      "000101" when "0101110010011111", -- t[23711] = 5
      "000101" when "0101110010100000", -- t[23712] = 5
      "000101" when "0101110010100001", -- t[23713] = 5
      "000101" when "0101110010100010", -- t[23714] = 5
      "000101" when "0101110010100011", -- t[23715] = 5
      "000101" when "0101110010100100", -- t[23716] = 5
      "000101" when "0101110010100101", -- t[23717] = 5
      "000101" when "0101110010100110", -- t[23718] = 5
      "000101" when "0101110010100111", -- t[23719] = 5
      "000101" when "0101110010101000", -- t[23720] = 5
      "000101" when "0101110010101001", -- t[23721] = 5
      "000101" when "0101110010101010", -- t[23722] = 5
      "000101" when "0101110010101011", -- t[23723] = 5
      "000101" when "0101110010101100", -- t[23724] = 5
      "000101" when "0101110010101101", -- t[23725] = 5
      "000101" when "0101110010101110", -- t[23726] = 5
      "000101" when "0101110010101111", -- t[23727] = 5
      "000101" when "0101110010110000", -- t[23728] = 5
      "000101" when "0101110010110001", -- t[23729] = 5
      "000101" when "0101110010110010", -- t[23730] = 5
      "000101" when "0101110010110011", -- t[23731] = 5
      "000101" when "0101110010110100", -- t[23732] = 5
      "000101" when "0101110010110101", -- t[23733] = 5
      "000101" when "0101110010110110", -- t[23734] = 5
      "000101" when "0101110010110111", -- t[23735] = 5
      "000101" when "0101110010111000", -- t[23736] = 5
      "000101" when "0101110010111001", -- t[23737] = 5
      "000101" when "0101110010111010", -- t[23738] = 5
      "000101" when "0101110010111011", -- t[23739] = 5
      "000101" when "0101110010111100", -- t[23740] = 5
      "000101" when "0101110010111101", -- t[23741] = 5
      "000101" when "0101110010111110", -- t[23742] = 5
      "000101" when "0101110010111111", -- t[23743] = 5
      "000101" when "0101110011000000", -- t[23744] = 5
      "000101" when "0101110011000001", -- t[23745] = 5
      "000101" when "0101110011000010", -- t[23746] = 5
      "000101" when "0101110011000011", -- t[23747] = 5
      "000101" when "0101110011000100", -- t[23748] = 5
      "000101" when "0101110011000101", -- t[23749] = 5
      "000101" when "0101110011000110", -- t[23750] = 5
      "000101" when "0101110011000111", -- t[23751] = 5
      "000101" when "0101110011001000", -- t[23752] = 5
      "000101" when "0101110011001001", -- t[23753] = 5
      "000101" when "0101110011001010", -- t[23754] = 5
      "000101" when "0101110011001011", -- t[23755] = 5
      "000101" when "0101110011001100", -- t[23756] = 5
      "000101" when "0101110011001101", -- t[23757] = 5
      "000101" when "0101110011001110", -- t[23758] = 5
      "000101" when "0101110011001111", -- t[23759] = 5
      "000101" when "0101110011010000", -- t[23760] = 5
      "000101" when "0101110011010001", -- t[23761] = 5
      "000101" when "0101110011010010", -- t[23762] = 5
      "000101" when "0101110011010011", -- t[23763] = 5
      "000101" when "0101110011010100", -- t[23764] = 5
      "000101" when "0101110011010101", -- t[23765] = 5
      "000101" when "0101110011010110", -- t[23766] = 5
      "000101" when "0101110011010111", -- t[23767] = 5
      "000101" when "0101110011011000", -- t[23768] = 5
      "000101" when "0101110011011001", -- t[23769] = 5
      "000101" when "0101110011011010", -- t[23770] = 5
      "000101" when "0101110011011011", -- t[23771] = 5
      "000101" when "0101110011011100", -- t[23772] = 5
      "000101" when "0101110011011101", -- t[23773] = 5
      "000101" when "0101110011011110", -- t[23774] = 5
      "000101" when "0101110011011111", -- t[23775] = 5
      "000101" when "0101110011100000", -- t[23776] = 5
      "000101" when "0101110011100001", -- t[23777] = 5
      "000101" when "0101110011100010", -- t[23778] = 5
      "000101" when "0101110011100011", -- t[23779] = 5
      "000101" when "0101110011100100", -- t[23780] = 5
      "000101" when "0101110011100101", -- t[23781] = 5
      "000101" when "0101110011100110", -- t[23782] = 5
      "000101" when "0101110011100111", -- t[23783] = 5
      "000101" when "0101110011101000", -- t[23784] = 5
      "000101" when "0101110011101001", -- t[23785] = 5
      "000101" when "0101110011101010", -- t[23786] = 5
      "000101" when "0101110011101011", -- t[23787] = 5
      "000101" when "0101110011101100", -- t[23788] = 5
      "000101" when "0101110011101101", -- t[23789] = 5
      "000101" when "0101110011101110", -- t[23790] = 5
      "000101" when "0101110011101111", -- t[23791] = 5
      "000101" when "0101110011110000", -- t[23792] = 5
      "000101" when "0101110011110001", -- t[23793] = 5
      "000101" when "0101110011110010", -- t[23794] = 5
      "000101" when "0101110011110011", -- t[23795] = 5
      "000101" when "0101110011110100", -- t[23796] = 5
      "000101" when "0101110011110101", -- t[23797] = 5
      "000101" when "0101110011110110", -- t[23798] = 5
      "000101" when "0101110011110111", -- t[23799] = 5
      "000101" when "0101110011111000", -- t[23800] = 5
      "000101" when "0101110011111001", -- t[23801] = 5
      "000101" when "0101110011111010", -- t[23802] = 5
      "000101" when "0101110011111011", -- t[23803] = 5
      "000101" when "0101110011111100", -- t[23804] = 5
      "000101" when "0101110011111101", -- t[23805] = 5
      "000101" when "0101110011111110", -- t[23806] = 5
      "000101" when "0101110011111111", -- t[23807] = 5
      "000101" when "0101110100000000", -- t[23808] = 5
      "000101" when "0101110100000001", -- t[23809] = 5
      "000101" when "0101110100000010", -- t[23810] = 5
      "000101" when "0101110100000011", -- t[23811] = 5
      "000101" when "0101110100000100", -- t[23812] = 5
      "000101" when "0101110100000101", -- t[23813] = 5
      "000101" when "0101110100000110", -- t[23814] = 5
      "000101" when "0101110100000111", -- t[23815] = 5
      "000101" when "0101110100001000", -- t[23816] = 5
      "000101" when "0101110100001001", -- t[23817] = 5
      "000101" when "0101110100001010", -- t[23818] = 5
      "000101" when "0101110100001011", -- t[23819] = 5
      "000101" when "0101110100001100", -- t[23820] = 5
      "000101" when "0101110100001101", -- t[23821] = 5
      "000101" when "0101110100001110", -- t[23822] = 5
      "000101" when "0101110100001111", -- t[23823] = 5
      "000101" when "0101110100010000", -- t[23824] = 5
      "000101" when "0101110100010001", -- t[23825] = 5
      "000101" when "0101110100010010", -- t[23826] = 5
      "000101" when "0101110100010011", -- t[23827] = 5
      "000101" when "0101110100010100", -- t[23828] = 5
      "000101" when "0101110100010101", -- t[23829] = 5
      "000101" when "0101110100010110", -- t[23830] = 5
      "000101" when "0101110100010111", -- t[23831] = 5
      "000101" when "0101110100011000", -- t[23832] = 5
      "000101" when "0101110100011001", -- t[23833] = 5
      "000101" when "0101110100011010", -- t[23834] = 5
      "000101" when "0101110100011011", -- t[23835] = 5
      "000101" when "0101110100011100", -- t[23836] = 5
      "000101" when "0101110100011101", -- t[23837] = 5
      "000101" when "0101110100011110", -- t[23838] = 5
      "000101" when "0101110100011111", -- t[23839] = 5
      "000101" when "0101110100100000", -- t[23840] = 5
      "000101" when "0101110100100001", -- t[23841] = 5
      "000101" when "0101110100100010", -- t[23842] = 5
      "000101" when "0101110100100011", -- t[23843] = 5
      "000101" when "0101110100100100", -- t[23844] = 5
      "000101" when "0101110100100101", -- t[23845] = 5
      "000101" when "0101110100100110", -- t[23846] = 5
      "000101" when "0101110100100111", -- t[23847] = 5
      "000101" when "0101110100101000", -- t[23848] = 5
      "000101" when "0101110100101001", -- t[23849] = 5
      "000101" when "0101110100101010", -- t[23850] = 5
      "000101" when "0101110100101011", -- t[23851] = 5
      "000101" when "0101110100101100", -- t[23852] = 5
      "000101" when "0101110100101101", -- t[23853] = 5
      "000101" when "0101110100101110", -- t[23854] = 5
      "000101" when "0101110100101111", -- t[23855] = 5
      "000101" when "0101110100110000", -- t[23856] = 5
      "000101" when "0101110100110001", -- t[23857] = 5
      "000101" when "0101110100110010", -- t[23858] = 5
      "000101" when "0101110100110011", -- t[23859] = 5
      "000101" when "0101110100110100", -- t[23860] = 5
      "000101" when "0101110100110101", -- t[23861] = 5
      "000101" when "0101110100110110", -- t[23862] = 5
      "000101" when "0101110100110111", -- t[23863] = 5
      "000101" when "0101110100111000", -- t[23864] = 5
      "000101" when "0101110100111001", -- t[23865] = 5
      "000101" when "0101110100111010", -- t[23866] = 5
      "000101" when "0101110100111011", -- t[23867] = 5
      "000101" when "0101110100111100", -- t[23868] = 5
      "000101" when "0101110100111101", -- t[23869] = 5
      "000101" when "0101110100111110", -- t[23870] = 5
      "000101" when "0101110100111111", -- t[23871] = 5
      "000101" when "0101110101000000", -- t[23872] = 5
      "000101" when "0101110101000001", -- t[23873] = 5
      "000101" when "0101110101000010", -- t[23874] = 5
      "000101" when "0101110101000011", -- t[23875] = 5
      "000101" when "0101110101000100", -- t[23876] = 5
      "000101" when "0101110101000101", -- t[23877] = 5
      "000101" when "0101110101000110", -- t[23878] = 5
      "000101" when "0101110101000111", -- t[23879] = 5
      "000101" when "0101110101001000", -- t[23880] = 5
      "000101" when "0101110101001001", -- t[23881] = 5
      "000101" when "0101110101001010", -- t[23882] = 5
      "000101" when "0101110101001011", -- t[23883] = 5
      "000101" when "0101110101001100", -- t[23884] = 5
      "000101" when "0101110101001101", -- t[23885] = 5
      "000101" when "0101110101001110", -- t[23886] = 5
      "000101" when "0101110101001111", -- t[23887] = 5
      "000101" when "0101110101010000", -- t[23888] = 5
      "000101" when "0101110101010001", -- t[23889] = 5
      "000101" when "0101110101010010", -- t[23890] = 5
      "000101" when "0101110101010011", -- t[23891] = 5
      "000101" when "0101110101010100", -- t[23892] = 5
      "000101" when "0101110101010101", -- t[23893] = 5
      "000101" when "0101110101010110", -- t[23894] = 5
      "000101" when "0101110101010111", -- t[23895] = 5
      "000101" when "0101110101011000", -- t[23896] = 5
      "000101" when "0101110101011001", -- t[23897] = 5
      "000101" when "0101110101011010", -- t[23898] = 5
      "000101" when "0101110101011011", -- t[23899] = 5
      "000101" when "0101110101011100", -- t[23900] = 5
      "000101" when "0101110101011101", -- t[23901] = 5
      "000101" when "0101110101011110", -- t[23902] = 5
      "000101" when "0101110101011111", -- t[23903] = 5
      "000101" when "0101110101100000", -- t[23904] = 5
      "000101" when "0101110101100001", -- t[23905] = 5
      "000101" when "0101110101100010", -- t[23906] = 5
      "000101" when "0101110101100011", -- t[23907] = 5
      "000101" when "0101110101100100", -- t[23908] = 5
      "000101" when "0101110101100101", -- t[23909] = 5
      "000101" when "0101110101100110", -- t[23910] = 5
      "000101" when "0101110101100111", -- t[23911] = 5
      "000101" when "0101110101101000", -- t[23912] = 5
      "000101" when "0101110101101001", -- t[23913] = 5
      "000101" when "0101110101101010", -- t[23914] = 5
      "000101" when "0101110101101011", -- t[23915] = 5
      "000101" when "0101110101101100", -- t[23916] = 5
      "000101" when "0101110101101101", -- t[23917] = 5
      "000101" when "0101110101101110", -- t[23918] = 5
      "000101" when "0101110101101111", -- t[23919] = 5
      "000101" when "0101110101110000", -- t[23920] = 5
      "000101" when "0101110101110001", -- t[23921] = 5
      "000101" when "0101110101110010", -- t[23922] = 5
      "000101" when "0101110101110011", -- t[23923] = 5
      "000101" when "0101110101110100", -- t[23924] = 5
      "000101" when "0101110101110101", -- t[23925] = 5
      "000101" when "0101110101110110", -- t[23926] = 5
      "000101" when "0101110101110111", -- t[23927] = 5
      "000101" when "0101110101111000", -- t[23928] = 5
      "000101" when "0101110101111001", -- t[23929] = 5
      "000101" when "0101110101111010", -- t[23930] = 5
      "000101" when "0101110101111011", -- t[23931] = 5
      "000101" when "0101110101111100", -- t[23932] = 5
      "000101" when "0101110101111101", -- t[23933] = 5
      "000101" when "0101110101111110", -- t[23934] = 5
      "000101" when "0101110101111111", -- t[23935] = 5
      "000101" when "0101110110000000", -- t[23936] = 5
      "000101" when "0101110110000001", -- t[23937] = 5
      "000101" when "0101110110000010", -- t[23938] = 5
      "000101" when "0101110110000011", -- t[23939] = 5
      "000101" when "0101110110000100", -- t[23940] = 5
      "000101" when "0101110110000101", -- t[23941] = 5
      "000101" when "0101110110000110", -- t[23942] = 5
      "000101" when "0101110110000111", -- t[23943] = 5
      "000101" when "0101110110001000", -- t[23944] = 5
      "000101" when "0101110110001001", -- t[23945] = 5
      "000101" when "0101110110001010", -- t[23946] = 5
      "000101" when "0101110110001011", -- t[23947] = 5
      "000101" when "0101110110001100", -- t[23948] = 5
      "000101" when "0101110110001101", -- t[23949] = 5
      "000101" when "0101110110001110", -- t[23950] = 5
      "000101" when "0101110110001111", -- t[23951] = 5
      "000101" when "0101110110010000", -- t[23952] = 5
      "000101" when "0101110110010001", -- t[23953] = 5
      "000101" when "0101110110010010", -- t[23954] = 5
      "000101" when "0101110110010011", -- t[23955] = 5
      "000101" when "0101110110010100", -- t[23956] = 5
      "000101" when "0101110110010101", -- t[23957] = 5
      "000101" when "0101110110010110", -- t[23958] = 5
      "000101" when "0101110110010111", -- t[23959] = 5
      "000101" when "0101110110011000", -- t[23960] = 5
      "000101" when "0101110110011001", -- t[23961] = 5
      "000101" when "0101110110011010", -- t[23962] = 5
      "000101" when "0101110110011011", -- t[23963] = 5
      "000101" when "0101110110011100", -- t[23964] = 5
      "000101" when "0101110110011101", -- t[23965] = 5
      "000101" when "0101110110011110", -- t[23966] = 5
      "000101" when "0101110110011111", -- t[23967] = 5
      "000101" when "0101110110100000", -- t[23968] = 5
      "000101" when "0101110110100001", -- t[23969] = 5
      "000101" when "0101110110100010", -- t[23970] = 5
      "000101" when "0101110110100011", -- t[23971] = 5
      "000101" when "0101110110100100", -- t[23972] = 5
      "000101" when "0101110110100101", -- t[23973] = 5
      "000101" when "0101110110100110", -- t[23974] = 5
      "000101" when "0101110110100111", -- t[23975] = 5
      "000101" when "0101110110101000", -- t[23976] = 5
      "000101" when "0101110110101001", -- t[23977] = 5
      "000101" when "0101110110101010", -- t[23978] = 5
      "000101" when "0101110110101011", -- t[23979] = 5
      "000101" when "0101110110101100", -- t[23980] = 5
      "000101" when "0101110110101101", -- t[23981] = 5
      "000101" when "0101110110101110", -- t[23982] = 5
      "000101" when "0101110110101111", -- t[23983] = 5
      "000101" when "0101110110110000", -- t[23984] = 5
      "000101" when "0101110110110001", -- t[23985] = 5
      "000101" when "0101110110110010", -- t[23986] = 5
      "000101" when "0101110110110011", -- t[23987] = 5
      "000101" when "0101110110110100", -- t[23988] = 5
      "000101" when "0101110110110101", -- t[23989] = 5
      "000101" when "0101110110110110", -- t[23990] = 5
      "000101" when "0101110110110111", -- t[23991] = 5
      "000101" when "0101110110111000", -- t[23992] = 5
      "000101" when "0101110110111001", -- t[23993] = 5
      "000101" when "0101110110111010", -- t[23994] = 5
      "000101" when "0101110110111011", -- t[23995] = 5
      "000101" when "0101110110111100", -- t[23996] = 5
      "000101" when "0101110110111101", -- t[23997] = 5
      "000101" when "0101110110111110", -- t[23998] = 5
      "000101" when "0101110110111111", -- t[23999] = 5
      "000101" when "0101110111000000", -- t[24000] = 5
      "000101" when "0101110111000001", -- t[24001] = 5
      "000101" when "0101110111000010", -- t[24002] = 5
      "000101" when "0101110111000011", -- t[24003] = 5
      "000101" when "0101110111000100", -- t[24004] = 5
      "000101" when "0101110111000101", -- t[24005] = 5
      "000101" when "0101110111000110", -- t[24006] = 5
      "000101" when "0101110111000111", -- t[24007] = 5
      "000101" when "0101110111001000", -- t[24008] = 5
      "000101" when "0101110111001001", -- t[24009] = 5
      "000101" when "0101110111001010", -- t[24010] = 5
      "000101" when "0101110111001011", -- t[24011] = 5
      "000101" when "0101110111001100", -- t[24012] = 5
      "000101" when "0101110111001101", -- t[24013] = 5
      "000101" when "0101110111001110", -- t[24014] = 5
      "000101" when "0101110111001111", -- t[24015] = 5
      "000101" when "0101110111010000", -- t[24016] = 5
      "000101" when "0101110111010001", -- t[24017] = 5
      "000101" when "0101110111010010", -- t[24018] = 5
      "000101" when "0101110111010011", -- t[24019] = 5
      "000101" when "0101110111010100", -- t[24020] = 5
      "000101" when "0101110111010101", -- t[24021] = 5
      "000101" when "0101110111010110", -- t[24022] = 5
      "000101" when "0101110111010111", -- t[24023] = 5
      "000101" when "0101110111011000", -- t[24024] = 5
      "000101" when "0101110111011001", -- t[24025] = 5
      "000101" when "0101110111011010", -- t[24026] = 5
      "000101" when "0101110111011011", -- t[24027] = 5
      "000101" when "0101110111011100", -- t[24028] = 5
      "000101" when "0101110111011101", -- t[24029] = 5
      "000101" when "0101110111011110", -- t[24030] = 5
      "000101" when "0101110111011111", -- t[24031] = 5
      "000101" when "0101110111100000", -- t[24032] = 5
      "000101" when "0101110111100001", -- t[24033] = 5
      "000101" when "0101110111100010", -- t[24034] = 5
      "000101" when "0101110111100011", -- t[24035] = 5
      "000101" when "0101110111100100", -- t[24036] = 5
      "000101" when "0101110111100101", -- t[24037] = 5
      "000101" when "0101110111100110", -- t[24038] = 5
      "000101" when "0101110111100111", -- t[24039] = 5
      "000101" when "0101110111101000", -- t[24040] = 5
      "000101" when "0101110111101001", -- t[24041] = 5
      "000101" when "0101110111101010", -- t[24042] = 5
      "000101" when "0101110111101011", -- t[24043] = 5
      "000101" when "0101110111101100", -- t[24044] = 5
      "000101" when "0101110111101101", -- t[24045] = 5
      "000101" when "0101110111101110", -- t[24046] = 5
      "000101" when "0101110111101111", -- t[24047] = 5
      "000101" when "0101110111110000", -- t[24048] = 5
      "000101" when "0101110111110001", -- t[24049] = 5
      "000101" when "0101110111110010", -- t[24050] = 5
      "000101" when "0101110111110011", -- t[24051] = 5
      "000101" when "0101110111110100", -- t[24052] = 5
      "000101" when "0101110111110101", -- t[24053] = 5
      "000101" when "0101110111110110", -- t[24054] = 5
      "000101" when "0101110111110111", -- t[24055] = 5
      "000101" when "0101110111111000", -- t[24056] = 5
      "000101" when "0101110111111001", -- t[24057] = 5
      "000101" when "0101110111111010", -- t[24058] = 5
      "000101" when "0101110111111011", -- t[24059] = 5
      "000101" when "0101110111111100", -- t[24060] = 5
      "000101" when "0101110111111101", -- t[24061] = 5
      "000101" when "0101110111111110", -- t[24062] = 5
      "000101" when "0101110111111111", -- t[24063] = 5
      "000101" when "0101111000000000", -- t[24064] = 5
      "000101" when "0101111000000001", -- t[24065] = 5
      "000101" when "0101111000000010", -- t[24066] = 5
      "000101" when "0101111000000011", -- t[24067] = 5
      "000101" when "0101111000000100", -- t[24068] = 5
      "000101" when "0101111000000101", -- t[24069] = 5
      "000101" when "0101111000000110", -- t[24070] = 5
      "000101" when "0101111000000111", -- t[24071] = 5
      "000101" when "0101111000001000", -- t[24072] = 5
      "000101" when "0101111000001001", -- t[24073] = 5
      "000101" when "0101111000001010", -- t[24074] = 5
      "000101" when "0101111000001011", -- t[24075] = 5
      "000101" when "0101111000001100", -- t[24076] = 5
      "000101" when "0101111000001101", -- t[24077] = 5
      "000101" when "0101111000001110", -- t[24078] = 5
      "000101" when "0101111000001111", -- t[24079] = 5
      "000101" when "0101111000010000", -- t[24080] = 5
      "000101" when "0101111000010001", -- t[24081] = 5
      "000101" when "0101111000010010", -- t[24082] = 5
      "000101" when "0101111000010011", -- t[24083] = 5
      "000101" when "0101111000010100", -- t[24084] = 5
      "000101" when "0101111000010101", -- t[24085] = 5
      "000101" when "0101111000010110", -- t[24086] = 5
      "000101" when "0101111000010111", -- t[24087] = 5
      "000101" when "0101111000011000", -- t[24088] = 5
      "000101" when "0101111000011001", -- t[24089] = 5
      "000101" when "0101111000011010", -- t[24090] = 5
      "000101" when "0101111000011011", -- t[24091] = 5
      "000101" when "0101111000011100", -- t[24092] = 5
      "000101" when "0101111000011101", -- t[24093] = 5
      "000101" when "0101111000011110", -- t[24094] = 5
      "000101" when "0101111000011111", -- t[24095] = 5
      "000101" when "0101111000100000", -- t[24096] = 5
      "000101" when "0101111000100001", -- t[24097] = 5
      "000101" when "0101111000100010", -- t[24098] = 5
      "000101" when "0101111000100011", -- t[24099] = 5
      "000101" when "0101111000100100", -- t[24100] = 5
      "000101" when "0101111000100101", -- t[24101] = 5
      "000101" when "0101111000100110", -- t[24102] = 5
      "000101" when "0101111000100111", -- t[24103] = 5
      "000101" when "0101111000101000", -- t[24104] = 5
      "000101" when "0101111000101001", -- t[24105] = 5
      "000101" when "0101111000101010", -- t[24106] = 5
      "000101" when "0101111000101011", -- t[24107] = 5
      "000101" when "0101111000101100", -- t[24108] = 5
      "000101" when "0101111000101101", -- t[24109] = 5
      "000101" when "0101111000101110", -- t[24110] = 5
      "000101" when "0101111000101111", -- t[24111] = 5
      "000101" when "0101111000110000", -- t[24112] = 5
      "000101" when "0101111000110001", -- t[24113] = 5
      "000101" when "0101111000110010", -- t[24114] = 5
      "000101" when "0101111000110011", -- t[24115] = 5
      "000101" when "0101111000110100", -- t[24116] = 5
      "000101" when "0101111000110101", -- t[24117] = 5
      "000101" when "0101111000110110", -- t[24118] = 5
      "000101" when "0101111000110111", -- t[24119] = 5
      "000101" when "0101111000111000", -- t[24120] = 5
      "000101" when "0101111000111001", -- t[24121] = 5
      "000101" when "0101111000111010", -- t[24122] = 5
      "000101" when "0101111000111011", -- t[24123] = 5
      "000101" when "0101111000111100", -- t[24124] = 5
      "000101" when "0101111000111101", -- t[24125] = 5
      "000101" when "0101111000111110", -- t[24126] = 5
      "000101" when "0101111000111111", -- t[24127] = 5
      "000101" when "0101111001000000", -- t[24128] = 5
      "000101" when "0101111001000001", -- t[24129] = 5
      "000101" when "0101111001000010", -- t[24130] = 5
      "000101" when "0101111001000011", -- t[24131] = 5
      "000101" when "0101111001000100", -- t[24132] = 5
      "000101" when "0101111001000101", -- t[24133] = 5
      "000101" when "0101111001000110", -- t[24134] = 5
      "000101" when "0101111001000111", -- t[24135] = 5
      "000101" when "0101111001001000", -- t[24136] = 5
      "000101" when "0101111001001001", -- t[24137] = 5
      "000101" when "0101111001001010", -- t[24138] = 5
      "000101" when "0101111001001011", -- t[24139] = 5
      "000101" when "0101111001001100", -- t[24140] = 5
      "000101" when "0101111001001101", -- t[24141] = 5
      "000101" when "0101111001001110", -- t[24142] = 5
      "000101" when "0101111001001111", -- t[24143] = 5
      "000101" when "0101111001010000", -- t[24144] = 5
      "000101" when "0101111001010001", -- t[24145] = 5
      "000101" when "0101111001010010", -- t[24146] = 5
      "000101" when "0101111001010011", -- t[24147] = 5
      "000101" when "0101111001010100", -- t[24148] = 5
      "000101" when "0101111001010101", -- t[24149] = 5
      "000101" when "0101111001010110", -- t[24150] = 5
      "000101" when "0101111001010111", -- t[24151] = 5
      "000101" when "0101111001011000", -- t[24152] = 5
      "000101" when "0101111001011001", -- t[24153] = 5
      "000101" when "0101111001011010", -- t[24154] = 5
      "000101" when "0101111001011011", -- t[24155] = 5
      "000101" when "0101111001011100", -- t[24156] = 5
      "000101" when "0101111001011101", -- t[24157] = 5
      "000101" when "0101111001011110", -- t[24158] = 5
      "000101" when "0101111001011111", -- t[24159] = 5
      "000101" when "0101111001100000", -- t[24160] = 5
      "000101" when "0101111001100001", -- t[24161] = 5
      "000101" when "0101111001100010", -- t[24162] = 5
      "000101" when "0101111001100011", -- t[24163] = 5
      "000101" when "0101111001100100", -- t[24164] = 5
      "000101" when "0101111001100101", -- t[24165] = 5
      "000101" when "0101111001100110", -- t[24166] = 5
      "000101" when "0101111001100111", -- t[24167] = 5
      "000101" when "0101111001101000", -- t[24168] = 5
      "000101" when "0101111001101001", -- t[24169] = 5
      "000101" when "0101111001101010", -- t[24170] = 5
      "000101" when "0101111001101011", -- t[24171] = 5
      "000101" when "0101111001101100", -- t[24172] = 5
      "000101" when "0101111001101101", -- t[24173] = 5
      "000101" when "0101111001101110", -- t[24174] = 5
      "000101" when "0101111001101111", -- t[24175] = 5
      "000101" when "0101111001110000", -- t[24176] = 5
      "000101" when "0101111001110001", -- t[24177] = 5
      "000101" when "0101111001110010", -- t[24178] = 5
      "000101" when "0101111001110011", -- t[24179] = 5
      "000101" when "0101111001110100", -- t[24180] = 5
      "000101" when "0101111001110101", -- t[24181] = 5
      "000101" when "0101111001110110", -- t[24182] = 5
      "000101" when "0101111001110111", -- t[24183] = 5
      "000101" when "0101111001111000", -- t[24184] = 5
      "000101" when "0101111001111001", -- t[24185] = 5
      "000101" when "0101111001111010", -- t[24186] = 5
      "000101" when "0101111001111011", -- t[24187] = 5
      "000101" when "0101111001111100", -- t[24188] = 5
      "000101" when "0101111001111101", -- t[24189] = 5
      "000101" when "0101111001111110", -- t[24190] = 5
      "000101" when "0101111001111111", -- t[24191] = 5
      "000101" when "0101111010000000", -- t[24192] = 5
      "000101" when "0101111010000001", -- t[24193] = 5
      "000101" when "0101111010000010", -- t[24194] = 5
      "000101" when "0101111010000011", -- t[24195] = 5
      "000101" when "0101111010000100", -- t[24196] = 5
      "000101" when "0101111010000101", -- t[24197] = 5
      "000101" when "0101111010000110", -- t[24198] = 5
      "000101" when "0101111010000111", -- t[24199] = 5
      "000101" when "0101111010001000", -- t[24200] = 5
      "000101" when "0101111010001001", -- t[24201] = 5
      "000101" when "0101111010001010", -- t[24202] = 5
      "000101" when "0101111010001011", -- t[24203] = 5
      "000101" when "0101111010001100", -- t[24204] = 5
      "000101" when "0101111010001101", -- t[24205] = 5
      "000101" when "0101111010001110", -- t[24206] = 5
      "000101" when "0101111010001111", -- t[24207] = 5
      "000101" when "0101111010010000", -- t[24208] = 5
      "000101" when "0101111010010001", -- t[24209] = 5
      "000101" when "0101111010010010", -- t[24210] = 5
      "000101" when "0101111010010011", -- t[24211] = 5
      "000101" when "0101111010010100", -- t[24212] = 5
      "000101" when "0101111010010101", -- t[24213] = 5
      "000101" when "0101111010010110", -- t[24214] = 5
      "000101" when "0101111010010111", -- t[24215] = 5
      "000101" when "0101111010011000", -- t[24216] = 5
      "000101" when "0101111010011001", -- t[24217] = 5
      "000101" when "0101111010011010", -- t[24218] = 5
      "000101" when "0101111010011011", -- t[24219] = 5
      "000101" when "0101111010011100", -- t[24220] = 5
      "000101" when "0101111010011101", -- t[24221] = 5
      "000101" when "0101111010011110", -- t[24222] = 5
      "000101" when "0101111010011111", -- t[24223] = 5
      "000101" when "0101111010100000", -- t[24224] = 5
      "000101" when "0101111010100001", -- t[24225] = 5
      "000101" when "0101111010100010", -- t[24226] = 5
      "000101" when "0101111010100011", -- t[24227] = 5
      "000101" when "0101111010100100", -- t[24228] = 5
      "000101" when "0101111010100101", -- t[24229] = 5
      "000101" when "0101111010100110", -- t[24230] = 5
      "000101" when "0101111010100111", -- t[24231] = 5
      "000101" when "0101111010101000", -- t[24232] = 5
      "000101" when "0101111010101001", -- t[24233] = 5
      "000101" when "0101111010101010", -- t[24234] = 5
      "000101" when "0101111010101011", -- t[24235] = 5
      "000101" when "0101111010101100", -- t[24236] = 5
      "000101" when "0101111010101101", -- t[24237] = 5
      "000101" when "0101111010101110", -- t[24238] = 5
      "000101" when "0101111010101111", -- t[24239] = 5
      "000101" when "0101111010110000", -- t[24240] = 5
      "000101" when "0101111010110001", -- t[24241] = 5
      "000101" when "0101111010110010", -- t[24242] = 5
      "000101" when "0101111010110011", -- t[24243] = 5
      "000101" when "0101111010110100", -- t[24244] = 5
      "000101" when "0101111010110101", -- t[24245] = 5
      "000101" when "0101111010110110", -- t[24246] = 5
      "000101" when "0101111010110111", -- t[24247] = 5
      "000101" when "0101111010111000", -- t[24248] = 5
      "000101" when "0101111010111001", -- t[24249] = 5
      "000101" when "0101111010111010", -- t[24250] = 5
      "000101" when "0101111010111011", -- t[24251] = 5
      "000101" when "0101111010111100", -- t[24252] = 5
      "000101" when "0101111010111101", -- t[24253] = 5
      "000101" when "0101111010111110", -- t[24254] = 5
      "000101" when "0101111010111111", -- t[24255] = 5
      "000101" when "0101111011000000", -- t[24256] = 5
      "000101" when "0101111011000001", -- t[24257] = 5
      "000101" when "0101111011000010", -- t[24258] = 5
      "000101" when "0101111011000011", -- t[24259] = 5
      "000101" when "0101111011000100", -- t[24260] = 5
      "000101" when "0101111011000101", -- t[24261] = 5
      "000101" when "0101111011000110", -- t[24262] = 5
      "000101" when "0101111011000111", -- t[24263] = 5
      "000101" when "0101111011001000", -- t[24264] = 5
      "000101" when "0101111011001001", -- t[24265] = 5
      "000101" when "0101111011001010", -- t[24266] = 5
      "000101" when "0101111011001011", -- t[24267] = 5
      "000101" when "0101111011001100", -- t[24268] = 5
      "000101" when "0101111011001101", -- t[24269] = 5
      "000101" when "0101111011001110", -- t[24270] = 5
      "000101" when "0101111011001111", -- t[24271] = 5
      "000101" when "0101111011010000", -- t[24272] = 5
      "000101" when "0101111011010001", -- t[24273] = 5
      "000101" when "0101111011010010", -- t[24274] = 5
      "000101" when "0101111011010011", -- t[24275] = 5
      "000101" when "0101111011010100", -- t[24276] = 5
      "000101" when "0101111011010101", -- t[24277] = 5
      "000101" when "0101111011010110", -- t[24278] = 5
      "000101" when "0101111011010111", -- t[24279] = 5
      "000101" when "0101111011011000", -- t[24280] = 5
      "000101" when "0101111011011001", -- t[24281] = 5
      "000101" when "0101111011011010", -- t[24282] = 5
      "000101" when "0101111011011011", -- t[24283] = 5
      "000101" when "0101111011011100", -- t[24284] = 5
      "000101" when "0101111011011101", -- t[24285] = 5
      "000101" when "0101111011011110", -- t[24286] = 5
      "000101" when "0101111011011111", -- t[24287] = 5
      "000101" when "0101111011100000", -- t[24288] = 5
      "000101" when "0101111011100001", -- t[24289] = 5
      "000110" when "0101111011100010", -- t[24290] = 6
      "000110" when "0101111011100011", -- t[24291] = 6
      "000110" when "0101111011100100", -- t[24292] = 6
      "000110" when "0101111011100101", -- t[24293] = 6
      "000110" when "0101111011100110", -- t[24294] = 6
      "000110" when "0101111011100111", -- t[24295] = 6
      "000110" when "0101111011101000", -- t[24296] = 6
      "000110" when "0101111011101001", -- t[24297] = 6
      "000110" when "0101111011101010", -- t[24298] = 6
      "000110" when "0101111011101011", -- t[24299] = 6
      "000110" when "0101111011101100", -- t[24300] = 6
      "000110" when "0101111011101101", -- t[24301] = 6
      "000110" when "0101111011101110", -- t[24302] = 6
      "000110" when "0101111011101111", -- t[24303] = 6
      "000110" when "0101111011110000", -- t[24304] = 6
      "000110" when "0101111011110001", -- t[24305] = 6
      "000110" when "0101111011110010", -- t[24306] = 6
      "000110" when "0101111011110011", -- t[24307] = 6
      "000110" when "0101111011110100", -- t[24308] = 6
      "000110" when "0101111011110101", -- t[24309] = 6
      "000110" when "0101111011110110", -- t[24310] = 6
      "000110" when "0101111011110111", -- t[24311] = 6
      "000110" when "0101111011111000", -- t[24312] = 6
      "000110" when "0101111011111001", -- t[24313] = 6
      "000110" when "0101111011111010", -- t[24314] = 6
      "000110" when "0101111011111011", -- t[24315] = 6
      "000110" when "0101111011111100", -- t[24316] = 6
      "000110" when "0101111011111101", -- t[24317] = 6
      "000110" when "0101111011111110", -- t[24318] = 6
      "000110" when "0101111011111111", -- t[24319] = 6
      "000110" when "0101111100000000", -- t[24320] = 6
      "000110" when "0101111100000001", -- t[24321] = 6
      "000110" when "0101111100000010", -- t[24322] = 6
      "000110" when "0101111100000011", -- t[24323] = 6
      "000110" when "0101111100000100", -- t[24324] = 6
      "000110" when "0101111100000101", -- t[24325] = 6
      "000110" when "0101111100000110", -- t[24326] = 6
      "000110" when "0101111100000111", -- t[24327] = 6
      "000110" when "0101111100001000", -- t[24328] = 6
      "000110" when "0101111100001001", -- t[24329] = 6
      "000110" when "0101111100001010", -- t[24330] = 6
      "000110" when "0101111100001011", -- t[24331] = 6
      "000110" when "0101111100001100", -- t[24332] = 6
      "000110" when "0101111100001101", -- t[24333] = 6
      "000110" when "0101111100001110", -- t[24334] = 6
      "000110" when "0101111100001111", -- t[24335] = 6
      "000110" when "0101111100010000", -- t[24336] = 6
      "000110" when "0101111100010001", -- t[24337] = 6
      "000110" when "0101111100010010", -- t[24338] = 6
      "000110" when "0101111100010011", -- t[24339] = 6
      "000110" when "0101111100010100", -- t[24340] = 6
      "000110" when "0101111100010101", -- t[24341] = 6
      "000110" when "0101111100010110", -- t[24342] = 6
      "000110" when "0101111100010111", -- t[24343] = 6
      "000110" when "0101111100011000", -- t[24344] = 6
      "000110" when "0101111100011001", -- t[24345] = 6
      "000110" when "0101111100011010", -- t[24346] = 6
      "000110" when "0101111100011011", -- t[24347] = 6
      "000110" when "0101111100011100", -- t[24348] = 6
      "000110" when "0101111100011101", -- t[24349] = 6
      "000110" when "0101111100011110", -- t[24350] = 6
      "000110" when "0101111100011111", -- t[24351] = 6
      "000110" when "0101111100100000", -- t[24352] = 6
      "000110" when "0101111100100001", -- t[24353] = 6
      "000110" when "0101111100100010", -- t[24354] = 6
      "000110" when "0101111100100011", -- t[24355] = 6
      "000110" when "0101111100100100", -- t[24356] = 6
      "000110" when "0101111100100101", -- t[24357] = 6
      "000110" when "0101111100100110", -- t[24358] = 6
      "000110" when "0101111100100111", -- t[24359] = 6
      "000110" when "0101111100101000", -- t[24360] = 6
      "000110" when "0101111100101001", -- t[24361] = 6
      "000110" when "0101111100101010", -- t[24362] = 6
      "000110" when "0101111100101011", -- t[24363] = 6
      "000110" when "0101111100101100", -- t[24364] = 6
      "000110" when "0101111100101101", -- t[24365] = 6
      "000110" when "0101111100101110", -- t[24366] = 6
      "000110" when "0101111100101111", -- t[24367] = 6
      "000110" when "0101111100110000", -- t[24368] = 6
      "000110" when "0101111100110001", -- t[24369] = 6
      "000110" when "0101111100110010", -- t[24370] = 6
      "000110" when "0101111100110011", -- t[24371] = 6
      "000110" when "0101111100110100", -- t[24372] = 6
      "000110" when "0101111100110101", -- t[24373] = 6
      "000110" when "0101111100110110", -- t[24374] = 6
      "000110" when "0101111100110111", -- t[24375] = 6
      "000110" when "0101111100111000", -- t[24376] = 6
      "000110" when "0101111100111001", -- t[24377] = 6
      "000110" when "0101111100111010", -- t[24378] = 6
      "000110" when "0101111100111011", -- t[24379] = 6
      "000110" when "0101111100111100", -- t[24380] = 6
      "000110" when "0101111100111101", -- t[24381] = 6
      "000110" when "0101111100111110", -- t[24382] = 6
      "000110" when "0101111100111111", -- t[24383] = 6
      "000110" when "0101111101000000", -- t[24384] = 6
      "000110" when "0101111101000001", -- t[24385] = 6
      "000110" when "0101111101000010", -- t[24386] = 6
      "000110" when "0101111101000011", -- t[24387] = 6
      "000110" when "0101111101000100", -- t[24388] = 6
      "000110" when "0101111101000101", -- t[24389] = 6
      "000110" when "0101111101000110", -- t[24390] = 6
      "000110" when "0101111101000111", -- t[24391] = 6
      "000110" when "0101111101001000", -- t[24392] = 6
      "000110" when "0101111101001001", -- t[24393] = 6
      "000110" when "0101111101001010", -- t[24394] = 6
      "000110" when "0101111101001011", -- t[24395] = 6
      "000110" when "0101111101001100", -- t[24396] = 6
      "000110" when "0101111101001101", -- t[24397] = 6
      "000110" when "0101111101001110", -- t[24398] = 6
      "000110" when "0101111101001111", -- t[24399] = 6
      "000110" when "0101111101010000", -- t[24400] = 6
      "000110" when "0101111101010001", -- t[24401] = 6
      "000110" when "0101111101010010", -- t[24402] = 6
      "000110" when "0101111101010011", -- t[24403] = 6
      "000110" when "0101111101010100", -- t[24404] = 6
      "000110" when "0101111101010101", -- t[24405] = 6
      "000110" when "0101111101010110", -- t[24406] = 6
      "000110" when "0101111101010111", -- t[24407] = 6
      "000110" when "0101111101011000", -- t[24408] = 6
      "000110" when "0101111101011001", -- t[24409] = 6
      "000110" when "0101111101011010", -- t[24410] = 6
      "000110" when "0101111101011011", -- t[24411] = 6
      "000110" when "0101111101011100", -- t[24412] = 6
      "000110" when "0101111101011101", -- t[24413] = 6
      "000110" when "0101111101011110", -- t[24414] = 6
      "000110" when "0101111101011111", -- t[24415] = 6
      "000110" when "0101111101100000", -- t[24416] = 6
      "000110" when "0101111101100001", -- t[24417] = 6
      "000110" when "0101111101100010", -- t[24418] = 6
      "000110" when "0101111101100011", -- t[24419] = 6
      "000110" when "0101111101100100", -- t[24420] = 6
      "000110" when "0101111101100101", -- t[24421] = 6
      "000110" when "0101111101100110", -- t[24422] = 6
      "000110" when "0101111101100111", -- t[24423] = 6
      "000110" when "0101111101101000", -- t[24424] = 6
      "000110" when "0101111101101001", -- t[24425] = 6
      "000110" when "0101111101101010", -- t[24426] = 6
      "000110" when "0101111101101011", -- t[24427] = 6
      "000110" when "0101111101101100", -- t[24428] = 6
      "000110" when "0101111101101101", -- t[24429] = 6
      "000110" when "0101111101101110", -- t[24430] = 6
      "000110" when "0101111101101111", -- t[24431] = 6
      "000110" when "0101111101110000", -- t[24432] = 6
      "000110" when "0101111101110001", -- t[24433] = 6
      "000110" when "0101111101110010", -- t[24434] = 6
      "000110" when "0101111101110011", -- t[24435] = 6
      "000110" when "0101111101110100", -- t[24436] = 6
      "000110" when "0101111101110101", -- t[24437] = 6
      "000110" when "0101111101110110", -- t[24438] = 6
      "000110" when "0101111101110111", -- t[24439] = 6
      "000110" when "0101111101111000", -- t[24440] = 6
      "000110" when "0101111101111001", -- t[24441] = 6
      "000110" when "0101111101111010", -- t[24442] = 6
      "000110" when "0101111101111011", -- t[24443] = 6
      "000110" when "0101111101111100", -- t[24444] = 6
      "000110" when "0101111101111101", -- t[24445] = 6
      "000110" when "0101111101111110", -- t[24446] = 6
      "000110" when "0101111101111111", -- t[24447] = 6
      "000110" when "0101111110000000", -- t[24448] = 6
      "000110" when "0101111110000001", -- t[24449] = 6
      "000110" when "0101111110000010", -- t[24450] = 6
      "000110" when "0101111110000011", -- t[24451] = 6
      "000110" when "0101111110000100", -- t[24452] = 6
      "000110" when "0101111110000101", -- t[24453] = 6
      "000110" when "0101111110000110", -- t[24454] = 6
      "000110" when "0101111110000111", -- t[24455] = 6
      "000110" when "0101111110001000", -- t[24456] = 6
      "000110" when "0101111110001001", -- t[24457] = 6
      "000110" when "0101111110001010", -- t[24458] = 6
      "000110" when "0101111110001011", -- t[24459] = 6
      "000110" when "0101111110001100", -- t[24460] = 6
      "000110" when "0101111110001101", -- t[24461] = 6
      "000110" when "0101111110001110", -- t[24462] = 6
      "000110" when "0101111110001111", -- t[24463] = 6
      "000110" when "0101111110010000", -- t[24464] = 6
      "000110" when "0101111110010001", -- t[24465] = 6
      "000110" when "0101111110010010", -- t[24466] = 6
      "000110" when "0101111110010011", -- t[24467] = 6
      "000110" when "0101111110010100", -- t[24468] = 6
      "000110" when "0101111110010101", -- t[24469] = 6
      "000110" when "0101111110010110", -- t[24470] = 6
      "000110" when "0101111110010111", -- t[24471] = 6
      "000110" when "0101111110011000", -- t[24472] = 6
      "000110" when "0101111110011001", -- t[24473] = 6
      "000110" when "0101111110011010", -- t[24474] = 6
      "000110" when "0101111110011011", -- t[24475] = 6
      "000110" when "0101111110011100", -- t[24476] = 6
      "000110" when "0101111110011101", -- t[24477] = 6
      "000110" when "0101111110011110", -- t[24478] = 6
      "000110" when "0101111110011111", -- t[24479] = 6
      "000110" when "0101111110100000", -- t[24480] = 6
      "000110" when "0101111110100001", -- t[24481] = 6
      "000110" when "0101111110100010", -- t[24482] = 6
      "000110" when "0101111110100011", -- t[24483] = 6
      "000110" when "0101111110100100", -- t[24484] = 6
      "000110" when "0101111110100101", -- t[24485] = 6
      "000110" when "0101111110100110", -- t[24486] = 6
      "000110" when "0101111110100111", -- t[24487] = 6
      "000110" when "0101111110101000", -- t[24488] = 6
      "000110" when "0101111110101001", -- t[24489] = 6
      "000110" when "0101111110101010", -- t[24490] = 6
      "000110" when "0101111110101011", -- t[24491] = 6
      "000110" when "0101111110101100", -- t[24492] = 6
      "000110" when "0101111110101101", -- t[24493] = 6
      "000110" when "0101111110101110", -- t[24494] = 6
      "000110" when "0101111110101111", -- t[24495] = 6
      "000110" when "0101111110110000", -- t[24496] = 6
      "000110" when "0101111110110001", -- t[24497] = 6
      "000110" when "0101111110110010", -- t[24498] = 6
      "000110" when "0101111110110011", -- t[24499] = 6
      "000110" when "0101111110110100", -- t[24500] = 6
      "000110" when "0101111110110101", -- t[24501] = 6
      "000110" when "0101111110110110", -- t[24502] = 6
      "000110" when "0101111110110111", -- t[24503] = 6
      "000110" when "0101111110111000", -- t[24504] = 6
      "000110" when "0101111110111001", -- t[24505] = 6
      "000110" when "0101111110111010", -- t[24506] = 6
      "000110" when "0101111110111011", -- t[24507] = 6
      "000110" when "0101111110111100", -- t[24508] = 6
      "000110" when "0101111110111101", -- t[24509] = 6
      "000110" when "0101111110111110", -- t[24510] = 6
      "000110" when "0101111110111111", -- t[24511] = 6
      "000110" when "0101111111000000", -- t[24512] = 6
      "000110" when "0101111111000001", -- t[24513] = 6
      "000110" when "0101111111000010", -- t[24514] = 6
      "000110" when "0101111111000011", -- t[24515] = 6
      "000110" when "0101111111000100", -- t[24516] = 6
      "000110" when "0101111111000101", -- t[24517] = 6
      "000110" when "0101111111000110", -- t[24518] = 6
      "000110" when "0101111111000111", -- t[24519] = 6
      "000110" when "0101111111001000", -- t[24520] = 6
      "000110" when "0101111111001001", -- t[24521] = 6
      "000110" when "0101111111001010", -- t[24522] = 6
      "000110" when "0101111111001011", -- t[24523] = 6
      "000110" when "0101111111001100", -- t[24524] = 6
      "000110" when "0101111111001101", -- t[24525] = 6
      "000110" when "0101111111001110", -- t[24526] = 6
      "000110" when "0101111111001111", -- t[24527] = 6
      "000110" when "0101111111010000", -- t[24528] = 6
      "000110" when "0101111111010001", -- t[24529] = 6
      "000110" when "0101111111010010", -- t[24530] = 6
      "000110" when "0101111111010011", -- t[24531] = 6
      "000110" when "0101111111010100", -- t[24532] = 6
      "000110" when "0101111111010101", -- t[24533] = 6
      "000110" when "0101111111010110", -- t[24534] = 6
      "000110" when "0101111111010111", -- t[24535] = 6
      "000110" when "0101111111011000", -- t[24536] = 6
      "000110" when "0101111111011001", -- t[24537] = 6
      "000110" when "0101111111011010", -- t[24538] = 6
      "000110" when "0101111111011011", -- t[24539] = 6
      "000110" when "0101111111011100", -- t[24540] = 6
      "000110" when "0101111111011101", -- t[24541] = 6
      "000110" when "0101111111011110", -- t[24542] = 6
      "000110" when "0101111111011111", -- t[24543] = 6
      "000110" when "0101111111100000", -- t[24544] = 6
      "000110" when "0101111111100001", -- t[24545] = 6
      "000110" when "0101111111100010", -- t[24546] = 6
      "000110" when "0101111111100011", -- t[24547] = 6
      "000110" when "0101111111100100", -- t[24548] = 6
      "000110" when "0101111111100101", -- t[24549] = 6
      "000110" when "0101111111100110", -- t[24550] = 6
      "000110" when "0101111111100111", -- t[24551] = 6
      "000110" when "0101111111101000", -- t[24552] = 6
      "000110" when "0101111111101001", -- t[24553] = 6
      "000110" when "0101111111101010", -- t[24554] = 6
      "000110" when "0101111111101011", -- t[24555] = 6
      "000110" when "0101111111101100", -- t[24556] = 6
      "000110" when "0101111111101101", -- t[24557] = 6
      "000110" when "0101111111101110", -- t[24558] = 6
      "000110" when "0101111111101111", -- t[24559] = 6
      "000110" when "0101111111110000", -- t[24560] = 6
      "000110" when "0101111111110001", -- t[24561] = 6
      "000110" when "0101111111110010", -- t[24562] = 6
      "000110" when "0101111111110011", -- t[24563] = 6
      "000110" when "0101111111110100", -- t[24564] = 6
      "000110" when "0101111111110101", -- t[24565] = 6
      "000110" when "0101111111110110", -- t[24566] = 6
      "000110" when "0101111111110111", -- t[24567] = 6
      "000110" when "0101111111111000", -- t[24568] = 6
      "000110" when "0101111111111001", -- t[24569] = 6
      "000110" when "0101111111111010", -- t[24570] = 6
      "000110" when "0101111111111011", -- t[24571] = 6
      "000110" when "0101111111111100", -- t[24572] = 6
      "000110" when "0101111111111101", -- t[24573] = 6
      "000110" when "0101111111111110", -- t[24574] = 6
      "000110" when "0101111111111111", -- t[24575] = 6
      "000110" when "0110000000000000", -- t[24576] = 6
      "000110" when "0110000000000001", -- t[24577] = 6
      "000110" when "0110000000000010", -- t[24578] = 6
      "000110" when "0110000000000011", -- t[24579] = 6
      "000110" when "0110000000000100", -- t[24580] = 6
      "000110" when "0110000000000101", -- t[24581] = 6
      "000110" when "0110000000000110", -- t[24582] = 6
      "000110" when "0110000000000111", -- t[24583] = 6
      "000110" when "0110000000001000", -- t[24584] = 6
      "000110" when "0110000000001001", -- t[24585] = 6
      "000110" when "0110000000001010", -- t[24586] = 6
      "000110" when "0110000000001011", -- t[24587] = 6
      "000110" when "0110000000001100", -- t[24588] = 6
      "000110" when "0110000000001101", -- t[24589] = 6
      "000110" when "0110000000001110", -- t[24590] = 6
      "000110" when "0110000000001111", -- t[24591] = 6
      "000110" when "0110000000010000", -- t[24592] = 6
      "000110" when "0110000000010001", -- t[24593] = 6
      "000110" when "0110000000010010", -- t[24594] = 6
      "000110" when "0110000000010011", -- t[24595] = 6
      "000110" when "0110000000010100", -- t[24596] = 6
      "000110" when "0110000000010101", -- t[24597] = 6
      "000110" when "0110000000010110", -- t[24598] = 6
      "000110" when "0110000000010111", -- t[24599] = 6
      "000110" when "0110000000011000", -- t[24600] = 6
      "000110" when "0110000000011001", -- t[24601] = 6
      "000110" when "0110000000011010", -- t[24602] = 6
      "000110" when "0110000000011011", -- t[24603] = 6
      "000110" when "0110000000011100", -- t[24604] = 6
      "000110" when "0110000000011101", -- t[24605] = 6
      "000110" when "0110000000011110", -- t[24606] = 6
      "000110" when "0110000000011111", -- t[24607] = 6
      "000110" when "0110000000100000", -- t[24608] = 6
      "000110" when "0110000000100001", -- t[24609] = 6
      "000110" when "0110000000100010", -- t[24610] = 6
      "000110" when "0110000000100011", -- t[24611] = 6
      "000110" when "0110000000100100", -- t[24612] = 6
      "000110" when "0110000000100101", -- t[24613] = 6
      "000110" when "0110000000100110", -- t[24614] = 6
      "000110" when "0110000000100111", -- t[24615] = 6
      "000110" when "0110000000101000", -- t[24616] = 6
      "000110" when "0110000000101001", -- t[24617] = 6
      "000110" when "0110000000101010", -- t[24618] = 6
      "000110" when "0110000000101011", -- t[24619] = 6
      "000110" when "0110000000101100", -- t[24620] = 6
      "000110" when "0110000000101101", -- t[24621] = 6
      "000110" when "0110000000101110", -- t[24622] = 6
      "000110" when "0110000000101111", -- t[24623] = 6
      "000110" when "0110000000110000", -- t[24624] = 6
      "000110" when "0110000000110001", -- t[24625] = 6
      "000110" when "0110000000110010", -- t[24626] = 6
      "000110" when "0110000000110011", -- t[24627] = 6
      "000110" when "0110000000110100", -- t[24628] = 6
      "000110" when "0110000000110101", -- t[24629] = 6
      "000110" when "0110000000110110", -- t[24630] = 6
      "000110" when "0110000000110111", -- t[24631] = 6
      "000110" when "0110000000111000", -- t[24632] = 6
      "000110" when "0110000000111001", -- t[24633] = 6
      "000110" when "0110000000111010", -- t[24634] = 6
      "000110" when "0110000000111011", -- t[24635] = 6
      "000110" when "0110000000111100", -- t[24636] = 6
      "000110" when "0110000000111101", -- t[24637] = 6
      "000110" when "0110000000111110", -- t[24638] = 6
      "000110" when "0110000000111111", -- t[24639] = 6
      "000110" when "0110000001000000", -- t[24640] = 6
      "000110" when "0110000001000001", -- t[24641] = 6
      "000110" when "0110000001000010", -- t[24642] = 6
      "000110" when "0110000001000011", -- t[24643] = 6
      "000110" when "0110000001000100", -- t[24644] = 6
      "000110" when "0110000001000101", -- t[24645] = 6
      "000110" when "0110000001000110", -- t[24646] = 6
      "000110" when "0110000001000111", -- t[24647] = 6
      "000110" when "0110000001001000", -- t[24648] = 6
      "000110" when "0110000001001001", -- t[24649] = 6
      "000110" when "0110000001001010", -- t[24650] = 6
      "000110" when "0110000001001011", -- t[24651] = 6
      "000110" when "0110000001001100", -- t[24652] = 6
      "000110" when "0110000001001101", -- t[24653] = 6
      "000110" when "0110000001001110", -- t[24654] = 6
      "000110" when "0110000001001111", -- t[24655] = 6
      "000110" when "0110000001010000", -- t[24656] = 6
      "000110" when "0110000001010001", -- t[24657] = 6
      "000110" when "0110000001010010", -- t[24658] = 6
      "000110" when "0110000001010011", -- t[24659] = 6
      "000110" when "0110000001010100", -- t[24660] = 6
      "000110" when "0110000001010101", -- t[24661] = 6
      "000110" when "0110000001010110", -- t[24662] = 6
      "000110" when "0110000001010111", -- t[24663] = 6
      "000110" when "0110000001011000", -- t[24664] = 6
      "000110" when "0110000001011001", -- t[24665] = 6
      "000110" when "0110000001011010", -- t[24666] = 6
      "000110" when "0110000001011011", -- t[24667] = 6
      "000110" when "0110000001011100", -- t[24668] = 6
      "000110" when "0110000001011101", -- t[24669] = 6
      "000110" when "0110000001011110", -- t[24670] = 6
      "000110" when "0110000001011111", -- t[24671] = 6
      "000110" when "0110000001100000", -- t[24672] = 6
      "000110" when "0110000001100001", -- t[24673] = 6
      "000110" when "0110000001100010", -- t[24674] = 6
      "000110" when "0110000001100011", -- t[24675] = 6
      "000110" when "0110000001100100", -- t[24676] = 6
      "000110" when "0110000001100101", -- t[24677] = 6
      "000110" when "0110000001100110", -- t[24678] = 6
      "000110" when "0110000001100111", -- t[24679] = 6
      "000110" when "0110000001101000", -- t[24680] = 6
      "000110" when "0110000001101001", -- t[24681] = 6
      "000110" when "0110000001101010", -- t[24682] = 6
      "000110" when "0110000001101011", -- t[24683] = 6
      "000110" when "0110000001101100", -- t[24684] = 6
      "000110" when "0110000001101101", -- t[24685] = 6
      "000110" when "0110000001101110", -- t[24686] = 6
      "000110" when "0110000001101111", -- t[24687] = 6
      "000110" when "0110000001110000", -- t[24688] = 6
      "000110" when "0110000001110001", -- t[24689] = 6
      "000110" when "0110000001110010", -- t[24690] = 6
      "000110" when "0110000001110011", -- t[24691] = 6
      "000110" when "0110000001110100", -- t[24692] = 6
      "000110" when "0110000001110101", -- t[24693] = 6
      "000110" when "0110000001110110", -- t[24694] = 6
      "000110" when "0110000001110111", -- t[24695] = 6
      "000110" when "0110000001111000", -- t[24696] = 6
      "000110" when "0110000001111001", -- t[24697] = 6
      "000110" when "0110000001111010", -- t[24698] = 6
      "000110" when "0110000001111011", -- t[24699] = 6
      "000110" when "0110000001111100", -- t[24700] = 6
      "000110" when "0110000001111101", -- t[24701] = 6
      "000110" when "0110000001111110", -- t[24702] = 6
      "000110" when "0110000001111111", -- t[24703] = 6
      "000110" when "0110000010000000", -- t[24704] = 6
      "000110" when "0110000010000001", -- t[24705] = 6
      "000110" when "0110000010000010", -- t[24706] = 6
      "000110" when "0110000010000011", -- t[24707] = 6
      "000110" when "0110000010000100", -- t[24708] = 6
      "000110" when "0110000010000101", -- t[24709] = 6
      "000110" when "0110000010000110", -- t[24710] = 6
      "000110" when "0110000010000111", -- t[24711] = 6
      "000110" when "0110000010001000", -- t[24712] = 6
      "000110" when "0110000010001001", -- t[24713] = 6
      "000110" when "0110000010001010", -- t[24714] = 6
      "000110" when "0110000010001011", -- t[24715] = 6
      "000110" when "0110000010001100", -- t[24716] = 6
      "000110" when "0110000010001101", -- t[24717] = 6
      "000110" when "0110000010001110", -- t[24718] = 6
      "000110" when "0110000010001111", -- t[24719] = 6
      "000110" when "0110000010010000", -- t[24720] = 6
      "000110" when "0110000010010001", -- t[24721] = 6
      "000110" when "0110000010010010", -- t[24722] = 6
      "000110" when "0110000010010011", -- t[24723] = 6
      "000110" when "0110000010010100", -- t[24724] = 6
      "000110" when "0110000010010101", -- t[24725] = 6
      "000110" when "0110000010010110", -- t[24726] = 6
      "000110" when "0110000010010111", -- t[24727] = 6
      "000110" when "0110000010011000", -- t[24728] = 6
      "000110" when "0110000010011001", -- t[24729] = 6
      "000110" when "0110000010011010", -- t[24730] = 6
      "000110" when "0110000010011011", -- t[24731] = 6
      "000110" when "0110000010011100", -- t[24732] = 6
      "000110" when "0110000010011101", -- t[24733] = 6
      "000110" when "0110000010011110", -- t[24734] = 6
      "000110" when "0110000010011111", -- t[24735] = 6
      "000110" when "0110000010100000", -- t[24736] = 6
      "000110" when "0110000010100001", -- t[24737] = 6
      "000110" when "0110000010100010", -- t[24738] = 6
      "000110" when "0110000010100011", -- t[24739] = 6
      "000110" when "0110000010100100", -- t[24740] = 6
      "000110" when "0110000010100101", -- t[24741] = 6
      "000110" when "0110000010100110", -- t[24742] = 6
      "000110" when "0110000010100111", -- t[24743] = 6
      "000110" when "0110000010101000", -- t[24744] = 6
      "000110" when "0110000010101001", -- t[24745] = 6
      "000110" when "0110000010101010", -- t[24746] = 6
      "000110" when "0110000010101011", -- t[24747] = 6
      "000110" when "0110000010101100", -- t[24748] = 6
      "000110" when "0110000010101101", -- t[24749] = 6
      "000110" when "0110000010101110", -- t[24750] = 6
      "000110" when "0110000010101111", -- t[24751] = 6
      "000110" when "0110000010110000", -- t[24752] = 6
      "000110" when "0110000010110001", -- t[24753] = 6
      "000110" when "0110000010110010", -- t[24754] = 6
      "000110" when "0110000010110011", -- t[24755] = 6
      "000110" when "0110000010110100", -- t[24756] = 6
      "000110" when "0110000010110101", -- t[24757] = 6
      "000110" when "0110000010110110", -- t[24758] = 6
      "000110" when "0110000010110111", -- t[24759] = 6
      "000110" when "0110000010111000", -- t[24760] = 6
      "000110" when "0110000010111001", -- t[24761] = 6
      "000110" when "0110000010111010", -- t[24762] = 6
      "000110" when "0110000010111011", -- t[24763] = 6
      "000110" when "0110000010111100", -- t[24764] = 6
      "000110" when "0110000010111101", -- t[24765] = 6
      "000110" when "0110000010111110", -- t[24766] = 6
      "000110" when "0110000010111111", -- t[24767] = 6
      "000110" when "0110000011000000", -- t[24768] = 6
      "000110" when "0110000011000001", -- t[24769] = 6
      "000110" when "0110000011000010", -- t[24770] = 6
      "000110" when "0110000011000011", -- t[24771] = 6
      "000110" when "0110000011000100", -- t[24772] = 6
      "000110" when "0110000011000101", -- t[24773] = 6
      "000110" when "0110000011000110", -- t[24774] = 6
      "000110" when "0110000011000111", -- t[24775] = 6
      "000110" when "0110000011001000", -- t[24776] = 6
      "000110" when "0110000011001001", -- t[24777] = 6
      "000110" when "0110000011001010", -- t[24778] = 6
      "000110" when "0110000011001011", -- t[24779] = 6
      "000110" when "0110000011001100", -- t[24780] = 6
      "000110" when "0110000011001101", -- t[24781] = 6
      "000110" when "0110000011001110", -- t[24782] = 6
      "000110" when "0110000011001111", -- t[24783] = 6
      "000110" when "0110000011010000", -- t[24784] = 6
      "000110" when "0110000011010001", -- t[24785] = 6
      "000110" when "0110000011010010", -- t[24786] = 6
      "000110" when "0110000011010011", -- t[24787] = 6
      "000110" when "0110000011010100", -- t[24788] = 6
      "000110" when "0110000011010101", -- t[24789] = 6
      "000110" when "0110000011010110", -- t[24790] = 6
      "000110" when "0110000011010111", -- t[24791] = 6
      "000110" when "0110000011011000", -- t[24792] = 6
      "000110" when "0110000011011001", -- t[24793] = 6
      "000110" when "0110000011011010", -- t[24794] = 6
      "000110" when "0110000011011011", -- t[24795] = 6
      "000110" when "0110000011011100", -- t[24796] = 6
      "000110" when "0110000011011101", -- t[24797] = 6
      "000110" when "0110000011011110", -- t[24798] = 6
      "000110" when "0110000011011111", -- t[24799] = 6
      "000110" when "0110000011100000", -- t[24800] = 6
      "000110" when "0110000011100001", -- t[24801] = 6
      "000110" when "0110000011100010", -- t[24802] = 6
      "000110" when "0110000011100011", -- t[24803] = 6
      "000110" when "0110000011100100", -- t[24804] = 6
      "000110" when "0110000011100101", -- t[24805] = 6
      "000110" when "0110000011100110", -- t[24806] = 6
      "000110" when "0110000011100111", -- t[24807] = 6
      "000110" when "0110000011101000", -- t[24808] = 6
      "000110" when "0110000011101001", -- t[24809] = 6
      "000110" when "0110000011101010", -- t[24810] = 6
      "000110" when "0110000011101011", -- t[24811] = 6
      "000110" when "0110000011101100", -- t[24812] = 6
      "000110" when "0110000011101101", -- t[24813] = 6
      "000110" when "0110000011101110", -- t[24814] = 6
      "000110" when "0110000011101111", -- t[24815] = 6
      "000110" when "0110000011110000", -- t[24816] = 6
      "000110" when "0110000011110001", -- t[24817] = 6
      "000110" when "0110000011110010", -- t[24818] = 6
      "000110" when "0110000011110011", -- t[24819] = 6
      "000110" when "0110000011110100", -- t[24820] = 6
      "000110" when "0110000011110101", -- t[24821] = 6
      "000110" when "0110000011110110", -- t[24822] = 6
      "000110" when "0110000011110111", -- t[24823] = 6
      "000110" when "0110000011111000", -- t[24824] = 6
      "000110" when "0110000011111001", -- t[24825] = 6
      "000110" when "0110000011111010", -- t[24826] = 6
      "000110" when "0110000011111011", -- t[24827] = 6
      "000110" when "0110000011111100", -- t[24828] = 6
      "000110" when "0110000011111101", -- t[24829] = 6
      "000110" when "0110000011111110", -- t[24830] = 6
      "000110" when "0110000011111111", -- t[24831] = 6
      "000110" when "0110000100000000", -- t[24832] = 6
      "000110" when "0110000100000001", -- t[24833] = 6
      "000110" when "0110000100000010", -- t[24834] = 6
      "000110" when "0110000100000011", -- t[24835] = 6
      "000110" when "0110000100000100", -- t[24836] = 6
      "000110" when "0110000100000101", -- t[24837] = 6
      "000110" when "0110000100000110", -- t[24838] = 6
      "000110" when "0110000100000111", -- t[24839] = 6
      "000110" when "0110000100001000", -- t[24840] = 6
      "000110" when "0110000100001001", -- t[24841] = 6
      "000110" when "0110000100001010", -- t[24842] = 6
      "000110" when "0110000100001011", -- t[24843] = 6
      "000110" when "0110000100001100", -- t[24844] = 6
      "000110" when "0110000100001101", -- t[24845] = 6
      "000110" when "0110000100001110", -- t[24846] = 6
      "000110" when "0110000100001111", -- t[24847] = 6
      "000110" when "0110000100010000", -- t[24848] = 6
      "000110" when "0110000100010001", -- t[24849] = 6
      "000110" when "0110000100010010", -- t[24850] = 6
      "000110" when "0110000100010011", -- t[24851] = 6
      "000110" when "0110000100010100", -- t[24852] = 6
      "000110" when "0110000100010101", -- t[24853] = 6
      "000110" when "0110000100010110", -- t[24854] = 6
      "000110" when "0110000100010111", -- t[24855] = 6
      "000110" when "0110000100011000", -- t[24856] = 6
      "000110" when "0110000100011001", -- t[24857] = 6
      "000110" when "0110000100011010", -- t[24858] = 6
      "000110" when "0110000100011011", -- t[24859] = 6
      "000110" when "0110000100011100", -- t[24860] = 6
      "000110" when "0110000100011101", -- t[24861] = 6
      "000110" when "0110000100011110", -- t[24862] = 6
      "000110" when "0110000100011111", -- t[24863] = 6
      "000110" when "0110000100100000", -- t[24864] = 6
      "000110" when "0110000100100001", -- t[24865] = 6
      "000110" when "0110000100100010", -- t[24866] = 6
      "000110" when "0110000100100011", -- t[24867] = 6
      "000110" when "0110000100100100", -- t[24868] = 6
      "000110" when "0110000100100101", -- t[24869] = 6
      "000110" when "0110000100100110", -- t[24870] = 6
      "000110" when "0110000100100111", -- t[24871] = 6
      "000110" when "0110000100101000", -- t[24872] = 6
      "000110" when "0110000100101001", -- t[24873] = 6
      "000110" when "0110000100101010", -- t[24874] = 6
      "000110" when "0110000100101011", -- t[24875] = 6
      "000110" when "0110000100101100", -- t[24876] = 6
      "000110" when "0110000100101101", -- t[24877] = 6
      "000110" when "0110000100101110", -- t[24878] = 6
      "000110" when "0110000100101111", -- t[24879] = 6
      "000110" when "0110000100110000", -- t[24880] = 6
      "000110" when "0110000100110001", -- t[24881] = 6
      "000110" when "0110000100110010", -- t[24882] = 6
      "000110" when "0110000100110011", -- t[24883] = 6
      "000110" when "0110000100110100", -- t[24884] = 6
      "000110" when "0110000100110101", -- t[24885] = 6
      "000110" when "0110000100110110", -- t[24886] = 6
      "000110" when "0110000100110111", -- t[24887] = 6
      "000110" when "0110000100111000", -- t[24888] = 6
      "000110" when "0110000100111001", -- t[24889] = 6
      "000110" when "0110000100111010", -- t[24890] = 6
      "000110" when "0110000100111011", -- t[24891] = 6
      "000110" when "0110000100111100", -- t[24892] = 6
      "000110" when "0110000100111101", -- t[24893] = 6
      "000110" when "0110000100111110", -- t[24894] = 6
      "000110" when "0110000100111111", -- t[24895] = 6
      "000110" when "0110000101000000", -- t[24896] = 6
      "000110" when "0110000101000001", -- t[24897] = 6
      "000110" when "0110000101000010", -- t[24898] = 6
      "000110" when "0110000101000011", -- t[24899] = 6
      "000110" when "0110000101000100", -- t[24900] = 6
      "000110" when "0110000101000101", -- t[24901] = 6
      "000110" when "0110000101000110", -- t[24902] = 6
      "000110" when "0110000101000111", -- t[24903] = 6
      "000110" when "0110000101001000", -- t[24904] = 6
      "000110" when "0110000101001001", -- t[24905] = 6
      "000110" when "0110000101001010", -- t[24906] = 6
      "000110" when "0110000101001011", -- t[24907] = 6
      "000110" when "0110000101001100", -- t[24908] = 6
      "000110" when "0110000101001101", -- t[24909] = 6
      "000110" when "0110000101001110", -- t[24910] = 6
      "000110" when "0110000101001111", -- t[24911] = 6
      "000110" when "0110000101010000", -- t[24912] = 6
      "000110" when "0110000101010001", -- t[24913] = 6
      "000110" when "0110000101010010", -- t[24914] = 6
      "000110" when "0110000101010011", -- t[24915] = 6
      "000110" when "0110000101010100", -- t[24916] = 6
      "000110" when "0110000101010101", -- t[24917] = 6
      "000110" when "0110000101010110", -- t[24918] = 6
      "000110" when "0110000101010111", -- t[24919] = 6
      "000110" when "0110000101011000", -- t[24920] = 6
      "000110" when "0110000101011001", -- t[24921] = 6
      "000110" when "0110000101011010", -- t[24922] = 6
      "000110" when "0110000101011011", -- t[24923] = 6
      "000110" when "0110000101011100", -- t[24924] = 6
      "000110" when "0110000101011101", -- t[24925] = 6
      "000110" when "0110000101011110", -- t[24926] = 6
      "000110" when "0110000101011111", -- t[24927] = 6
      "000110" when "0110000101100000", -- t[24928] = 6
      "000110" when "0110000101100001", -- t[24929] = 6
      "000110" when "0110000101100010", -- t[24930] = 6
      "000110" when "0110000101100011", -- t[24931] = 6
      "000110" when "0110000101100100", -- t[24932] = 6
      "000110" when "0110000101100101", -- t[24933] = 6
      "000110" when "0110000101100110", -- t[24934] = 6
      "000110" when "0110000101100111", -- t[24935] = 6
      "000110" when "0110000101101000", -- t[24936] = 6
      "000110" when "0110000101101001", -- t[24937] = 6
      "000110" when "0110000101101010", -- t[24938] = 6
      "000110" when "0110000101101011", -- t[24939] = 6
      "000110" when "0110000101101100", -- t[24940] = 6
      "000110" when "0110000101101101", -- t[24941] = 6
      "000110" when "0110000101101110", -- t[24942] = 6
      "000110" when "0110000101101111", -- t[24943] = 6
      "000110" when "0110000101110000", -- t[24944] = 6
      "000110" when "0110000101110001", -- t[24945] = 6
      "000110" when "0110000101110010", -- t[24946] = 6
      "000110" when "0110000101110011", -- t[24947] = 6
      "000110" when "0110000101110100", -- t[24948] = 6
      "000110" when "0110000101110101", -- t[24949] = 6
      "000110" when "0110000101110110", -- t[24950] = 6
      "000110" when "0110000101110111", -- t[24951] = 6
      "000110" when "0110000101111000", -- t[24952] = 6
      "000110" when "0110000101111001", -- t[24953] = 6
      "000110" when "0110000101111010", -- t[24954] = 6
      "000110" when "0110000101111011", -- t[24955] = 6
      "000110" when "0110000101111100", -- t[24956] = 6
      "000110" when "0110000101111101", -- t[24957] = 6
      "000110" when "0110000101111110", -- t[24958] = 6
      "000110" when "0110000101111111", -- t[24959] = 6
      "000110" when "0110000110000000", -- t[24960] = 6
      "000110" when "0110000110000001", -- t[24961] = 6
      "000110" when "0110000110000010", -- t[24962] = 6
      "000110" when "0110000110000011", -- t[24963] = 6
      "000110" when "0110000110000100", -- t[24964] = 6
      "000110" when "0110000110000101", -- t[24965] = 6
      "000110" when "0110000110000110", -- t[24966] = 6
      "000110" when "0110000110000111", -- t[24967] = 6
      "000110" when "0110000110001000", -- t[24968] = 6
      "000110" when "0110000110001001", -- t[24969] = 6
      "000110" when "0110000110001010", -- t[24970] = 6
      "000110" when "0110000110001011", -- t[24971] = 6
      "000110" when "0110000110001100", -- t[24972] = 6
      "000110" when "0110000110001101", -- t[24973] = 6
      "000110" when "0110000110001110", -- t[24974] = 6
      "000110" when "0110000110001111", -- t[24975] = 6
      "000110" when "0110000110010000", -- t[24976] = 6
      "000110" when "0110000110010001", -- t[24977] = 6
      "000110" when "0110000110010010", -- t[24978] = 6
      "000110" when "0110000110010011", -- t[24979] = 6
      "000110" when "0110000110010100", -- t[24980] = 6
      "000110" when "0110000110010101", -- t[24981] = 6
      "000110" when "0110000110010110", -- t[24982] = 6
      "000110" when "0110000110010111", -- t[24983] = 6
      "000110" when "0110000110011000", -- t[24984] = 6
      "000110" when "0110000110011001", -- t[24985] = 6
      "000110" when "0110000110011010", -- t[24986] = 6
      "000110" when "0110000110011011", -- t[24987] = 6
      "000110" when "0110000110011100", -- t[24988] = 6
      "000110" when "0110000110011101", -- t[24989] = 6
      "000110" when "0110000110011110", -- t[24990] = 6
      "000110" when "0110000110011111", -- t[24991] = 6
      "000110" when "0110000110100000", -- t[24992] = 6
      "000110" when "0110000110100001", -- t[24993] = 6
      "000110" when "0110000110100010", -- t[24994] = 6
      "000110" when "0110000110100011", -- t[24995] = 6
      "000110" when "0110000110100100", -- t[24996] = 6
      "000110" when "0110000110100101", -- t[24997] = 6
      "000110" when "0110000110100110", -- t[24998] = 6
      "000110" when "0110000110100111", -- t[24999] = 6
      "000110" when "0110000110101000", -- t[25000] = 6
      "000110" when "0110000110101001", -- t[25001] = 6
      "000110" when "0110000110101010", -- t[25002] = 6
      "000110" when "0110000110101011", -- t[25003] = 6
      "000110" when "0110000110101100", -- t[25004] = 6
      "000110" when "0110000110101101", -- t[25005] = 6
      "000110" when "0110000110101110", -- t[25006] = 6
      "000110" when "0110000110101111", -- t[25007] = 6
      "000110" when "0110000110110000", -- t[25008] = 6
      "000110" when "0110000110110001", -- t[25009] = 6
      "000110" when "0110000110110010", -- t[25010] = 6
      "000110" when "0110000110110011", -- t[25011] = 6
      "000110" when "0110000110110100", -- t[25012] = 6
      "000110" when "0110000110110101", -- t[25013] = 6
      "000110" when "0110000110110110", -- t[25014] = 6
      "000110" when "0110000110110111", -- t[25015] = 6
      "000110" when "0110000110111000", -- t[25016] = 6
      "000110" when "0110000110111001", -- t[25017] = 6
      "000110" when "0110000110111010", -- t[25018] = 6
      "000110" when "0110000110111011", -- t[25019] = 6
      "000110" when "0110000110111100", -- t[25020] = 6
      "000110" when "0110000110111101", -- t[25021] = 6
      "000110" when "0110000110111110", -- t[25022] = 6
      "000110" when "0110000110111111", -- t[25023] = 6
      "000110" when "0110000111000000", -- t[25024] = 6
      "000110" when "0110000111000001", -- t[25025] = 6
      "000110" when "0110000111000010", -- t[25026] = 6
      "000110" when "0110000111000011", -- t[25027] = 6
      "000110" when "0110000111000100", -- t[25028] = 6
      "000110" when "0110000111000101", -- t[25029] = 6
      "000110" when "0110000111000110", -- t[25030] = 6
      "000110" when "0110000111000111", -- t[25031] = 6
      "000110" when "0110000111001000", -- t[25032] = 6
      "000110" when "0110000111001001", -- t[25033] = 6
      "000110" when "0110000111001010", -- t[25034] = 6
      "000110" when "0110000111001011", -- t[25035] = 6
      "000110" when "0110000111001100", -- t[25036] = 6
      "000110" when "0110000111001101", -- t[25037] = 6
      "000110" when "0110000111001110", -- t[25038] = 6
      "000110" when "0110000111001111", -- t[25039] = 6
      "000110" when "0110000111010000", -- t[25040] = 6
      "000110" when "0110000111010001", -- t[25041] = 6
      "000110" when "0110000111010010", -- t[25042] = 6
      "000110" when "0110000111010011", -- t[25043] = 6
      "000110" when "0110000111010100", -- t[25044] = 6
      "000110" when "0110000111010101", -- t[25045] = 6
      "000110" when "0110000111010110", -- t[25046] = 6
      "000110" when "0110000111010111", -- t[25047] = 6
      "000110" when "0110000111011000", -- t[25048] = 6
      "000110" when "0110000111011001", -- t[25049] = 6
      "000110" when "0110000111011010", -- t[25050] = 6
      "000110" when "0110000111011011", -- t[25051] = 6
      "000110" when "0110000111011100", -- t[25052] = 6
      "000110" when "0110000111011101", -- t[25053] = 6
      "000110" when "0110000111011110", -- t[25054] = 6
      "000110" when "0110000111011111", -- t[25055] = 6
      "000110" when "0110000111100000", -- t[25056] = 6
      "000110" when "0110000111100001", -- t[25057] = 6
      "000110" when "0110000111100010", -- t[25058] = 6
      "000110" when "0110000111100011", -- t[25059] = 6
      "000110" when "0110000111100100", -- t[25060] = 6
      "000110" when "0110000111100101", -- t[25061] = 6
      "000110" when "0110000111100110", -- t[25062] = 6
      "000110" when "0110000111100111", -- t[25063] = 6
      "000110" when "0110000111101000", -- t[25064] = 6
      "000110" when "0110000111101001", -- t[25065] = 6
      "000110" when "0110000111101010", -- t[25066] = 6
      "000110" when "0110000111101011", -- t[25067] = 6
      "000110" when "0110000111101100", -- t[25068] = 6
      "000110" when "0110000111101101", -- t[25069] = 6
      "000110" when "0110000111101110", -- t[25070] = 6
      "000110" when "0110000111101111", -- t[25071] = 6
      "000110" when "0110000111110000", -- t[25072] = 6
      "000110" when "0110000111110001", -- t[25073] = 6
      "000110" when "0110000111110010", -- t[25074] = 6
      "000110" when "0110000111110011", -- t[25075] = 6
      "000110" when "0110000111110100", -- t[25076] = 6
      "000110" when "0110000111110101", -- t[25077] = 6
      "000110" when "0110000111110110", -- t[25078] = 6
      "000110" when "0110000111110111", -- t[25079] = 6
      "000110" when "0110000111111000", -- t[25080] = 6
      "000110" when "0110000111111001", -- t[25081] = 6
      "000110" when "0110000111111010", -- t[25082] = 6
      "000110" when "0110000111111011", -- t[25083] = 6
      "000110" when "0110000111111100", -- t[25084] = 6
      "000110" when "0110000111111101", -- t[25085] = 6
      "000110" when "0110000111111110", -- t[25086] = 6
      "000110" when "0110000111111111", -- t[25087] = 6
      "000110" when "0110001000000000", -- t[25088] = 6
      "000110" when "0110001000000001", -- t[25089] = 6
      "000110" when "0110001000000010", -- t[25090] = 6
      "000110" when "0110001000000011", -- t[25091] = 6
      "000110" when "0110001000000100", -- t[25092] = 6
      "000110" when "0110001000000101", -- t[25093] = 6
      "000110" when "0110001000000110", -- t[25094] = 6
      "000110" when "0110001000000111", -- t[25095] = 6
      "000110" when "0110001000001000", -- t[25096] = 6
      "000110" when "0110001000001001", -- t[25097] = 6
      "000110" when "0110001000001010", -- t[25098] = 6
      "000110" when "0110001000001011", -- t[25099] = 6
      "000110" when "0110001000001100", -- t[25100] = 6
      "000110" when "0110001000001101", -- t[25101] = 6
      "000110" when "0110001000001110", -- t[25102] = 6
      "000110" when "0110001000001111", -- t[25103] = 6
      "000110" when "0110001000010000", -- t[25104] = 6
      "000110" when "0110001000010001", -- t[25105] = 6
      "000110" when "0110001000010010", -- t[25106] = 6
      "000110" when "0110001000010011", -- t[25107] = 6
      "000110" when "0110001000010100", -- t[25108] = 6
      "000110" when "0110001000010101", -- t[25109] = 6
      "000110" when "0110001000010110", -- t[25110] = 6
      "000110" when "0110001000010111", -- t[25111] = 6
      "000110" when "0110001000011000", -- t[25112] = 6
      "000110" when "0110001000011001", -- t[25113] = 6
      "000110" when "0110001000011010", -- t[25114] = 6
      "000110" when "0110001000011011", -- t[25115] = 6
      "000110" when "0110001000011100", -- t[25116] = 6
      "000110" when "0110001000011101", -- t[25117] = 6
      "000110" when "0110001000011110", -- t[25118] = 6
      "000110" when "0110001000011111", -- t[25119] = 6
      "000110" when "0110001000100000", -- t[25120] = 6
      "000110" when "0110001000100001", -- t[25121] = 6
      "000110" when "0110001000100010", -- t[25122] = 6
      "000110" when "0110001000100011", -- t[25123] = 6
      "000110" when "0110001000100100", -- t[25124] = 6
      "000110" when "0110001000100101", -- t[25125] = 6
      "000110" when "0110001000100110", -- t[25126] = 6
      "000110" when "0110001000100111", -- t[25127] = 6
      "000110" when "0110001000101000", -- t[25128] = 6
      "000110" when "0110001000101001", -- t[25129] = 6
      "000110" when "0110001000101010", -- t[25130] = 6
      "000110" when "0110001000101011", -- t[25131] = 6
      "000110" when "0110001000101100", -- t[25132] = 6
      "000110" when "0110001000101101", -- t[25133] = 6
      "000110" when "0110001000101110", -- t[25134] = 6
      "000110" when "0110001000101111", -- t[25135] = 6
      "000110" when "0110001000110000", -- t[25136] = 6
      "000110" when "0110001000110001", -- t[25137] = 6
      "000110" when "0110001000110010", -- t[25138] = 6
      "000110" when "0110001000110011", -- t[25139] = 6
      "000110" when "0110001000110100", -- t[25140] = 6
      "000110" when "0110001000110101", -- t[25141] = 6
      "000110" when "0110001000110110", -- t[25142] = 6
      "000110" when "0110001000110111", -- t[25143] = 6
      "000110" when "0110001000111000", -- t[25144] = 6
      "000110" when "0110001000111001", -- t[25145] = 6
      "000110" when "0110001000111010", -- t[25146] = 6
      "000110" when "0110001000111011", -- t[25147] = 6
      "000110" when "0110001000111100", -- t[25148] = 6
      "000110" when "0110001000111101", -- t[25149] = 6
      "000110" when "0110001000111110", -- t[25150] = 6
      "000110" when "0110001000111111", -- t[25151] = 6
      "000110" when "0110001001000000", -- t[25152] = 6
      "000110" when "0110001001000001", -- t[25153] = 6
      "000110" when "0110001001000010", -- t[25154] = 6
      "000110" when "0110001001000011", -- t[25155] = 6
      "000110" when "0110001001000100", -- t[25156] = 6
      "000110" when "0110001001000101", -- t[25157] = 6
      "000110" when "0110001001000110", -- t[25158] = 6
      "000110" when "0110001001000111", -- t[25159] = 6
      "000110" when "0110001001001000", -- t[25160] = 6
      "000110" when "0110001001001001", -- t[25161] = 6
      "000110" when "0110001001001010", -- t[25162] = 6
      "000110" when "0110001001001011", -- t[25163] = 6
      "000110" when "0110001001001100", -- t[25164] = 6
      "000110" when "0110001001001101", -- t[25165] = 6
      "000110" when "0110001001001110", -- t[25166] = 6
      "000110" when "0110001001001111", -- t[25167] = 6
      "000110" when "0110001001010000", -- t[25168] = 6
      "000110" when "0110001001010001", -- t[25169] = 6
      "000110" when "0110001001010010", -- t[25170] = 6
      "000110" when "0110001001010011", -- t[25171] = 6
      "000110" when "0110001001010100", -- t[25172] = 6
      "000110" when "0110001001010101", -- t[25173] = 6
      "000110" when "0110001001010110", -- t[25174] = 6
      "000110" when "0110001001010111", -- t[25175] = 6
      "000110" when "0110001001011000", -- t[25176] = 6
      "000110" when "0110001001011001", -- t[25177] = 6
      "000110" when "0110001001011010", -- t[25178] = 6
      "000110" when "0110001001011011", -- t[25179] = 6
      "000110" when "0110001001011100", -- t[25180] = 6
      "000110" when "0110001001011101", -- t[25181] = 6
      "000110" when "0110001001011110", -- t[25182] = 6
      "000110" when "0110001001011111", -- t[25183] = 6
      "000110" when "0110001001100000", -- t[25184] = 6
      "000110" when "0110001001100001", -- t[25185] = 6
      "000110" when "0110001001100010", -- t[25186] = 6
      "000110" when "0110001001100011", -- t[25187] = 6
      "000110" when "0110001001100100", -- t[25188] = 6
      "000110" when "0110001001100101", -- t[25189] = 6
      "000110" when "0110001001100110", -- t[25190] = 6
      "000110" when "0110001001100111", -- t[25191] = 6
      "000110" when "0110001001101000", -- t[25192] = 6
      "000110" when "0110001001101001", -- t[25193] = 6
      "000110" when "0110001001101010", -- t[25194] = 6
      "000110" when "0110001001101011", -- t[25195] = 6
      "000110" when "0110001001101100", -- t[25196] = 6
      "000110" when "0110001001101101", -- t[25197] = 6
      "000110" when "0110001001101110", -- t[25198] = 6
      "000110" when "0110001001101111", -- t[25199] = 6
      "000110" when "0110001001110000", -- t[25200] = 6
      "000110" when "0110001001110001", -- t[25201] = 6
      "000110" when "0110001001110010", -- t[25202] = 6
      "000110" when "0110001001110011", -- t[25203] = 6
      "000110" when "0110001001110100", -- t[25204] = 6
      "000110" when "0110001001110101", -- t[25205] = 6
      "000110" when "0110001001110110", -- t[25206] = 6
      "000110" when "0110001001110111", -- t[25207] = 6
      "000110" when "0110001001111000", -- t[25208] = 6
      "000110" when "0110001001111001", -- t[25209] = 6
      "000110" when "0110001001111010", -- t[25210] = 6
      "000110" when "0110001001111011", -- t[25211] = 6
      "000110" when "0110001001111100", -- t[25212] = 6
      "000110" when "0110001001111101", -- t[25213] = 6
      "000110" when "0110001001111110", -- t[25214] = 6
      "000110" when "0110001001111111", -- t[25215] = 6
      "000110" when "0110001010000000", -- t[25216] = 6
      "000110" when "0110001010000001", -- t[25217] = 6
      "000110" when "0110001010000010", -- t[25218] = 6
      "000110" when "0110001010000011", -- t[25219] = 6
      "000110" when "0110001010000100", -- t[25220] = 6
      "000110" when "0110001010000101", -- t[25221] = 6
      "000110" when "0110001010000110", -- t[25222] = 6
      "000110" when "0110001010000111", -- t[25223] = 6
      "000110" when "0110001010001000", -- t[25224] = 6
      "000110" when "0110001010001001", -- t[25225] = 6
      "000110" when "0110001010001010", -- t[25226] = 6
      "000110" when "0110001010001011", -- t[25227] = 6
      "000110" when "0110001010001100", -- t[25228] = 6
      "000110" when "0110001010001101", -- t[25229] = 6
      "000110" when "0110001010001110", -- t[25230] = 6
      "000110" when "0110001010001111", -- t[25231] = 6
      "000110" when "0110001010010000", -- t[25232] = 6
      "000110" when "0110001010010001", -- t[25233] = 6
      "000110" when "0110001010010010", -- t[25234] = 6
      "000110" when "0110001010010011", -- t[25235] = 6
      "000110" when "0110001010010100", -- t[25236] = 6
      "000110" when "0110001010010101", -- t[25237] = 6
      "000110" when "0110001010010110", -- t[25238] = 6
      "000110" when "0110001010010111", -- t[25239] = 6
      "000110" when "0110001010011000", -- t[25240] = 6
      "000110" when "0110001010011001", -- t[25241] = 6
      "000110" when "0110001010011010", -- t[25242] = 6
      "000110" when "0110001010011011", -- t[25243] = 6
      "000110" when "0110001010011100", -- t[25244] = 6
      "000110" when "0110001010011101", -- t[25245] = 6
      "000110" when "0110001010011110", -- t[25246] = 6
      "000110" when "0110001010011111", -- t[25247] = 6
      "000110" when "0110001010100000", -- t[25248] = 6
      "000110" when "0110001010100001", -- t[25249] = 6
      "000110" when "0110001010100010", -- t[25250] = 6
      "000110" when "0110001010100011", -- t[25251] = 6
      "000110" when "0110001010100100", -- t[25252] = 6
      "000110" when "0110001010100101", -- t[25253] = 6
      "000110" when "0110001010100110", -- t[25254] = 6
      "000110" when "0110001010100111", -- t[25255] = 6
      "000110" when "0110001010101000", -- t[25256] = 6
      "000110" when "0110001010101001", -- t[25257] = 6
      "000110" when "0110001010101010", -- t[25258] = 6
      "000110" when "0110001010101011", -- t[25259] = 6
      "000110" when "0110001010101100", -- t[25260] = 6
      "000110" when "0110001010101101", -- t[25261] = 6
      "000110" when "0110001010101110", -- t[25262] = 6
      "000110" when "0110001010101111", -- t[25263] = 6
      "000110" when "0110001010110000", -- t[25264] = 6
      "000110" when "0110001010110001", -- t[25265] = 6
      "000110" when "0110001010110010", -- t[25266] = 6
      "000110" when "0110001010110011", -- t[25267] = 6
      "000110" when "0110001010110100", -- t[25268] = 6
      "000110" when "0110001010110101", -- t[25269] = 6
      "000110" when "0110001010110110", -- t[25270] = 6
      "000110" when "0110001010110111", -- t[25271] = 6
      "000110" when "0110001010111000", -- t[25272] = 6
      "000110" when "0110001010111001", -- t[25273] = 6
      "000110" when "0110001010111010", -- t[25274] = 6
      "000110" when "0110001010111011", -- t[25275] = 6
      "000111" when "0110001010111100", -- t[25276] = 7
      "000111" when "0110001010111101", -- t[25277] = 7
      "000111" when "0110001010111110", -- t[25278] = 7
      "000111" when "0110001010111111", -- t[25279] = 7
      "000111" when "0110001011000000", -- t[25280] = 7
      "000111" when "0110001011000001", -- t[25281] = 7
      "000111" when "0110001011000010", -- t[25282] = 7
      "000111" when "0110001011000011", -- t[25283] = 7
      "000111" when "0110001011000100", -- t[25284] = 7
      "000111" when "0110001011000101", -- t[25285] = 7
      "000111" when "0110001011000110", -- t[25286] = 7
      "000111" when "0110001011000111", -- t[25287] = 7
      "000111" when "0110001011001000", -- t[25288] = 7
      "000111" when "0110001011001001", -- t[25289] = 7
      "000111" when "0110001011001010", -- t[25290] = 7
      "000111" when "0110001011001011", -- t[25291] = 7
      "000111" when "0110001011001100", -- t[25292] = 7
      "000111" when "0110001011001101", -- t[25293] = 7
      "000111" when "0110001011001110", -- t[25294] = 7
      "000111" when "0110001011001111", -- t[25295] = 7
      "000111" when "0110001011010000", -- t[25296] = 7
      "000111" when "0110001011010001", -- t[25297] = 7
      "000111" when "0110001011010010", -- t[25298] = 7
      "000111" when "0110001011010011", -- t[25299] = 7
      "000111" when "0110001011010100", -- t[25300] = 7
      "000111" when "0110001011010101", -- t[25301] = 7
      "000111" when "0110001011010110", -- t[25302] = 7
      "000111" when "0110001011010111", -- t[25303] = 7
      "000111" when "0110001011011000", -- t[25304] = 7
      "000111" when "0110001011011001", -- t[25305] = 7
      "000111" when "0110001011011010", -- t[25306] = 7
      "000111" when "0110001011011011", -- t[25307] = 7
      "000111" when "0110001011011100", -- t[25308] = 7
      "000111" when "0110001011011101", -- t[25309] = 7
      "000111" when "0110001011011110", -- t[25310] = 7
      "000111" when "0110001011011111", -- t[25311] = 7
      "000111" when "0110001011100000", -- t[25312] = 7
      "000111" when "0110001011100001", -- t[25313] = 7
      "000111" when "0110001011100010", -- t[25314] = 7
      "000111" when "0110001011100011", -- t[25315] = 7
      "000111" when "0110001011100100", -- t[25316] = 7
      "000111" when "0110001011100101", -- t[25317] = 7
      "000111" when "0110001011100110", -- t[25318] = 7
      "000111" when "0110001011100111", -- t[25319] = 7
      "000111" when "0110001011101000", -- t[25320] = 7
      "000111" when "0110001011101001", -- t[25321] = 7
      "000111" when "0110001011101010", -- t[25322] = 7
      "000111" when "0110001011101011", -- t[25323] = 7
      "000111" when "0110001011101100", -- t[25324] = 7
      "000111" when "0110001011101101", -- t[25325] = 7
      "000111" when "0110001011101110", -- t[25326] = 7
      "000111" when "0110001011101111", -- t[25327] = 7
      "000111" when "0110001011110000", -- t[25328] = 7
      "000111" when "0110001011110001", -- t[25329] = 7
      "000111" when "0110001011110010", -- t[25330] = 7
      "000111" when "0110001011110011", -- t[25331] = 7
      "000111" when "0110001011110100", -- t[25332] = 7
      "000111" when "0110001011110101", -- t[25333] = 7
      "000111" when "0110001011110110", -- t[25334] = 7
      "000111" when "0110001011110111", -- t[25335] = 7
      "000111" when "0110001011111000", -- t[25336] = 7
      "000111" when "0110001011111001", -- t[25337] = 7
      "000111" when "0110001011111010", -- t[25338] = 7
      "000111" when "0110001011111011", -- t[25339] = 7
      "000111" when "0110001011111100", -- t[25340] = 7
      "000111" when "0110001011111101", -- t[25341] = 7
      "000111" when "0110001011111110", -- t[25342] = 7
      "000111" when "0110001011111111", -- t[25343] = 7
      "000111" when "0110001100000000", -- t[25344] = 7
      "000111" when "0110001100000001", -- t[25345] = 7
      "000111" when "0110001100000010", -- t[25346] = 7
      "000111" when "0110001100000011", -- t[25347] = 7
      "000111" when "0110001100000100", -- t[25348] = 7
      "000111" when "0110001100000101", -- t[25349] = 7
      "000111" when "0110001100000110", -- t[25350] = 7
      "000111" when "0110001100000111", -- t[25351] = 7
      "000111" when "0110001100001000", -- t[25352] = 7
      "000111" when "0110001100001001", -- t[25353] = 7
      "000111" when "0110001100001010", -- t[25354] = 7
      "000111" when "0110001100001011", -- t[25355] = 7
      "000111" when "0110001100001100", -- t[25356] = 7
      "000111" when "0110001100001101", -- t[25357] = 7
      "000111" when "0110001100001110", -- t[25358] = 7
      "000111" when "0110001100001111", -- t[25359] = 7
      "000111" when "0110001100010000", -- t[25360] = 7
      "000111" when "0110001100010001", -- t[25361] = 7
      "000111" when "0110001100010010", -- t[25362] = 7
      "000111" when "0110001100010011", -- t[25363] = 7
      "000111" when "0110001100010100", -- t[25364] = 7
      "000111" when "0110001100010101", -- t[25365] = 7
      "000111" when "0110001100010110", -- t[25366] = 7
      "000111" when "0110001100010111", -- t[25367] = 7
      "000111" when "0110001100011000", -- t[25368] = 7
      "000111" when "0110001100011001", -- t[25369] = 7
      "000111" when "0110001100011010", -- t[25370] = 7
      "000111" when "0110001100011011", -- t[25371] = 7
      "000111" when "0110001100011100", -- t[25372] = 7
      "000111" when "0110001100011101", -- t[25373] = 7
      "000111" when "0110001100011110", -- t[25374] = 7
      "000111" when "0110001100011111", -- t[25375] = 7
      "000111" when "0110001100100000", -- t[25376] = 7
      "000111" when "0110001100100001", -- t[25377] = 7
      "000111" when "0110001100100010", -- t[25378] = 7
      "000111" when "0110001100100011", -- t[25379] = 7
      "000111" when "0110001100100100", -- t[25380] = 7
      "000111" when "0110001100100101", -- t[25381] = 7
      "000111" when "0110001100100110", -- t[25382] = 7
      "000111" when "0110001100100111", -- t[25383] = 7
      "000111" when "0110001100101000", -- t[25384] = 7
      "000111" when "0110001100101001", -- t[25385] = 7
      "000111" when "0110001100101010", -- t[25386] = 7
      "000111" when "0110001100101011", -- t[25387] = 7
      "000111" when "0110001100101100", -- t[25388] = 7
      "000111" when "0110001100101101", -- t[25389] = 7
      "000111" when "0110001100101110", -- t[25390] = 7
      "000111" when "0110001100101111", -- t[25391] = 7
      "000111" when "0110001100110000", -- t[25392] = 7
      "000111" when "0110001100110001", -- t[25393] = 7
      "000111" when "0110001100110010", -- t[25394] = 7
      "000111" when "0110001100110011", -- t[25395] = 7
      "000111" when "0110001100110100", -- t[25396] = 7
      "000111" when "0110001100110101", -- t[25397] = 7
      "000111" when "0110001100110110", -- t[25398] = 7
      "000111" when "0110001100110111", -- t[25399] = 7
      "000111" when "0110001100111000", -- t[25400] = 7
      "000111" when "0110001100111001", -- t[25401] = 7
      "000111" when "0110001100111010", -- t[25402] = 7
      "000111" when "0110001100111011", -- t[25403] = 7
      "000111" when "0110001100111100", -- t[25404] = 7
      "000111" when "0110001100111101", -- t[25405] = 7
      "000111" when "0110001100111110", -- t[25406] = 7
      "000111" when "0110001100111111", -- t[25407] = 7
      "000111" when "0110001101000000", -- t[25408] = 7
      "000111" when "0110001101000001", -- t[25409] = 7
      "000111" when "0110001101000010", -- t[25410] = 7
      "000111" when "0110001101000011", -- t[25411] = 7
      "000111" when "0110001101000100", -- t[25412] = 7
      "000111" when "0110001101000101", -- t[25413] = 7
      "000111" when "0110001101000110", -- t[25414] = 7
      "000111" when "0110001101000111", -- t[25415] = 7
      "000111" when "0110001101001000", -- t[25416] = 7
      "000111" when "0110001101001001", -- t[25417] = 7
      "000111" when "0110001101001010", -- t[25418] = 7
      "000111" when "0110001101001011", -- t[25419] = 7
      "000111" when "0110001101001100", -- t[25420] = 7
      "000111" when "0110001101001101", -- t[25421] = 7
      "000111" when "0110001101001110", -- t[25422] = 7
      "000111" when "0110001101001111", -- t[25423] = 7
      "000111" when "0110001101010000", -- t[25424] = 7
      "000111" when "0110001101010001", -- t[25425] = 7
      "000111" when "0110001101010010", -- t[25426] = 7
      "000111" when "0110001101010011", -- t[25427] = 7
      "000111" when "0110001101010100", -- t[25428] = 7
      "000111" when "0110001101010101", -- t[25429] = 7
      "000111" when "0110001101010110", -- t[25430] = 7
      "000111" when "0110001101010111", -- t[25431] = 7
      "000111" when "0110001101011000", -- t[25432] = 7
      "000111" when "0110001101011001", -- t[25433] = 7
      "000111" when "0110001101011010", -- t[25434] = 7
      "000111" when "0110001101011011", -- t[25435] = 7
      "000111" when "0110001101011100", -- t[25436] = 7
      "000111" when "0110001101011101", -- t[25437] = 7
      "000111" when "0110001101011110", -- t[25438] = 7
      "000111" when "0110001101011111", -- t[25439] = 7
      "000111" when "0110001101100000", -- t[25440] = 7
      "000111" when "0110001101100001", -- t[25441] = 7
      "000111" when "0110001101100010", -- t[25442] = 7
      "000111" when "0110001101100011", -- t[25443] = 7
      "000111" when "0110001101100100", -- t[25444] = 7
      "000111" when "0110001101100101", -- t[25445] = 7
      "000111" when "0110001101100110", -- t[25446] = 7
      "000111" when "0110001101100111", -- t[25447] = 7
      "000111" when "0110001101101000", -- t[25448] = 7
      "000111" when "0110001101101001", -- t[25449] = 7
      "000111" when "0110001101101010", -- t[25450] = 7
      "000111" when "0110001101101011", -- t[25451] = 7
      "000111" when "0110001101101100", -- t[25452] = 7
      "000111" when "0110001101101101", -- t[25453] = 7
      "000111" when "0110001101101110", -- t[25454] = 7
      "000111" when "0110001101101111", -- t[25455] = 7
      "000111" when "0110001101110000", -- t[25456] = 7
      "000111" when "0110001101110001", -- t[25457] = 7
      "000111" when "0110001101110010", -- t[25458] = 7
      "000111" when "0110001101110011", -- t[25459] = 7
      "000111" when "0110001101110100", -- t[25460] = 7
      "000111" when "0110001101110101", -- t[25461] = 7
      "000111" when "0110001101110110", -- t[25462] = 7
      "000111" when "0110001101110111", -- t[25463] = 7
      "000111" when "0110001101111000", -- t[25464] = 7
      "000111" when "0110001101111001", -- t[25465] = 7
      "000111" when "0110001101111010", -- t[25466] = 7
      "000111" when "0110001101111011", -- t[25467] = 7
      "000111" when "0110001101111100", -- t[25468] = 7
      "000111" when "0110001101111101", -- t[25469] = 7
      "000111" when "0110001101111110", -- t[25470] = 7
      "000111" when "0110001101111111", -- t[25471] = 7
      "000111" when "0110001110000000", -- t[25472] = 7
      "000111" when "0110001110000001", -- t[25473] = 7
      "000111" when "0110001110000010", -- t[25474] = 7
      "000111" when "0110001110000011", -- t[25475] = 7
      "000111" when "0110001110000100", -- t[25476] = 7
      "000111" when "0110001110000101", -- t[25477] = 7
      "000111" when "0110001110000110", -- t[25478] = 7
      "000111" when "0110001110000111", -- t[25479] = 7
      "000111" when "0110001110001000", -- t[25480] = 7
      "000111" when "0110001110001001", -- t[25481] = 7
      "000111" when "0110001110001010", -- t[25482] = 7
      "000111" when "0110001110001011", -- t[25483] = 7
      "000111" when "0110001110001100", -- t[25484] = 7
      "000111" when "0110001110001101", -- t[25485] = 7
      "000111" when "0110001110001110", -- t[25486] = 7
      "000111" when "0110001110001111", -- t[25487] = 7
      "000111" when "0110001110010000", -- t[25488] = 7
      "000111" when "0110001110010001", -- t[25489] = 7
      "000111" when "0110001110010010", -- t[25490] = 7
      "000111" when "0110001110010011", -- t[25491] = 7
      "000111" when "0110001110010100", -- t[25492] = 7
      "000111" when "0110001110010101", -- t[25493] = 7
      "000111" when "0110001110010110", -- t[25494] = 7
      "000111" when "0110001110010111", -- t[25495] = 7
      "000111" when "0110001110011000", -- t[25496] = 7
      "000111" when "0110001110011001", -- t[25497] = 7
      "000111" when "0110001110011010", -- t[25498] = 7
      "000111" when "0110001110011011", -- t[25499] = 7
      "000111" when "0110001110011100", -- t[25500] = 7
      "000111" when "0110001110011101", -- t[25501] = 7
      "000111" when "0110001110011110", -- t[25502] = 7
      "000111" when "0110001110011111", -- t[25503] = 7
      "000111" when "0110001110100000", -- t[25504] = 7
      "000111" when "0110001110100001", -- t[25505] = 7
      "000111" when "0110001110100010", -- t[25506] = 7
      "000111" when "0110001110100011", -- t[25507] = 7
      "000111" when "0110001110100100", -- t[25508] = 7
      "000111" when "0110001110100101", -- t[25509] = 7
      "000111" when "0110001110100110", -- t[25510] = 7
      "000111" when "0110001110100111", -- t[25511] = 7
      "000111" when "0110001110101000", -- t[25512] = 7
      "000111" when "0110001110101001", -- t[25513] = 7
      "000111" when "0110001110101010", -- t[25514] = 7
      "000111" when "0110001110101011", -- t[25515] = 7
      "000111" when "0110001110101100", -- t[25516] = 7
      "000111" when "0110001110101101", -- t[25517] = 7
      "000111" when "0110001110101110", -- t[25518] = 7
      "000111" when "0110001110101111", -- t[25519] = 7
      "000111" when "0110001110110000", -- t[25520] = 7
      "000111" when "0110001110110001", -- t[25521] = 7
      "000111" when "0110001110110010", -- t[25522] = 7
      "000111" when "0110001110110011", -- t[25523] = 7
      "000111" when "0110001110110100", -- t[25524] = 7
      "000111" when "0110001110110101", -- t[25525] = 7
      "000111" when "0110001110110110", -- t[25526] = 7
      "000111" when "0110001110110111", -- t[25527] = 7
      "000111" when "0110001110111000", -- t[25528] = 7
      "000111" when "0110001110111001", -- t[25529] = 7
      "000111" when "0110001110111010", -- t[25530] = 7
      "000111" when "0110001110111011", -- t[25531] = 7
      "000111" when "0110001110111100", -- t[25532] = 7
      "000111" when "0110001110111101", -- t[25533] = 7
      "000111" when "0110001110111110", -- t[25534] = 7
      "000111" when "0110001110111111", -- t[25535] = 7
      "000111" when "0110001111000000", -- t[25536] = 7
      "000111" when "0110001111000001", -- t[25537] = 7
      "000111" when "0110001111000010", -- t[25538] = 7
      "000111" when "0110001111000011", -- t[25539] = 7
      "000111" when "0110001111000100", -- t[25540] = 7
      "000111" when "0110001111000101", -- t[25541] = 7
      "000111" when "0110001111000110", -- t[25542] = 7
      "000111" when "0110001111000111", -- t[25543] = 7
      "000111" when "0110001111001000", -- t[25544] = 7
      "000111" when "0110001111001001", -- t[25545] = 7
      "000111" when "0110001111001010", -- t[25546] = 7
      "000111" when "0110001111001011", -- t[25547] = 7
      "000111" when "0110001111001100", -- t[25548] = 7
      "000111" when "0110001111001101", -- t[25549] = 7
      "000111" when "0110001111001110", -- t[25550] = 7
      "000111" when "0110001111001111", -- t[25551] = 7
      "000111" when "0110001111010000", -- t[25552] = 7
      "000111" when "0110001111010001", -- t[25553] = 7
      "000111" when "0110001111010010", -- t[25554] = 7
      "000111" when "0110001111010011", -- t[25555] = 7
      "000111" when "0110001111010100", -- t[25556] = 7
      "000111" when "0110001111010101", -- t[25557] = 7
      "000111" when "0110001111010110", -- t[25558] = 7
      "000111" when "0110001111010111", -- t[25559] = 7
      "000111" when "0110001111011000", -- t[25560] = 7
      "000111" when "0110001111011001", -- t[25561] = 7
      "000111" when "0110001111011010", -- t[25562] = 7
      "000111" when "0110001111011011", -- t[25563] = 7
      "000111" when "0110001111011100", -- t[25564] = 7
      "000111" when "0110001111011101", -- t[25565] = 7
      "000111" when "0110001111011110", -- t[25566] = 7
      "000111" when "0110001111011111", -- t[25567] = 7
      "000111" when "0110001111100000", -- t[25568] = 7
      "000111" when "0110001111100001", -- t[25569] = 7
      "000111" when "0110001111100010", -- t[25570] = 7
      "000111" when "0110001111100011", -- t[25571] = 7
      "000111" when "0110001111100100", -- t[25572] = 7
      "000111" when "0110001111100101", -- t[25573] = 7
      "000111" when "0110001111100110", -- t[25574] = 7
      "000111" when "0110001111100111", -- t[25575] = 7
      "000111" when "0110001111101000", -- t[25576] = 7
      "000111" when "0110001111101001", -- t[25577] = 7
      "000111" when "0110001111101010", -- t[25578] = 7
      "000111" when "0110001111101011", -- t[25579] = 7
      "000111" when "0110001111101100", -- t[25580] = 7
      "000111" when "0110001111101101", -- t[25581] = 7
      "000111" when "0110001111101110", -- t[25582] = 7
      "000111" when "0110001111101111", -- t[25583] = 7
      "000111" when "0110001111110000", -- t[25584] = 7
      "000111" when "0110001111110001", -- t[25585] = 7
      "000111" when "0110001111110010", -- t[25586] = 7
      "000111" when "0110001111110011", -- t[25587] = 7
      "000111" when "0110001111110100", -- t[25588] = 7
      "000111" when "0110001111110101", -- t[25589] = 7
      "000111" when "0110001111110110", -- t[25590] = 7
      "000111" when "0110001111110111", -- t[25591] = 7
      "000111" when "0110001111111000", -- t[25592] = 7
      "000111" when "0110001111111001", -- t[25593] = 7
      "000111" when "0110001111111010", -- t[25594] = 7
      "000111" when "0110001111111011", -- t[25595] = 7
      "000111" when "0110001111111100", -- t[25596] = 7
      "000111" when "0110001111111101", -- t[25597] = 7
      "000111" when "0110001111111110", -- t[25598] = 7
      "000111" when "0110001111111111", -- t[25599] = 7
      "000111" when "0110010000000000", -- t[25600] = 7
      "000111" when "0110010000000001", -- t[25601] = 7
      "000111" when "0110010000000010", -- t[25602] = 7
      "000111" when "0110010000000011", -- t[25603] = 7
      "000111" when "0110010000000100", -- t[25604] = 7
      "000111" when "0110010000000101", -- t[25605] = 7
      "000111" when "0110010000000110", -- t[25606] = 7
      "000111" when "0110010000000111", -- t[25607] = 7
      "000111" when "0110010000001000", -- t[25608] = 7
      "000111" when "0110010000001001", -- t[25609] = 7
      "000111" when "0110010000001010", -- t[25610] = 7
      "000111" when "0110010000001011", -- t[25611] = 7
      "000111" when "0110010000001100", -- t[25612] = 7
      "000111" when "0110010000001101", -- t[25613] = 7
      "000111" when "0110010000001110", -- t[25614] = 7
      "000111" when "0110010000001111", -- t[25615] = 7
      "000111" when "0110010000010000", -- t[25616] = 7
      "000111" when "0110010000010001", -- t[25617] = 7
      "000111" when "0110010000010010", -- t[25618] = 7
      "000111" when "0110010000010011", -- t[25619] = 7
      "000111" when "0110010000010100", -- t[25620] = 7
      "000111" when "0110010000010101", -- t[25621] = 7
      "000111" when "0110010000010110", -- t[25622] = 7
      "000111" when "0110010000010111", -- t[25623] = 7
      "000111" when "0110010000011000", -- t[25624] = 7
      "000111" when "0110010000011001", -- t[25625] = 7
      "000111" when "0110010000011010", -- t[25626] = 7
      "000111" when "0110010000011011", -- t[25627] = 7
      "000111" when "0110010000011100", -- t[25628] = 7
      "000111" when "0110010000011101", -- t[25629] = 7
      "000111" when "0110010000011110", -- t[25630] = 7
      "000111" when "0110010000011111", -- t[25631] = 7
      "000111" when "0110010000100000", -- t[25632] = 7
      "000111" when "0110010000100001", -- t[25633] = 7
      "000111" when "0110010000100010", -- t[25634] = 7
      "000111" when "0110010000100011", -- t[25635] = 7
      "000111" when "0110010000100100", -- t[25636] = 7
      "000111" when "0110010000100101", -- t[25637] = 7
      "000111" when "0110010000100110", -- t[25638] = 7
      "000111" when "0110010000100111", -- t[25639] = 7
      "000111" when "0110010000101000", -- t[25640] = 7
      "000111" when "0110010000101001", -- t[25641] = 7
      "000111" when "0110010000101010", -- t[25642] = 7
      "000111" when "0110010000101011", -- t[25643] = 7
      "000111" when "0110010000101100", -- t[25644] = 7
      "000111" when "0110010000101101", -- t[25645] = 7
      "000111" when "0110010000101110", -- t[25646] = 7
      "000111" when "0110010000101111", -- t[25647] = 7
      "000111" when "0110010000110000", -- t[25648] = 7
      "000111" when "0110010000110001", -- t[25649] = 7
      "000111" when "0110010000110010", -- t[25650] = 7
      "000111" when "0110010000110011", -- t[25651] = 7
      "000111" when "0110010000110100", -- t[25652] = 7
      "000111" when "0110010000110101", -- t[25653] = 7
      "000111" when "0110010000110110", -- t[25654] = 7
      "000111" when "0110010000110111", -- t[25655] = 7
      "000111" when "0110010000111000", -- t[25656] = 7
      "000111" when "0110010000111001", -- t[25657] = 7
      "000111" when "0110010000111010", -- t[25658] = 7
      "000111" when "0110010000111011", -- t[25659] = 7
      "000111" when "0110010000111100", -- t[25660] = 7
      "000111" when "0110010000111101", -- t[25661] = 7
      "000111" when "0110010000111110", -- t[25662] = 7
      "000111" when "0110010000111111", -- t[25663] = 7
      "000111" when "0110010001000000", -- t[25664] = 7
      "000111" when "0110010001000001", -- t[25665] = 7
      "000111" when "0110010001000010", -- t[25666] = 7
      "000111" when "0110010001000011", -- t[25667] = 7
      "000111" when "0110010001000100", -- t[25668] = 7
      "000111" when "0110010001000101", -- t[25669] = 7
      "000111" when "0110010001000110", -- t[25670] = 7
      "000111" when "0110010001000111", -- t[25671] = 7
      "000111" when "0110010001001000", -- t[25672] = 7
      "000111" when "0110010001001001", -- t[25673] = 7
      "000111" when "0110010001001010", -- t[25674] = 7
      "000111" when "0110010001001011", -- t[25675] = 7
      "000111" when "0110010001001100", -- t[25676] = 7
      "000111" when "0110010001001101", -- t[25677] = 7
      "000111" when "0110010001001110", -- t[25678] = 7
      "000111" when "0110010001001111", -- t[25679] = 7
      "000111" when "0110010001010000", -- t[25680] = 7
      "000111" when "0110010001010001", -- t[25681] = 7
      "000111" when "0110010001010010", -- t[25682] = 7
      "000111" when "0110010001010011", -- t[25683] = 7
      "000111" when "0110010001010100", -- t[25684] = 7
      "000111" when "0110010001010101", -- t[25685] = 7
      "000111" when "0110010001010110", -- t[25686] = 7
      "000111" when "0110010001010111", -- t[25687] = 7
      "000111" when "0110010001011000", -- t[25688] = 7
      "000111" when "0110010001011001", -- t[25689] = 7
      "000111" when "0110010001011010", -- t[25690] = 7
      "000111" when "0110010001011011", -- t[25691] = 7
      "000111" when "0110010001011100", -- t[25692] = 7
      "000111" when "0110010001011101", -- t[25693] = 7
      "000111" when "0110010001011110", -- t[25694] = 7
      "000111" when "0110010001011111", -- t[25695] = 7
      "000111" when "0110010001100000", -- t[25696] = 7
      "000111" when "0110010001100001", -- t[25697] = 7
      "000111" when "0110010001100010", -- t[25698] = 7
      "000111" when "0110010001100011", -- t[25699] = 7
      "000111" when "0110010001100100", -- t[25700] = 7
      "000111" when "0110010001100101", -- t[25701] = 7
      "000111" when "0110010001100110", -- t[25702] = 7
      "000111" when "0110010001100111", -- t[25703] = 7
      "000111" when "0110010001101000", -- t[25704] = 7
      "000111" when "0110010001101001", -- t[25705] = 7
      "000111" when "0110010001101010", -- t[25706] = 7
      "000111" when "0110010001101011", -- t[25707] = 7
      "000111" when "0110010001101100", -- t[25708] = 7
      "000111" when "0110010001101101", -- t[25709] = 7
      "000111" when "0110010001101110", -- t[25710] = 7
      "000111" when "0110010001101111", -- t[25711] = 7
      "000111" when "0110010001110000", -- t[25712] = 7
      "000111" when "0110010001110001", -- t[25713] = 7
      "000111" when "0110010001110010", -- t[25714] = 7
      "000111" when "0110010001110011", -- t[25715] = 7
      "000111" when "0110010001110100", -- t[25716] = 7
      "000111" when "0110010001110101", -- t[25717] = 7
      "000111" when "0110010001110110", -- t[25718] = 7
      "000111" when "0110010001110111", -- t[25719] = 7
      "000111" when "0110010001111000", -- t[25720] = 7
      "000111" when "0110010001111001", -- t[25721] = 7
      "000111" when "0110010001111010", -- t[25722] = 7
      "000111" when "0110010001111011", -- t[25723] = 7
      "000111" when "0110010001111100", -- t[25724] = 7
      "000111" when "0110010001111101", -- t[25725] = 7
      "000111" when "0110010001111110", -- t[25726] = 7
      "000111" when "0110010001111111", -- t[25727] = 7
      "000111" when "0110010010000000", -- t[25728] = 7
      "000111" when "0110010010000001", -- t[25729] = 7
      "000111" when "0110010010000010", -- t[25730] = 7
      "000111" when "0110010010000011", -- t[25731] = 7
      "000111" when "0110010010000100", -- t[25732] = 7
      "000111" when "0110010010000101", -- t[25733] = 7
      "000111" when "0110010010000110", -- t[25734] = 7
      "000111" when "0110010010000111", -- t[25735] = 7
      "000111" when "0110010010001000", -- t[25736] = 7
      "000111" when "0110010010001001", -- t[25737] = 7
      "000111" when "0110010010001010", -- t[25738] = 7
      "000111" when "0110010010001011", -- t[25739] = 7
      "000111" when "0110010010001100", -- t[25740] = 7
      "000111" when "0110010010001101", -- t[25741] = 7
      "000111" when "0110010010001110", -- t[25742] = 7
      "000111" when "0110010010001111", -- t[25743] = 7
      "000111" when "0110010010010000", -- t[25744] = 7
      "000111" when "0110010010010001", -- t[25745] = 7
      "000111" when "0110010010010010", -- t[25746] = 7
      "000111" when "0110010010010011", -- t[25747] = 7
      "000111" when "0110010010010100", -- t[25748] = 7
      "000111" when "0110010010010101", -- t[25749] = 7
      "000111" when "0110010010010110", -- t[25750] = 7
      "000111" when "0110010010010111", -- t[25751] = 7
      "000111" when "0110010010011000", -- t[25752] = 7
      "000111" when "0110010010011001", -- t[25753] = 7
      "000111" when "0110010010011010", -- t[25754] = 7
      "000111" when "0110010010011011", -- t[25755] = 7
      "000111" when "0110010010011100", -- t[25756] = 7
      "000111" when "0110010010011101", -- t[25757] = 7
      "000111" when "0110010010011110", -- t[25758] = 7
      "000111" when "0110010010011111", -- t[25759] = 7
      "000111" when "0110010010100000", -- t[25760] = 7
      "000111" when "0110010010100001", -- t[25761] = 7
      "000111" when "0110010010100010", -- t[25762] = 7
      "000111" when "0110010010100011", -- t[25763] = 7
      "000111" when "0110010010100100", -- t[25764] = 7
      "000111" when "0110010010100101", -- t[25765] = 7
      "000111" when "0110010010100110", -- t[25766] = 7
      "000111" when "0110010010100111", -- t[25767] = 7
      "000111" when "0110010010101000", -- t[25768] = 7
      "000111" when "0110010010101001", -- t[25769] = 7
      "000111" when "0110010010101010", -- t[25770] = 7
      "000111" when "0110010010101011", -- t[25771] = 7
      "000111" when "0110010010101100", -- t[25772] = 7
      "000111" when "0110010010101101", -- t[25773] = 7
      "000111" when "0110010010101110", -- t[25774] = 7
      "000111" when "0110010010101111", -- t[25775] = 7
      "000111" when "0110010010110000", -- t[25776] = 7
      "000111" when "0110010010110001", -- t[25777] = 7
      "000111" when "0110010010110010", -- t[25778] = 7
      "000111" when "0110010010110011", -- t[25779] = 7
      "000111" when "0110010010110100", -- t[25780] = 7
      "000111" when "0110010010110101", -- t[25781] = 7
      "000111" when "0110010010110110", -- t[25782] = 7
      "000111" when "0110010010110111", -- t[25783] = 7
      "000111" when "0110010010111000", -- t[25784] = 7
      "000111" when "0110010010111001", -- t[25785] = 7
      "000111" when "0110010010111010", -- t[25786] = 7
      "000111" when "0110010010111011", -- t[25787] = 7
      "000111" when "0110010010111100", -- t[25788] = 7
      "000111" when "0110010010111101", -- t[25789] = 7
      "000111" when "0110010010111110", -- t[25790] = 7
      "000111" when "0110010010111111", -- t[25791] = 7
      "000111" when "0110010011000000", -- t[25792] = 7
      "000111" when "0110010011000001", -- t[25793] = 7
      "000111" when "0110010011000010", -- t[25794] = 7
      "000111" when "0110010011000011", -- t[25795] = 7
      "000111" when "0110010011000100", -- t[25796] = 7
      "000111" when "0110010011000101", -- t[25797] = 7
      "000111" when "0110010011000110", -- t[25798] = 7
      "000111" when "0110010011000111", -- t[25799] = 7
      "000111" when "0110010011001000", -- t[25800] = 7
      "000111" when "0110010011001001", -- t[25801] = 7
      "000111" when "0110010011001010", -- t[25802] = 7
      "000111" when "0110010011001011", -- t[25803] = 7
      "000111" when "0110010011001100", -- t[25804] = 7
      "000111" when "0110010011001101", -- t[25805] = 7
      "000111" when "0110010011001110", -- t[25806] = 7
      "000111" when "0110010011001111", -- t[25807] = 7
      "000111" when "0110010011010000", -- t[25808] = 7
      "000111" when "0110010011010001", -- t[25809] = 7
      "000111" when "0110010011010010", -- t[25810] = 7
      "000111" when "0110010011010011", -- t[25811] = 7
      "000111" when "0110010011010100", -- t[25812] = 7
      "000111" when "0110010011010101", -- t[25813] = 7
      "000111" when "0110010011010110", -- t[25814] = 7
      "000111" when "0110010011010111", -- t[25815] = 7
      "000111" when "0110010011011000", -- t[25816] = 7
      "000111" when "0110010011011001", -- t[25817] = 7
      "000111" when "0110010011011010", -- t[25818] = 7
      "000111" when "0110010011011011", -- t[25819] = 7
      "000111" when "0110010011011100", -- t[25820] = 7
      "000111" when "0110010011011101", -- t[25821] = 7
      "000111" when "0110010011011110", -- t[25822] = 7
      "000111" when "0110010011011111", -- t[25823] = 7
      "000111" when "0110010011100000", -- t[25824] = 7
      "000111" when "0110010011100001", -- t[25825] = 7
      "000111" when "0110010011100010", -- t[25826] = 7
      "000111" when "0110010011100011", -- t[25827] = 7
      "000111" when "0110010011100100", -- t[25828] = 7
      "000111" when "0110010011100101", -- t[25829] = 7
      "000111" when "0110010011100110", -- t[25830] = 7
      "000111" when "0110010011100111", -- t[25831] = 7
      "000111" when "0110010011101000", -- t[25832] = 7
      "000111" when "0110010011101001", -- t[25833] = 7
      "000111" when "0110010011101010", -- t[25834] = 7
      "000111" when "0110010011101011", -- t[25835] = 7
      "000111" when "0110010011101100", -- t[25836] = 7
      "000111" when "0110010011101101", -- t[25837] = 7
      "000111" when "0110010011101110", -- t[25838] = 7
      "000111" when "0110010011101111", -- t[25839] = 7
      "000111" when "0110010011110000", -- t[25840] = 7
      "000111" when "0110010011110001", -- t[25841] = 7
      "000111" when "0110010011110010", -- t[25842] = 7
      "000111" when "0110010011110011", -- t[25843] = 7
      "000111" when "0110010011110100", -- t[25844] = 7
      "000111" when "0110010011110101", -- t[25845] = 7
      "000111" when "0110010011110110", -- t[25846] = 7
      "000111" when "0110010011110111", -- t[25847] = 7
      "000111" when "0110010011111000", -- t[25848] = 7
      "000111" when "0110010011111001", -- t[25849] = 7
      "000111" when "0110010011111010", -- t[25850] = 7
      "000111" when "0110010011111011", -- t[25851] = 7
      "000111" when "0110010011111100", -- t[25852] = 7
      "000111" when "0110010011111101", -- t[25853] = 7
      "000111" when "0110010011111110", -- t[25854] = 7
      "000111" when "0110010011111111", -- t[25855] = 7
      "000111" when "0110010100000000", -- t[25856] = 7
      "000111" when "0110010100000001", -- t[25857] = 7
      "000111" when "0110010100000010", -- t[25858] = 7
      "000111" when "0110010100000011", -- t[25859] = 7
      "000111" when "0110010100000100", -- t[25860] = 7
      "000111" when "0110010100000101", -- t[25861] = 7
      "000111" when "0110010100000110", -- t[25862] = 7
      "000111" when "0110010100000111", -- t[25863] = 7
      "000111" when "0110010100001000", -- t[25864] = 7
      "000111" when "0110010100001001", -- t[25865] = 7
      "000111" when "0110010100001010", -- t[25866] = 7
      "000111" when "0110010100001011", -- t[25867] = 7
      "000111" when "0110010100001100", -- t[25868] = 7
      "000111" when "0110010100001101", -- t[25869] = 7
      "000111" when "0110010100001110", -- t[25870] = 7
      "000111" when "0110010100001111", -- t[25871] = 7
      "000111" when "0110010100010000", -- t[25872] = 7
      "000111" when "0110010100010001", -- t[25873] = 7
      "000111" when "0110010100010010", -- t[25874] = 7
      "000111" when "0110010100010011", -- t[25875] = 7
      "000111" when "0110010100010100", -- t[25876] = 7
      "000111" when "0110010100010101", -- t[25877] = 7
      "000111" when "0110010100010110", -- t[25878] = 7
      "000111" when "0110010100010111", -- t[25879] = 7
      "000111" when "0110010100011000", -- t[25880] = 7
      "000111" when "0110010100011001", -- t[25881] = 7
      "000111" when "0110010100011010", -- t[25882] = 7
      "000111" when "0110010100011011", -- t[25883] = 7
      "000111" when "0110010100011100", -- t[25884] = 7
      "000111" when "0110010100011101", -- t[25885] = 7
      "000111" when "0110010100011110", -- t[25886] = 7
      "000111" when "0110010100011111", -- t[25887] = 7
      "000111" when "0110010100100000", -- t[25888] = 7
      "000111" when "0110010100100001", -- t[25889] = 7
      "000111" when "0110010100100010", -- t[25890] = 7
      "000111" when "0110010100100011", -- t[25891] = 7
      "000111" when "0110010100100100", -- t[25892] = 7
      "000111" when "0110010100100101", -- t[25893] = 7
      "000111" when "0110010100100110", -- t[25894] = 7
      "000111" when "0110010100100111", -- t[25895] = 7
      "000111" when "0110010100101000", -- t[25896] = 7
      "000111" when "0110010100101001", -- t[25897] = 7
      "000111" when "0110010100101010", -- t[25898] = 7
      "000111" when "0110010100101011", -- t[25899] = 7
      "000111" when "0110010100101100", -- t[25900] = 7
      "000111" when "0110010100101101", -- t[25901] = 7
      "000111" when "0110010100101110", -- t[25902] = 7
      "000111" when "0110010100101111", -- t[25903] = 7
      "000111" when "0110010100110000", -- t[25904] = 7
      "000111" when "0110010100110001", -- t[25905] = 7
      "000111" when "0110010100110010", -- t[25906] = 7
      "000111" when "0110010100110011", -- t[25907] = 7
      "000111" when "0110010100110100", -- t[25908] = 7
      "000111" when "0110010100110101", -- t[25909] = 7
      "000111" when "0110010100110110", -- t[25910] = 7
      "000111" when "0110010100110111", -- t[25911] = 7
      "000111" when "0110010100111000", -- t[25912] = 7
      "000111" when "0110010100111001", -- t[25913] = 7
      "000111" when "0110010100111010", -- t[25914] = 7
      "000111" when "0110010100111011", -- t[25915] = 7
      "000111" when "0110010100111100", -- t[25916] = 7
      "000111" when "0110010100111101", -- t[25917] = 7
      "000111" when "0110010100111110", -- t[25918] = 7
      "000111" when "0110010100111111", -- t[25919] = 7
      "000111" when "0110010101000000", -- t[25920] = 7
      "000111" when "0110010101000001", -- t[25921] = 7
      "000111" when "0110010101000010", -- t[25922] = 7
      "000111" when "0110010101000011", -- t[25923] = 7
      "000111" when "0110010101000100", -- t[25924] = 7
      "000111" when "0110010101000101", -- t[25925] = 7
      "000111" when "0110010101000110", -- t[25926] = 7
      "000111" when "0110010101000111", -- t[25927] = 7
      "000111" when "0110010101001000", -- t[25928] = 7
      "000111" when "0110010101001001", -- t[25929] = 7
      "000111" when "0110010101001010", -- t[25930] = 7
      "000111" when "0110010101001011", -- t[25931] = 7
      "000111" when "0110010101001100", -- t[25932] = 7
      "000111" when "0110010101001101", -- t[25933] = 7
      "000111" when "0110010101001110", -- t[25934] = 7
      "000111" when "0110010101001111", -- t[25935] = 7
      "000111" when "0110010101010000", -- t[25936] = 7
      "000111" when "0110010101010001", -- t[25937] = 7
      "000111" when "0110010101010010", -- t[25938] = 7
      "000111" when "0110010101010011", -- t[25939] = 7
      "000111" when "0110010101010100", -- t[25940] = 7
      "000111" when "0110010101010101", -- t[25941] = 7
      "000111" when "0110010101010110", -- t[25942] = 7
      "000111" when "0110010101010111", -- t[25943] = 7
      "000111" when "0110010101011000", -- t[25944] = 7
      "000111" when "0110010101011001", -- t[25945] = 7
      "000111" when "0110010101011010", -- t[25946] = 7
      "000111" when "0110010101011011", -- t[25947] = 7
      "000111" when "0110010101011100", -- t[25948] = 7
      "000111" when "0110010101011101", -- t[25949] = 7
      "000111" when "0110010101011110", -- t[25950] = 7
      "000111" when "0110010101011111", -- t[25951] = 7
      "000111" when "0110010101100000", -- t[25952] = 7
      "000111" when "0110010101100001", -- t[25953] = 7
      "000111" when "0110010101100010", -- t[25954] = 7
      "000111" when "0110010101100011", -- t[25955] = 7
      "000111" when "0110010101100100", -- t[25956] = 7
      "000111" when "0110010101100101", -- t[25957] = 7
      "000111" when "0110010101100110", -- t[25958] = 7
      "000111" when "0110010101100111", -- t[25959] = 7
      "000111" when "0110010101101000", -- t[25960] = 7
      "000111" when "0110010101101001", -- t[25961] = 7
      "000111" when "0110010101101010", -- t[25962] = 7
      "000111" when "0110010101101011", -- t[25963] = 7
      "000111" when "0110010101101100", -- t[25964] = 7
      "000111" when "0110010101101101", -- t[25965] = 7
      "000111" when "0110010101101110", -- t[25966] = 7
      "000111" when "0110010101101111", -- t[25967] = 7
      "000111" when "0110010101110000", -- t[25968] = 7
      "000111" when "0110010101110001", -- t[25969] = 7
      "000111" when "0110010101110010", -- t[25970] = 7
      "000111" when "0110010101110011", -- t[25971] = 7
      "000111" when "0110010101110100", -- t[25972] = 7
      "000111" when "0110010101110101", -- t[25973] = 7
      "000111" when "0110010101110110", -- t[25974] = 7
      "000111" when "0110010101110111", -- t[25975] = 7
      "000111" when "0110010101111000", -- t[25976] = 7
      "000111" when "0110010101111001", -- t[25977] = 7
      "000111" when "0110010101111010", -- t[25978] = 7
      "000111" when "0110010101111011", -- t[25979] = 7
      "000111" when "0110010101111100", -- t[25980] = 7
      "000111" when "0110010101111101", -- t[25981] = 7
      "000111" when "0110010101111110", -- t[25982] = 7
      "000111" when "0110010101111111", -- t[25983] = 7
      "000111" when "0110010110000000", -- t[25984] = 7
      "000111" when "0110010110000001", -- t[25985] = 7
      "000111" when "0110010110000010", -- t[25986] = 7
      "000111" when "0110010110000011", -- t[25987] = 7
      "000111" when "0110010110000100", -- t[25988] = 7
      "000111" when "0110010110000101", -- t[25989] = 7
      "000111" when "0110010110000110", -- t[25990] = 7
      "000111" when "0110010110000111", -- t[25991] = 7
      "000111" when "0110010110001000", -- t[25992] = 7
      "000111" when "0110010110001001", -- t[25993] = 7
      "000111" when "0110010110001010", -- t[25994] = 7
      "000111" when "0110010110001011", -- t[25995] = 7
      "000111" when "0110010110001100", -- t[25996] = 7
      "000111" when "0110010110001101", -- t[25997] = 7
      "000111" when "0110010110001110", -- t[25998] = 7
      "000111" when "0110010110001111", -- t[25999] = 7
      "000111" when "0110010110010000", -- t[26000] = 7
      "000111" when "0110010110010001", -- t[26001] = 7
      "000111" when "0110010110010010", -- t[26002] = 7
      "000111" when "0110010110010011", -- t[26003] = 7
      "000111" when "0110010110010100", -- t[26004] = 7
      "000111" when "0110010110010101", -- t[26005] = 7
      "000111" when "0110010110010110", -- t[26006] = 7
      "000111" when "0110010110010111", -- t[26007] = 7
      "000111" when "0110010110011000", -- t[26008] = 7
      "000111" when "0110010110011001", -- t[26009] = 7
      "000111" when "0110010110011010", -- t[26010] = 7
      "000111" when "0110010110011011", -- t[26011] = 7
      "000111" when "0110010110011100", -- t[26012] = 7
      "000111" when "0110010110011101", -- t[26013] = 7
      "000111" when "0110010110011110", -- t[26014] = 7
      "000111" when "0110010110011111", -- t[26015] = 7
      "000111" when "0110010110100000", -- t[26016] = 7
      "000111" when "0110010110100001", -- t[26017] = 7
      "000111" when "0110010110100010", -- t[26018] = 7
      "000111" when "0110010110100011", -- t[26019] = 7
      "000111" when "0110010110100100", -- t[26020] = 7
      "000111" when "0110010110100101", -- t[26021] = 7
      "000111" when "0110010110100110", -- t[26022] = 7
      "000111" when "0110010110100111", -- t[26023] = 7
      "000111" when "0110010110101000", -- t[26024] = 7
      "000111" when "0110010110101001", -- t[26025] = 7
      "000111" when "0110010110101010", -- t[26026] = 7
      "000111" when "0110010110101011", -- t[26027] = 7
      "000111" when "0110010110101100", -- t[26028] = 7
      "000111" when "0110010110101101", -- t[26029] = 7
      "000111" when "0110010110101110", -- t[26030] = 7
      "000111" when "0110010110101111", -- t[26031] = 7
      "000111" when "0110010110110000", -- t[26032] = 7
      "000111" when "0110010110110001", -- t[26033] = 7
      "000111" when "0110010110110010", -- t[26034] = 7
      "000111" when "0110010110110011", -- t[26035] = 7
      "000111" when "0110010110110100", -- t[26036] = 7
      "000111" when "0110010110110101", -- t[26037] = 7
      "000111" when "0110010110110110", -- t[26038] = 7
      "000111" when "0110010110110111", -- t[26039] = 7
      "000111" when "0110010110111000", -- t[26040] = 7
      "000111" when "0110010110111001", -- t[26041] = 7
      "000111" when "0110010110111010", -- t[26042] = 7
      "000111" when "0110010110111011", -- t[26043] = 7
      "000111" when "0110010110111100", -- t[26044] = 7
      "000111" when "0110010110111101", -- t[26045] = 7
      "000111" when "0110010110111110", -- t[26046] = 7
      "000111" when "0110010110111111", -- t[26047] = 7
      "000111" when "0110010111000000", -- t[26048] = 7
      "000111" when "0110010111000001", -- t[26049] = 7
      "000111" when "0110010111000010", -- t[26050] = 7
      "000111" when "0110010111000011", -- t[26051] = 7
      "000111" when "0110010111000100", -- t[26052] = 7
      "000111" when "0110010111000101", -- t[26053] = 7
      "000111" when "0110010111000110", -- t[26054] = 7
      "000111" when "0110010111000111", -- t[26055] = 7
      "000111" when "0110010111001000", -- t[26056] = 7
      "000111" when "0110010111001001", -- t[26057] = 7
      "000111" when "0110010111001010", -- t[26058] = 7
      "000111" when "0110010111001011", -- t[26059] = 7
      "000111" when "0110010111001100", -- t[26060] = 7
      "000111" when "0110010111001101", -- t[26061] = 7
      "000111" when "0110010111001110", -- t[26062] = 7
      "000111" when "0110010111001111", -- t[26063] = 7
      "000111" when "0110010111010000", -- t[26064] = 7
      "000111" when "0110010111010001", -- t[26065] = 7
      "000111" when "0110010111010010", -- t[26066] = 7
      "000111" when "0110010111010011", -- t[26067] = 7
      "000111" when "0110010111010100", -- t[26068] = 7
      "000111" when "0110010111010101", -- t[26069] = 7
      "000111" when "0110010111010110", -- t[26070] = 7
      "000111" when "0110010111010111", -- t[26071] = 7
      "000111" when "0110010111011000", -- t[26072] = 7
      "000111" when "0110010111011001", -- t[26073] = 7
      "000111" when "0110010111011010", -- t[26074] = 7
      "000111" when "0110010111011011", -- t[26075] = 7
      "000111" when "0110010111011100", -- t[26076] = 7
      "000111" when "0110010111011101", -- t[26077] = 7
      "000111" when "0110010111011110", -- t[26078] = 7
      "000111" when "0110010111011111", -- t[26079] = 7
      "000111" when "0110010111100000", -- t[26080] = 7
      "000111" when "0110010111100001", -- t[26081] = 7
      "000111" when "0110010111100010", -- t[26082] = 7
      "000111" when "0110010111100011", -- t[26083] = 7
      "000111" when "0110010111100100", -- t[26084] = 7
      "000111" when "0110010111100101", -- t[26085] = 7
      "000111" when "0110010111100110", -- t[26086] = 7
      "000111" when "0110010111100111", -- t[26087] = 7
      "000111" when "0110010111101000", -- t[26088] = 7
      "000111" when "0110010111101001", -- t[26089] = 7
      "000111" when "0110010111101010", -- t[26090] = 7
      "000111" when "0110010111101011", -- t[26091] = 7
      "000111" when "0110010111101100", -- t[26092] = 7
      "000111" when "0110010111101101", -- t[26093] = 7
      "000111" when "0110010111101110", -- t[26094] = 7
      "000111" when "0110010111101111", -- t[26095] = 7
      "000111" when "0110010111110000", -- t[26096] = 7
      "000111" when "0110010111110001", -- t[26097] = 7
      "000111" when "0110010111110010", -- t[26098] = 7
      "000111" when "0110010111110011", -- t[26099] = 7
      "000111" when "0110010111110100", -- t[26100] = 7
      "000111" when "0110010111110101", -- t[26101] = 7
      "000111" when "0110010111110110", -- t[26102] = 7
      "000111" when "0110010111110111", -- t[26103] = 7
      "000111" when "0110010111111000", -- t[26104] = 7
      "000111" when "0110010111111001", -- t[26105] = 7
      "000111" when "0110010111111010", -- t[26106] = 7
      "000111" when "0110010111111011", -- t[26107] = 7
      "000111" when "0110010111111100", -- t[26108] = 7
      "000111" when "0110010111111101", -- t[26109] = 7
      "000111" when "0110010111111110", -- t[26110] = 7
      "000111" when "0110010111111111", -- t[26111] = 7
      "000111" when "0110011000000000", -- t[26112] = 7
      "000111" when "0110011000000001", -- t[26113] = 7
      "000111" when "0110011000000010", -- t[26114] = 7
      "000111" when "0110011000000011", -- t[26115] = 7
      "000111" when "0110011000000100", -- t[26116] = 7
      "000111" when "0110011000000101", -- t[26117] = 7
      "000111" when "0110011000000110", -- t[26118] = 7
      "000111" when "0110011000000111", -- t[26119] = 7
      "000111" when "0110011000001000", -- t[26120] = 7
      "000111" when "0110011000001001", -- t[26121] = 7
      "001000" when "0110011000001010", -- t[26122] = 8
      "001000" when "0110011000001011", -- t[26123] = 8
      "001000" when "0110011000001100", -- t[26124] = 8
      "001000" when "0110011000001101", -- t[26125] = 8
      "001000" when "0110011000001110", -- t[26126] = 8
      "001000" when "0110011000001111", -- t[26127] = 8
      "001000" when "0110011000010000", -- t[26128] = 8
      "001000" when "0110011000010001", -- t[26129] = 8
      "001000" when "0110011000010010", -- t[26130] = 8
      "001000" when "0110011000010011", -- t[26131] = 8
      "001000" when "0110011000010100", -- t[26132] = 8
      "001000" when "0110011000010101", -- t[26133] = 8
      "001000" when "0110011000010110", -- t[26134] = 8
      "001000" when "0110011000010111", -- t[26135] = 8
      "001000" when "0110011000011000", -- t[26136] = 8
      "001000" when "0110011000011001", -- t[26137] = 8
      "001000" when "0110011000011010", -- t[26138] = 8
      "001000" when "0110011000011011", -- t[26139] = 8
      "001000" when "0110011000011100", -- t[26140] = 8
      "001000" when "0110011000011101", -- t[26141] = 8
      "001000" when "0110011000011110", -- t[26142] = 8
      "001000" when "0110011000011111", -- t[26143] = 8
      "001000" when "0110011000100000", -- t[26144] = 8
      "001000" when "0110011000100001", -- t[26145] = 8
      "001000" when "0110011000100010", -- t[26146] = 8
      "001000" when "0110011000100011", -- t[26147] = 8
      "001000" when "0110011000100100", -- t[26148] = 8
      "001000" when "0110011000100101", -- t[26149] = 8
      "001000" when "0110011000100110", -- t[26150] = 8
      "001000" when "0110011000100111", -- t[26151] = 8
      "001000" when "0110011000101000", -- t[26152] = 8
      "001000" when "0110011000101001", -- t[26153] = 8
      "001000" when "0110011000101010", -- t[26154] = 8
      "001000" when "0110011000101011", -- t[26155] = 8
      "001000" when "0110011000101100", -- t[26156] = 8
      "001000" when "0110011000101101", -- t[26157] = 8
      "001000" when "0110011000101110", -- t[26158] = 8
      "001000" when "0110011000101111", -- t[26159] = 8
      "001000" when "0110011000110000", -- t[26160] = 8
      "001000" when "0110011000110001", -- t[26161] = 8
      "001000" when "0110011000110010", -- t[26162] = 8
      "001000" when "0110011000110011", -- t[26163] = 8
      "001000" when "0110011000110100", -- t[26164] = 8
      "001000" when "0110011000110101", -- t[26165] = 8
      "001000" when "0110011000110110", -- t[26166] = 8
      "001000" when "0110011000110111", -- t[26167] = 8
      "001000" when "0110011000111000", -- t[26168] = 8
      "001000" when "0110011000111001", -- t[26169] = 8
      "001000" when "0110011000111010", -- t[26170] = 8
      "001000" when "0110011000111011", -- t[26171] = 8
      "001000" when "0110011000111100", -- t[26172] = 8
      "001000" when "0110011000111101", -- t[26173] = 8
      "001000" when "0110011000111110", -- t[26174] = 8
      "001000" when "0110011000111111", -- t[26175] = 8
      "001000" when "0110011001000000", -- t[26176] = 8
      "001000" when "0110011001000001", -- t[26177] = 8
      "001000" when "0110011001000010", -- t[26178] = 8
      "001000" when "0110011001000011", -- t[26179] = 8
      "001000" when "0110011001000100", -- t[26180] = 8
      "001000" when "0110011001000101", -- t[26181] = 8
      "001000" when "0110011001000110", -- t[26182] = 8
      "001000" when "0110011001000111", -- t[26183] = 8
      "001000" when "0110011001001000", -- t[26184] = 8
      "001000" when "0110011001001001", -- t[26185] = 8
      "001000" when "0110011001001010", -- t[26186] = 8
      "001000" when "0110011001001011", -- t[26187] = 8
      "001000" when "0110011001001100", -- t[26188] = 8
      "001000" when "0110011001001101", -- t[26189] = 8
      "001000" when "0110011001001110", -- t[26190] = 8
      "001000" when "0110011001001111", -- t[26191] = 8
      "001000" when "0110011001010000", -- t[26192] = 8
      "001000" when "0110011001010001", -- t[26193] = 8
      "001000" when "0110011001010010", -- t[26194] = 8
      "001000" when "0110011001010011", -- t[26195] = 8
      "001000" when "0110011001010100", -- t[26196] = 8
      "001000" when "0110011001010101", -- t[26197] = 8
      "001000" when "0110011001010110", -- t[26198] = 8
      "001000" when "0110011001010111", -- t[26199] = 8
      "001000" when "0110011001011000", -- t[26200] = 8
      "001000" when "0110011001011001", -- t[26201] = 8
      "001000" when "0110011001011010", -- t[26202] = 8
      "001000" when "0110011001011011", -- t[26203] = 8
      "001000" when "0110011001011100", -- t[26204] = 8
      "001000" when "0110011001011101", -- t[26205] = 8
      "001000" when "0110011001011110", -- t[26206] = 8
      "001000" when "0110011001011111", -- t[26207] = 8
      "001000" when "0110011001100000", -- t[26208] = 8
      "001000" when "0110011001100001", -- t[26209] = 8
      "001000" when "0110011001100010", -- t[26210] = 8
      "001000" when "0110011001100011", -- t[26211] = 8
      "001000" when "0110011001100100", -- t[26212] = 8
      "001000" when "0110011001100101", -- t[26213] = 8
      "001000" when "0110011001100110", -- t[26214] = 8
      "001000" when "0110011001100111", -- t[26215] = 8
      "001000" when "0110011001101000", -- t[26216] = 8
      "001000" when "0110011001101001", -- t[26217] = 8
      "001000" when "0110011001101010", -- t[26218] = 8
      "001000" when "0110011001101011", -- t[26219] = 8
      "001000" when "0110011001101100", -- t[26220] = 8
      "001000" when "0110011001101101", -- t[26221] = 8
      "001000" when "0110011001101110", -- t[26222] = 8
      "001000" when "0110011001101111", -- t[26223] = 8
      "001000" when "0110011001110000", -- t[26224] = 8
      "001000" when "0110011001110001", -- t[26225] = 8
      "001000" when "0110011001110010", -- t[26226] = 8
      "001000" when "0110011001110011", -- t[26227] = 8
      "001000" when "0110011001110100", -- t[26228] = 8
      "001000" when "0110011001110101", -- t[26229] = 8
      "001000" when "0110011001110110", -- t[26230] = 8
      "001000" when "0110011001110111", -- t[26231] = 8
      "001000" when "0110011001111000", -- t[26232] = 8
      "001000" when "0110011001111001", -- t[26233] = 8
      "001000" when "0110011001111010", -- t[26234] = 8
      "001000" when "0110011001111011", -- t[26235] = 8
      "001000" when "0110011001111100", -- t[26236] = 8
      "001000" when "0110011001111101", -- t[26237] = 8
      "001000" when "0110011001111110", -- t[26238] = 8
      "001000" when "0110011001111111", -- t[26239] = 8
      "001000" when "0110011010000000", -- t[26240] = 8
      "001000" when "0110011010000001", -- t[26241] = 8
      "001000" when "0110011010000010", -- t[26242] = 8
      "001000" when "0110011010000011", -- t[26243] = 8
      "001000" when "0110011010000100", -- t[26244] = 8
      "001000" when "0110011010000101", -- t[26245] = 8
      "001000" when "0110011010000110", -- t[26246] = 8
      "001000" when "0110011010000111", -- t[26247] = 8
      "001000" when "0110011010001000", -- t[26248] = 8
      "001000" when "0110011010001001", -- t[26249] = 8
      "001000" when "0110011010001010", -- t[26250] = 8
      "001000" when "0110011010001011", -- t[26251] = 8
      "001000" when "0110011010001100", -- t[26252] = 8
      "001000" when "0110011010001101", -- t[26253] = 8
      "001000" when "0110011010001110", -- t[26254] = 8
      "001000" when "0110011010001111", -- t[26255] = 8
      "001000" when "0110011010010000", -- t[26256] = 8
      "001000" when "0110011010010001", -- t[26257] = 8
      "001000" when "0110011010010010", -- t[26258] = 8
      "001000" when "0110011010010011", -- t[26259] = 8
      "001000" when "0110011010010100", -- t[26260] = 8
      "001000" when "0110011010010101", -- t[26261] = 8
      "001000" when "0110011010010110", -- t[26262] = 8
      "001000" when "0110011010010111", -- t[26263] = 8
      "001000" when "0110011010011000", -- t[26264] = 8
      "001000" when "0110011010011001", -- t[26265] = 8
      "001000" when "0110011010011010", -- t[26266] = 8
      "001000" when "0110011010011011", -- t[26267] = 8
      "001000" when "0110011010011100", -- t[26268] = 8
      "001000" when "0110011010011101", -- t[26269] = 8
      "001000" when "0110011010011110", -- t[26270] = 8
      "001000" when "0110011010011111", -- t[26271] = 8
      "001000" when "0110011010100000", -- t[26272] = 8
      "001000" when "0110011010100001", -- t[26273] = 8
      "001000" when "0110011010100010", -- t[26274] = 8
      "001000" when "0110011010100011", -- t[26275] = 8
      "001000" when "0110011010100100", -- t[26276] = 8
      "001000" when "0110011010100101", -- t[26277] = 8
      "001000" when "0110011010100110", -- t[26278] = 8
      "001000" when "0110011010100111", -- t[26279] = 8
      "001000" when "0110011010101000", -- t[26280] = 8
      "001000" when "0110011010101001", -- t[26281] = 8
      "001000" when "0110011010101010", -- t[26282] = 8
      "001000" when "0110011010101011", -- t[26283] = 8
      "001000" when "0110011010101100", -- t[26284] = 8
      "001000" when "0110011010101101", -- t[26285] = 8
      "001000" when "0110011010101110", -- t[26286] = 8
      "001000" when "0110011010101111", -- t[26287] = 8
      "001000" when "0110011010110000", -- t[26288] = 8
      "001000" when "0110011010110001", -- t[26289] = 8
      "001000" when "0110011010110010", -- t[26290] = 8
      "001000" when "0110011010110011", -- t[26291] = 8
      "001000" when "0110011010110100", -- t[26292] = 8
      "001000" when "0110011010110101", -- t[26293] = 8
      "001000" when "0110011010110110", -- t[26294] = 8
      "001000" when "0110011010110111", -- t[26295] = 8
      "001000" when "0110011010111000", -- t[26296] = 8
      "001000" when "0110011010111001", -- t[26297] = 8
      "001000" when "0110011010111010", -- t[26298] = 8
      "001000" when "0110011010111011", -- t[26299] = 8
      "001000" when "0110011010111100", -- t[26300] = 8
      "001000" when "0110011010111101", -- t[26301] = 8
      "001000" when "0110011010111110", -- t[26302] = 8
      "001000" when "0110011010111111", -- t[26303] = 8
      "001000" when "0110011011000000", -- t[26304] = 8
      "001000" when "0110011011000001", -- t[26305] = 8
      "001000" when "0110011011000010", -- t[26306] = 8
      "001000" when "0110011011000011", -- t[26307] = 8
      "001000" when "0110011011000100", -- t[26308] = 8
      "001000" when "0110011011000101", -- t[26309] = 8
      "001000" when "0110011011000110", -- t[26310] = 8
      "001000" when "0110011011000111", -- t[26311] = 8
      "001000" when "0110011011001000", -- t[26312] = 8
      "001000" when "0110011011001001", -- t[26313] = 8
      "001000" when "0110011011001010", -- t[26314] = 8
      "001000" when "0110011011001011", -- t[26315] = 8
      "001000" when "0110011011001100", -- t[26316] = 8
      "001000" when "0110011011001101", -- t[26317] = 8
      "001000" when "0110011011001110", -- t[26318] = 8
      "001000" when "0110011011001111", -- t[26319] = 8
      "001000" when "0110011011010000", -- t[26320] = 8
      "001000" when "0110011011010001", -- t[26321] = 8
      "001000" when "0110011011010010", -- t[26322] = 8
      "001000" when "0110011011010011", -- t[26323] = 8
      "001000" when "0110011011010100", -- t[26324] = 8
      "001000" when "0110011011010101", -- t[26325] = 8
      "001000" when "0110011011010110", -- t[26326] = 8
      "001000" when "0110011011010111", -- t[26327] = 8
      "001000" when "0110011011011000", -- t[26328] = 8
      "001000" when "0110011011011001", -- t[26329] = 8
      "001000" when "0110011011011010", -- t[26330] = 8
      "001000" when "0110011011011011", -- t[26331] = 8
      "001000" when "0110011011011100", -- t[26332] = 8
      "001000" when "0110011011011101", -- t[26333] = 8
      "001000" when "0110011011011110", -- t[26334] = 8
      "001000" when "0110011011011111", -- t[26335] = 8
      "001000" when "0110011011100000", -- t[26336] = 8
      "001000" when "0110011011100001", -- t[26337] = 8
      "001000" when "0110011011100010", -- t[26338] = 8
      "001000" when "0110011011100011", -- t[26339] = 8
      "001000" when "0110011011100100", -- t[26340] = 8
      "001000" when "0110011011100101", -- t[26341] = 8
      "001000" when "0110011011100110", -- t[26342] = 8
      "001000" when "0110011011100111", -- t[26343] = 8
      "001000" when "0110011011101000", -- t[26344] = 8
      "001000" when "0110011011101001", -- t[26345] = 8
      "001000" when "0110011011101010", -- t[26346] = 8
      "001000" when "0110011011101011", -- t[26347] = 8
      "001000" when "0110011011101100", -- t[26348] = 8
      "001000" when "0110011011101101", -- t[26349] = 8
      "001000" when "0110011011101110", -- t[26350] = 8
      "001000" when "0110011011101111", -- t[26351] = 8
      "001000" when "0110011011110000", -- t[26352] = 8
      "001000" when "0110011011110001", -- t[26353] = 8
      "001000" when "0110011011110010", -- t[26354] = 8
      "001000" when "0110011011110011", -- t[26355] = 8
      "001000" when "0110011011110100", -- t[26356] = 8
      "001000" when "0110011011110101", -- t[26357] = 8
      "001000" when "0110011011110110", -- t[26358] = 8
      "001000" when "0110011011110111", -- t[26359] = 8
      "001000" when "0110011011111000", -- t[26360] = 8
      "001000" when "0110011011111001", -- t[26361] = 8
      "001000" when "0110011011111010", -- t[26362] = 8
      "001000" when "0110011011111011", -- t[26363] = 8
      "001000" when "0110011011111100", -- t[26364] = 8
      "001000" when "0110011011111101", -- t[26365] = 8
      "001000" when "0110011011111110", -- t[26366] = 8
      "001000" when "0110011011111111", -- t[26367] = 8
      "001000" when "0110011100000000", -- t[26368] = 8
      "001000" when "0110011100000001", -- t[26369] = 8
      "001000" when "0110011100000010", -- t[26370] = 8
      "001000" when "0110011100000011", -- t[26371] = 8
      "001000" when "0110011100000100", -- t[26372] = 8
      "001000" when "0110011100000101", -- t[26373] = 8
      "001000" when "0110011100000110", -- t[26374] = 8
      "001000" when "0110011100000111", -- t[26375] = 8
      "001000" when "0110011100001000", -- t[26376] = 8
      "001000" when "0110011100001001", -- t[26377] = 8
      "001000" when "0110011100001010", -- t[26378] = 8
      "001000" when "0110011100001011", -- t[26379] = 8
      "001000" when "0110011100001100", -- t[26380] = 8
      "001000" when "0110011100001101", -- t[26381] = 8
      "001000" when "0110011100001110", -- t[26382] = 8
      "001000" when "0110011100001111", -- t[26383] = 8
      "001000" when "0110011100010000", -- t[26384] = 8
      "001000" when "0110011100010001", -- t[26385] = 8
      "001000" when "0110011100010010", -- t[26386] = 8
      "001000" when "0110011100010011", -- t[26387] = 8
      "001000" when "0110011100010100", -- t[26388] = 8
      "001000" when "0110011100010101", -- t[26389] = 8
      "001000" when "0110011100010110", -- t[26390] = 8
      "001000" when "0110011100010111", -- t[26391] = 8
      "001000" when "0110011100011000", -- t[26392] = 8
      "001000" when "0110011100011001", -- t[26393] = 8
      "001000" when "0110011100011010", -- t[26394] = 8
      "001000" when "0110011100011011", -- t[26395] = 8
      "001000" when "0110011100011100", -- t[26396] = 8
      "001000" when "0110011100011101", -- t[26397] = 8
      "001000" when "0110011100011110", -- t[26398] = 8
      "001000" when "0110011100011111", -- t[26399] = 8
      "001000" when "0110011100100000", -- t[26400] = 8
      "001000" when "0110011100100001", -- t[26401] = 8
      "001000" when "0110011100100010", -- t[26402] = 8
      "001000" when "0110011100100011", -- t[26403] = 8
      "001000" when "0110011100100100", -- t[26404] = 8
      "001000" when "0110011100100101", -- t[26405] = 8
      "001000" when "0110011100100110", -- t[26406] = 8
      "001000" when "0110011100100111", -- t[26407] = 8
      "001000" when "0110011100101000", -- t[26408] = 8
      "001000" when "0110011100101001", -- t[26409] = 8
      "001000" when "0110011100101010", -- t[26410] = 8
      "001000" when "0110011100101011", -- t[26411] = 8
      "001000" when "0110011100101100", -- t[26412] = 8
      "001000" when "0110011100101101", -- t[26413] = 8
      "001000" when "0110011100101110", -- t[26414] = 8
      "001000" when "0110011100101111", -- t[26415] = 8
      "001000" when "0110011100110000", -- t[26416] = 8
      "001000" when "0110011100110001", -- t[26417] = 8
      "001000" when "0110011100110010", -- t[26418] = 8
      "001000" when "0110011100110011", -- t[26419] = 8
      "001000" when "0110011100110100", -- t[26420] = 8
      "001000" when "0110011100110101", -- t[26421] = 8
      "001000" when "0110011100110110", -- t[26422] = 8
      "001000" when "0110011100110111", -- t[26423] = 8
      "001000" when "0110011100111000", -- t[26424] = 8
      "001000" when "0110011100111001", -- t[26425] = 8
      "001000" when "0110011100111010", -- t[26426] = 8
      "001000" when "0110011100111011", -- t[26427] = 8
      "001000" when "0110011100111100", -- t[26428] = 8
      "001000" when "0110011100111101", -- t[26429] = 8
      "001000" when "0110011100111110", -- t[26430] = 8
      "001000" when "0110011100111111", -- t[26431] = 8
      "001000" when "0110011101000000", -- t[26432] = 8
      "001000" when "0110011101000001", -- t[26433] = 8
      "001000" when "0110011101000010", -- t[26434] = 8
      "001000" when "0110011101000011", -- t[26435] = 8
      "001000" when "0110011101000100", -- t[26436] = 8
      "001000" when "0110011101000101", -- t[26437] = 8
      "001000" when "0110011101000110", -- t[26438] = 8
      "001000" when "0110011101000111", -- t[26439] = 8
      "001000" when "0110011101001000", -- t[26440] = 8
      "001000" when "0110011101001001", -- t[26441] = 8
      "001000" when "0110011101001010", -- t[26442] = 8
      "001000" when "0110011101001011", -- t[26443] = 8
      "001000" when "0110011101001100", -- t[26444] = 8
      "001000" when "0110011101001101", -- t[26445] = 8
      "001000" when "0110011101001110", -- t[26446] = 8
      "001000" when "0110011101001111", -- t[26447] = 8
      "001000" when "0110011101010000", -- t[26448] = 8
      "001000" when "0110011101010001", -- t[26449] = 8
      "001000" when "0110011101010010", -- t[26450] = 8
      "001000" when "0110011101010011", -- t[26451] = 8
      "001000" when "0110011101010100", -- t[26452] = 8
      "001000" when "0110011101010101", -- t[26453] = 8
      "001000" when "0110011101010110", -- t[26454] = 8
      "001000" when "0110011101010111", -- t[26455] = 8
      "001000" when "0110011101011000", -- t[26456] = 8
      "001000" when "0110011101011001", -- t[26457] = 8
      "001000" when "0110011101011010", -- t[26458] = 8
      "001000" when "0110011101011011", -- t[26459] = 8
      "001000" when "0110011101011100", -- t[26460] = 8
      "001000" when "0110011101011101", -- t[26461] = 8
      "001000" when "0110011101011110", -- t[26462] = 8
      "001000" when "0110011101011111", -- t[26463] = 8
      "001000" when "0110011101100000", -- t[26464] = 8
      "001000" when "0110011101100001", -- t[26465] = 8
      "001000" when "0110011101100010", -- t[26466] = 8
      "001000" when "0110011101100011", -- t[26467] = 8
      "001000" when "0110011101100100", -- t[26468] = 8
      "001000" when "0110011101100101", -- t[26469] = 8
      "001000" when "0110011101100110", -- t[26470] = 8
      "001000" when "0110011101100111", -- t[26471] = 8
      "001000" when "0110011101101000", -- t[26472] = 8
      "001000" when "0110011101101001", -- t[26473] = 8
      "001000" when "0110011101101010", -- t[26474] = 8
      "001000" when "0110011101101011", -- t[26475] = 8
      "001000" when "0110011101101100", -- t[26476] = 8
      "001000" when "0110011101101101", -- t[26477] = 8
      "001000" when "0110011101101110", -- t[26478] = 8
      "001000" when "0110011101101111", -- t[26479] = 8
      "001000" when "0110011101110000", -- t[26480] = 8
      "001000" when "0110011101110001", -- t[26481] = 8
      "001000" when "0110011101110010", -- t[26482] = 8
      "001000" when "0110011101110011", -- t[26483] = 8
      "001000" when "0110011101110100", -- t[26484] = 8
      "001000" when "0110011101110101", -- t[26485] = 8
      "001000" when "0110011101110110", -- t[26486] = 8
      "001000" when "0110011101110111", -- t[26487] = 8
      "001000" when "0110011101111000", -- t[26488] = 8
      "001000" when "0110011101111001", -- t[26489] = 8
      "001000" when "0110011101111010", -- t[26490] = 8
      "001000" when "0110011101111011", -- t[26491] = 8
      "001000" when "0110011101111100", -- t[26492] = 8
      "001000" when "0110011101111101", -- t[26493] = 8
      "001000" when "0110011101111110", -- t[26494] = 8
      "001000" when "0110011101111111", -- t[26495] = 8
      "001000" when "0110011110000000", -- t[26496] = 8
      "001000" when "0110011110000001", -- t[26497] = 8
      "001000" when "0110011110000010", -- t[26498] = 8
      "001000" when "0110011110000011", -- t[26499] = 8
      "001000" when "0110011110000100", -- t[26500] = 8
      "001000" when "0110011110000101", -- t[26501] = 8
      "001000" when "0110011110000110", -- t[26502] = 8
      "001000" when "0110011110000111", -- t[26503] = 8
      "001000" when "0110011110001000", -- t[26504] = 8
      "001000" when "0110011110001001", -- t[26505] = 8
      "001000" when "0110011110001010", -- t[26506] = 8
      "001000" when "0110011110001011", -- t[26507] = 8
      "001000" when "0110011110001100", -- t[26508] = 8
      "001000" when "0110011110001101", -- t[26509] = 8
      "001000" when "0110011110001110", -- t[26510] = 8
      "001000" when "0110011110001111", -- t[26511] = 8
      "001000" when "0110011110010000", -- t[26512] = 8
      "001000" when "0110011110010001", -- t[26513] = 8
      "001000" when "0110011110010010", -- t[26514] = 8
      "001000" when "0110011110010011", -- t[26515] = 8
      "001000" when "0110011110010100", -- t[26516] = 8
      "001000" when "0110011110010101", -- t[26517] = 8
      "001000" when "0110011110010110", -- t[26518] = 8
      "001000" when "0110011110010111", -- t[26519] = 8
      "001000" when "0110011110011000", -- t[26520] = 8
      "001000" when "0110011110011001", -- t[26521] = 8
      "001000" when "0110011110011010", -- t[26522] = 8
      "001000" when "0110011110011011", -- t[26523] = 8
      "001000" when "0110011110011100", -- t[26524] = 8
      "001000" when "0110011110011101", -- t[26525] = 8
      "001000" when "0110011110011110", -- t[26526] = 8
      "001000" when "0110011110011111", -- t[26527] = 8
      "001000" when "0110011110100000", -- t[26528] = 8
      "001000" when "0110011110100001", -- t[26529] = 8
      "001000" when "0110011110100010", -- t[26530] = 8
      "001000" when "0110011110100011", -- t[26531] = 8
      "001000" when "0110011110100100", -- t[26532] = 8
      "001000" when "0110011110100101", -- t[26533] = 8
      "001000" when "0110011110100110", -- t[26534] = 8
      "001000" when "0110011110100111", -- t[26535] = 8
      "001000" when "0110011110101000", -- t[26536] = 8
      "001000" when "0110011110101001", -- t[26537] = 8
      "001000" when "0110011110101010", -- t[26538] = 8
      "001000" when "0110011110101011", -- t[26539] = 8
      "001000" when "0110011110101100", -- t[26540] = 8
      "001000" when "0110011110101101", -- t[26541] = 8
      "001000" when "0110011110101110", -- t[26542] = 8
      "001000" when "0110011110101111", -- t[26543] = 8
      "001000" when "0110011110110000", -- t[26544] = 8
      "001000" when "0110011110110001", -- t[26545] = 8
      "001000" when "0110011110110010", -- t[26546] = 8
      "001000" when "0110011110110011", -- t[26547] = 8
      "001000" when "0110011110110100", -- t[26548] = 8
      "001000" when "0110011110110101", -- t[26549] = 8
      "001000" when "0110011110110110", -- t[26550] = 8
      "001000" when "0110011110110111", -- t[26551] = 8
      "001000" when "0110011110111000", -- t[26552] = 8
      "001000" when "0110011110111001", -- t[26553] = 8
      "001000" when "0110011110111010", -- t[26554] = 8
      "001000" when "0110011110111011", -- t[26555] = 8
      "001000" when "0110011110111100", -- t[26556] = 8
      "001000" when "0110011110111101", -- t[26557] = 8
      "001000" when "0110011110111110", -- t[26558] = 8
      "001000" when "0110011110111111", -- t[26559] = 8
      "001000" when "0110011111000000", -- t[26560] = 8
      "001000" when "0110011111000001", -- t[26561] = 8
      "001000" when "0110011111000010", -- t[26562] = 8
      "001000" when "0110011111000011", -- t[26563] = 8
      "001000" when "0110011111000100", -- t[26564] = 8
      "001000" when "0110011111000101", -- t[26565] = 8
      "001000" when "0110011111000110", -- t[26566] = 8
      "001000" when "0110011111000111", -- t[26567] = 8
      "001000" when "0110011111001000", -- t[26568] = 8
      "001000" when "0110011111001001", -- t[26569] = 8
      "001000" when "0110011111001010", -- t[26570] = 8
      "001000" when "0110011111001011", -- t[26571] = 8
      "001000" when "0110011111001100", -- t[26572] = 8
      "001000" when "0110011111001101", -- t[26573] = 8
      "001000" when "0110011111001110", -- t[26574] = 8
      "001000" when "0110011111001111", -- t[26575] = 8
      "001000" when "0110011111010000", -- t[26576] = 8
      "001000" when "0110011111010001", -- t[26577] = 8
      "001000" when "0110011111010010", -- t[26578] = 8
      "001000" when "0110011111010011", -- t[26579] = 8
      "001000" when "0110011111010100", -- t[26580] = 8
      "001000" when "0110011111010101", -- t[26581] = 8
      "001000" when "0110011111010110", -- t[26582] = 8
      "001000" when "0110011111010111", -- t[26583] = 8
      "001000" when "0110011111011000", -- t[26584] = 8
      "001000" when "0110011111011001", -- t[26585] = 8
      "001000" when "0110011111011010", -- t[26586] = 8
      "001000" when "0110011111011011", -- t[26587] = 8
      "001000" when "0110011111011100", -- t[26588] = 8
      "001000" when "0110011111011101", -- t[26589] = 8
      "001000" when "0110011111011110", -- t[26590] = 8
      "001000" when "0110011111011111", -- t[26591] = 8
      "001000" when "0110011111100000", -- t[26592] = 8
      "001000" when "0110011111100001", -- t[26593] = 8
      "001000" when "0110011111100010", -- t[26594] = 8
      "001000" when "0110011111100011", -- t[26595] = 8
      "001000" when "0110011111100100", -- t[26596] = 8
      "001000" when "0110011111100101", -- t[26597] = 8
      "001000" when "0110011111100110", -- t[26598] = 8
      "001000" when "0110011111100111", -- t[26599] = 8
      "001000" when "0110011111101000", -- t[26600] = 8
      "001000" when "0110011111101001", -- t[26601] = 8
      "001000" when "0110011111101010", -- t[26602] = 8
      "001000" when "0110011111101011", -- t[26603] = 8
      "001000" when "0110011111101100", -- t[26604] = 8
      "001000" when "0110011111101101", -- t[26605] = 8
      "001000" when "0110011111101110", -- t[26606] = 8
      "001000" when "0110011111101111", -- t[26607] = 8
      "001000" when "0110011111110000", -- t[26608] = 8
      "001000" when "0110011111110001", -- t[26609] = 8
      "001000" when "0110011111110010", -- t[26610] = 8
      "001000" when "0110011111110011", -- t[26611] = 8
      "001000" when "0110011111110100", -- t[26612] = 8
      "001000" when "0110011111110101", -- t[26613] = 8
      "001000" when "0110011111110110", -- t[26614] = 8
      "001000" when "0110011111110111", -- t[26615] = 8
      "001000" when "0110011111111000", -- t[26616] = 8
      "001000" when "0110011111111001", -- t[26617] = 8
      "001000" when "0110011111111010", -- t[26618] = 8
      "001000" when "0110011111111011", -- t[26619] = 8
      "001000" when "0110011111111100", -- t[26620] = 8
      "001000" when "0110011111111101", -- t[26621] = 8
      "001000" when "0110011111111110", -- t[26622] = 8
      "001000" when "0110011111111111", -- t[26623] = 8
      "001000" when "0110100000000000", -- t[26624] = 8
      "001000" when "0110100000000001", -- t[26625] = 8
      "001000" when "0110100000000010", -- t[26626] = 8
      "001000" when "0110100000000011", -- t[26627] = 8
      "001000" when "0110100000000100", -- t[26628] = 8
      "001000" when "0110100000000101", -- t[26629] = 8
      "001000" when "0110100000000110", -- t[26630] = 8
      "001000" when "0110100000000111", -- t[26631] = 8
      "001000" when "0110100000001000", -- t[26632] = 8
      "001000" when "0110100000001001", -- t[26633] = 8
      "001000" when "0110100000001010", -- t[26634] = 8
      "001000" when "0110100000001011", -- t[26635] = 8
      "001000" when "0110100000001100", -- t[26636] = 8
      "001000" when "0110100000001101", -- t[26637] = 8
      "001000" when "0110100000001110", -- t[26638] = 8
      "001000" when "0110100000001111", -- t[26639] = 8
      "001000" when "0110100000010000", -- t[26640] = 8
      "001000" when "0110100000010001", -- t[26641] = 8
      "001000" when "0110100000010010", -- t[26642] = 8
      "001000" when "0110100000010011", -- t[26643] = 8
      "001000" when "0110100000010100", -- t[26644] = 8
      "001000" when "0110100000010101", -- t[26645] = 8
      "001000" when "0110100000010110", -- t[26646] = 8
      "001000" when "0110100000010111", -- t[26647] = 8
      "001000" when "0110100000011000", -- t[26648] = 8
      "001000" when "0110100000011001", -- t[26649] = 8
      "001000" when "0110100000011010", -- t[26650] = 8
      "001000" when "0110100000011011", -- t[26651] = 8
      "001000" when "0110100000011100", -- t[26652] = 8
      "001000" when "0110100000011101", -- t[26653] = 8
      "001000" when "0110100000011110", -- t[26654] = 8
      "001000" when "0110100000011111", -- t[26655] = 8
      "001000" when "0110100000100000", -- t[26656] = 8
      "001000" when "0110100000100001", -- t[26657] = 8
      "001000" when "0110100000100010", -- t[26658] = 8
      "001000" when "0110100000100011", -- t[26659] = 8
      "001000" when "0110100000100100", -- t[26660] = 8
      "001000" when "0110100000100101", -- t[26661] = 8
      "001000" when "0110100000100110", -- t[26662] = 8
      "001000" when "0110100000100111", -- t[26663] = 8
      "001000" when "0110100000101000", -- t[26664] = 8
      "001000" when "0110100000101001", -- t[26665] = 8
      "001000" when "0110100000101010", -- t[26666] = 8
      "001000" when "0110100000101011", -- t[26667] = 8
      "001000" when "0110100000101100", -- t[26668] = 8
      "001000" when "0110100000101101", -- t[26669] = 8
      "001000" when "0110100000101110", -- t[26670] = 8
      "001000" when "0110100000101111", -- t[26671] = 8
      "001000" when "0110100000110000", -- t[26672] = 8
      "001000" when "0110100000110001", -- t[26673] = 8
      "001000" when "0110100000110010", -- t[26674] = 8
      "001000" when "0110100000110011", -- t[26675] = 8
      "001000" when "0110100000110100", -- t[26676] = 8
      "001000" when "0110100000110101", -- t[26677] = 8
      "001000" when "0110100000110110", -- t[26678] = 8
      "001000" when "0110100000110111", -- t[26679] = 8
      "001000" when "0110100000111000", -- t[26680] = 8
      "001000" when "0110100000111001", -- t[26681] = 8
      "001000" when "0110100000111010", -- t[26682] = 8
      "001000" when "0110100000111011", -- t[26683] = 8
      "001000" when "0110100000111100", -- t[26684] = 8
      "001000" when "0110100000111101", -- t[26685] = 8
      "001000" when "0110100000111110", -- t[26686] = 8
      "001000" when "0110100000111111", -- t[26687] = 8
      "001000" when "0110100001000000", -- t[26688] = 8
      "001000" when "0110100001000001", -- t[26689] = 8
      "001000" when "0110100001000010", -- t[26690] = 8
      "001000" when "0110100001000011", -- t[26691] = 8
      "001000" when "0110100001000100", -- t[26692] = 8
      "001000" when "0110100001000101", -- t[26693] = 8
      "001000" when "0110100001000110", -- t[26694] = 8
      "001000" when "0110100001000111", -- t[26695] = 8
      "001000" when "0110100001001000", -- t[26696] = 8
      "001000" when "0110100001001001", -- t[26697] = 8
      "001000" when "0110100001001010", -- t[26698] = 8
      "001000" when "0110100001001011", -- t[26699] = 8
      "001000" when "0110100001001100", -- t[26700] = 8
      "001000" when "0110100001001101", -- t[26701] = 8
      "001000" when "0110100001001110", -- t[26702] = 8
      "001000" when "0110100001001111", -- t[26703] = 8
      "001000" when "0110100001010000", -- t[26704] = 8
      "001000" when "0110100001010001", -- t[26705] = 8
      "001000" when "0110100001010010", -- t[26706] = 8
      "001000" when "0110100001010011", -- t[26707] = 8
      "001000" when "0110100001010100", -- t[26708] = 8
      "001000" when "0110100001010101", -- t[26709] = 8
      "001000" when "0110100001010110", -- t[26710] = 8
      "001000" when "0110100001010111", -- t[26711] = 8
      "001000" when "0110100001011000", -- t[26712] = 8
      "001000" when "0110100001011001", -- t[26713] = 8
      "001000" when "0110100001011010", -- t[26714] = 8
      "001000" when "0110100001011011", -- t[26715] = 8
      "001000" when "0110100001011100", -- t[26716] = 8
      "001000" when "0110100001011101", -- t[26717] = 8
      "001000" when "0110100001011110", -- t[26718] = 8
      "001000" when "0110100001011111", -- t[26719] = 8
      "001000" when "0110100001100000", -- t[26720] = 8
      "001000" when "0110100001100001", -- t[26721] = 8
      "001000" when "0110100001100010", -- t[26722] = 8
      "001000" when "0110100001100011", -- t[26723] = 8
      "001000" when "0110100001100100", -- t[26724] = 8
      "001000" when "0110100001100101", -- t[26725] = 8
      "001000" when "0110100001100110", -- t[26726] = 8
      "001000" when "0110100001100111", -- t[26727] = 8
      "001000" when "0110100001101000", -- t[26728] = 8
      "001000" when "0110100001101001", -- t[26729] = 8
      "001000" when "0110100001101010", -- t[26730] = 8
      "001000" when "0110100001101011", -- t[26731] = 8
      "001000" when "0110100001101100", -- t[26732] = 8
      "001000" when "0110100001101101", -- t[26733] = 8
      "001000" when "0110100001101110", -- t[26734] = 8
      "001000" when "0110100001101111", -- t[26735] = 8
      "001000" when "0110100001110000", -- t[26736] = 8
      "001000" when "0110100001110001", -- t[26737] = 8
      "001000" when "0110100001110010", -- t[26738] = 8
      "001000" when "0110100001110011", -- t[26739] = 8
      "001000" when "0110100001110100", -- t[26740] = 8
      "001000" when "0110100001110101", -- t[26741] = 8
      "001000" when "0110100001110110", -- t[26742] = 8
      "001000" when "0110100001110111", -- t[26743] = 8
      "001000" when "0110100001111000", -- t[26744] = 8
      "001000" when "0110100001111001", -- t[26745] = 8
      "001000" when "0110100001111010", -- t[26746] = 8
      "001000" when "0110100001111011", -- t[26747] = 8
      "001000" when "0110100001111100", -- t[26748] = 8
      "001000" when "0110100001111101", -- t[26749] = 8
      "001000" when "0110100001111110", -- t[26750] = 8
      "001000" when "0110100001111111", -- t[26751] = 8
      "001000" when "0110100010000000", -- t[26752] = 8
      "001000" when "0110100010000001", -- t[26753] = 8
      "001000" when "0110100010000010", -- t[26754] = 8
      "001000" when "0110100010000011", -- t[26755] = 8
      "001000" when "0110100010000100", -- t[26756] = 8
      "001000" when "0110100010000101", -- t[26757] = 8
      "001000" when "0110100010000110", -- t[26758] = 8
      "001000" when "0110100010000111", -- t[26759] = 8
      "001000" when "0110100010001000", -- t[26760] = 8
      "001000" when "0110100010001001", -- t[26761] = 8
      "001000" when "0110100010001010", -- t[26762] = 8
      "001000" when "0110100010001011", -- t[26763] = 8
      "001000" when "0110100010001100", -- t[26764] = 8
      "001000" when "0110100010001101", -- t[26765] = 8
      "001000" when "0110100010001110", -- t[26766] = 8
      "001000" when "0110100010001111", -- t[26767] = 8
      "001000" when "0110100010010000", -- t[26768] = 8
      "001000" when "0110100010010001", -- t[26769] = 8
      "001000" when "0110100010010010", -- t[26770] = 8
      "001000" when "0110100010010011", -- t[26771] = 8
      "001000" when "0110100010010100", -- t[26772] = 8
      "001000" when "0110100010010101", -- t[26773] = 8
      "001000" when "0110100010010110", -- t[26774] = 8
      "001000" when "0110100010010111", -- t[26775] = 8
      "001000" when "0110100010011000", -- t[26776] = 8
      "001000" when "0110100010011001", -- t[26777] = 8
      "001000" when "0110100010011010", -- t[26778] = 8
      "001000" when "0110100010011011", -- t[26779] = 8
      "001000" when "0110100010011100", -- t[26780] = 8
      "001000" when "0110100010011101", -- t[26781] = 8
      "001000" when "0110100010011110", -- t[26782] = 8
      "001000" when "0110100010011111", -- t[26783] = 8
      "001000" when "0110100010100000", -- t[26784] = 8
      "001000" when "0110100010100001", -- t[26785] = 8
      "001000" when "0110100010100010", -- t[26786] = 8
      "001000" when "0110100010100011", -- t[26787] = 8
      "001000" when "0110100010100100", -- t[26788] = 8
      "001000" when "0110100010100101", -- t[26789] = 8
      "001000" when "0110100010100110", -- t[26790] = 8
      "001000" when "0110100010100111", -- t[26791] = 8
      "001000" when "0110100010101000", -- t[26792] = 8
      "001000" when "0110100010101001", -- t[26793] = 8
      "001000" when "0110100010101010", -- t[26794] = 8
      "001000" when "0110100010101011", -- t[26795] = 8
      "001000" when "0110100010101100", -- t[26796] = 8
      "001000" when "0110100010101101", -- t[26797] = 8
      "001000" when "0110100010101110", -- t[26798] = 8
      "001000" when "0110100010101111", -- t[26799] = 8
      "001000" when "0110100010110000", -- t[26800] = 8
      "001000" when "0110100010110001", -- t[26801] = 8
      "001000" when "0110100010110010", -- t[26802] = 8
      "001000" when "0110100010110011", -- t[26803] = 8
      "001000" when "0110100010110100", -- t[26804] = 8
      "001000" when "0110100010110101", -- t[26805] = 8
      "001000" when "0110100010110110", -- t[26806] = 8
      "001000" when "0110100010110111", -- t[26807] = 8
      "001000" when "0110100010111000", -- t[26808] = 8
      "001000" when "0110100010111001", -- t[26809] = 8
      "001000" when "0110100010111010", -- t[26810] = 8
      "001000" when "0110100010111011", -- t[26811] = 8
      "001000" when "0110100010111100", -- t[26812] = 8
      "001000" when "0110100010111101", -- t[26813] = 8
      "001000" when "0110100010111110", -- t[26814] = 8
      "001000" when "0110100010111111", -- t[26815] = 8
      "001000" when "0110100011000000", -- t[26816] = 8
      "001000" when "0110100011000001", -- t[26817] = 8
      "001000" when "0110100011000010", -- t[26818] = 8
      "001000" when "0110100011000011", -- t[26819] = 8
      "001000" when "0110100011000100", -- t[26820] = 8
      "001000" when "0110100011000101", -- t[26821] = 8
      "001000" when "0110100011000110", -- t[26822] = 8
      "001000" when "0110100011000111", -- t[26823] = 8
      "001000" when "0110100011001000", -- t[26824] = 8
      "001000" when "0110100011001001", -- t[26825] = 8
      "001000" when "0110100011001010", -- t[26826] = 8
      "001000" when "0110100011001011", -- t[26827] = 8
      "001000" when "0110100011001100", -- t[26828] = 8
      "001000" when "0110100011001101", -- t[26829] = 8
      "001000" when "0110100011001110", -- t[26830] = 8
      "001000" when "0110100011001111", -- t[26831] = 8
      "001000" when "0110100011010000", -- t[26832] = 8
      "001000" when "0110100011010001", -- t[26833] = 8
      "001000" when "0110100011010010", -- t[26834] = 8
      "001000" when "0110100011010011", -- t[26835] = 8
      "001000" when "0110100011010100", -- t[26836] = 8
      "001000" when "0110100011010101", -- t[26837] = 8
      "001000" when "0110100011010110", -- t[26838] = 8
      "001000" when "0110100011010111", -- t[26839] = 8
      "001000" when "0110100011011000", -- t[26840] = 8
      "001000" when "0110100011011001", -- t[26841] = 8
      "001000" when "0110100011011010", -- t[26842] = 8
      "001000" when "0110100011011011", -- t[26843] = 8
      "001000" when "0110100011011100", -- t[26844] = 8
      "001000" when "0110100011011101", -- t[26845] = 8
      "001000" when "0110100011011110", -- t[26846] = 8
      "001000" when "0110100011011111", -- t[26847] = 8
      "001000" when "0110100011100000", -- t[26848] = 8
      "001000" when "0110100011100001", -- t[26849] = 8
      "001000" when "0110100011100010", -- t[26850] = 8
      "001000" when "0110100011100011", -- t[26851] = 8
      "001000" when "0110100011100100", -- t[26852] = 8
      "001000" when "0110100011100101", -- t[26853] = 8
      "001000" when "0110100011100110", -- t[26854] = 8
      "001000" when "0110100011100111", -- t[26855] = 8
      "001000" when "0110100011101000", -- t[26856] = 8
      "001000" when "0110100011101001", -- t[26857] = 8
      "001000" when "0110100011101010", -- t[26858] = 8
      "001000" when "0110100011101011", -- t[26859] = 8
      "001000" when "0110100011101100", -- t[26860] = 8
      "001001" when "0110100011101101", -- t[26861] = 9
      "001001" when "0110100011101110", -- t[26862] = 9
      "001001" when "0110100011101111", -- t[26863] = 9
      "001001" when "0110100011110000", -- t[26864] = 9
      "001001" when "0110100011110001", -- t[26865] = 9
      "001001" when "0110100011110010", -- t[26866] = 9
      "001001" when "0110100011110011", -- t[26867] = 9
      "001001" when "0110100011110100", -- t[26868] = 9
      "001001" when "0110100011110101", -- t[26869] = 9
      "001001" when "0110100011110110", -- t[26870] = 9
      "001001" when "0110100011110111", -- t[26871] = 9
      "001001" when "0110100011111000", -- t[26872] = 9
      "001001" when "0110100011111001", -- t[26873] = 9
      "001001" when "0110100011111010", -- t[26874] = 9
      "001001" when "0110100011111011", -- t[26875] = 9
      "001001" when "0110100011111100", -- t[26876] = 9
      "001001" when "0110100011111101", -- t[26877] = 9
      "001001" when "0110100011111110", -- t[26878] = 9
      "001001" when "0110100011111111", -- t[26879] = 9
      "001001" when "0110100100000000", -- t[26880] = 9
      "001001" when "0110100100000001", -- t[26881] = 9
      "001001" when "0110100100000010", -- t[26882] = 9
      "001001" when "0110100100000011", -- t[26883] = 9
      "001001" when "0110100100000100", -- t[26884] = 9
      "001001" when "0110100100000101", -- t[26885] = 9
      "001001" when "0110100100000110", -- t[26886] = 9
      "001001" when "0110100100000111", -- t[26887] = 9
      "001001" when "0110100100001000", -- t[26888] = 9
      "001001" when "0110100100001001", -- t[26889] = 9
      "001001" when "0110100100001010", -- t[26890] = 9
      "001001" when "0110100100001011", -- t[26891] = 9
      "001001" when "0110100100001100", -- t[26892] = 9
      "001001" when "0110100100001101", -- t[26893] = 9
      "001001" when "0110100100001110", -- t[26894] = 9
      "001001" when "0110100100001111", -- t[26895] = 9
      "001001" when "0110100100010000", -- t[26896] = 9
      "001001" when "0110100100010001", -- t[26897] = 9
      "001001" when "0110100100010010", -- t[26898] = 9
      "001001" when "0110100100010011", -- t[26899] = 9
      "001001" when "0110100100010100", -- t[26900] = 9
      "001001" when "0110100100010101", -- t[26901] = 9
      "001001" when "0110100100010110", -- t[26902] = 9
      "001001" when "0110100100010111", -- t[26903] = 9
      "001001" when "0110100100011000", -- t[26904] = 9
      "001001" when "0110100100011001", -- t[26905] = 9
      "001001" when "0110100100011010", -- t[26906] = 9
      "001001" when "0110100100011011", -- t[26907] = 9
      "001001" when "0110100100011100", -- t[26908] = 9
      "001001" when "0110100100011101", -- t[26909] = 9
      "001001" when "0110100100011110", -- t[26910] = 9
      "001001" when "0110100100011111", -- t[26911] = 9
      "001001" when "0110100100100000", -- t[26912] = 9
      "001001" when "0110100100100001", -- t[26913] = 9
      "001001" when "0110100100100010", -- t[26914] = 9
      "001001" when "0110100100100011", -- t[26915] = 9
      "001001" when "0110100100100100", -- t[26916] = 9
      "001001" when "0110100100100101", -- t[26917] = 9
      "001001" when "0110100100100110", -- t[26918] = 9
      "001001" when "0110100100100111", -- t[26919] = 9
      "001001" when "0110100100101000", -- t[26920] = 9
      "001001" when "0110100100101001", -- t[26921] = 9
      "001001" when "0110100100101010", -- t[26922] = 9
      "001001" when "0110100100101011", -- t[26923] = 9
      "001001" when "0110100100101100", -- t[26924] = 9
      "001001" when "0110100100101101", -- t[26925] = 9
      "001001" when "0110100100101110", -- t[26926] = 9
      "001001" when "0110100100101111", -- t[26927] = 9
      "001001" when "0110100100110000", -- t[26928] = 9
      "001001" when "0110100100110001", -- t[26929] = 9
      "001001" when "0110100100110010", -- t[26930] = 9
      "001001" when "0110100100110011", -- t[26931] = 9
      "001001" when "0110100100110100", -- t[26932] = 9
      "001001" when "0110100100110101", -- t[26933] = 9
      "001001" when "0110100100110110", -- t[26934] = 9
      "001001" when "0110100100110111", -- t[26935] = 9
      "001001" when "0110100100111000", -- t[26936] = 9
      "001001" when "0110100100111001", -- t[26937] = 9
      "001001" when "0110100100111010", -- t[26938] = 9
      "001001" when "0110100100111011", -- t[26939] = 9
      "001001" when "0110100100111100", -- t[26940] = 9
      "001001" when "0110100100111101", -- t[26941] = 9
      "001001" when "0110100100111110", -- t[26942] = 9
      "001001" when "0110100100111111", -- t[26943] = 9
      "001001" when "0110100101000000", -- t[26944] = 9
      "001001" when "0110100101000001", -- t[26945] = 9
      "001001" when "0110100101000010", -- t[26946] = 9
      "001001" when "0110100101000011", -- t[26947] = 9
      "001001" when "0110100101000100", -- t[26948] = 9
      "001001" when "0110100101000101", -- t[26949] = 9
      "001001" when "0110100101000110", -- t[26950] = 9
      "001001" when "0110100101000111", -- t[26951] = 9
      "001001" when "0110100101001000", -- t[26952] = 9
      "001001" when "0110100101001001", -- t[26953] = 9
      "001001" when "0110100101001010", -- t[26954] = 9
      "001001" when "0110100101001011", -- t[26955] = 9
      "001001" when "0110100101001100", -- t[26956] = 9
      "001001" when "0110100101001101", -- t[26957] = 9
      "001001" when "0110100101001110", -- t[26958] = 9
      "001001" when "0110100101001111", -- t[26959] = 9
      "001001" when "0110100101010000", -- t[26960] = 9
      "001001" when "0110100101010001", -- t[26961] = 9
      "001001" when "0110100101010010", -- t[26962] = 9
      "001001" when "0110100101010011", -- t[26963] = 9
      "001001" when "0110100101010100", -- t[26964] = 9
      "001001" when "0110100101010101", -- t[26965] = 9
      "001001" when "0110100101010110", -- t[26966] = 9
      "001001" when "0110100101010111", -- t[26967] = 9
      "001001" when "0110100101011000", -- t[26968] = 9
      "001001" when "0110100101011001", -- t[26969] = 9
      "001001" when "0110100101011010", -- t[26970] = 9
      "001001" when "0110100101011011", -- t[26971] = 9
      "001001" when "0110100101011100", -- t[26972] = 9
      "001001" when "0110100101011101", -- t[26973] = 9
      "001001" when "0110100101011110", -- t[26974] = 9
      "001001" when "0110100101011111", -- t[26975] = 9
      "001001" when "0110100101100000", -- t[26976] = 9
      "001001" when "0110100101100001", -- t[26977] = 9
      "001001" when "0110100101100010", -- t[26978] = 9
      "001001" when "0110100101100011", -- t[26979] = 9
      "001001" when "0110100101100100", -- t[26980] = 9
      "001001" when "0110100101100101", -- t[26981] = 9
      "001001" when "0110100101100110", -- t[26982] = 9
      "001001" when "0110100101100111", -- t[26983] = 9
      "001001" when "0110100101101000", -- t[26984] = 9
      "001001" when "0110100101101001", -- t[26985] = 9
      "001001" when "0110100101101010", -- t[26986] = 9
      "001001" when "0110100101101011", -- t[26987] = 9
      "001001" when "0110100101101100", -- t[26988] = 9
      "001001" when "0110100101101101", -- t[26989] = 9
      "001001" when "0110100101101110", -- t[26990] = 9
      "001001" when "0110100101101111", -- t[26991] = 9
      "001001" when "0110100101110000", -- t[26992] = 9
      "001001" when "0110100101110001", -- t[26993] = 9
      "001001" when "0110100101110010", -- t[26994] = 9
      "001001" when "0110100101110011", -- t[26995] = 9
      "001001" when "0110100101110100", -- t[26996] = 9
      "001001" when "0110100101110101", -- t[26997] = 9
      "001001" when "0110100101110110", -- t[26998] = 9
      "001001" when "0110100101110111", -- t[26999] = 9
      "001001" when "0110100101111000", -- t[27000] = 9
      "001001" when "0110100101111001", -- t[27001] = 9
      "001001" when "0110100101111010", -- t[27002] = 9
      "001001" when "0110100101111011", -- t[27003] = 9
      "001001" when "0110100101111100", -- t[27004] = 9
      "001001" when "0110100101111101", -- t[27005] = 9
      "001001" when "0110100101111110", -- t[27006] = 9
      "001001" when "0110100101111111", -- t[27007] = 9
      "001001" when "0110100110000000", -- t[27008] = 9
      "001001" when "0110100110000001", -- t[27009] = 9
      "001001" when "0110100110000010", -- t[27010] = 9
      "001001" when "0110100110000011", -- t[27011] = 9
      "001001" when "0110100110000100", -- t[27012] = 9
      "001001" when "0110100110000101", -- t[27013] = 9
      "001001" when "0110100110000110", -- t[27014] = 9
      "001001" when "0110100110000111", -- t[27015] = 9
      "001001" when "0110100110001000", -- t[27016] = 9
      "001001" when "0110100110001001", -- t[27017] = 9
      "001001" when "0110100110001010", -- t[27018] = 9
      "001001" when "0110100110001011", -- t[27019] = 9
      "001001" when "0110100110001100", -- t[27020] = 9
      "001001" when "0110100110001101", -- t[27021] = 9
      "001001" when "0110100110001110", -- t[27022] = 9
      "001001" when "0110100110001111", -- t[27023] = 9
      "001001" when "0110100110010000", -- t[27024] = 9
      "001001" when "0110100110010001", -- t[27025] = 9
      "001001" when "0110100110010010", -- t[27026] = 9
      "001001" when "0110100110010011", -- t[27027] = 9
      "001001" when "0110100110010100", -- t[27028] = 9
      "001001" when "0110100110010101", -- t[27029] = 9
      "001001" when "0110100110010110", -- t[27030] = 9
      "001001" when "0110100110010111", -- t[27031] = 9
      "001001" when "0110100110011000", -- t[27032] = 9
      "001001" when "0110100110011001", -- t[27033] = 9
      "001001" when "0110100110011010", -- t[27034] = 9
      "001001" when "0110100110011011", -- t[27035] = 9
      "001001" when "0110100110011100", -- t[27036] = 9
      "001001" when "0110100110011101", -- t[27037] = 9
      "001001" when "0110100110011110", -- t[27038] = 9
      "001001" when "0110100110011111", -- t[27039] = 9
      "001001" when "0110100110100000", -- t[27040] = 9
      "001001" when "0110100110100001", -- t[27041] = 9
      "001001" when "0110100110100010", -- t[27042] = 9
      "001001" when "0110100110100011", -- t[27043] = 9
      "001001" when "0110100110100100", -- t[27044] = 9
      "001001" when "0110100110100101", -- t[27045] = 9
      "001001" when "0110100110100110", -- t[27046] = 9
      "001001" when "0110100110100111", -- t[27047] = 9
      "001001" when "0110100110101000", -- t[27048] = 9
      "001001" when "0110100110101001", -- t[27049] = 9
      "001001" when "0110100110101010", -- t[27050] = 9
      "001001" when "0110100110101011", -- t[27051] = 9
      "001001" when "0110100110101100", -- t[27052] = 9
      "001001" when "0110100110101101", -- t[27053] = 9
      "001001" when "0110100110101110", -- t[27054] = 9
      "001001" when "0110100110101111", -- t[27055] = 9
      "001001" when "0110100110110000", -- t[27056] = 9
      "001001" when "0110100110110001", -- t[27057] = 9
      "001001" when "0110100110110010", -- t[27058] = 9
      "001001" when "0110100110110011", -- t[27059] = 9
      "001001" when "0110100110110100", -- t[27060] = 9
      "001001" when "0110100110110101", -- t[27061] = 9
      "001001" when "0110100110110110", -- t[27062] = 9
      "001001" when "0110100110110111", -- t[27063] = 9
      "001001" when "0110100110111000", -- t[27064] = 9
      "001001" when "0110100110111001", -- t[27065] = 9
      "001001" when "0110100110111010", -- t[27066] = 9
      "001001" when "0110100110111011", -- t[27067] = 9
      "001001" when "0110100110111100", -- t[27068] = 9
      "001001" when "0110100110111101", -- t[27069] = 9
      "001001" when "0110100110111110", -- t[27070] = 9
      "001001" when "0110100110111111", -- t[27071] = 9
      "001001" when "0110100111000000", -- t[27072] = 9
      "001001" when "0110100111000001", -- t[27073] = 9
      "001001" when "0110100111000010", -- t[27074] = 9
      "001001" when "0110100111000011", -- t[27075] = 9
      "001001" when "0110100111000100", -- t[27076] = 9
      "001001" when "0110100111000101", -- t[27077] = 9
      "001001" when "0110100111000110", -- t[27078] = 9
      "001001" when "0110100111000111", -- t[27079] = 9
      "001001" when "0110100111001000", -- t[27080] = 9
      "001001" when "0110100111001001", -- t[27081] = 9
      "001001" when "0110100111001010", -- t[27082] = 9
      "001001" when "0110100111001011", -- t[27083] = 9
      "001001" when "0110100111001100", -- t[27084] = 9
      "001001" when "0110100111001101", -- t[27085] = 9
      "001001" when "0110100111001110", -- t[27086] = 9
      "001001" when "0110100111001111", -- t[27087] = 9
      "001001" when "0110100111010000", -- t[27088] = 9
      "001001" when "0110100111010001", -- t[27089] = 9
      "001001" when "0110100111010010", -- t[27090] = 9
      "001001" when "0110100111010011", -- t[27091] = 9
      "001001" when "0110100111010100", -- t[27092] = 9
      "001001" when "0110100111010101", -- t[27093] = 9
      "001001" when "0110100111010110", -- t[27094] = 9
      "001001" when "0110100111010111", -- t[27095] = 9
      "001001" when "0110100111011000", -- t[27096] = 9
      "001001" when "0110100111011001", -- t[27097] = 9
      "001001" when "0110100111011010", -- t[27098] = 9
      "001001" when "0110100111011011", -- t[27099] = 9
      "001001" when "0110100111011100", -- t[27100] = 9
      "001001" when "0110100111011101", -- t[27101] = 9
      "001001" when "0110100111011110", -- t[27102] = 9
      "001001" when "0110100111011111", -- t[27103] = 9
      "001001" when "0110100111100000", -- t[27104] = 9
      "001001" when "0110100111100001", -- t[27105] = 9
      "001001" when "0110100111100010", -- t[27106] = 9
      "001001" when "0110100111100011", -- t[27107] = 9
      "001001" when "0110100111100100", -- t[27108] = 9
      "001001" when "0110100111100101", -- t[27109] = 9
      "001001" when "0110100111100110", -- t[27110] = 9
      "001001" when "0110100111100111", -- t[27111] = 9
      "001001" when "0110100111101000", -- t[27112] = 9
      "001001" when "0110100111101001", -- t[27113] = 9
      "001001" when "0110100111101010", -- t[27114] = 9
      "001001" when "0110100111101011", -- t[27115] = 9
      "001001" when "0110100111101100", -- t[27116] = 9
      "001001" when "0110100111101101", -- t[27117] = 9
      "001001" when "0110100111101110", -- t[27118] = 9
      "001001" when "0110100111101111", -- t[27119] = 9
      "001001" when "0110100111110000", -- t[27120] = 9
      "001001" when "0110100111110001", -- t[27121] = 9
      "001001" when "0110100111110010", -- t[27122] = 9
      "001001" when "0110100111110011", -- t[27123] = 9
      "001001" when "0110100111110100", -- t[27124] = 9
      "001001" when "0110100111110101", -- t[27125] = 9
      "001001" when "0110100111110110", -- t[27126] = 9
      "001001" when "0110100111110111", -- t[27127] = 9
      "001001" when "0110100111111000", -- t[27128] = 9
      "001001" when "0110100111111001", -- t[27129] = 9
      "001001" when "0110100111111010", -- t[27130] = 9
      "001001" when "0110100111111011", -- t[27131] = 9
      "001001" when "0110100111111100", -- t[27132] = 9
      "001001" when "0110100111111101", -- t[27133] = 9
      "001001" when "0110100111111110", -- t[27134] = 9
      "001001" when "0110100111111111", -- t[27135] = 9
      "001001" when "0110101000000000", -- t[27136] = 9
      "001001" when "0110101000000001", -- t[27137] = 9
      "001001" when "0110101000000010", -- t[27138] = 9
      "001001" when "0110101000000011", -- t[27139] = 9
      "001001" when "0110101000000100", -- t[27140] = 9
      "001001" when "0110101000000101", -- t[27141] = 9
      "001001" when "0110101000000110", -- t[27142] = 9
      "001001" when "0110101000000111", -- t[27143] = 9
      "001001" when "0110101000001000", -- t[27144] = 9
      "001001" when "0110101000001001", -- t[27145] = 9
      "001001" when "0110101000001010", -- t[27146] = 9
      "001001" when "0110101000001011", -- t[27147] = 9
      "001001" when "0110101000001100", -- t[27148] = 9
      "001001" when "0110101000001101", -- t[27149] = 9
      "001001" when "0110101000001110", -- t[27150] = 9
      "001001" when "0110101000001111", -- t[27151] = 9
      "001001" when "0110101000010000", -- t[27152] = 9
      "001001" when "0110101000010001", -- t[27153] = 9
      "001001" when "0110101000010010", -- t[27154] = 9
      "001001" when "0110101000010011", -- t[27155] = 9
      "001001" when "0110101000010100", -- t[27156] = 9
      "001001" when "0110101000010101", -- t[27157] = 9
      "001001" when "0110101000010110", -- t[27158] = 9
      "001001" when "0110101000010111", -- t[27159] = 9
      "001001" when "0110101000011000", -- t[27160] = 9
      "001001" when "0110101000011001", -- t[27161] = 9
      "001001" when "0110101000011010", -- t[27162] = 9
      "001001" when "0110101000011011", -- t[27163] = 9
      "001001" when "0110101000011100", -- t[27164] = 9
      "001001" when "0110101000011101", -- t[27165] = 9
      "001001" when "0110101000011110", -- t[27166] = 9
      "001001" when "0110101000011111", -- t[27167] = 9
      "001001" when "0110101000100000", -- t[27168] = 9
      "001001" when "0110101000100001", -- t[27169] = 9
      "001001" when "0110101000100010", -- t[27170] = 9
      "001001" when "0110101000100011", -- t[27171] = 9
      "001001" when "0110101000100100", -- t[27172] = 9
      "001001" when "0110101000100101", -- t[27173] = 9
      "001001" when "0110101000100110", -- t[27174] = 9
      "001001" when "0110101000100111", -- t[27175] = 9
      "001001" when "0110101000101000", -- t[27176] = 9
      "001001" when "0110101000101001", -- t[27177] = 9
      "001001" when "0110101000101010", -- t[27178] = 9
      "001001" when "0110101000101011", -- t[27179] = 9
      "001001" when "0110101000101100", -- t[27180] = 9
      "001001" when "0110101000101101", -- t[27181] = 9
      "001001" when "0110101000101110", -- t[27182] = 9
      "001001" when "0110101000101111", -- t[27183] = 9
      "001001" when "0110101000110000", -- t[27184] = 9
      "001001" when "0110101000110001", -- t[27185] = 9
      "001001" when "0110101000110010", -- t[27186] = 9
      "001001" when "0110101000110011", -- t[27187] = 9
      "001001" when "0110101000110100", -- t[27188] = 9
      "001001" when "0110101000110101", -- t[27189] = 9
      "001001" when "0110101000110110", -- t[27190] = 9
      "001001" when "0110101000110111", -- t[27191] = 9
      "001001" when "0110101000111000", -- t[27192] = 9
      "001001" when "0110101000111001", -- t[27193] = 9
      "001001" when "0110101000111010", -- t[27194] = 9
      "001001" when "0110101000111011", -- t[27195] = 9
      "001001" when "0110101000111100", -- t[27196] = 9
      "001001" when "0110101000111101", -- t[27197] = 9
      "001001" when "0110101000111110", -- t[27198] = 9
      "001001" when "0110101000111111", -- t[27199] = 9
      "001001" when "0110101001000000", -- t[27200] = 9
      "001001" when "0110101001000001", -- t[27201] = 9
      "001001" when "0110101001000010", -- t[27202] = 9
      "001001" when "0110101001000011", -- t[27203] = 9
      "001001" when "0110101001000100", -- t[27204] = 9
      "001001" when "0110101001000101", -- t[27205] = 9
      "001001" when "0110101001000110", -- t[27206] = 9
      "001001" when "0110101001000111", -- t[27207] = 9
      "001001" when "0110101001001000", -- t[27208] = 9
      "001001" when "0110101001001001", -- t[27209] = 9
      "001001" when "0110101001001010", -- t[27210] = 9
      "001001" when "0110101001001011", -- t[27211] = 9
      "001001" when "0110101001001100", -- t[27212] = 9
      "001001" when "0110101001001101", -- t[27213] = 9
      "001001" when "0110101001001110", -- t[27214] = 9
      "001001" when "0110101001001111", -- t[27215] = 9
      "001001" when "0110101001010000", -- t[27216] = 9
      "001001" when "0110101001010001", -- t[27217] = 9
      "001001" when "0110101001010010", -- t[27218] = 9
      "001001" when "0110101001010011", -- t[27219] = 9
      "001001" when "0110101001010100", -- t[27220] = 9
      "001001" when "0110101001010101", -- t[27221] = 9
      "001001" when "0110101001010110", -- t[27222] = 9
      "001001" when "0110101001010111", -- t[27223] = 9
      "001001" when "0110101001011000", -- t[27224] = 9
      "001001" when "0110101001011001", -- t[27225] = 9
      "001001" when "0110101001011010", -- t[27226] = 9
      "001001" when "0110101001011011", -- t[27227] = 9
      "001001" when "0110101001011100", -- t[27228] = 9
      "001001" when "0110101001011101", -- t[27229] = 9
      "001001" when "0110101001011110", -- t[27230] = 9
      "001001" when "0110101001011111", -- t[27231] = 9
      "001001" when "0110101001100000", -- t[27232] = 9
      "001001" when "0110101001100001", -- t[27233] = 9
      "001001" when "0110101001100010", -- t[27234] = 9
      "001001" when "0110101001100011", -- t[27235] = 9
      "001001" when "0110101001100100", -- t[27236] = 9
      "001001" when "0110101001100101", -- t[27237] = 9
      "001001" when "0110101001100110", -- t[27238] = 9
      "001001" when "0110101001100111", -- t[27239] = 9
      "001001" when "0110101001101000", -- t[27240] = 9
      "001001" when "0110101001101001", -- t[27241] = 9
      "001001" when "0110101001101010", -- t[27242] = 9
      "001001" when "0110101001101011", -- t[27243] = 9
      "001001" when "0110101001101100", -- t[27244] = 9
      "001001" when "0110101001101101", -- t[27245] = 9
      "001001" when "0110101001101110", -- t[27246] = 9
      "001001" when "0110101001101111", -- t[27247] = 9
      "001001" when "0110101001110000", -- t[27248] = 9
      "001001" when "0110101001110001", -- t[27249] = 9
      "001001" when "0110101001110010", -- t[27250] = 9
      "001001" when "0110101001110011", -- t[27251] = 9
      "001001" when "0110101001110100", -- t[27252] = 9
      "001001" when "0110101001110101", -- t[27253] = 9
      "001001" when "0110101001110110", -- t[27254] = 9
      "001001" when "0110101001110111", -- t[27255] = 9
      "001001" when "0110101001111000", -- t[27256] = 9
      "001001" when "0110101001111001", -- t[27257] = 9
      "001001" when "0110101001111010", -- t[27258] = 9
      "001001" when "0110101001111011", -- t[27259] = 9
      "001001" when "0110101001111100", -- t[27260] = 9
      "001001" when "0110101001111101", -- t[27261] = 9
      "001001" when "0110101001111110", -- t[27262] = 9
      "001001" when "0110101001111111", -- t[27263] = 9
      "001001" when "0110101010000000", -- t[27264] = 9
      "001001" when "0110101010000001", -- t[27265] = 9
      "001001" when "0110101010000010", -- t[27266] = 9
      "001001" when "0110101010000011", -- t[27267] = 9
      "001001" when "0110101010000100", -- t[27268] = 9
      "001001" when "0110101010000101", -- t[27269] = 9
      "001001" when "0110101010000110", -- t[27270] = 9
      "001001" when "0110101010000111", -- t[27271] = 9
      "001001" when "0110101010001000", -- t[27272] = 9
      "001001" when "0110101010001001", -- t[27273] = 9
      "001001" when "0110101010001010", -- t[27274] = 9
      "001001" when "0110101010001011", -- t[27275] = 9
      "001001" when "0110101010001100", -- t[27276] = 9
      "001001" when "0110101010001101", -- t[27277] = 9
      "001001" when "0110101010001110", -- t[27278] = 9
      "001001" when "0110101010001111", -- t[27279] = 9
      "001001" when "0110101010010000", -- t[27280] = 9
      "001001" when "0110101010010001", -- t[27281] = 9
      "001001" when "0110101010010010", -- t[27282] = 9
      "001001" when "0110101010010011", -- t[27283] = 9
      "001001" when "0110101010010100", -- t[27284] = 9
      "001001" when "0110101010010101", -- t[27285] = 9
      "001001" when "0110101010010110", -- t[27286] = 9
      "001001" when "0110101010010111", -- t[27287] = 9
      "001001" when "0110101010011000", -- t[27288] = 9
      "001001" when "0110101010011001", -- t[27289] = 9
      "001001" when "0110101010011010", -- t[27290] = 9
      "001001" when "0110101010011011", -- t[27291] = 9
      "001001" when "0110101010011100", -- t[27292] = 9
      "001001" when "0110101010011101", -- t[27293] = 9
      "001001" when "0110101010011110", -- t[27294] = 9
      "001001" when "0110101010011111", -- t[27295] = 9
      "001001" when "0110101010100000", -- t[27296] = 9
      "001001" when "0110101010100001", -- t[27297] = 9
      "001001" when "0110101010100010", -- t[27298] = 9
      "001001" when "0110101010100011", -- t[27299] = 9
      "001001" when "0110101010100100", -- t[27300] = 9
      "001001" when "0110101010100101", -- t[27301] = 9
      "001001" when "0110101010100110", -- t[27302] = 9
      "001001" when "0110101010100111", -- t[27303] = 9
      "001001" when "0110101010101000", -- t[27304] = 9
      "001001" when "0110101010101001", -- t[27305] = 9
      "001001" when "0110101010101010", -- t[27306] = 9
      "001001" when "0110101010101011", -- t[27307] = 9
      "001001" when "0110101010101100", -- t[27308] = 9
      "001001" when "0110101010101101", -- t[27309] = 9
      "001001" when "0110101010101110", -- t[27310] = 9
      "001001" when "0110101010101111", -- t[27311] = 9
      "001001" when "0110101010110000", -- t[27312] = 9
      "001001" when "0110101010110001", -- t[27313] = 9
      "001001" when "0110101010110010", -- t[27314] = 9
      "001001" when "0110101010110011", -- t[27315] = 9
      "001001" when "0110101010110100", -- t[27316] = 9
      "001001" when "0110101010110101", -- t[27317] = 9
      "001001" when "0110101010110110", -- t[27318] = 9
      "001001" when "0110101010110111", -- t[27319] = 9
      "001001" when "0110101010111000", -- t[27320] = 9
      "001001" when "0110101010111001", -- t[27321] = 9
      "001001" when "0110101010111010", -- t[27322] = 9
      "001001" when "0110101010111011", -- t[27323] = 9
      "001001" when "0110101010111100", -- t[27324] = 9
      "001001" when "0110101010111101", -- t[27325] = 9
      "001001" when "0110101010111110", -- t[27326] = 9
      "001001" when "0110101010111111", -- t[27327] = 9
      "001001" when "0110101011000000", -- t[27328] = 9
      "001001" when "0110101011000001", -- t[27329] = 9
      "001001" when "0110101011000010", -- t[27330] = 9
      "001001" when "0110101011000011", -- t[27331] = 9
      "001001" when "0110101011000100", -- t[27332] = 9
      "001001" when "0110101011000101", -- t[27333] = 9
      "001001" when "0110101011000110", -- t[27334] = 9
      "001001" when "0110101011000111", -- t[27335] = 9
      "001001" when "0110101011001000", -- t[27336] = 9
      "001001" when "0110101011001001", -- t[27337] = 9
      "001001" when "0110101011001010", -- t[27338] = 9
      "001001" when "0110101011001011", -- t[27339] = 9
      "001001" when "0110101011001100", -- t[27340] = 9
      "001001" when "0110101011001101", -- t[27341] = 9
      "001001" when "0110101011001110", -- t[27342] = 9
      "001001" when "0110101011001111", -- t[27343] = 9
      "001001" when "0110101011010000", -- t[27344] = 9
      "001001" when "0110101011010001", -- t[27345] = 9
      "001001" when "0110101011010010", -- t[27346] = 9
      "001001" when "0110101011010011", -- t[27347] = 9
      "001001" when "0110101011010100", -- t[27348] = 9
      "001001" when "0110101011010101", -- t[27349] = 9
      "001001" when "0110101011010110", -- t[27350] = 9
      "001001" when "0110101011010111", -- t[27351] = 9
      "001001" when "0110101011011000", -- t[27352] = 9
      "001001" when "0110101011011001", -- t[27353] = 9
      "001001" when "0110101011011010", -- t[27354] = 9
      "001001" when "0110101011011011", -- t[27355] = 9
      "001001" when "0110101011011100", -- t[27356] = 9
      "001001" when "0110101011011101", -- t[27357] = 9
      "001001" when "0110101011011110", -- t[27358] = 9
      "001001" when "0110101011011111", -- t[27359] = 9
      "001001" when "0110101011100000", -- t[27360] = 9
      "001001" when "0110101011100001", -- t[27361] = 9
      "001001" when "0110101011100010", -- t[27362] = 9
      "001001" when "0110101011100011", -- t[27363] = 9
      "001001" when "0110101011100100", -- t[27364] = 9
      "001001" when "0110101011100101", -- t[27365] = 9
      "001001" when "0110101011100110", -- t[27366] = 9
      "001001" when "0110101011100111", -- t[27367] = 9
      "001001" when "0110101011101000", -- t[27368] = 9
      "001001" when "0110101011101001", -- t[27369] = 9
      "001001" when "0110101011101010", -- t[27370] = 9
      "001001" when "0110101011101011", -- t[27371] = 9
      "001001" when "0110101011101100", -- t[27372] = 9
      "001001" when "0110101011101101", -- t[27373] = 9
      "001001" when "0110101011101110", -- t[27374] = 9
      "001001" when "0110101011101111", -- t[27375] = 9
      "001001" when "0110101011110000", -- t[27376] = 9
      "001001" when "0110101011110001", -- t[27377] = 9
      "001001" when "0110101011110010", -- t[27378] = 9
      "001001" when "0110101011110011", -- t[27379] = 9
      "001001" when "0110101011110100", -- t[27380] = 9
      "001001" when "0110101011110101", -- t[27381] = 9
      "001001" when "0110101011110110", -- t[27382] = 9
      "001001" when "0110101011110111", -- t[27383] = 9
      "001001" when "0110101011111000", -- t[27384] = 9
      "001001" when "0110101011111001", -- t[27385] = 9
      "001001" when "0110101011111010", -- t[27386] = 9
      "001001" when "0110101011111011", -- t[27387] = 9
      "001001" when "0110101011111100", -- t[27388] = 9
      "001001" when "0110101011111101", -- t[27389] = 9
      "001001" when "0110101011111110", -- t[27390] = 9
      "001001" when "0110101011111111", -- t[27391] = 9
      "001001" when "0110101100000000", -- t[27392] = 9
      "001001" when "0110101100000001", -- t[27393] = 9
      "001001" when "0110101100000010", -- t[27394] = 9
      "001001" when "0110101100000011", -- t[27395] = 9
      "001001" when "0110101100000100", -- t[27396] = 9
      "001001" when "0110101100000101", -- t[27397] = 9
      "001001" when "0110101100000110", -- t[27398] = 9
      "001001" when "0110101100000111", -- t[27399] = 9
      "001001" when "0110101100001000", -- t[27400] = 9
      "001001" when "0110101100001001", -- t[27401] = 9
      "001001" when "0110101100001010", -- t[27402] = 9
      "001001" when "0110101100001011", -- t[27403] = 9
      "001001" when "0110101100001100", -- t[27404] = 9
      "001001" when "0110101100001101", -- t[27405] = 9
      "001001" when "0110101100001110", -- t[27406] = 9
      "001001" when "0110101100001111", -- t[27407] = 9
      "001001" when "0110101100010000", -- t[27408] = 9
      "001001" when "0110101100010001", -- t[27409] = 9
      "001001" when "0110101100010010", -- t[27410] = 9
      "001001" when "0110101100010011", -- t[27411] = 9
      "001001" when "0110101100010100", -- t[27412] = 9
      "001001" when "0110101100010101", -- t[27413] = 9
      "001001" when "0110101100010110", -- t[27414] = 9
      "001001" when "0110101100010111", -- t[27415] = 9
      "001001" when "0110101100011000", -- t[27416] = 9
      "001001" when "0110101100011001", -- t[27417] = 9
      "001001" when "0110101100011010", -- t[27418] = 9
      "001001" when "0110101100011011", -- t[27419] = 9
      "001001" when "0110101100011100", -- t[27420] = 9
      "001001" when "0110101100011101", -- t[27421] = 9
      "001001" when "0110101100011110", -- t[27422] = 9
      "001001" when "0110101100011111", -- t[27423] = 9
      "001001" when "0110101100100000", -- t[27424] = 9
      "001001" when "0110101100100001", -- t[27425] = 9
      "001001" when "0110101100100010", -- t[27426] = 9
      "001001" when "0110101100100011", -- t[27427] = 9
      "001001" when "0110101100100100", -- t[27428] = 9
      "001001" when "0110101100100101", -- t[27429] = 9
      "001001" when "0110101100100110", -- t[27430] = 9
      "001001" when "0110101100100111", -- t[27431] = 9
      "001001" when "0110101100101000", -- t[27432] = 9
      "001001" when "0110101100101001", -- t[27433] = 9
      "001001" when "0110101100101010", -- t[27434] = 9
      "001001" when "0110101100101011", -- t[27435] = 9
      "001001" when "0110101100101100", -- t[27436] = 9
      "001001" when "0110101100101101", -- t[27437] = 9
      "001001" when "0110101100101110", -- t[27438] = 9
      "001001" when "0110101100101111", -- t[27439] = 9
      "001001" when "0110101100110000", -- t[27440] = 9
      "001001" when "0110101100110001", -- t[27441] = 9
      "001001" when "0110101100110010", -- t[27442] = 9
      "001001" when "0110101100110011", -- t[27443] = 9
      "001001" when "0110101100110100", -- t[27444] = 9
      "001001" when "0110101100110101", -- t[27445] = 9
      "001001" when "0110101100110110", -- t[27446] = 9
      "001001" when "0110101100110111", -- t[27447] = 9
      "001001" when "0110101100111000", -- t[27448] = 9
      "001001" when "0110101100111001", -- t[27449] = 9
      "001001" when "0110101100111010", -- t[27450] = 9
      "001001" when "0110101100111011", -- t[27451] = 9
      "001001" when "0110101100111100", -- t[27452] = 9
      "001001" when "0110101100111101", -- t[27453] = 9
      "001001" when "0110101100111110", -- t[27454] = 9
      "001001" when "0110101100111111", -- t[27455] = 9
      "001001" when "0110101101000000", -- t[27456] = 9
      "001001" when "0110101101000001", -- t[27457] = 9
      "001001" when "0110101101000010", -- t[27458] = 9
      "001001" when "0110101101000011", -- t[27459] = 9
      "001001" when "0110101101000100", -- t[27460] = 9
      "001001" when "0110101101000101", -- t[27461] = 9
      "001001" when "0110101101000110", -- t[27462] = 9
      "001001" when "0110101101000111", -- t[27463] = 9
      "001001" when "0110101101001000", -- t[27464] = 9
      "001001" when "0110101101001001", -- t[27465] = 9
      "001001" when "0110101101001010", -- t[27466] = 9
      "001001" when "0110101101001011", -- t[27467] = 9
      "001001" when "0110101101001100", -- t[27468] = 9
      "001001" when "0110101101001101", -- t[27469] = 9
      "001001" when "0110101101001110", -- t[27470] = 9
      "001001" when "0110101101001111", -- t[27471] = 9
      "001001" when "0110101101010000", -- t[27472] = 9
      "001001" when "0110101101010001", -- t[27473] = 9
      "001001" when "0110101101010010", -- t[27474] = 9
      "001001" when "0110101101010011", -- t[27475] = 9
      "001001" when "0110101101010100", -- t[27476] = 9
      "001001" when "0110101101010101", -- t[27477] = 9
      "001001" when "0110101101010110", -- t[27478] = 9
      "001001" when "0110101101010111", -- t[27479] = 9
      "001001" when "0110101101011000", -- t[27480] = 9
      "001001" when "0110101101011001", -- t[27481] = 9
      "001001" when "0110101101011010", -- t[27482] = 9
      "001001" when "0110101101011011", -- t[27483] = 9
      "001001" when "0110101101011100", -- t[27484] = 9
      "001001" when "0110101101011101", -- t[27485] = 9
      "001001" when "0110101101011110", -- t[27486] = 9
      "001001" when "0110101101011111", -- t[27487] = 9
      "001001" when "0110101101100000", -- t[27488] = 9
      "001001" when "0110101101100001", -- t[27489] = 9
      "001001" when "0110101101100010", -- t[27490] = 9
      "001001" when "0110101101100011", -- t[27491] = 9
      "001001" when "0110101101100100", -- t[27492] = 9
      "001001" when "0110101101100101", -- t[27493] = 9
      "001001" when "0110101101100110", -- t[27494] = 9
      "001001" when "0110101101100111", -- t[27495] = 9
      "001001" when "0110101101101000", -- t[27496] = 9
      "001001" when "0110101101101001", -- t[27497] = 9
      "001001" when "0110101101101010", -- t[27498] = 9
      "001001" when "0110101101101011", -- t[27499] = 9
      "001001" when "0110101101101100", -- t[27500] = 9
      "001001" when "0110101101101101", -- t[27501] = 9
      "001001" when "0110101101101110", -- t[27502] = 9
      "001001" when "0110101101101111", -- t[27503] = 9
      "001001" when "0110101101110000", -- t[27504] = 9
      "001001" when "0110101101110001", -- t[27505] = 9
      "001001" when "0110101101110010", -- t[27506] = 9
      "001001" when "0110101101110011", -- t[27507] = 9
      "001001" when "0110101101110100", -- t[27508] = 9
      "001001" when "0110101101110101", -- t[27509] = 9
      "001001" when "0110101101110110", -- t[27510] = 9
      "001001" when "0110101101110111", -- t[27511] = 9
      "001001" when "0110101101111000", -- t[27512] = 9
      "001001" when "0110101101111001", -- t[27513] = 9
      "001001" when "0110101101111010", -- t[27514] = 9
      "001001" when "0110101101111011", -- t[27515] = 9
      "001001" when "0110101101111100", -- t[27516] = 9
      "001010" when "0110101101111101", -- t[27517] = 10
      "001010" when "0110101101111110", -- t[27518] = 10
      "001010" when "0110101101111111", -- t[27519] = 10
      "001010" when "0110101110000000", -- t[27520] = 10
      "001010" when "0110101110000001", -- t[27521] = 10
      "001010" when "0110101110000010", -- t[27522] = 10
      "001010" when "0110101110000011", -- t[27523] = 10
      "001010" when "0110101110000100", -- t[27524] = 10
      "001010" when "0110101110000101", -- t[27525] = 10
      "001010" when "0110101110000110", -- t[27526] = 10
      "001010" when "0110101110000111", -- t[27527] = 10
      "001010" when "0110101110001000", -- t[27528] = 10
      "001010" when "0110101110001001", -- t[27529] = 10
      "001010" when "0110101110001010", -- t[27530] = 10
      "001010" when "0110101110001011", -- t[27531] = 10
      "001010" when "0110101110001100", -- t[27532] = 10
      "001010" when "0110101110001101", -- t[27533] = 10
      "001010" when "0110101110001110", -- t[27534] = 10
      "001010" when "0110101110001111", -- t[27535] = 10
      "001010" when "0110101110010000", -- t[27536] = 10
      "001010" when "0110101110010001", -- t[27537] = 10
      "001010" when "0110101110010010", -- t[27538] = 10
      "001010" when "0110101110010011", -- t[27539] = 10
      "001010" when "0110101110010100", -- t[27540] = 10
      "001010" when "0110101110010101", -- t[27541] = 10
      "001010" when "0110101110010110", -- t[27542] = 10
      "001010" when "0110101110010111", -- t[27543] = 10
      "001010" when "0110101110011000", -- t[27544] = 10
      "001010" when "0110101110011001", -- t[27545] = 10
      "001010" when "0110101110011010", -- t[27546] = 10
      "001010" when "0110101110011011", -- t[27547] = 10
      "001010" when "0110101110011100", -- t[27548] = 10
      "001010" when "0110101110011101", -- t[27549] = 10
      "001010" when "0110101110011110", -- t[27550] = 10
      "001010" when "0110101110011111", -- t[27551] = 10
      "001010" when "0110101110100000", -- t[27552] = 10
      "001010" when "0110101110100001", -- t[27553] = 10
      "001010" when "0110101110100010", -- t[27554] = 10
      "001010" when "0110101110100011", -- t[27555] = 10
      "001010" when "0110101110100100", -- t[27556] = 10
      "001010" when "0110101110100101", -- t[27557] = 10
      "001010" when "0110101110100110", -- t[27558] = 10
      "001010" when "0110101110100111", -- t[27559] = 10
      "001010" when "0110101110101000", -- t[27560] = 10
      "001010" when "0110101110101001", -- t[27561] = 10
      "001010" when "0110101110101010", -- t[27562] = 10
      "001010" when "0110101110101011", -- t[27563] = 10
      "001010" when "0110101110101100", -- t[27564] = 10
      "001010" when "0110101110101101", -- t[27565] = 10
      "001010" when "0110101110101110", -- t[27566] = 10
      "001010" when "0110101110101111", -- t[27567] = 10
      "001010" when "0110101110110000", -- t[27568] = 10
      "001010" when "0110101110110001", -- t[27569] = 10
      "001010" when "0110101110110010", -- t[27570] = 10
      "001010" when "0110101110110011", -- t[27571] = 10
      "001010" when "0110101110110100", -- t[27572] = 10
      "001010" when "0110101110110101", -- t[27573] = 10
      "001010" when "0110101110110110", -- t[27574] = 10
      "001010" when "0110101110110111", -- t[27575] = 10
      "001010" when "0110101110111000", -- t[27576] = 10
      "001010" when "0110101110111001", -- t[27577] = 10
      "001010" when "0110101110111010", -- t[27578] = 10
      "001010" when "0110101110111011", -- t[27579] = 10
      "001010" when "0110101110111100", -- t[27580] = 10
      "001010" when "0110101110111101", -- t[27581] = 10
      "001010" when "0110101110111110", -- t[27582] = 10
      "001010" when "0110101110111111", -- t[27583] = 10
      "001010" when "0110101111000000", -- t[27584] = 10
      "001010" when "0110101111000001", -- t[27585] = 10
      "001010" when "0110101111000010", -- t[27586] = 10
      "001010" when "0110101111000011", -- t[27587] = 10
      "001010" when "0110101111000100", -- t[27588] = 10
      "001010" when "0110101111000101", -- t[27589] = 10
      "001010" when "0110101111000110", -- t[27590] = 10
      "001010" when "0110101111000111", -- t[27591] = 10
      "001010" when "0110101111001000", -- t[27592] = 10
      "001010" when "0110101111001001", -- t[27593] = 10
      "001010" when "0110101111001010", -- t[27594] = 10
      "001010" when "0110101111001011", -- t[27595] = 10
      "001010" when "0110101111001100", -- t[27596] = 10
      "001010" when "0110101111001101", -- t[27597] = 10
      "001010" when "0110101111001110", -- t[27598] = 10
      "001010" when "0110101111001111", -- t[27599] = 10
      "001010" when "0110101111010000", -- t[27600] = 10
      "001010" when "0110101111010001", -- t[27601] = 10
      "001010" when "0110101111010010", -- t[27602] = 10
      "001010" when "0110101111010011", -- t[27603] = 10
      "001010" when "0110101111010100", -- t[27604] = 10
      "001010" when "0110101111010101", -- t[27605] = 10
      "001010" when "0110101111010110", -- t[27606] = 10
      "001010" when "0110101111010111", -- t[27607] = 10
      "001010" when "0110101111011000", -- t[27608] = 10
      "001010" when "0110101111011001", -- t[27609] = 10
      "001010" when "0110101111011010", -- t[27610] = 10
      "001010" when "0110101111011011", -- t[27611] = 10
      "001010" when "0110101111011100", -- t[27612] = 10
      "001010" when "0110101111011101", -- t[27613] = 10
      "001010" when "0110101111011110", -- t[27614] = 10
      "001010" when "0110101111011111", -- t[27615] = 10
      "001010" when "0110101111100000", -- t[27616] = 10
      "001010" when "0110101111100001", -- t[27617] = 10
      "001010" when "0110101111100010", -- t[27618] = 10
      "001010" when "0110101111100011", -- t[27619] = 10
      "001010" when "0110101111100100", -- t[27620] = 10
      "001010" when "0110101111100101", -- t[27621] = 10
      "001010" when "0110101111100110", -- t[27622] = 10
      "001010" when "0110101111100111", -- t[27623] = 10
      "001010" when "0110101111101000", -- t[27624] = 10
      "001010" when "0110101111101001", -- t[27625] = 10
      "001010" when "0110101111101010", -- t[27626] = 10
      "001010" when "0110101111101011", -- t[27627] = 10
      "001010" when "0110101111101100", -- t[27628] = 10
      "001010" when "0110101111101101", -- t[27629] = 10
      "001010" when "0110101111101110", -- t[27630] = 10
      "001010" when "0110101111101111", -- t[27631] = 10
      "001010" when "0110101111110000", -- t[27632] = 10
      "001010" when "0110101111110001", -- t[27633] = 10
      "001010" when "0110101111110010", -- t[27634] = 10
      "001010" when "0110101111110011", -- t[27635] = 10
      "001010" when "0110101111110100", -- t[27636] = 10
      "001010" when "0110101111110101", -- t[27637] = 10
      "001010" when "0110101111110110", -- t[27638] = 10
      "001010" when "0110101111110111", -- t[27639] = 10
      "001010" when "0110101111111000", -- t[27640] = 10
      "001010" when "0110101111111001", -- t[27641] = 10
      "001010" when "0110101111111010", -- t[27642] = 10
      "001010" when "0110101111111011", -- t[27643] = 10
      "001010" when "0110101111111100", -- t[27644] = 10
      "001010" when "0110101111111101", -- t[27645] = 10
      "001010" when "0110101111111110", -- t[27646] = 10
      "001010" when "0110101111111111", -- t[27647] = 10
      "001010" when "0110110000000000", -- t[27648] = 10
      "001010" when "0110110000000001", -- t[27649] = 10
      "001010" when "0110110000000010", -- t[27650] = 10
      "001010" when "0110110000000011", -- t[27651] = 10
      "001010" when "0110110000000100", -- t[27652] = 10
      "001010" when "0110110000000101", -- t[27653] = 10
      "001010" when "0110110000000110", -- t[27654] = 10
      "001010" when "0110110000000111", -- t[27655] = 10
      "001010" when "0110110000001000", -- t[27656] = 10
      "001010" when "0110110000001001", -- t[27657] = 10
      "001010" when "0110110000001010", -- t[27658] = 10
      "001010" when "0110110000001011", -- t[27659] = 10
      "001010" when "0110110000001100", -- t[27660] = 10
      "001010" when "0110110000001101", -- t[27661] = 10
      "001010" when "0110110000001110", -- t[27662] = 10
      "001010" when "0110110000001111", -- t[27663] = 10
      "001010" when "0110110000010000", -- t[27664] = 10
      "001010" when "0110110000010001", -- t[27665] = 10
      "001010" when "0110110000010010", -- t[27666] = 10
      "001010" when "0110110000010011", -- t[27667] = 10
      "001010" when "0110110000010100", -- t[27668] = 10
      "001010" when "0110110000010101", -- t[27669] = 10
      "001010" when "0110110000010110", -- t[27670] = 10
      "001010" when "0110110000010111", -- t[27671] = 10
      "001010" when "0110110000011000", -- t[27672] = 10
      "001010" when "0110110000011001", -- t[27673] = 10
      "001010" when "0110110000011010", -- t[27674] = 10
      "001010" when "0110110000011011", -- t[27675] = 10
      "001010" when "0110110000011100", -- t[27676] = 10
      "001010" when "0110110000011101", -- t[27677] = 10
      "001010" when "0110110000011110", -- t[27678] = 10
      "001010" when "0110110000011111", -- t[27679] = 10
      "001010" when "0110110000100000", -- t[27680] = 10
      "001010" when "0110110000100001", -- t[27681] = 10
      "001010" when "0110110000100010", -- t[27682] = 10
      "001010" when "0110110000100011", -- t[27683] = 10
      "001010" when "0110110000100100", -- t[27684] = 10
      "001010" when "0110110000100101", -- t[27685] = 10
      "001010" when "0110110000100110", -- t[27686] = 10
      "001010" when "0110110000100111", -- t[27687] = 10
      "001010" when "0110110000101000", -- t[27688] = 10
      "001010" when "0110110000101001", -- t[27689] = 10
      "001010" when "0110110000101010", -- t[27690] = 10
      "001010" when "0110110000101011", -- t[27691] = 10
      "001010" when "0110110000101100", -- t[27692] = 10
      "001010" when "0110110000101101", -- t[27693] = 10
      "001010" when "0110110000101110", -- t[27694] = 10
      "001010" when "0110110000101111", -- t[27695] = 10
      "001010" when "0110110000110000", -- t[27696] = 10
      "001010" when "0110110000110001", -- t[27697] = 10
      "001010" when "0110110000110010", -- t[27698] = 10
      "001010" when "0110110000110011", -- t[27699] = 10
      "001010" when "0110110000110100", -- t[27700] = 10
      "001010" when "0110110000110101", -- t[27701] = 10
      "001010" when "0110110000110110", -- t[27702] = 10
      "001010" when "0110110000110111", -- t[27703] = 10
      "001010" when "0110110000111000", -- t[27704] = 10
      "001010" when "0110110000111001", -- t[27705] = 10
      "001010" when "0110110000111010", -- t[27706] = 10
      "001010" when "0110110000111011", -- t[27707] = 10
      "001010" when "0110110000111100", -- t[27708] = 10
      "001010" when "0110110000111101", -- t[27709] = 10
      "001010" when "0110110000111110", -- t[27710] = 10
      "001010" when "0110110000111111", -- t[27711] = 10
      "001010" when "0110110001000000", -- t[27712] = 10
      "001010" when "0110110001000001", -- t[27713] = 10
      "001010" when "0110110001000010", -- t[27714] = 10
      "001010" when "0110110001000011", -- t[27715] = 10
      "001010" when "0110110001000100", -- t[27716] = 10
      "001010" when "0110110001000101", -- t[27717] = 10
      "001010" when "0110110001000110", -- t[27718] = 10
      "001010" when "0110110001000111", -- t[27719] = 10
      "001010" when "0110110001001000", -- t[27720] = 10
      "001010" when "0110110001001001", -- t[27721] = 10
      "001010" when "0110110001001010", -- t[27722] = 10
      "001010" when "0110110001001011", -- t[27723] = 10
      "001010" when "0110110001001100", -- t[27724] = 10
      "001010" when "0110110001001101", -- t[27725] = 10
      "001010" when "0110110001001110", -- t[27726] = 10
      "001010" when "0110110001001111", -- t[27727] = 10
      "001010" when "0110110001010000", -- t[27728] = 10
      "001010" when "0110110001010001", -- t[27729] = 10
      "001010" when "0110110001010010", -- t[27730] = 10
      "001010" when "0110110001010011", -- t[27731] = 10
      "001010" when "0110110001010100", -- t[27732] = 10
      "001010" when "0110110001010101", -- t[27733] = 10
      "001010" when "0110110001010110", -- t[27734] = 10
      "001010" when "0110110001010111", -- t[27735] = 10
      "001010" when "0110110001011000", -- t[27736] = 10
      "001010" when "0110110001011001", -- t[27737] = 10
      "001010" when "0110110001011010", -- t[27738] = 10
      "001010" when "0110110001011011", -- t[27739] = 10
      "001010" when "0110110001011100", -- t[27740] = 10
      "001010" when "0110110001011101", -- t[27741] = 10
      "001010" when "0110110001011110", -- t[27742] = 10
      "001010" when "0110110001011111", -- t[27743] = 10
      "001010" when "0110110001100000", -- t[27744] = 10
      "001010" when "0110110001100001", -- t[27745] = 10
      "001010" when "0110110001100010", -- t[27746] = 10
      "001010" when "0110110001100011", -- t[27747] = 10
      "001010" when "0110110001100100", -- t[27748] = 10
      "001010" when "0110110001100101", -- t[27749] = 10
      "001010" when "0110110001100110", -- t[27750] = 10
      "001010" when "0110110001100111", -- t[27751] = 10
      "001010" when "0110110001101000", -- t[27752] = 10
      "001010" when "0110110001101001", -- t[27753] = 10
      "001010" when "0110110001101010", -- t[27754] = 10
      "001010" when "0110110001101011", -- t[27755] = 10
      "001010" when "0110110001101100", -- t[27756] = 10
      "001010" when "0110110001101101", -- t[27757] = 10
      "001010" when "0110110001101110", -- t[27758] = 10
      "001010" when "0110110001101111", -- t[27759] = 10
      "001010" when "0110110001110000", -- t[27760] = 10
      "001010" when "0110110001110001", -- t[27761] = 10
      "001010" when "0110110001110010", -- t[27762] = 10
      "001010" when "0110110001110011", -- t[27763] = 10
      "001010" when "0110110001110100", -- t[27764] = 10
      "001010" when "0110110001110101", -- t[27765] = 10
      "001010" when "0110110001110110", -- t[27766] = 10
      "001010" when "0110110001110111", -- t[27767] = 10
      "001010" when "0110110001111000", -- t[27768] = 10
      "001010" when "0110110001111001", -- t[27769] = 10
      "001010" when "0110110001111010", -- t[27770] = 10
      "001010" when "0110110001111011", -- t[27771] = 10
      "001010" when "0110110001111100", -- t[27772] = 10
      "001010" when "0110110001111101", -- t[27773] = 10
      "001010" when "0110110001111110", -- t[27774] = 10
      "001010" when "0110110001111111", -- t[27775] = 10
      "001010" when "0110110010000000", -- t[27776] = 10
      "001010" when "0110110010000001", -- t[27777] = 10
      "001010" when "0110110010000010", -- t[27778] = 10
      "001010" when "0110110010000011", -- t[27779] = 10
      "001010" when "0110110010000100", -- t[27780] = 10
      "001010" when "0110110010000101", -- t[27781] = 10
      "001010" when "0110110010000110", -- t[27782] = 10
      "001010" when "0110110010000111", -- t[27783] = 10
      "001010" when "0110110010001000", -- t[27784] = 10
      "001010" when "0110110010001001", -- t[27785] = 10
      "001010" when "0110110010001010", -- t[27786] = 10
      "001010" when "0110110010001011", -- t[27787] = 10
      "001010" when "0110110010001100", -- t[27788] = 10
      "001010" when "0110110010001101", -- t[27789] = 10
      "001010" when "0110110010001110", -- t[27790] = 10
      "001010" when "0110110010001111", -- t[27791] = 10
      "001010" when "0110110010010000", -- t[27792] = 10
      "001010" when "0110110010010001", -- t[27793] = 10
      "001010" when "0110110010010010", -- t[27794] = 10
      "001010" when "0110110010010011", -- t[27795] = 10
      "001010" when "0110110010010100", -- t[27796] = 10
      "001010" when "0110110010010101", -- t[27797] = 10
      "001010" when "0110110010010110", -- t[27798] = 10
      "001010" when "0110110010010111", -- t[27799] = 10
      "001010" when "0110110010011000", -- t[27800] = 10
      "001010" when "0110110010011001", -- t[27801] = 10
      "001010" when "0110110010011010", -- t[27802] = 10
      "001010" when "0110110010011011", -- t[27803] = 10
      "001010" when "0110110010011100", -- t[27804] = 10
      "001010" when "0110110010011101", -- t[27805] = 10
      "001010" when "0110110010011110", -- t[27806] = 10
      "001010" when "0110110010011111", -- t[27807] = 10
      "001010" when "0110110010100000", -- t[27808] = 10
      "001010" when "0110110010100001", -- t[27809] = 10
      "001010" when "0110110010100010", -- t[27810] = 10
      "001010" when "0110110010100011", -- t[27811] = 10
      "001010" when "0110110010100100", -- t[27812] = 10
      "001010" when "0110110010100101", -- t[27813] = 10
      "001010" when "0110110010100110", -- t[27814] = 10
      "001010" when "0110110010100111", -- t[27815] = 10
      "001010" when "0110110010101000", -- t[27816] = 10
      "001010" when "0110110010101001", -- t[27817] = 10
      "001010" when "0110110010101010", -- t[27818] = 10
      "001010" when "0110110010101011", -- t[27819] = 10
      "001010" when "0110110010101100", -- t[27820] = 10
      "001010" when "0110110010101101", -- t[27821] = 10
      "001010" when "0110110010101110", -- t[27822] = 10
      "001010" when "0110110010101111", -- t[27823] = 10
      "001010" when "0110110010110000", -- t[27824] = 10
      "001010" when "0110110010110001", -- t[27825] = 10
      "001010" when "0110110010110010", -- t[27826] = 10
      "001010" when "0110110010110011", -- t[27827] = 10
      "001010" when "0110110010110100", -- t[27828] = 10
      "001010" when "0110110010110101", -- t[27829] = 10
      "001010" when "0110110010110110", -- t[27830] = 10
      "001010" when "0110110010110111", -- t[27831] = 10
      "001010" when "0110110010111000", -- t[27832] = 10
      "001010" when "0110110010111001", -- t[27833] = 10
      "001010" when "0110110010111010", -- t[27834] = 10
      "001010" when "0110110010111011", -- t[27835] = 10
      "001010" when "0110110010111100", -- t[27836] = 10
      "001010" when "0110110010111101", -- t[27837] = 10
      "001010" when "0110110010111110", -- t[27838] = 10
      "001010" when "0110110010111111", -- t[27839] = 10
      "001010" when "0110110011000000", -- t[27840] = 10
      "001010" when "0110110011000001", -- t[27841] = 10
      "001010" when "0110110011000010", -- t[27842] = 10
      "001010" when "0110110011000011", -- t[27843] = 10
      "001010" when "0110110011000100", -- t[27844] = 10
      "001010" when "0110110011000101", -- t[27845] = 10
      "001010" when "0110110011000110", -- t[27846] = 10
      "001010" when "0110110011000111", -- t[27847] = 10
      "001010" when "0110110011001000", -- t[27848] = 10
      "001010" when "0110110011001001", -- t[27849] = 10
      "001010" when "0110110011001010", -- t[27850] = 10
      "001010" when "0110110011001011", -- t[27851] = 10
      "001010" when "0110110011001100", -- t[27852] = 10
      "001010" when "0110110011001101", -- t[27853] = 10
      "001010" when "0110110011001110", -- t[27854] = 10
      "001010" when "0110110011001111", -- t[27855] = 10
      "001010" when "0110110011010000", -- t[27856] = 10
      "001010" when "0110110011010001", -- t[27857] = 10
      "001010" when "0110110011010010", -- t[27858] = 10
      "001010" when "0110110011010011", -- t[27859] = 10
      "001010" when "0110110011010100", -- t[27860] = 10
      "001010" when "0110110011010101", -- t[27861] = 10
      "001010" when "0110110011010110", -- t[27862] = 10
      "001010" when "0110110011010111", -- t[27863] = 10
      "001010" when "0110110011011000", -- t[27864] = 10
      "001010" when "0110110011011001", -- t[27865] = 10
      "001010" when "0110110011011010", -- t[27866] = 10
      "001010" when "0110110011011011", -- t[27867] = 10
      "001010" when "0110110011011100", -- t[27868] = 10
      "001010" when "0110110011011101", -- t[27869] = 10
      "001010" when "0110110011011110", -- t[27870] = 10
      "001010" when "0110110011011111", -- t[27871] = 10
      "001010" when "0110110011100000", -- t[27872] = 10
      "001010" when "0110110011100001", -- t[27873] = 10
      "001010" when "0110110011100010", -- t[27874] = 10
      "001010" when "0110110011100011", -- t[27875] = 10
      "001010" when "0110110011100100", -- t[27876] = 10
      "001010" when "0110110011100101", -- t[27877] = 10
      "001010" when "0110110011100110", -- t[27878] = 10
      "001010" when "0110110011100111", -- t[27879] = 10
      "001010" when "0110110011101000", -- t[27880] = 10
      "001010" when "0110110011101001", -- t[27881] = 10
      "001010" when "0110110011101010", -- t[27882] = 10
      "001010" when "0110110011101011", -- t[27883] = 10
      "001010" when "0110110011101100", -- t[27884] = 10
      "001010" when "0110110011101101", -- t[27885] = 10
      "001010" when "0110110011101110", -- t[27886] = 10
      "001010" when "0110110011101111", -- t[27887] = 10
      "001010" when "0110110011110000", -- t[27888] = 10
      "001010" when "0110110011110001", -- t[27889] = 10
      "001010" when "0110110011110010", -- t[27890] = 10
      "001010" when "0110110011110011", -- t[27891] = 10
      "001010" when "0110110011110100", -- t[27892] = 10
      "001010" when "0110110011110101", -- t[27893] = 10
      "001010" when "0110110011110110", -- t[27894] = 10
      "001010" when "0110110011110111", -- t[27895] = 10
      "001010" when "0110110011111000", -- t[27896] = 10
      "001010" when "0110110011111001", -- t[27897] = 10
      "001010" when "0110110011111010", -- t[27898] = 10
      "001010" when "0110110011111011", -- t[27899] = 10
      "001010" when "0110110011111100", -- t[27900] = 10
      "001010" when "0110110011111101", -- t[27901] = 10
      "001010" when "0110110011111110", -- t[27902] = 10
      "001010" when "0110110011111111", -- t[27903] = 10
      "001010" when "0110110100000000", -- t[27904] = 10
      "001010" when "0110110100000001", -- t[27905] = 10
      "001010" when "0110110100000010", -- t[27906] = 10
      "001010" when "0110110100000011", -- t[27907] = 10
      "001010" when "0110110100000100", -- t[27908] = 10
      "001010" when "0110110100000101", -- t[27909] = 10
      "001010" when "0110110100000110", -- t[27910] = 10
      "001010" when "0110110100000111", -- t[27911] = 10
      "001010" when "0110110100001000", -- t[27912] = 10
      "001010" when "0110110100001001", -- t[27913] = 10
      "001010" when "0110110100001010", -- t[27914] = 10
      "001010" when "0110110100001011", -- t[27915] = 10
      "001010" when "0110110100001100", -- t[27916] = 10
      "001010" when "0110110100001101", -- t[27917] = 10
      "001010" when "0110110100001110", -- t[27918] = 10
      "001010" when "0110110100001111", -- t[27919] = 10
      "001010" when "0110110100010000", -- t[27920] = 10
      "001010" when "0110110100010001", -- t[27921] = 10
      "001010" when "0110110100010010", -- t[27922] = 10
      "001010" when "0110110100010011", -- t[27923] = 10
      "001010" when "0110110100010100", -- t[27924] = 10
      "001010" when "0110110100010101", -- t[27925] = 10
      "001010" when "0110110100010110", -- t[27926] = 10
      "001010" when "0110110100010111", -- t[27927] = 10
      "001010" when "0110110100011000", -- t[27928] = 10
      "001010" when "0110110100011001", -- t[27929] = 10
      "001010" when "0110110100011010", -- t[27930] = 10
      "001010" when "0110110100011011", -- t[27931] = 10
      "001010" when "0110110100011100", -- t[27932] = 10
      "001010" when "0110110100011101", -- t[27933] = 10
      "001010" when "0110110100011110", -- t[27934] = 10
      "001010" when "0110110100011111", -- t[27935] = 10
      "001010" when "0110110100100000", -- t[27936] = 10
      "001010" when "0110110100100001", -- t[27937] = 10
      "001010" when "0110110100100010", -- t[27938] = 10
      "001010" when "0110110100100011", -- t[27939] = 10
      "001010" when "0110110100100100", -- t[27940] = 10
      "001010" when "0110110100100101", -- t[27941] = 10
      "001010" when "0110110100100110", -- t[27942] = 10
      "001010" when "0110110100100111", -- t[27943] = 10
      "001010" when "0110110100101000", -- t[27944] = 10
      "001010" when "0110110100101001", -- t[27945] = 10
      "001010" when "0110110100101010", -- t[27946] = 10
      "001010" when "0110110100101011", -- t[27947] = 10
      "001010" when "0110110100101100", -- t[27948] = 10
      "001010" when "0110110100101101", -- t[27949] = 10
      "001010" when "0110110100101110", -- t[27950] = 10
      "001010" when "0110110100101111", -- t[27951] = 10
      "001010" when "0110110100110000", -- t[27952] = 10
      "001010" when "0110110100110001", -- t[27953] = 10
      "001010" when "0110110100110010", -- t[27954] = 10
      "001010" when "0110110100110011", -- t[27955] = 10
      "001010" when "0110110100110100", -- t[27956] = 10
      "001010" when "0110110100110101", -- t[27957] = 10
      "001010" when "0110110100110110", -- t[27958] = 10
      "001010" when "0110110100110111", -- t[27959] = 10
      "001010" when "0110110100111000", -- t[27960] = 10
      "001010" when "0110110100111001", -- t[27961] = 10
      "001010" when "0110110100111010", -- t[27962] = 10
      "001010" when "0110110100111011", -- t[27963] = 10
      "001010" when "0110110100111100", -- t[27964] = 10
      "001010" when "0110110100111101", -- t[27965] = 10
      "001010" when "0110110100111110", -- t[27966] = 10
      "001010" when "0110110100111111", -- t[27967] = 10
      "001010" when "0110110101000000", -- t[27968] = 10
      "001010" when "0110110101000001", -- t[27969] = 10
      "001010" when "0110110101000010", -- t[27970] = 10
      "001010" when "0110110101000011", -- t[27971] = 10
      "001010" when "0110110101000100", -- t[27972] = 10
      "001010" when "0110110101000101", -- t[27973] = 10
      "001010" when "0110110101000110", -- t[27974] = 10
      "001010" when "0110110101000111", -- t[27975] = 10
      "001010" when "0110110101001000", -- t[27976] = 10
      "001010" when "0110110101001001", -- t[27977] = 10
      "001010" when "0110110101001010", -- t[27978] = 10
      "001010" when "0110110101001011", -- t[27979] = 10
      "001010" when "0110110101001100", -- t[27980] = 10
      "001010" when "0110110101001101", -- t[27981] = 10
      "001010" when "0110110101001110", -- t[27982] = 10
      "001010" when "0110110101001111", -- t[27983] = 10
      "001010" when "0110110101010000", -- t[27984] = 10
      "001010" when "0110110101010001", -- t[27985] = 10
      "001010" when "0110110101010010", -- t[27986] = 10
      "001010" when "0110110101010011", -- t[27987] = 10
      "001010" when "0110110101010100", -- t[27988] = 10
      "001010" when "0110110101010101", -- t[27989] = 10
      "001010" when "0110110101010110", -- t[27990] = 10
      "001010" when "0110110101010111", -- t[27991] = 10
      "001010" when "0110110101011000", -- t[27992] = 10
      "001010" when "0110110101011001", -- t[27993] = 10
      "001010" when "0110110101011010", -- t[27994] = 10
      "001010" when "0110110101011011", -- t[27995] = 10
      "001010" when "0110110101011100", -- t[27996] = 10
      "001010" when "0110110101011101", -- t[27997] = 10
      "001010" when "0110110101011110", -- t[27998] = 10
      "001010" when "0110110101011111", -- t[27999] = 10
      "001010" when "0110110101100000", -- t[28000] = 10
      "001010" when "0110110101100001", -- t[28001] = 10
      "001010" when "0110110101100010", -- t[28002] = 10
      "001010" when "0110110101100011", -- t[28003] = 10
      "001010" when "0110110101100100", -- t[28004] = 10
      "001010" when "0110110101100101", -- t[28005] = 10
      "001010" when "0110110101100110", -- t[28006] = 10
      "001010" when "0110110101100111", -- t[28007] = 10
      "001010" when "0110110101101000", -- t[28008] = 10
      "001010" when "0110110101101001", -- t[28009] = 10
      "001010" when "0110110101101010", -- t[28010] = 10
      "001010" when "0110110101101011", -- t[28011] = 10
      "001010" when "0110110101101100", -- t[28012] = 10
      "001010" when "0110110101101101", -- t[28013] = 10
      "001010" when "0110110101101110", -- t[28014] = 10
      "001010" when "0110110101101111", -- t[28015] = 10
      "001010" when "0110110101110000", -- t[28016] = 10
      "001010" when "0110110101110001", -- t[28017] = 10
      "001010" when "0110110101110010", -- t[28018] = 10
      "001010" when "0110110101110011", -- t[28019] = 10
      "001010" when "0110110101110100", -- t[28020] = 10
      "001010" when "0110110101110101", -- t[28021] = 10
      "001010" when "0110110101110110", -- t[28022] = 10
      "001010" when "0110110101110111", -- t[28023] = 10
      "001010" when "0110110101111000", -- t[28024] = 10
      "001010" when "0110110101111001", -- t[28025] = 10
      "001010" when "0110110101111010", -- t[28026] = 10
      "001010" when "0110110101111011", -- t[28027] = 10
      "001010" when "0110110101111100", -- t[28028] = 10
      "001010" when "0110110101111101", -- t[28029] = 10
      "001010" when "0110110101111110", -- t[28030] = 10
      "001010" when "0110110101111111", -- t[28031] = 10
      "001010" when "0110110110000000", -- t[28032] = 10
      "001010" when "0110110110000001", -- t[28033] = 10
      "001010" when "0110110110000010", -- t[28034] = 10
      "001010" when "0110110110000011", -- t[28035] = 10
      "001010" when "0110110110000100", -- t[28036] = 10
      "001010" when "0110110110000101", -- t[28037] = 10
      "001010" when "0110110110000110", -- t[28038] = 10
      "001010" when "0110110110000111", -- t[28039] = 10
      "001010" when "0110110110001000", -- t[28040] = 10
      "001010" when "0110110110001001", -- t[28041] = 10
      "001010" when "0110110110001010", -- t[28042] = 10
      "001010" when "0110110110001011", -- t[28043] = 10
      "001010" when "0110110110001100", -- t[28044] = 10
      "001010" when "0110110110001101", -- t[28045] = 10
      "001010" when "0110110110001110", -- t[28046] = 10
      "001010" when "0110110110001111", -- t[28047] = 10
      "001010" when "0110110110010000", -- t[28048] = 10
      "001010" when "0110110110010001", -- t[28049] = 10
      "001010" when "0110110110010010", -- t[28050] = 10
      "001010" when "0110110110010011", -- t[28051] = 10
      "001010" when "0110110110010100", -- t[28052] = 10
      "001010" when "0110110110010101", -- t[28053] = 10
      "001010" when "0110110110010110", -- t[28054] = 10
      "001010" when "0110110110010111", -- t[28055] = 10
      "001010" when "0110110110011000", -- t[28056] = 10
      "001010" when "0110110110011001", -- t[28057] = 10
      "001010" when "0110110110011010", -- t[28058] = 10
      "001010" when "0110110110011011", -- t[28059] = 10
      "001010" when "0110110110011100", -- t[28060] = 10
      "001010" when "0110110110011101", -- t[28061] = 10
      "001010" when "0110110110011110", -- t[28062] = 10
      "001010" when "0110110110011111", -- t[28063] = 10
      "001010" when "0110110110100000", -- t[28064] = 10
      "001010" when "0110110110100001", -- t[28065] = 10
      "001010" when "0110110110100010", -- t[28066] = 10
      "001010" when "0110110110100011", -- t[28067] = 10
      "001010" when "0110110110100100", -- t[28068] = 10
      "001010" when "0110110110100101", -- t[28069] = 10
      "001010" when "0110110110100110", -- t[28070] = 10
      "001010" when "0110110110100111", -- t[28071] = 10
      "001010" when "0110110110101000", -- t[28072] = 10
      "001010" when "0110110110101001", -- t[28073] = 10
      "001010" when "0110110110101010", -- t[28074] = 10
      "001010" when "0110110110101011", -- t[28075] = 10
      "001010" when "0110110110101100", -- t[28076] = 10
      "001010" when "0110110110101101", -- t[28077] = 10
      "001010" when "0110110110101110", -- t[28078] = 10
      "001010" when "0110110110101111", -- t[28079] = 10
      "001010" when "0110110110110000", -- t[28080] = 10
      "001010" when "0110110110110001", -- t[28081] = 10
      "001010" when "0110110110110010", -- t[28082] = 10
      "001010" when "0110110110110011", -- t[28083] = 10
      "001010" when "0110110110110100", -- t[28084] = 10
      "001010" when "0110110110110101", -- t[28085] = 10
      "001010" when "0110110110110110", -- t[28086] = 10
      "001010" when "0110110110110111", -- t[28087] = 10
      "001010" when "0110110110111000", -- t[28088] = 10
      "001010" when "0110110110111001", -- t[28089] = 10
      "001010" when "0110110110111010", -- t[28090] = 10
      "001010" when "0110110110111011", -- t[28091] = 10
      "001010" when "0110110110111100", -- t[28092] = 10
      "001010" when "0110110110111101", -- t[28093] = 10
      "001010" when "0110110110111110", -- t[28094] = 10
      "001010" when "0110110110111111", -- t[28095] = 10
      "001010" when "0110110111000000", -- t[28096] = 10
      "001010" when "0110110111000001", -- t[28097] = 10
      "001010" when "0110110111000010", -- t[28098] = 10
      "001010" when "0110110111000011", -- t[28099] = 10
      "001010" when "0110110111000100", -- t[28100] = 10
      "001010" when "0110110111000101", -- t[28101] = 10
      "001010" when "0110110111000110", -- t[28102] = 10
      "001010" when "0110110111000111", -- t[28103] = 10
      "001010" when "0110110111001000", -- t[28104] = 10
      "001010" when "0110110111001001", -- t[28105] = 10
      "001010" when "0110110111001010", -- t[28106] = 10
      "001010" when "0110110111001011", -- t[28107] = 10
      "001011" when "0110110111001100", -- t[28108] = 11
      "001011" when "0110110111001101", -- t[28109] = 11
      "001011" when "0110110111001110", -- t[28110] = 11
      "001011" when "0110110111001111", -- t[28111] = 11
      "001011" when "0110110111010000", -- t[28112] = 11
      "001011" when "0110110111010001", -- t[28113] = 11
      "001011" when "0110110111010010", -- t[28114] = 11
      "001011" when "0110110111010011", -- t[28115] = 11
      "001011" when "0110110111010100", -- t[28116] = 11
      "001011" when "0110110111010101", -- t[28117] = 11
      "001011" when "0110110111010110", -- t[28118] = 11
      "001011" when "0110110111010111", -- t[28119] = 11
      "001011" when "0110110111011000", -- t[28120] = 11
      "001011" when "0110110111011001", -- t[28121] = 11
      "001011" when "0110110111011010", -- t[28122] = 11
      "001011" when "0110110111011011", -- t[28123] = 11
      "001011" when "0110110111011100", -- t[28124] = 11
      "001011" when "0110110111011101", -- t[28125] = 11
      "001011" when "0110110111011110", -- t[28126] = 11
      "001011" when "0110110111011111", -- t[28127] = 11
      "001011" when "0110110111100000", -- t[28128] = 11
      "001011" when "0110110111100001", -- t[28129] = 11
      "001011" when "0110110111100010", -- t[28130] = 11
      "001011" when "0110110111100011", -- t[28131] = 11
      "001011" when "0110110111100100", -- t[28132] = 11
      "001011" when "0110110111100101", -- t[28133] = 11
      "001011" when "0110110111100110", -- t[28134] = 11
      "001011" when "0110110111100111", -- t[28135] = 11
      "001011" when "0110110111101000", -- t[28136] = 11
      "001011" when "0110110111101001", -- t[28137] = 11
      "001011" when "0110110111101010", -- t[28138] = 11
      "001011" when "0110110111101011", -- t[28139] = 11
      "001011" when "0110110111101100", -- t[28140] = 11
      "001011" when "0110110111101101", -- t[28141] = 11
      "001011" when "0110110111101110", -- t[28142] = 11
      "001011" when "0110110111101111", -- t[28143] = 11
      "001011" when "0110110111110000", -- t[28144] = 11
      "001011" when "0110110111110001", -- t[28145] = 11
      "001011" when "0110110111110010", -- t[28146] = 11
      "001011" when "0110110111110011", -- t[28147] = 11
      "001011" when "0110110111110100", -- t[28148] = 11
      "001011" when "0110110111110101", -- t[28149] = 11
      "001011" when "0110110111110110", -- t[28150] = 11
      "001011" when "0110110111110111", -- t[28151] = 11
      "001011" when "0110110111111000", -- t[28152] = 11
      "001011" when "0110110111111001", -- t[28153] = 11
      "001011" when "0110110111111010", -- t[28154] = 11
      "001011" when "0110110111111011", -- t[28155] = 11
      "001011" when "0110110111111100", -- t[28156] = 11
      "001011" when "0110110111111101", -- t[28157] = 11
      "001011" when "0110110111111110", -- t[28158] = 11
      "001011" when "0110110111111111", -- t[28159] = 11
      "001011" when "0110111000000000", -- t[28160] = 11
      "001011" when "0110111000000001", -- t[28161] = 11
      "001011" when "0110111000000010", -- t[28162] = 11
      "001011" when "0110111000000011", -- t[28163] = 11
      "001011" when "0110111000000100", -- t[28164] = 11
      "001011" when "0110111000000101", -- t[28165] = 11
      "001011" when "0110111000000110", -- t[28166] = 11
      "001011" when "0110111000000111", -- t[28167] = 11
      "001011" when "0110111000001000", -- t[28168] = 11
      "001011" when "0110111000001001", -- t[28169] = 11
      "001011" when "0110111000001010", -- t[28170] = 11
      "001011" when "0110111000001011", -- t[28171] = 11
      "001011" when "0110111000001100", -- t[28172] = 11
      "001011" when "0110111000001101", -- t[28173] = 11
      "001011" when "0110111000001110", -- t[28174] = 11
      "001011" when "0110111000001111", -- t[28175] = 11
      "001011" when "0110111000010000", -- t[28176] = 11
      "001011" when "0110111000010001", -- t[28177] = 11
      "001011" when "0110111000010010", -- t[28178] = 11
      "001011" when "0110111000010011", -- t[28179] = 11
      "001011" when "0110111000010100", -- t[28180] = 11
      "001011" when "0110111000010101", -- t[28181] = 11
      "001011" when "0110111000010110", -- t[28182] = 11
      "001011" when "0110111000010111", -- t[28183] = 11
      "001011" when "0110111000011000", -- t[28184] = 11
      "001011" when "0110111000011001", -- t[28185] = 11
      "001011" when "0110111000011010", -- t[28186] = 11
      "001011" when "0110111000011011", -- t[28187] = 11
      "001011" when "0110111000011100", -- t[28188] = 11
      "001011" when "0110111000011101", -- t[28189] = 11
      "001011" when "0110111000011110", -- t[28190] = 11
      "001011" when "0110111000011111", -- t[28191] = 11
      "001011" when "0110111000100000", -- t[28192] = 11
      "001011" when "0110111000100001", -- t[28193] = 11
      "001011" when "0110111000100010", -- t[28194] = 11
      "001011" when "0110111000100011", -- t[28195] = 11
      "001011" when "0110111000100100", -- t[28196] = 11
      "001011" when "0110111000100101", -- t[28197] = 11
      "001011" when "0110111000100110", -- t[28198] = 11
      "001011" when "0110111000100111", -- t[28199] = 11
      "001011" when "0110111000101000", -- t[28200] = 11
      "001011" when "0110111000101001", -- t[28201] = 11
      "001011" when "0110111000101010", -- t[28202] = 11
      "001011" when "0110111000101011", -- t[28203] = 11
      "001011" when "0110111000101100", -- t[28204] = 11
      "001011" when "0110111000101101", -- t[28205] = 11
      "001011" when "0110111000101110", -- t[28206] = 11
      "001011" when "0110111000101111", -- t[28207] = 11
      "001011" when "0110111000110000", -- t[28208] = 11
      "001011" when "0110111000110001", -- t[28209] = 11
      "001011" when "0110111000110010", -- t[28210] = 11
      "001011" when "0110111000110011", -- t[28211] = 11
      "001011" when "0110111000110100", -- t[28212] = 11
      "001011" when "0110111000110101", -- t[28213] = 11
      "001011" when "0110111000110110", -- t[28214] = 11
      "001011" when "0110111000110111", -- t[28215] = 11
      "001011" when "0110111000111000", -- t[28216] = 11
      "001011" when "0110111000111001", -- t[28217] = 11
      "001011" when "0110111000111010", -- t[28218] = 11
      "001011" when "0110111000111011", -- t[28219] = 11
      "001011" when "0110111000111100", -- t[28220] = 11
      "001011" when "0110111000111101", -- t[28221] = 11
      "001011" when "0110111000111110", -- t[28222] = 11
      "001011" when "0110111000111111", -- t[28223] = 11
      "001011" when "0110111001000000", -- t[28224] = 11
      "001011" when "0110111001000001", -- t[28225] = 11
      "001011" when "0110111001000010", -- t[28226] = 11
      "001011" when "0110111001000011", -- t[28227] = 11
      "001011" when "0110111001000100", -- t[28228] = 11
      "001011" when "0110111001000101", -- t[28229] = 11
      "001011" when "0110111001000110", -- t[28230] = 11
      "001011" when "0110111001000111", -- t[28231] = 11
      "001011" when "0110111001001000", -- t[28232] = 11
      "001011" when "0110111001001001", -- t[28233] = 11
      "001011" when "0110111001001010", -- t[28234] = 11
      "001011" when "0110111001001011", -- t[28235] = 11
      "001011" when "0110111001001100", -- t[28236] = 11
      "001011" when "0110111001001101", -- t[28237] = 11
      "001011" when "0110111001001110", -- t[28238] = 11
      "001011" when "0110111001001111", -- t[28239] = 11
      "001011" when "0110111001010000", -- t[28240] = 11
      "001011" when "0110111001010001", -- t[28241] = 11
      "001011" when "0110111001010010", -- t[28242] = 11
      "001011" when "0110111001010011", -- t[28243] = 11
      "001011" when "0110111001010100", -- t[28244] = 11
      "001011" when "0110111001010101", -- t[28245] = 11
      "001011" when "0110111001010110", -- t[28246] = 11
      "001011" when "0110111001010111", -- t[28247] = 11
      "001011" when "0110111001011000", -- t[28248] = 11
      "001011" when "0110111001011001", -- t[28249] = 11
      "001011" when "0110111001011010", -- t[28250] = 11
      "001011" when "0110111001011011", -- t[28251] = 11
      "001011" when "0110111001011100", -- t[28252] = 11
      "001011" when "0110111001011101", -- t[28253] = 11
      "001011" when "0110111001011110", -- t[28254] = 11
      "001011" when "0110111001011111", -- t[28255] = 11
      "001011" when "0110111001100000", -- t[28256] = 11
      "001011" when "0110111001100001", -- t[28257] = 11
      "001011" when "0110111001100010", -- t[28258] = 11
      "001011" when "0110111001100011", -- t[28259] = 11
      "001011" when "0110111001100100", -- t[28260] = 11
      "001011" when "0110111001100101", -- t[28261] = 11
      "001011" when "0110111001100110", -- t[28262] = 11
      "001011" when "0110111001100111", -- t[28263] = 11
      "001011" when "0110111001101000", -- t[28264] = 11
      "001011" when "0110111001101001", -- t[28265] = 11
      "001011" when "0110111001101010", -- t[28266] = 11
      "001011" when "0110111001101011", -- t[28267] = 11
      "001011" when "0110111001101100", -- t[28268] = 11
      "001011" when "0110111001101101", -- t[28269] = 11
      "001011" when "0110111001101110", -- t[28270] = 11
      "001011" when "0110111001101111", -- t[28271] = 11
      "001011" when "0110111001110000", -- t[28272] = 11
      "001011" when "0110111001110001", -- t[28273] = 11
      "001011" when "0110111001110010", -- t[28274] = 11
      "001011" when "0110111001110011", -- t[28275] = 11
      "001011" when "0110111001110100", -- t[28276] = 11
      "001011" when "0110111001110101", -- t[28277] = 11
      "001011" when "0110111001110110", -- t[28278] = 11
      "001011" when "0110111001110111", -- t[28279] = 11
      "001011" when "0110111001111000", -- t[28280] = 11
      "001011" when "0110111001111001", -- t[28281] = 11
      "001011" when "0110111001111010", -- t[28282] = 11
      "001011" when "0110111001111011", -- t[28283] = 11
      "001011" when "0110111001111100", -- t[28284] = 11
      "001011" when "0110111001111101", -- t[28285] = 11
      "001011" when "0110111001111110", -- t[28286] = 11
      "001011" when "0110111001111111", -- t[28287] = 11
      "001011" when "0110111010000000", -- t[28288] = 11
      "001011" when "0110111010000001", -- t[28289] = 11
      "001011" when "0110111010000010", -- t[28290] = 11
      "001011" when "0110111010000011", -- t[28291] = 11
      "001011" when "0110111010000100", -- t[28292] = 11
      "001011" when "0110111010000101", -- t[28293] = 11
      "001011" when "0110111010000110", -- t[28294] = 11
      "001011" when "0110111010000111", -- t[28295] = 11
      "001011" when "0110111010001000", -- t[28296] = 11
      "001011" when "0110111010001001", -- t[28297] = 11
      "001011" when "0110111010001010", -- t[28298] = 11
      "001011" when "0110111010001011", -- t[28299] = 11
      "001011" when "0110111010001100", -- t[28300] = 11
      "001011" when "0110111010001101", -- t[28301] = 11
      "001011" when "0110111010001110", -- t[28302] = 11
      "001011" when "0110111010001111", -- t[28303] = 11
      "001011" when "0110111010010000", -- t[28304] = 11
      "001011" when "0110111010010001", -- t[28305] = 11
      "001011" when "0110111010010010", -- t[28306] = 11
      "001011" when "0110111010010011", -- t[28307] = 11
      "001011" when "0110111010010100", -- t[28308] = 11
      "001011" when "0110111010010101", -- t[28309] = 11
      "001011" when "0110111010010110", -- t[28310] = 11
      "001011" when "0110111010010111", -- t[28311] = 11
      "001011" when "0110111010011000", -- t[28312] = 11
      "001011" when "0110111010011001", -- t[28313] = 11
      "001011" when "0110111010011010", -- t[28314] = 11
      "001011" when "0110111010011011", -- t[28315] = 11
      "001011" when "0110111010011100", -- t[28316] = 11
      "001011" when "0110111010011101", -- t[28317] = 11
      "001011" when "0110111010011110", -- t[28318] = 11
      "001011" when "0110111010011111", -- t[28319] = 11
      "001011" when "0110111010100000", -- t[28320] = 11
      "001011" when "0110111010100001", -- t[28321] = 11
      "001011" when "0110111010100010", -- t[28322] = 11
      "001011" when "0110111010100011", -- t[28323] = 11
      "001011" when "0110111010100100", -- t[28324] = 11
      "001011" when "0110111010100101", -- t[28325] = 11
      "001011" when "0110111010100110", -- t[28326] = 11
      "001011" when "0110111010100111", -- t[28327] = 11
      "001011" when "0110111010101000", -- t[28328] = 11
      "001011" when "0110111010101001", -- t[28329] = 11
      "001011" when "0110111010101010", -- t[28330] = 11
      "001011" when "0110111010101011", -- t[28331] = 11
      "001011" when "0110111010101100", -- t[28332] = 11
      "001011" when "0110111010101101", -- t[28333] = 11
      "001011" when "0110111010101110", -- t[28334] = 11
      "001011" when "0110111010101111", -- t[28335] = 11
      "001011" when "0110111010110000", -- t[28336] = 11
      "001011" when "0110111010110001", -- t[28337] = 11
      "001011" when "0110111010110010", -- t[28338] = 11
      "001011" when "0110111010110011", -- t[28339] = 11
      "001011" when "0110111010110100", -- t[28340] = 11
      "001011" when "0110111010110101", -- t[28341] = 11
      "001011" when "0110111010110110", -- t[28342] = 11
      "001011" when "0110111010110111", -- t[28343] = 11
      "001011" when "0110111010111000", -- t[28344] = 11
      "001011" when "0110111010111001", -- t[28345] = 11
      "001011" when "0110111010111010", -- t[28346] = 11
      "001011" when "0110111010111011", -- t[28347] = 11
      "001011" when "0110111010111100", -- t[28348] = 11
      "001011" when "0110111010111101", -- t[28349] = 11
      "001011" when "0110111010111110", -- t[28350] = 11
      "001011" when "0110111010111111", -- t[28351] = 11
      "001011" when "0110111011000000", -- t[28352] = 11
      "001011" when "0110111011000001", -- t[28353] = 11
      "001011" when "0110111011000010", -- t[28354] = 11
      "001011" when "0110111011000011", -- t[28355] = 11
      "001011" when "0110111011000100", -- t[28356] = 11
      "001011" when "0110111011000101", -- t[28357] = 11
      "001011" when "0110111011000110", -- t[28358] = 11
      "001011" when "0110111011000111", -- t[28359] = 11
      "001011" when "0110111011001000", -- t[28360] = 11
      "001011" when "0110111011001001", -- t[28361] = 11
      "001011" when "0110111011001010", -- t[28362] = 11
      "001011" when "0110111011001011", -- t[28363] = 11
      "001011" when "0110111011001100", -- t[28364] = 11
      "001011" when "0110111011001101", -- t[28365] = 11
      "001011" when "0110111011001110", -- t[28366] = 11
      "001011" when "0110111011001111", -- t[28367] = 11
      "001011" when "0110111011010000", -- t[28368] = 11
      "001011" when "0110111011010001", -- t[28369] = 11
      "001011" when "0110111011010010", -- t[28370] = 11
      "001011" when "0110111011010011", -- t[28371] = 11
      "001011" when "0110111011010100", -- t[28372] = 11
      "001011" when "0110111011010101", -- t[28373] = 11
      "001011" when "0110111011010110", -- t[28374] = 11
      "001011" when "0110111011010111", -- t[28375] = 11
      "001011" when "0110111011011000", -- t[28376] = 11
      "001011" when "0110111011011001", -- t[28377] = 11
      "001011" when "0110111011011010", -- t[28378] = 11
      "001011" when "0110111011011011", -- t[28379] = 11
      "001011" when "0110111011011100", -- t[28380] = 11
      "001011" when "0110111011011101", -- t[28381] = 11
      "001011" when "0110111011011110", -- t[28382] = 11
      "001011" when "0110111011011111", -- t[28383] = 11
      "001011" when "0110111011100000", -- t[28384] = 11
      "001011" when "0110111011100001", -- t[28385] = 11
      "001011" when "0110111011100010", -- t[28386] = 11
      "001011" when "0110111011100011", -- t[28387] = 11
      "001011" when "0110111011100100", -- t[28388] = 11
      "001011" when "0110111011100101", -- t[28389] = 11
      "001011" when "0110111011100110", -- t[28390] = 11
      "001011" when "0110111011100111", -- t[28391] = 11
      "001011" when "0110111011101000", -- t[28392] = 11
      "001011" when "0110111011101001", -- t[28393] = 11
      "001011" when "0110111011101010", -- t[28394] = 11
      "001011" when "0110111011101011", -- t[28395] = 11
      "001011" when "0110111011101100", -- t[28396] = 11
      "001011" when "0110111011101101", -- t[28397] = 11
      "001011" when "0110111011101110", -- t[28398] = 11
      "001011" when "0110111011101111", -- t[28399] = 11
      "001011" when "0110111011110000", -- t[28400] = 11
      "001011" when "0110111011110001", -- t[28401] = 11
      "001011" when "0110111011110010", -- t[28402] = 11
      "001011" when "0110111011110011", -- t[28403] = 11
      "001011" when "0110111011110100", -- t[28404] = 11
      "001011" when "0110111011110101", -- t[28405] = 11
      "001011" when "0110111011110110", -- t[28406] = 11
      "001011" when "0110111011110111", -- t[28407] = 11
      "001011" when "0110111011111000", -- t[28408] = 11
      "001011" when "0110111011111001", -- t[28409] = 11
      "001011" when "0110111011111010", -- t[28410] = 11
      "001011" when "0110111011111011", -- t[28411] = 11
      "001011" when "0110111011111100", -- t[28412] = 11
      "001011" when "0110111011111101", -- t[28413] = 11
      "001011" when "0110111011111110", -- t[28414] = 11
      "001011" when "0110111011111111", -- t[28415] = 11
      "001011" when "0110111100000000", -- t[28416] = 11
      "001011" when "0110111100000001", -- t[28417] = 11
      "001011" when "0110111100000010", -- t[28418] = 11
      "001011" when "0110111100000011", -- t[28419] = 11
      "001011" when "0110111100000100", -- t[28420] = 11
      "001011" when "0110111100000101", -- t[28421] = 11
      "001011" when "0110111100000110", -- t[28422] = 11
      "001011" when "0110111100000111", -- t[28423] = 11
      "001011" when "0110111100001000", -- t[28424] = 11
      "001011" when "0110111100001001", -- t[28425] = 11
      "001011" when "0110111100001010", -- t[28426] = 11
      "001011" when "0110111100001011", -- t[28427] = 11
      "001011" when "0110111100001100", -- t[28428] = 11
      "001011" when "0110111100001101", -- t[28429] = 11
      "001011" when "0110111100001110", -- t[28430] = 11
      "001011" when "0110111100001111", -- t[28431] = 11
      "001011" when "0110111100010000", -- t[28432] = 11
      "001011" when "0110111100010001", -- t[28433] = 11
      "001011" when "0110111100010010", -- t[28434] = 11
      "001011" when "0110111100010011", -- t[28435] = 11
      "001011" when "0110111100010100", -- t[28436] = 11
      "001011" when "0110111100010101", -- t[28437] = 11
      "001011" when "0110111100010110", -- t[28438] = 11
      "001011" when "0110111100010111", -- t[28439] = 11
      "001011" when "0110111100011000", -- t[28440] = 11
      "001011" when "0110111100011001", -- t[28441] = 11
      "001011" when "0110111100011010", -- t[28442] = 11
      "001011" when "0110111100011011", -- t[28443] = 11
      "001011" when "0110111100011100", -- t[28444] = 11
      "001011" when "0110111100011101", -- t[28445] = 11
      "001011" when "0110111100011110", -- t[28446] = 11
      "001011" when "0110111100011111", -- t[28447] = 11
      "001011" when "0110111100100000", -- t[28448] = 11
      "001011" when "0110111100100001", -- t[28449] = 11
      "001011" when "0110111100100010", -- t[28450] = 11
      "001011" when "0110111100100011", -- t[28451] = 11
      "001011" when "0110111100100100", -- t[28452] = 11
      "001011" when "0110111100100101", -- t[28453] = 11
      "001011" when "0110111100100110", -- t[28454] = 11
      "001011" when "0110111100100111", -- t[28455] = 11
      "001011" when "0110111100101000", -- t[28456] = 11
      "001011" when "0110111100101001", -- t[28457] = 11
      "001011" when "0110111100101010", -- t[28458] = 11
      "001011" when "0110111100101011", -- t[28459] = 11
      "001011" when "0110111100101100", -- t[28460] = 11
      "001011" when "0110111100101101", -- t[28461] = 11
      "001011" when "0110111100101110", -- t[28462] = 11
      "001011" when "0110111100101111", -- t[28463] = 11
      "001011" when "0110111100110000", -- t[28464] = 11
      "001011" when "0110111100110001", -- t[28465] = 11
      "001011" when "0110111100110010", -- t[28466] = 11
      "001011" when "0110111100110011", -- t[28467] = 11
      "001011" when "0110111100110100", -- t[28468] = 11
      "001011" when "0110111100110101", -- t[28469] = 11
      "001011" when "0110111100110110", -- t[28470] = 11
      "001011" when "0110111100110111", -- t[28471] = 11
      "001011" when "0110111100111000", -- t[28472] = 11
      "001011" when "0110111100111001", -- t[28473] = 11
      "001011" when "0110111100111010", -- t[28474] = 11
      "001011" when "0110111100111011", -- t[28475] = 11
      "001011" when "0110111100111100", -- t[28476] = 11
      "001011" when "0110111100111101", -- t[28477] = 11
      "001011" when "0110111100111110", -- t[28478] = 11
      "001011" when "0110111100111111", -- t[28479] = 11
      "001011" when "0110111101000000", -- t[28480] = 11
      "001011" when "0110111101000001", -- t[28481] = 11
      "001011" when "0110111101000010", -- t[28482] = 11
      "001011" when "0110111101000011", -- t[28483] = 11
      "001011" when "0110111101000100", -- t[28484] = 11
      "001011" when "0110111101000101", -- t[28485] = 11
      "001011" when "0110111101000110", -- t[28486] = 11
      "001011" when "0110111101000111", -- t[28487] = 11
      "001011" when "0110111101001000", -- t[28488] = 11
      "001011" when "0110111101001001", -- t[28489] = 11
      "001011" when "0110111101001010", -- t[28490] = 11
      "001011" when "0110111101001011", -- t[28491] = 11
      "001011" when "0110111101001100", -- t[28492] = 11
      "001011" when "0110111101001101", -- t[28493] = 11
      "001011" when "0110111101001110", -- t[28494] = 11
      "001011" when "0110111101001111", -- t[28495] = 11
      "001011" when "0110111101010000", -- t[28496] = 11
      "001011" when "0110111101010001", -- t[28497] = 11
      "001011" when "0110111101010010", -- t[28498] = 11
      "001011" when "0110111101010011", -- t[28499] = 11
      "001011" when "0110111101010100", -- t[28500] = 11
      "001011" when "0110111101010101", -- t[28501] = 11
      "001011" when "0110111101010110", -- t[28502] = 11
      "001011" when "0110111101010111", -- t[28503] = 11
      "001011" when "0110111101011000", -- t[28504] = 11
      "001011" when "0110111101011001", -- t[28505] = 11
      "001011" when "0110111101011010", -- t[28506] = 11
      "001011" when "0110111101011011", -- t[28507] = 11
      "001011" when "0110111101011100", -- t[28508] = 11
      "001011" when "0110111101011101", -- t[28509] = 11
      "001011" when "0110111101011110", -- t[28510] = 11
      "001011" when "0110111101011111", -- t[28511] = 11
      "001011" when "0110111101100000", -- t[28512] = 11
      "001011" when "0110111101100001", -- t[28513] = 11
      "001011" when "0110111101100010", -- t[28514] = 11
      "001011" when "0110111101100011", -- t[28515] = 11
      "001011" when "0110111101100100", -- t[28516] = 11
      "001011" when "0110111101100101", -- t[28517] = 11
      "001011" when "0110111101100110", -- t[28518] = 11
      "001011" when "0110111101100111", -- t[28519] = 11
      "001011" when "0110111101101000", -- t[28520] = 11
      "001011" when "0110111101101001", -- t[28521] = 11
      "001011" when "0110111101101010", -- t[28522] = 11
      "001011" when "0110111101101011", -- t[28523] = 11
      "001011" when "0110111101101100", -- t[28524] = 11
      "001011" when "0110111101101101", -- t[28525] = 11
      "001011" when "0110111101101110", -- t[28526] = 11
      "001011" when "0110111101101111", -- t[28527] = 11
      "001011" when "0110111101110000", -- t[28528] = 11
      "001011" when "0110111101110001", -- t[28529] = 11
      "001011" when "0110111101110010", -- t[28530] = 11
      "001011" when "0110111101110011", -- t[28531] = 11
      "001011" when "0110111101110100", -- t[28532] = 11
      "001011" when "0110111101110101", -- t[28533] = 11
      "001011" when "0110111101110110", -- t[28534] = 11
      "001011" when "0110111101110111", -- t[28535] = 11
      "001011" when "0110111101111000", -- t[28536] = 11
      "001011" when "0110111101111001", -- t[28537] = 11
      "001011" when "0110111101111010", -- t[28538] = 11
      "001011" when "0110111101111011", -- t[28539] = 11
      "001011" when "0110111101111100", -- t[28540] = 11
      "001011" when "0110111101111101", -- t[28541] = 11
      "001011" when "0110111101111110", -- t[28542] = 11
      "001011" when "0110111101111111", -- t[28543] = 11
      "001011" when "0110111110000000", -- t[28544] = 11
      "001011" when "0110111110000001", -- t[28545] = 11
      "001011" when "0110111110000010", -- t[28546] = 11
      "001011" when "0110111110000011", -- t[28547] = 11
      "001011" when "0110111110000100", -- t[28548] = 11
      "001011" when "0110111110000101", -- t[28549] = 11
      "001011" when "0110111110000110", -- t[28550] = 11
      "001011" when "0110111110000111", -- t[28551] = 11
      "001011" when "0110111110001000", -- t[28552] = 11
      "001011" when "0110111110001001", -- t[28553] = 11
      "001011" when "0110111110001010", -- t[28554] = 11
      "001011" when "0110111110001011", -- t[28555] = 11
      "001011" when "0110111110001100", -- t[28556] = 11
      "001011" when "0110111110001101", -- t[28557] = 11
      "001011" when "0110111110001110", -- t[28558] = 11
      "001011" when "0110111110001111", -- t[28559] = 11
      "001011" when "0110111110010000", -- t[28560] = 11
      "001011" when "0110111110010001", -- t[28561] = 11
      "001011" when "0110111110010010", -- t[28562] = 11
      "001011" when "0110111110010011", -- t[28563] = 11
      "001011" when "0110111110010100", -- t[28564] = 11
      "001011" when "0110111110010101", -- t[28565] = 11
      "001011" when "0110111110010110", -- t[28566] = 11
      "001011" when "0110111110010111", -- t[28567] = 11
      "001011" when "0110111110011000", -- t[28568] = 11
      "001011" when "0110111110011001", -- t[28569] = 11
      "001011" when "0110111110011010", -- t[28570] = 11
      "001011" when "0110111110011011", -- t[28571] = 11
      "001011" when "0110111110011100", -- t[28572] = 11
      "001011" when "0110111110011101", -- t[28573] = 11
      "001011" when "0110111110011110", -- t[28574] = 11
      "001011" when "0110111110011111", -- t[28575] = 11
      "001011" when "0110111110100000", -- t[28576] = 11
      "001011" when "0110111110100001", -- t[28577] = 11
      "001011" when "0110111110100010", -- t[28578] = 11
      "001011" when "0110111110100011", -- t[28579] = 11
      "001011" when "0110111110100100", -- t[28580] = 11
      "001011" when "0110111110100101", -- t[28581] = 11
      "001011" when "0110111110100110", -- t[28582] = 11
      "001011" when "0110111110100111", -- t[28583] = 11
      "001011" when "0110111110101000", -- t[28584] = 11
      "001011" when "0110111110101001", -- t[28585] = 11
      "001011" when "0110111110101010", -- t[28586] = 11
      "001011" when "0110111110101011", -- t[28587] = 11
      "001011" when "0110111110101100", -- t[28588] = 11
      "001011" when "0110111110101101", -- t[28589] = 11
      "001011" when "0110111110101110", -- t[28590] = 11
      "001011" when "0110111110101111", -- t[28591] = 11
      "001011" when "0110111110110000", -- t[28592] = 11
      "001011" when "0110111110110001", -- t[28593] = 11
      "001011" when "0110111110110010", -- t[28594] = 11
      "001011" when "0110111110110011", -- t[28595] = 11
      "001011" when "0110111110110100", -- t[28596] = 11
      "001011" when "0110111110110101", -- t[28597] = 11
      "001011" when "0110111110110110", -- t[28598] = 11
      "001011" when "0110111110110111", -- t[28599] = 11
      "001011" when "0110111110111000", -- t[28600] = 11
      "001011" when "0110111110111001", -- t[28601] = 11
      "001011" when "0110111110111010", -- t[28602] = 11
      "001011" when "0110111110111011", -- t[28603] = 11
      "001011" when "0110111110111100", -- t[28604] = 11
      "001011" when "0110111110111101", -- t[28605] = 11
      "001011" when "0110111110111110", -- t[28606] = 11
      "001011" when "0110111110111111", -- t[28607] = 11
      "001011" when "0110111111000000", -- t[28608] = 11
      "001011" when "0110111111000001", -- t[28609] = 11
      "001011" when "0110111111000010", -- t[28610] = 11
      "001011" when "0110111111000011", -- t[28611] = 11
      "001011" when "0110111111000100", -- t[28612] = 11
      "001011" when "0110111111000101", -- t[28613] = 11
      "001011" when "0110111111000110", -- t[28614] = 11
      "001011" when "0110111111000111", -- t[28615] = 11
      "001011" when "0110111111001000", -- t[28616] = 11
      "001011" when "0110111111001001", -- t[28617] = 11
      "001011" when "0110111111001010", -- t[28618] = 11
      "001011" when "0110111111001011", -- t[28619] = 11
      "001011" when "0110111111001100", -- t[28620] = 11
      "001011" when "0110111111001101", -- t[28621] = 11
      "001011" when "0110111111001110", -- t[28622] = 11
      "001011" when "0110111111001111", -- t[28623] = 11
      "001011" when "0110111111010000", -- t[28624] = 11
      "001011" when "0110111111010001", -- t[28625] = 11
      "001011" when "0110111111010010", -- t[28626] = 11
      "001011" when "0110111111010011", -- t[28627] = 11
      "001011" when "0110111111010100", -- t[28628] = 11
      "001011" when "0110111111010101", -- t[28629] = 11
      "001011" when "0110111111010110", -- t[28630] = 11
      "001011" when "0110111111010111", -- t[28631] = 11
      "001011" when "0110111111011000", -- t[28632] = 11
      "001011" when "0110111111011001", -- t[28633] = 11
      "001011" when "0110111111011010", -- t[28634] = 11
      "001011" when "0110111111011011", -- t[28635] = 11
      "001011" when "0110111111011100", -- t[28636] = 11
      "001011" when "0110111111011101", -- t[28637] = 11
      "001011" when "0110111111011110", -- t[28638] = 11
      "001011" when "0110111111011111", -- t[28639] = 11
      "001011" when "0110111111100000", -- t[28640] = 11
      "001011" when "0110111111100001", -- t[28641] = 11
      "001011" when "0110111111100010", -- t[28642] = 11
      "001011" when "0110111111100011", -- t[28643] = 11
      "001011" when "0110111111100100", -- t[28644] = 11
      "001100" when "0110111111100101", -- t[28645] = 12
      "001100" when "0110111111100110", -- t[28646] = 12
      "001100" when "0110111111100111", -- t[28647] = 12
      "001100" when "0110111111101000", -- t[28648] = 12
      "001100" when "0110111111101001", -- t[28649] = 12
      "001100" when "0110111111101010", -- t[28650] = 12
      "001100" when "0110111111101011", -- t[28651] = 12
      "001100" when "0110111111101100", -- t[28652] = 12
      "001100" when "0110111111101101", -- t[28653] = 12
      "001100" when "0110111111101110", -- t[28654] = 12
      "001100" when "0110111111101111", -- t[28655] = 12
      "001100" when "0110111111110000", -- t[28656] = 12
      "001100" when "0110111111110001", -- t[28657] = 12
      "001100" when "0110111111110010", -- t[28658] = 12
      "001100" when "0110111111110011", -- t[28659] = 12
      "001100" when "0110111111110100", -- t[28660] = 12
      "001100" when "0110111111110101", -- t[28661] = 12
      "001100" when "0110111111110110", -- t[28662] = 12
      "001100" when "0110111111110111", -- t[28663] = 12
      "001100" when "0110111111111000", -- t[28664] = 12
      "001100" when "0110111111111001", -- t[28665] = 12
      "001100" when "0110111111111010", -- t[28666] = 12
      "001100" when "0110111111111011", -- t[28667] = 12
      "001100" when "0110111111111100", -- t[28668] = 12
      "001100" when "0110111111111101", -- t[28669] = 12
      "001100" when "0110111111111110", -- t[28670] = 12
      "001100" when "0110111111111111", -- t[28671] = 12
      "001100" when "0111000000000000", -- t[28672] = 12
      "001100" when "0111000000000001", -- t[28673] = 12
      "001100" when "0111000000000010", -- t[28674] = 12
      "001100" when "0111000000000011", -- t[28675] = 12
      "001100" when "0111000000000100", -- t[28676] = 12
      "001100" when "0111000000000101", -- t[28677] = 12
      "001100" when "0111000000000110", -- t[28678] = 12
      "001100" when "0111000000000111", -- t[28679] = 12
      "001100" when "0111000000001000", -- t[28680] = 12
      "001100" when "0111000000001001", -- t[28681] = 12
      "001100" when "0111000000001010", -- t[28682] = 12
      "001100" when "0111000000001011", -- t[28683] = 12
      "001100" when "0111000000001100", -- t[28684] = 12
      "001100" when "0111000000001101", -- t[28685] = 12
      "001100" when "0111000000001110", -- t[28686] = 12
      "001100" when "0111000000001111", -- t[28687] = 12
      "001100" when "0111000000010000", -- t[28688] = 12
      "001100" when "0111000000010001", -- t[28689] = 12
      "001100" when "0111000000010010", -- t[28690] = 12
      "001100" when "0111000000010011", -- t[28691] = 12
      "001100" when "0111000000010100", -- t[28692] = 12
      "001100" when "0111000000010101", -- t[28693] = 12
      "001100" when "0111000000010110", -- t[28694] = 12
      "001100" when "0111000000010111", -- t[28695] = 12
      "001100" when "0111000000011000", -- t[28696] = 12
      "001100" when "0111000000011001", -- t[28697] = 12
      "001100" when "0111000000011010", -- t[28698] = 12
      "001100" when "0111000000011011", -- t[28699] = 12
      "001100" when "0111000000011100", -- t[28700] = 12
      "001100" when "0111000000011101", -- t[28701] = 12
      "001100" when "0111000000011110", -- t[28702] = 12
      "001100" when "0111000000011111", -- t[28703] = 12
      "001100" when "0111000000100000", -- t[28704] = 12
      "001100" when "0111000000100001", -- t[28705] = 12
      "001100" when "0111000000100010", -- t[28706] = 12
      "001100" when "0111000000100011", -- t[28707] = 12
      "001100" when "0111000000100100", -- t[28708] = 12
      "001100" when "0111000000100101", -- t[28709] = 12
      "001100" when "0111000000100110", -- t[28710] = 12
      "001100" when "0111000000100111", -- t[28711] = 12
      "001100" when "0111000000101000", -- t[28712] = 12
      "001100" when "0111000000101001", -- t[28713] = 12
      "001100" when "0111000000101010", -- t[28714] = 12
      "001100" when "0111000000101011", -- t[28715] = 12
      "001100" when "0111000000101100", -- t[28716] = 12
      "001100" when "0111000000101101", -- t[28717] = 12
      "001100" when "0111000000101110", -- t[28718] = 12
      "001100" when "0111000000101111", -- t[28719] = 12
      "001100" when "0111000000110000", -- t[28720] = 12
      "001100" when "0111000000110001", -- t[28721] = 12
      "001100" when "0111000000110010", -- t[28722] = 12
      "001100" when "0111000000110011", -- t[28723] = 12
      "001100" when "0111000000110100", -- t[28724] = 12
      "001100" when "0111000000110101", -- t[28725] = 12
      "001100" when "0111000000110110", -- t[28726] = 12
      "001100" when "0111000000110111", -- t[28727] = 12
      "001100" when "0111000000111000", -- t[28728] = 12
      "001100" when "0111000000111001", -- t[28729] = 12
      "001100" when "0111000000111010", -- t[28730] = 12
      "001100" when "0111000000111011", -- t[28731] = 12
      "001100" when "0111000000111100", -- t[28732] = 12
      "001100" when "0111000000111101", -- t[28733] = 12
      "001100" when "0111000000111110", -- t[28734] = 12
      "001100" when "0111000000111111", -- t[28735] = 12
      "001100" when "0111000001000000", -- t[28736] = 12
      "001100" when "0111000001000001", -- t[28737] = 12
      "001100" when "0111000001000010", -- t[28738] = 12
      "001100" when "0111000001000011", -- t[28739] = 12
      "001100" when "0111000001000100", -- t[28740] = 12
      "001100" when "0111000001000101", -- t[28741] = 12
      "001100" when "0111000001000110", -- t[28742] = 12
      "001100" when "0111000001000111", -- t[28743] = 12
      "001100" when "0111000001001000", -- t[28744] = 12
      "001100" when "0111000001001001", -- t[28745] = 12
      "001100" when "0111000001001010", -- t[28746] = 12
      "001100" when "0111000001001011", -- t[28747] = 12
      "001100" when "0111000001001100", -- t[28748] = 12
      "001100" when "0111000001001101", -- t[28749] = 12
      "001100" when "0111000001001110", -- t[28750] = 12
      "001100" when "0111000001001111", -- t[28751] = 12
      "001100" when "0111000001010000", -- t[28752] = 12
      "001100" when "0111000001010001", -- t[28753] = 12
      "001100" when "0111000001010010", -- t[28754] = 12
      "001100" when "0111000001010011", -- t[28755] = 12
      "001100" when "0111000001010100", -- t[28756] = 12
      "001100" when "0111000001010101", -- t[28757] = 12
      "001100" when "0111000001010110", -- t[28758] = 12
      "001100" when "0111000001010111", -- t[28759] = 12
      "001100" when "0111000001011000", -- t[28760] = 12
      "001100" when "0111000001011001", -- t[28761] = 12
      "001100" when "0111000001011010", -- t[28762] = 12
      "001100" when "0111000001011011", -- t[28763] = 12
      "001100" when "0111000001011100", -- t[28764] = 12
      "001100" when "0111000001011101", -- t[28765] = 12
      "001100" when "0111000001011110", -- t[28766] = 12
      "001100" when "0111000001011111", -- t[28767] = 12
      "001100" when "0111000001100000", -- t[28768] = 12
      "001100" when "0111000001100001", -- t[28769] = 12
      "001100" when "0111000001100010", -- t[28770] = 12
      "001100" when "0111000001100011", -- t[28771] = 12
      "001100" when "0111000001100100", -- t[28772] = 12
      "001100" when "0111000001100101", -- t[28773] = 12
      "001100" when "0111000001100110", -- t[28774] = 12
      "001100" when "0111000001100111", -- t[28775] = 12
      "001100" when "0111000001101000", -- t[28776] = 12
      "001100" when "0111000001101001", -- t[28777] = 12
      "001100" when "0111000001101010", -- t[28778] = 12
      "001100" when "0111000001101011", -- t[28779] = 12
      "001100" when "0111000001101100", -- t[28780] = 12
      "001100" when "0111000001101101", -- t[28781] = 12
      "001100" when "0111000001101110", -- t[28782] = 12
      "001100" when "0111000001101111", -- t[28783] = 12
      "001100" when "0111000001110000", -- t[28784] = 12
      "001100" when "0111000001110001", -- t[28785] = 12
      "001100" when "0111000001110010", -- t[28786] = 12
      "001100" when "0111000001110011", -- t[28787] = 12
      "001100" when "0111000001110100", -- t[28788] = 12
      "001100" when "0111000001110101", -- t[28789] = 12
      "001100" when "0111000001110110", -- t[28790] = 12
      "001100" when "0111000001110111", -- t[28791] = 12
      "001100" when "0111000001111000", -- t[28792] = 12
      "001100" when "0111000001111001", -- t[28793] = 12
      "001100" when "0111000001111010", -- t[28794] = 12
      "001100" when "0111000001111011", -- t[28795] = 12
      "001100" when "0111000001111100", -- t[28796] = 12
      "001100" when "0111000001111101", -- t[28797] = 12
      "001100" when "0111000001111110", -- t[28798] = 12
      "001100" when "0111000001111111", -- t[28799] = 12
      "001100" when "0111000010000000", -- t[28800] = 12
      "001100" when "0111000010000001", -- t[28801] = 12
      "001100" when "0111000010000010", -- t[28802] = 12
      "001100" when "0111000010000011", -- t[28803] = 12
      "001100" when "0111000010000100", -- t[28804] = 12
      "001100" when "0111000010000101", -- t[28805] = 12
      "001100" when "0111000010000110", -- t[28806] = 12
      "001100" when "0111000010000111", -- t[28807] = 12
      "001100" when "0111000010001000", -- t[28808] = 12
      "001100" when "0111000010001001", -- t[28809] = 12
      "001100" when "0111000010001010", -- t[28810] = 12
      "001100" when "0111000010001011", -- t[28811] = 12
      "001100" when "0111000010001100", -- t[28812] = 12
      "001100" when "0111000010001101", -- t[28813] = 12
      "001100" when "0111000010001110", -- t[28814] = 12
      "001100" when "0111000010001111", -- t[28815] = 12
      "001100" when "0111000010010000", -- t[28816] = 12
      "001100" when "0111000010010001", -- t[28817] = 12
      "001100" when "0111000010010010", -- t[28818] = 12
      "001100" when "0111000010010011", -- t[28819] = 12
      "001100" when "0111000010010100", -- t[28820] = 12
      "001100" when "0111000010010101", -- t[28821] = 12
      "001100" when "0111000010010110", -- t[28822] = 12
      "001100" when "0111000010010111", -- t[28823] = 12
      "001100" when "0111000010011000", -- t[28824] = 12
      "001100" when "0111000010011001", -- t[28825] = 12
      "001100" when "0111000010011010", -- t[28826] = 12
      "001100" when "0111000010011011", -- t[28827] = 12
      "001100" when "0111000010011100", -- t[28828] = 12
      "001100" when "0111000010011101", -- t[28829] = 12
      "001100" when "0111000010011110", -- t[28830] = 12
      "001100" when "0111000010011111", -- t[28831] = 12
      "001100" when "0111000010100000", -- t[28832] = 12
      "001100" when "0111000010100001", -- t[28833] = 12
      "001100" when "0111000010100010", -- t[28834] = 12
      "001100" when "0111000010100011", -- t[28835] = 12
      "001100" when "0111000010100100", -- t[28836] = 12
      "001100" when "0111000010100101", -- t[28837] = 12
      "001100" when "0111000010100110", -- t[28838] = 12
      "001100" when "0111000010100111", -- t[28839] = 12
      "001100" when "0111000010101000", -- t[28840] = 12
      "001100" when "0111000010101001", -- t[28841] = 12
      "001100" when "0111000010101010", -- t[28842] = 12
      "001100" when "0111000010101011", -- t[28843] = 12
      "001100" when "0111000010101100", -- t[28844] = 12
      "001100" when "0111000010101101", -- t[28845] = 12
      "001100" when "0111000010101110", -- t[28846] = 12
      "001100" when "0111000010101111", -- t[28847] = 12
      "001100" when "0111000010110000", -- t[28848] = 12
      "001100" when "0111000010110001", -- t[28849] = 12
      "001100" when "0111000010110010", -- t[28850] = 12
      "001100" when "0111000010110011", -- t[28851] = 12
      "001100" when "0111000010110100", -- t[28852] = 12
      "001100" when "0111000010110101", -- t[28853] = 12
      "001100" when "0111000010110110", -- t[28854] = 12
      "001100" when "0111000010110111", -- t[28855] = 12
      "001100" when "0111000010111000", -- t[28856] = 12
      "001100" when "0111000010111001", -- t[28857] = 12
      "001100" when "0111000010111010", -- t[28858] = 12
      "001100" when "0111000010111011", -- t[28859] = 12
      "001100" when "0111000010111100", -- t[28860] = 12
      "001100" when "0111000010111101", -- t[28861] = 12
      "001100" when "0111000010111110", -- t[28862] = 12
      "001100" when "0111000010111111", -- t[28863] = 12
      "001100" when "0111000011000000", -- t[28864] = 12
      "001100" when "0111000011000001", -- t[28865] = 12
      "001100" when "0111000011000010", -- t[28866] = 12
      "001100" when "0111000011000011", -- t[28867] = 12
      "001100" when "0111000011000100", -- t[28868] = 12
      "001100" when "0111000011000101", -- t[28869] = 12
      "001100" when "0111000011000110", -- t[28870] = 12
      "001100" when "0111000011000111", -- t[28871] = 12
      "001100" when "0111000011001000", -- t[28872] = 12
      "001100" when "0111000011001001", -- t[28873] = 12
      "001100" when "0111000011001010", -- t[28874] = 12
      "001100" when "0111000011001011", -- t[28875] = 12
      "001100" when "0111000011001100", -- t[28876] = 12
      "001100" when "0111000011001101", -- t[28877] = 12
      "001100" when "0111000011001110", -- t[28878] = 12
      "001100" when "0111000011001111", -- t[28879] = 12
      "001100" when "0111000011010000", -- t[28880] = 12
      "001100" when "0111000011010001", -- t[28881] = 12
      "001100" when "0111000011010010", -- t[28882] = 12
      "001100" when "0111000011010011", -- t[28883] = 12
      "001100" when "0111000011010100", -- t[28884] = 12
      "001100" when "0111000011010101", -- t[28885] = 12
      "001100" when "0111000011010110", -- t[28886] = 12
      "001100" when "0111000011010111", -- t[28887] = 12
      "001100" when "0111000011011000", -- t[28888] = 12
      "001100" when "0111000011011001", -- t[28889] = 12
      "001100" when "0111000011011010", -- t[28890] = 12
      "001100" when "0111000011011011", -- t[28891] = 12
      "001100" when "0111000011011100", -- t[28892] = 12
      "001100" when "0111000011011101", -- t[28893] = 12
      "001100" when "0111000011011110", -- t[28894] = 12
      "001100" when "0111000011011111", -- t[28895] = 12
      "001100" when "0111000011100000", -- t[28896] = 12
      "001100" when "0111000011100001", -- t[28897] = 12
      "001100" when "0111000011100010", -- t[28898] = 12
      "001100" when "0111000011100011", -- t[28899] = 12
      "001100" when "0111000011100100", -- t[28900] = 12
      "001100" when "0111000011100101", -- t[28901] = 12
      "001100" when "0111000011100110", -- t[28902] = 12
      "001100" when "0111000011100111", -- t[28903] = 12
      "001100" when "0111000011101000", -- t[28904] = 12
      "001100" when "0111000011101001", -- t[28905] = 12
      "001100" when "0111000011101010", -- t[28906] = 12
      "001100" when "0111000011101011", -- t[28907] = 12
      "001100" when "0111000011101100", -- t[28908] = 12
      "001100" when "0111000011101101", -- t[28909] = 12
      "001100" when "0111000011101110", -- t[28910] = 12
      "001100" when "0111000011101111", -- t[28911] = 12
      "001100" when "0111000011110000", -- t[28912] = 12
      "001100" when "0111000011110001", -- t[28913] = 12
      "001100" when "0111000011110010", -- t[28914] = 12
      "001100" when "0111000011110011", -- t[28915] = 12
      "001100" when "0111000011110100", -- t[28916] = 12
      "001100" when "0111000011110101", -- t[28917] = 12
      "001100" when "0111000011110110", -- t[28918] = 12
      "001100" when "0111000011110111", -- t[28919] = 12
      "001100" when "0111000011111000", -- t[28920] = 12
      "001100" when "0111000011111001", -- t[28921] = 12
      "001100" when "0111000011111010", -- t[28922] = 12
      "001100" when "0111000011111011", -- t[28923] = 12
      "001100" when "0111000011111100", -- t[28924] = 12
      "001100" when "0111000011111101", -- t[28925] = 12
      "001100" when "0111000011111110", -- t[28926] = 12
      "001100" when "0111000011111111", -- t[28927] = 12
      "001100" when "0111000100000000", -- t[28928] = 12
      "001100" when "0111000100000001", -- t[28929] = 12
      "001100" when "0111000100000010", -- t[28930] = 12
      "001100" when "0111000100000011", -- t[28931] = 12
      "001100" when "0111000100000100", -- t[28932] = 12
      "001100" when "0111000100000101", -- t[28933] = 12
      "001100" when "0111000100000110", -- t[28934] = 12
      "001100" when "0111000100000111", -- t[28935] = 12
      "001100" when "0111000100001000", -- t[28936] = 12
      "001100" when "0111000100001001", -- t[28937] = 12
      "001100" when "0111000100001010", -- t[28938] = 12
      "001100" when "0111000100001011", -- t[28939] = 12
      "001100" when "0111000100001100", -- t[28940] = 12
      "001100" when "0111000100001101", -- t[28941] = 12
      "001100" when "0111000100001110", -- t[28942] = 12
      "001100" when "0111000100001111", -- t[28943] = 12
      "001100" when "0111000100010000", -- t[28944] = 12
      "001100" when "0111000100010001", -- t[28945] = 12
      "001100" when "0111000100010010", -- t[28946] = 12
      "001100" when "0111000100010011", -- t[28947] = 12
      "001100" when "0111000100010100", -- t[28948] = 12
      "001100" when "0111000100010101", -- t[28949] = 12
      "001100" when "0111000100010110", -- t[28950] = 12
      "001100" when "0111000100010111", -- t[28951] = 12
      "001100" when "0111000100011000", -- t[28952] = 12
      "001100" when "0111000100011001", -- t[28953] = 12
      "001100" when "0111000100011010", -- t[28954] = 12
      "001100" when "0111000100011011", -- t[28955] = 12
      "001100" when "0111000100011100", -- t[28956] = 12
      "001100" when "0111000100011101", -- t[28957] = 12
      "001100" when "0111000100011110", -- t[28958] = 12
      "001100" when "0111000100011111", -- t[28959] = 12
      "001100" when "0111000100100000", -- t[28960] = 12
      "001100" when "0111000100100001", -- t[28961] = 12
      "001100" when "0111000100100010", -- t[28962] = 12
      "001100" when "0111000100100011", -- t[28963] = 12
      "001100" when "0111000100100100", -- t[28964] = 12
      "001100" when "0111000100100101", -- t[28965] = 12
      "001100" when "0111000100100110", -- t[28966] = 12
      "001100" when "0111000100100111", -- t[28967] = 12
      "001100" when "0111000100101000", -- t[28968] = 12
      "001100" when "0111000100101001", -- t[28969] = 12
      "001100" when "0111000100101010", -- t[28970] = 12
      "001100" when "0111000100101011", -- t[28971] = 12
      "001100" when "0111000100101100", -- t[28972] = 12
      "001100" when "0111000100101101", -- t[28973] = 12
      "001100" when "0111000100101110", -- t[28974] = 12
      "001100" when "0111000100101111", -- t[28975] = 12
      "001100" when "0111000100110000", -- t[28976] = 12
      "001100" when "0111000100110001", -- t[28977] = 12
      "001100" when "0111000100110010", -- t[28978] = 12
      "001100" when "0111000100110011", -- t[28979] = 12
      "001100" when "0111000100110100", -- t[28980] = 12
      "001100" when "0111000100110101", -- t[28981] = 12
      "001100" when "0111000100110110", -- t[28982] = 12
      "001100" when "0111000100110111", -- t[28983] = 12
      "001100" when "0111000100111000", -- t[28984] = 12
      "001100" when "0111000100111001", -- t[28985] = 12
      "001100" when "0111000100111010", -- t[28986] = 12
      "001100" when "0111000100111011", -- t[28987] = 12
      "001100" when "0111000100111100", -- t[28988] = 12
      "001100" when "0111000100111101", -- t[28989] = 12
      "001100" when "0111000100111110", -- t[28990] = 12
      "001100" when "0111000100111111", -- t[28991] = 12
      "001100" when "0111000101000000", -- t[28992] = 12
      "001100" when "0111000101000001", -- t[28993] = 12
      "001100" when "0111000101000010", -- t[28994] = 12
      "001100" when "0111000101000011", -- t[28995] = 12
      "001100" when "0111000101000100", -- t[28996] = 12
      "001100" when "0111000101000101", -- t[28997] = 12
      "001100" when "0111000101000110", -- t[28998] = 12
      "001100" when "0111000101000111", -- t[28999] = 12
      "001100" when "0111000101001000", -- t[29000] = 12
      "001100" when "0111000101001001", -- t[29001] = 12
      "001100" when "0111000101001010", -- t[29002] = 12
      "001100" when "0111000101001011", -- t[29003] = 12
      "001100" when "0111000101001100", -- t[29004] = 12
      "001100" when "0111000101001101", -- t[29005] = 12
      "001100" when "0111000101001110", -- t[29006] = 12
      "001100" when "0111000101001111", -- t[29007] = 12
      "001100" when "0111000101010000", -- t[29008] = 12
      "001100" when "0111000101010001", -- t[29009] = 12
      "001100" when "0111000101010010", -- t[29010] = 12
      "001100" when "0111000101010011", -- t[29011] = 12
      "001100" when "0111000101010100", -- t[29012] = 12
      "001100" when "0111000101010101", -- t[29013] = 12
      "001100" when "0111000101010110", -- t[29014] = 12
      "001100" when "0111000101010111", -- t[29015] = 12
      "001100" when "0111000101011000", -- t[29016] = 12
      "001100" when "0111000101011001", -- t[29017] = 12
      "001100" when "0111000101011010", -- t[29018] = 12
      "001100" when "0111000101011011", -- t[29019] = 12
      "001100" when "0111000101011100", -- t[29020] = 12
      "001100" when "0111000101011101", -- t[29021] = 12
      "001100" when "0111000101011110", -- t[29022] = 12
      "001100" when "0111000101011111", -- t[29023] = 12
      "001100" when "0111000101100000", -- t[29024] = 12
      "001100" when "0111000101100001", -- t[29025] = 12
      "001100" when "0111000101100010", -- t[29026] = 12
      "001100" when "0111000101100011", -- t[29027] = 12
      "001100" when "0111000101100100", -- t[29028] = 12
      "001100" when "0111000101100101", -- t[29029] = 12
      "001100" when "0111000101100110", -- t[29030] = 12
      "001100" when "0111000101100111", -- t[29031] = 12
      "001100" when "0111000101101000", -- t[29032] = 12
      "001100" when "0111000101101001", -- t[29033] = 12
      "001100" when "0111000101101010", -- t[29034] = 12
      "001100" when "0111000101101011", -- t[29035] = 12
      "001100" when "0111000101101100", -- t[29036] = 12
      "001100" when "0111000101101101", -- t[29037] = 12
      "001100" when "0111000101101110", -- t[29038] = 12
      "001100" when "0111000101101111", -- t[29039] = 12
      "001100" when "0111000101110000", -- t[29040] = 12
      "001100" when "0111000101110001", -- t[29041] = 12
      "001100" when "0111000101110010", -- t[29042] = 12
      "001100" when "0111000101110011", -- t[29043] = 12
      "001100" when "0111000101110100", -- t[29044] = 12
      "001100" when "0111000101110101", -- t[29045] = 12
      "001100" when "0111000101110110", -- t[29046] = 12
      "001100" when "0111000101110111", -- t[29047] = 12
      "001100" when "0111000101111000", -- t[29048] = 12
      "001100" when "0111000101111001", -- t[29049] = 12
      "001100" when "0111000101111010", -- t[29050] = 12
      "001100" when "0111000101111011", -- t[29051] = 12
      "001100" when "0111000101111100", -- t[29052] = 12
      "001100" when "0111000101111101", -- t[29053] = 12
      "001100" when "0111000101111110", -- t[29054] = 12
      "001100" when "0111000101111111", -- t[29055] = 12
      "001100" when "0111000110000000", -- t[29056] = 12
      "001100" when "0111000110000001", -- t[29057] = 12
      "001100" when "0111000110000010", -- t[29058] = 12
      "001100" when "0111000110000011", -- t[29059] = 12
      "001100" when "0111000110000100", -- t[29060] = 12
      "001100" when "0111000110000101", -- t[29061] = 12
      "001100" when "0111000110000110", -- t[29062] = 12
      "001100" when "0111000110000111", -- t[29063] = 12
      "001100" when "0111000110001000", -- t[29064] = 12
      "001100" when "0111000110001001", -- t[29065] = 12
      "001100" when "0111000110001010", -- t[29066] = 12
      "001100" when "0111000110001011", -- t[29067] = 12
      "001100" when "0111000110001100", -- t[29068] = 12
      "001100" when "0111000110001101", -- t[29069] = 12
      "001100" when "0111000110001110", -- t[29070] = 12
      "001100" when "0111000110001111", -- t[29071] = 12
      "001100" when "0111000110010000", -- t[29072] = 12
      "001100" when "0111000110010001", -- t[29073] = 12
      "001100" when "0111000110010010", -- t[29074] = 12
      "001100" when "0111000110010011", -- t[29075] = 12
      "001100" when "0111000110010100", -- t[29076] = 12
      "001100" when "0111000110010101", -- t[29077] = 12
      "001100" when "0111000110010110", -- t[29078] = 12
      "001100" when "0111000110010111", -- t[29079] = 12
      "001100" when "0111000110011000", -- t[29080] = 12
      "001100" when "0111000110011001", -- t[29081] = 12
      "001100" when "0111000110011010", -- t[29082] = 12
      "001100" when "0111000110011011", -- t[29083] = 12
      "001100" when "0111000110011100", -- t[29084] = 12
      "001100" when "0111000110011101", -- t[29085] = 12
      "001100" when "0111000110011110", -- t[29086] = 12
      "001100" when "0111000110011111", -- t[29087] = 12
      "001100" when "0111000110100000", -- t[29088] = 12
      "001100" when "0111000110100001", -- t[29089] = 12
      "001100" when "0111000110100010", -- t[29090] = 12
      "001100" when "0111000110100011", -- t[29091] = 12
      "001100" when "0111000110100100", -- t[29092] = 12
      "001100" when "0111000110100101", -- t[29093] = 12
      "001100" when "0111000110100110", -- t[29094] = 12
      "001100" when "0111000110100111", -- t[29095] = 12
      "001100" when "0111000110101000", -- t[29096] = 12
      "001100" when "0111000110101001", -- t[29097] = 12
      "001100" when "0111000110101010", -- t[29098] = 12
      "001100" when "0111000110101011", -- t[29099] = 12
      "001100" when "0111000110101100", -- t[29100] = 12
      "001100" when "0111000110101101", -- t[29101] = 12
      "001100" when "0111000110101110", -- t[29102] = 12
      "001100" when "0111000110101111", -- t[29103] = 12
      "001100" when "0111000110110000", -- t[29104] = 12
      "001100" when "0111000110110001", -- t[29105] = 12
      "001100" when "0111000110110010", -- t[29106] = 12
      "001100" when "0111000110110011", -- t[29107] = 12
      "001100" when "0111000110110100", -- t[29108] = 12
      "001100" when "0111000110110101", -- t[29109] = 12
      "001100" when "0111000110110110", -- t[29110] = 12
      "001100" when "0111000110110111", -- t[29111] = 12
      "001100" when "0111000110111000", -- t[29112] = 12
      "001100" when "0111000110111001", -- t[29113] = 12
      "001100" when "0111000110111010", -- t[29114] = 12
      "001100" when "0111000110111011", -- t[29115] = 12
      "001100" when "0111000110111100", -- t[29116] = 12
      "001100" when "0111000110111101", -- t[29117] = 12
      "001100" when "0111000110111110", -- t[29118] = 12
      "001100" when "0111000110111111", -- t[29119] = 12
      "001100" when "0111000111000000", -- t[29120] = 12
      "001100" when "0111000111000001", -- t[29121] = 12
      "001100" when "0111000111000010", -- t[29122] = 12
      "001100" when "0111000111000011", -- t[29123] = 12
      "001100" when "0111000111000100", -- t[29124] = 12
      "001100" when "0111000111000101", -- t[29125] = 12
      "001100" when "0111000111000110", -- t[29126] = 12
      "001100" when "0111000111000111", -- t[29127] = 12
      "001100" when "0111000111001000", -- t[29128] = 12
      "001100" when "0111000111001001", -- t[29129] = 12
      "001100" when "0111000111001010", -- t[29130] = 12
      "001100" when "0111000111001011", -- t[29131] = 12
      "001100" when "0111000111001100", -- t[29132] = 12
      "001100" when "0111000111001101", -- t[29133] = 12
      "001100" when "0111000111001110", -- t[29134] = 12
      "001100" when "0111000111001111", -- t[29135] = 12
      "001100" when "0111000111010000", -- t[29136] = 12
      "001100" when "0111000111010001", -- t[29137] = 12
      "001101" when "0111000111010010", -- t[29138] = 13
      "001101" when "0111000111010011", -- t[29139] = 13
      "001101" when "0111000111010100", -- t[29140] = 13
      "001101" when "0111000111010101", -- t[29141] = 13
      "001101" when "0111000111010110", -- t[29142] = 13
      "001101" when "0111000111010111", -- t[29143] = 13
      "001101" when "0111000111011000", -- t[29144] = 13
      "001101" when "0111000111011001", -- t[29145] = 13
      "001101" when "0111000111011010", -- t[29146] = 13
      "001101" when "0111000111011011", -- t[29147] = 13
      "001101" when "0111000111011100", -- t[29148] = 13
      "001101" when "0111000111011101", -- t[29149] = 13
      "001101" when "0111000111011110", -- t[29150] = 13
      "001101" when "0111000111011111", -- t[29151] = 13
      "001101" when "0111000111100000", -- t[29152] = 13
      "001101" when "0111000111100001", -- t[29153] = 13
      "001101" when "0111000111100010", -- t[29154] = 13
      "001101" when "0111000111100011", -- t[29155] = 13
      "001101" when "0111000111100100", -- t[29156] = 13
      "001101" when "0111000111100101", -- t[29157] = 13
      "001101" when "0111000111100110", -- t[29158] = 13
      "001101" when "0111000111100111", -- t[29159] = 13
      "001101" when "0111000111101000", -- t[29160] = 13
      "001101" when "0111000111101001", -- t[29161] = 13
      "001101" when "0111000111101010", -- t[29162] = 13
      "001101" when "0111000111101011", -- t[29163] = 13
      "001101" when "0111000111101100", -- t[29164] = 13
      "001101" when "0111000111101101", -- t[29165] = 13
      "001101" when "0111000111101110", -- t[29166] = 13
      "001101" when "0111000111101111", -- t[29167] = 13
      "001101" when "0111000111110000", -- t[29168] = 13
      "001101" when "0111000111110001", -- t[29169] = 13
      "001101" when "0111000111110010", -- t[29170] = 13
      "001101" when "0111000111110011", -- t[29171] = 13
      "001101" when "0111000111110100", -- t[29172] = 13
      "001101" when "0111000111110101", -- t[29173] = 13
      "001101" when "0111000111110110", -- t[29174] = 13
      "001101" when "0111000111110111", -- t[29175] = 13
      "001101" when "0111000111111000", -- t[29176] = 13
      "001101" when "0111000111111001", -- t[29177] = 13
      "001101" when "0111000111111010", -- t[29178] = 13
      "001101" when "0111000111111011", -- t[29179] = 13
      "001101" when "0111000111111100", -- t[29180] = 13
      "001101" when "0111000111111101", -- t[29181] = 13
      "001101" when "0111000111111110", -- t[29182] = 13
      "001101" when "0111000111111111", -- t[29183] = 13
      "001101" when "0111001000000000", -- t[29184] = 13
      "001101" when "0111001000000001", -- t[29185] = 13
      "001101" when "0111001000000010", -- t[29186] = 13
      "001101" when "0111001000000011", -- t[29187] = 13
      "001101" when "0111001000000100", -- t[29188] = 13
      "001101" when "0111001000000101", -- t[29189] = 13
      "001101" when "0111001000000110", -- t[29190] = 13
      "001101" when "0111001000000111", -- t[29191] = 13
      "001101" when "0111001000001000", -- t[29192] = 13
      "001101" when "0111001000001001", -- t[29193] = 13
      "001101" when "0111001000001010", -- t[29194] = 13
      "001101" when "0111001000001011", -- t[29195] = 13
      "001101" when "0111001000001100", -- t[29196] = 13
      "001101" when "0111001000001101", -- t[29197] = 13
      "001101" when "0111001000001110", -- t[29198] = 13
      "001101" when "0111001000001111", -- t[29199] = 13
      "001101" when "0111001000010000", -- t[29200] = 13
      "001101" when "0111001000010001", -- t[29201] = 13
      "001101" when "0111001000010010", -- t[29202] = 13
      "001101" when "0111001000010011", -- t[29203] = 13
      "001101" when "0111001000010100", -- t[29204] = 13
      "001101" when "0111001000010101", -- t[29205] = 13
      "001101" when "0111001000010110", -- t[29206] = 13
      "001101" when "0111001000010111", -- t[29207] = 13
      "001101" when "0111001000011000", -- t[29208] = 13
      "001101" when "0111001000011001", -- t[29209] = 13
      "001101" when "0111001000011010", -- t[29210] = 13
      "001101" when "0111001000011011", -- t[29211] = 13
      "001101" when "0111001000011100", -- t[29212] = 13
      "001101" when "0111001000011101", -- t[29213] = 13
      "001101" when "0111001000011110", -- t[29214] = 13
      "001101" when "0111001000011111", -- t[29215] = 13
      "001101" when "0111001000100000", -- t[29216] = 13
      "001101" when "0111001000100001", -- t[29217] = 13
      "001101" when "0111001000100010", -- t[29218] = 13
      "001101" when "0111001000100011", -- t[29219] = 13
      "001101" when "0111001000100100", -- t[29220] = 13
      "001101" when "0111001000100101", -- t[29221] = 13
      "001101" when "0111001000100110", -- t[29222] = 13
      "001101" when "0111001000100111", -- t[29223] = 13
      "001101" when "0111001000101000", -- t[29224] = 13
      "001101" when "0111001000101001", -- t[29225] = 13
      "001101" when "0111001000101010", -- t[29226] = 13
      "001101" when "0111001000101011", -- t[29227] = 13
      "001101" when "0111001000101100", -- t[29228] = 13
      "001101" when "0111001000101101", -- t[29229] = 13
      "001101" when "0111001000101110", -- t[29230] = 13
      "001101" when "0111001000101111", -- t[29231] = 13
      "001101" when "0111001000110000", -- t[29232] = 13
      "001101" when "0111001000110001", -- t[29233] = 13
      "001101" when "0111001000110010", -- t[29234] = 13
      "001101" when "0111001000110011", -- t[29235] = 13
      "001101" when "0111001000110100", -- t[29236] = 13
      "001101" when "0111001000110101", -- t[29237] = 13
      "001101" when "0111001000110110", -- t[29238] = 13
      "001101" when "0111001000110111", -- t[29239] = 13
      "001101" when "0111001000111000", -- t[29240] = 13
      "001101" when "0111001000111001", -- t[29241] = 13
      "001101" when "0111001000111010", -- t[29242] = 13
      "001101" when "0111001000111011", -- t[29243] = 13
      "001101" when "0111001000111100", -- t[29244] = 13
      "001101" when "0111001000111101", -- t[29245] = 13
      "001101" when "0111001000111110", -- t[29246] = 13
      "001101" when "0111001000111111", -- t[29247] = 13
      "001101" when "0111001001000000", -- t[29248] = 13
      "001101" when "0111001001000001", -- t[29249] = 13
      "001101" when "0111001001000010", -- t[29250] = 13
      "001101" when "0111001001000011", -- t[29251] = 13
      "001101" when "0111001001000100", -- t[29252] = 13
      "001101" when "0111001001000101", -- t[29253] = 13
      "001101" when "0111001001000110", -- t[29254] = 13
      "001101" when "0111001001000111", -- t[29255] = 13
      "001101" when "0111001001001000", -- t[29256] = 13
      "001101" when "0111001001001001", -- t[29257] = 13
      "001101" when "0111001001001010", -- t[29258] = 13
      "001101" when "0111001001001011", -- t[29259] = 13
      "001101" when "0111001001001100", -- t[29260] = 13
      "001101" when "0111001001001101", -- t[29261] = 13
      "001101" when "0111001001001110", -- t[29262] = 13
      "001101" when "0111001001001111", -- t[29263] = 13
      "001101" when "0111001001010000", -- t[29264] = 13
      "001101" when "0111001001010001", -- t[29265] = 13
      "001101" when "0111001001010010", -- t[29266] = 13
      "001101" when "0111001001010011", -- t[29267] = 13
      "001101" when "0111001001010100", -- t[29268] = 13
      "001101" when "0111001001010101", -- t[29269] = 13
      "001101" when "0111001001010110", -- t[29270] = 13
      "001101" when "0111001001010111", -- t[29271] = 13
      "001101" when "0111001001011000", -- t[29272] = 13
      "001101" when "0111001001011001", -- t[29273] = 13
      "001101" when "0111001001011010", -- t[29274] = 13
      "001101" when "0111001001011011", -- t[29275] = 13
      "001101" when "0111001001011100", -- t[29276] = 13
      "001101" when "0111001001011101", -- t[29277] = 13
      "001101" when "0111001001011110", -- t[29278] = 13
      "001101" when "0111001001011111", -- t[29279] = 13
      "001101" when "0111001001100000", -- t[29280] = 13
      "001101" when "0111001001100001", -- t[29281] = 13
      "001101" when "0111001001100010", -- t[29282] = 13
      "001101" when "0111001001100011", -- t[29283] = 13
      "001101" when "0111001001100100", -- t[29284] = 13
      "001101" when "0111001001100101", -- t[29285] = 13
      "001101" when "0111001001100110", -- t[29286] = 13
      "001101" when "0111001001100111", -- t[29287] = 13
      "001101" when "0111001001101000", -- t[29288] = 13
      "001101" when "0111001001101001", -- t[29289] = 13
      "001101" when "0111001001101010", -- t[29290] = 13
      "001101" when "0111001001101011", -- t[29291] = 13
      "001101" when "0111001001101100", -- t[29292] = 13
      "001101" when "0111001001101101", -- t[29293] = 13
      "001101" when "0111001001101110", -- t[29294] = 13
      "001101" when "0111001001101111", -- t[29295] = 13
      "001101" when "0111001001110000", -- t[29296] = 13
      "001101" when "0111001001110001", -- t[29297] = 13
      "001101" when "0111001001110010", -- t[29298] = 13
      "001101" when "0111001001110011", -- t[29299] = 13
      "001101" when "0111001001110100", -- t[29300] = 13
      "001101" when "0111001001110101", -- t[29301] = 13
      "001101" when "0111001001110110", -- t[29302] = 13
      "001101" when "0111001001110111", -- t[29303] = 13
      "001101" when "0111001001111000", -- t[29304] = 13
      "001101" when "0111001001111001", -- t[29305] = 13
      "001101" when "0111001001111010", -- t[29306] = 13
      "001101" when "0111001001111011", -- t[29307] = 13
      "001101" when "0111001001111100", -- t[29308] = 13
      "001101" when "0111001001111101", -- t[29309] = 13
      "001101" when "0111001001111110", -- t[29310] = 13
      "001101" when "0111001001111111", -- t[29311] = 13
      "001101" when "0111001010000000", -- t[29312] = 13
      "001101" when "0111001010000001", -- t[29313] = 13
      "001101" when "0111001010000010", -- t[29314] = 13
      "001101" when "0111001010000011", -- t[29315] = 13
      "001101" when "0111001010000100", -- t[29316] = 13
      "001101" when "0111001010000101", -- t[29317] = 13
      "001101" when "0111001010000110", -- t[29318] = 13
      "001101" when "0111001010000111", -- t[29319] = 13
      "001101" when "0111001010001000", -- t[29320] = 13
      "001101" when "0111001010001001", -- t[29321] = 13
      "001101" when "0111001010001010", -- t[29322] = 13
      "001101" when "0111001010001011", -- t[29323] = 13
      "001101" when "0111001010001100", -- t[29324] = 13
      "001101" when "0111001010001101", -- t[29325] = 13
      "001101" when "0111001010001110", -- t[29326] = 13
      "001101" when "0111001010001111", -- t[29327] = 13
      "001101" when "0111001010010000", -- t[29328] = 13
      "001101" when "0111001010010001", -- t[29329] = 13
      "001101" when "0111001010010010", -- t[29330] = 13
      "001101" when "0111001010010011", -- t[29331] = 13
      "001101" when "0111001010010100", -- t[29332] = 13
      "001101" when "0111001010010101", -- t[29333] = 13
      "001101" when "0111001010010110", -- t[29334] = 13
      "001101" when "0111001010010111", -- t[29335] = 13
      "001101" when "0111001010011000", -- t[29336] = 13
      "001101" when "0111001010011001", -- t[29337] = 13
      "001101" when "0111001010011010", -- t[29338] = 13
      "001101" when "0111001010011011", -- t[29339] = 13
      "001101" when "0111001010011100", -- t[29340] = 13
      "001101" when "0111001010011101", -- t[29341] = 13
      "001101" when "0111001010011110", -- t[29342] = 13
      "001101" when "0111001010011111", -- t[29343] = 13
      "001101" when "0111001010100000", -- t[29344] = 13
      "001101" when "0111001010100001", -- t[29345] = 13
      "001101" when "0111001010100010", -- t[29346] = 13
      "001101" when "0111001010100011", -- t[29347] = 13
      "001101" when "0111001010100100", -- t[29348] = 13
      "001101" when "0111001010100101", -- t[29349] = 13
      "001101" when "0111001010100110", -- t[29350] = 13
      "001101" when "0111001010100111", -- t[29351] = 13
      "001101" when "0111001010101000", -- t[29352] = 13
      "001101" when "0111001010101001", -- t[29353] = 13
      "001101" when "0111001010101010", -- t[29354] = 13
      "001101" when "0111001010101011", -- t[29355] = 13
      "001101" when "0111001010101100", -- t[29356] = 13
      "001101" when "0111001010101101", -- t[29357] = 13
      "001101" when "0111001010101110", -- t[29358] = 13
      "001101" when "0111001010101111", -- t[29359] = 13
      "001101" when "0111001010110000", -- t[29360] = 13
      "001101" when "0111001010110001", -- t[29361] = 13
      "001101" when "0111001010110010", -- t[29362] = 13
      "001101" when "0111001010110011", -- t[29363] = 13
      "001101" when "0111001010110100", -- t[29364] = 13
      "001101" when "0111001010110101", -- t[29365] = 13
      "001101" when "0111001010110110", -- t[29366] = 13
      "001101" when "0111001010110111", -- t[29367] = 13
      "001101" when "0111001010111000", -- t[29368] = 13
      "001101" when "0111001010111001", -- t[29369] = 13
      "001101" when "0111001010111010", -- t[29370] = 13
      "001101" when "0111001010111011", -- t[29371] = 13
      "001101" when "0111001010111100", -- t[29372] = 13
      "001101" when "0111001010111101", -- t[29373] = 13
      "001101" when "0111001010111110", -- t[29374] = 13
      "001101" when "0111001010111111", -- t[29375] = 13
      "001101" when "0111001011000000", -- t[29376] = 13
      "001101" when "0111001011000001", -- t[29377] = 13
      "001101" when "0111001011000010", -- t[29378] = 13
      "001101" when "0111001011000011", -- t[29379] = 13
      "001101" when "0111001011000100", -- t[29380] = 13
      "001101" when "0111001011000101", -- t[29381] = 13
      "001101" when "0111001011000110", -- t[29382] = 13
      "001101" when "0111001011000111", -- t[29383] = 13
      "001101" when "0111001011001000", -- t[29384] = 13
      "001101" when "0111001011001001", -- t[29385] = 13
      "001101" when "0111001011001010", -- t[29386] = 13
      "001101" when "0111001011001011", -- t[29387] = 13
      "001101" when "0111001011001100", -- t[29388] = 13
      "001101" when "0111001011001101", -- t[29389] = 13
      "001101" when "0111001011001110", -- t[29390] = 13
      "001101" when "0111001011001111", -- t[29391] = 13
      "001101" when "0111001011010000", -- t[29392] = 13
      "001101" when "0111001011010001", -- t[29393] = 13
      "001101" when "0111001011010010", -- t[29394] = 13
      "001101" when "0111001011010011", -- t[29395] = 13
      "001101" when "0111001011010100", -- t[29396] = 13
      "001101" when "0111001011010101", -- t[29397] = 13
      "001101" when "0111001011010110", -- t[29398] = 13
      "001101" when "0111001011010111", -- t[29399] = 13
      "001101" when "0111001011011000", -- t[29400] = 13
      "001101" when "0111001011011001", -- t[29401] = 13
      "001101" when "0111001011011010", -- t[29402] = 13
      "001101" when "0111001011011011", -- t[29403] = 13
      "001101" when "0111001011011100", -- t[29404] = 13
      "001101" when "0111001011011101", -- t[29405] = 13
      "001101" when "0111001011011110", -- t[29406] = 13
      "001101" when "0111001011011111", -- t[29407] = 13
      "001101" when "0111001011100000", -- t[29408] = 13
      "001101" when "0111001011100001", -- t[29409] = 13
      "001101" when "0111001011100010", -- t[29410] = 13
      "001101" when "0111001011100011", -- t[29411] = 13
      "001101" when "0111001011100100", -- t[29412] = 13
      "001101" when "0111001011100101", -- t[29413] = 13
      "001101" when "0111001011100110", -- t[29414] = 13
      "001101" when "0111001011100111", -- t[29415] = 13
      "001101" when "0111001011101000", -- t[29416] = 13
      "001101" when "0111001011101001", -- t[29417] = 13
      "001101" when "0111001011101010", -- t[29418] = 13
      "001101" when "0111001011101011", -- t[29419] = 13
      "001101" when "0111001011101100", -- t[29420] = 13
      "001101" when "0111001011101101", -- t[29421] = 13
      "001101" when "0111001011101110", -- t[29422] = 13
      "001101" when "0111001011101111", -- t[29423] = 13
      "001101" when "0111001011110000", -- t[29424] = 13
      "001101" when "0111001011110001", -- t[29425] = 13
      "001101" when "0111001011110010", -- t[29426] = 13
      "001101" when "0111001011110011", -- t[29427] = 13
      "001101" when "0111001011110100", -- t[29428] = 13
      "001101" when "0111001011110101", -- t[29429] = 13
      "001101" when "0111001011110110", -- t[29430] = 13
      "001101" when "0111001011110111", -- t[29431] = 13
      "001101" when "0111001011111000", -- t[29432] = 13
      "001101" when "0111001011111001", -- t[29433] = 13
      "001101" when "0111001011111010", -- t[29434] = 13
      "001101" when "0111001011111011", -- t[29435] = 13
      "001101" when "0111001011111100", -- t[29436] = 13
      "001101" when "0111001011111101", -- t[29437] = 13
      "001101" when "0111001011111110", -- t[29438] = 13
      "001101" when "0111001011111111", -- t[29439] = 13
      "001101" when "0111001100000000", -- t[29440] = 13
      "001101" when "0111001100000001", -- t[29441] = 13
      "001101" when "0111001100000010", -- t[29442] = 13
      "001101" when "0111001100000011", -- t[29443] = 13
      "001101" when "0111001100000100", -- t[29444] = 13
      "001101" when "0111001100000101", -- t[29445] = 13
      "001101" when "0111001100000110", -- t[29446] = 13
      "001101" when "0111001100000111", -- t[29447] = 13
      "001101" when "0111001100001000", -- t[29448] = 13
      "001101" when "0111001100001001", -- t[29449] = 13
      "001101" when "0111001100001010", -- t[29450] = 13
      "001101" when "0111001100001011", -- t[29451] = 13
      "001101" when "0111001100001100", -- t[29452] = 13
      "001101" when "0111001100001101", -- t[29453] = 13
      "001101" when "0111001100001110", -- t[29454] = 13
      "001101" when "0111001100001111", -- t[29455] = 13
      "001101" when "0111001100010000", -- t[29456] = 13
      "001101" when "0111001100010001", -- t[29457] = 13
      "001101" when "0111001100010010", -- t[29458] = 13
      "001101" when "0111001100010011", -- t[29459] = 13
      "001101" when "0111001100010100", -- t[29460] = 13
      "001101" when "0111001100010101", -- t[29461] = 13
      "001101" when "0111001100010110", -- t[29462] = 13
      "001101" when "0111001100010111", -- t[29463] = 13
      "001101" when "0111001100011000", -- t[29464] = 13
      "001101" when "0111001100011001", -- t[29465] = 13
      "001101" when "0111001100011010", -- t[29466] = 13
      "001101" when "0111001100011011", -- t[29467] = 13
      "001101" when "0111001100011100", -- t[29468] = 13
      "001101" when "0111001100011101", -- t[29469] = 13
      "001101" when "0111001100011110", -- t[29470] = 13
      "001101" when "0111001100011111", -- t[29471] = 13
      "001101" when "0111001100100000", -- t[29472] = 13
      "001101" when "0111001100100001", -- t[29473] = 13
      "001101" when "0111001100100010", -- t[29474] = 13
      "001101" when "0111001100100011", -- t[29475] = 13
      "001101" when "0111001100100100", -- t[29476] = 13
      "001101" when "0111001100100101", -- t[29477] = 13
      "001101" when "0111001100100110", -- t[29478] = 13
      "001101" when "0111001100100111", -- t[29479] = 13
      "001101" when "0111001100101000", -- t[29480] = 13
      "001101" when "0111001100101001", -- t[29481] = 13
      "001101" when "0111001100101010", -- t[29482] = 13
      "001101" when "0111001100101011", -- t[29483] = 13
      "001101" when "0111001100101100", -- t[29484] = 13
      "001101" when "0111001100101101", -- t[29485] = 13
      "001101" when "0111001100101110", -- t[29486] = 13
      "001101" when "0111001100101111", -- t[29487] = 13
      "001101" when "0111001100110000", -- t[29488] = 13
      "001101" when "0111001100110001", -- t[29489] = 13
      "001101" when "0111001100110010", -- t[29490] = 13
      "001101" when "0111001100110011", -- t[29491] = 13
      "001101" when "0111001100110100", -- t[29492] = 13
      "001101" when "0111001100110101", -- t[29493] = 13
      "001101" when "0111001100110110", -- t[29494] = 13
      "001101" when "0111001100110111", -- t[29495] = 13
      "001101" when "0111001100111000", -- t[29496] = 13
      "001101" when "0111001100111001", -- t[29497] = 13
      "001101" when "0111001100111010", -- t[29498] = 13
      "001101" when "0111001100111011", -- t[29499] = 13
      "001101" when "0111001100111100", -- t[29500] = 13
      "001101" when "0111001100111101", -- t[29501] = 13
      "001101" when "0111001100111110", -- t[29502] = 13
      "001101" when "0111001100111111", -- t[29503] = 13
      "001101" when "0111001101000000", -- t[29504] = 13
      "001101" when "0111001101000001", -- t[29505] = 13
      "001101" when "0111001101000010", -- t[29506] = 13
      "001101" when "0111001101000011", -- t[29507] = 13
      "001101" when "0111001101000100", -- t[29508] = 13
      "001101" when "0111001101000101", -- t[29509] = 13
      "001101" when "0111001101000110", -- t[29510] = 13
      "001101" when "0111001101000111", -- t[29511] = 13
      "001101" when "0111001101001000", -- t[29512] = 13
      "001101" when "0111001101001001", -- t[29513] = 13
      "001101" when "0111001101001010", -- t[29514] = 13
      "001101" when "0111001101001011", -- t[29515] = 13
      "001101" when "0111001101001100", -- t[29516] = 13
      "001101" when "0111001101001101", -- t[29517] = 13
      "001101" when "0111001101001110", -- t[29518] = 13
      "001101" when "0111001101001111", -- t[29519] = 13
      "001101" when "0111001101010000", -- t[29520] = 13
      "001101" when "0111001101010001", -- t[29521] = 13
      "001101" when "0111001101010010", -- t[29522] = 13
      "001101" when "0111001101010011", -- t[29523] = 13
      "001101" when "0111001101010100", -- t[29524] = 13
      "001101" when "0111001101010101", -- t[29525] = 13
      "001101" when "0111001101010110", -- t[29526] = 13
      "001101" when "0111001101010111", -- t[29527] = 13
      "001101" when "0111001101011000", -- t[29528] = 13
      "001101" when "0111001101011001", -- t[29529] = 13
      "001101" when "0111001101011010", -- t[29530] = 13
      "001101" when "0111001101011011", -- t[29531] = 13
      "001101" when "0111001101011100", -- t[29532] = 13
      "001101" when "0111001101011101", -- t[29533] = 13
      "001101" when "0111001101011110", -- t[29534] = 13
      "001101" when "0111001101011111", -- t[29535] = 13
      "001101" when "0111001101100000", -- t[29536] = 13
      "001101" when "0111001101100001", -- t[29537] = 13
      "001101" when "0111001101100010", -- t[29538] = 13
      "001101" when "0111001101100011", -- t[29539] = 13
      "001101" when "0111001101100100", -- t[29540] = 13
      "001101" when "0111001101100101", -- t[29541] = 13
      "001101" when "0111001101100110", -- t[29542] = 13
      "001101" when "0111001101100111", -- t[29543] = 13
      "001101" when "0111001101101000", -- t[29544] = 13
      "001101" when "0111001101101001", -- t[29545] = 13
      "001101" when "0111001101101010", -- t[29546] = 13
      "001101" when "0111001101101011", -- t[29547] = 13
      "001101" when "0111001101101100", -- t[29548] = 13
      "001101" when "0111001101101101", -- t[29549] = 13
      "001101" when "0111001101101110", -- t[29550] = 13
      "001101" when "0111001101101111", -- t[29551] = 13
      "001101" when "0111001101110000", -- t[29552] = 13
      "001101" when "0111001101110001", -- t[29553] = 13
      "001101" when "0111001101110010", -- t[29554] = 13
      "001101" when "0111001101110011", -- t[29555] = 13
      "001101" when "0111001101110100", -- t[29556] = 13
      "001101" when "0111001101110101", -- t[29557] = 13
      "001101" when "0111001101110110", -- t[29558] = 13
      "001101" when "0111001101110111", -- t[29559] = 13
      "001101" when "0111001101111000", -- t[29560] = 13
      "001101" when "0111001101111001", -- t[29561] = 13
      "001101" when "0111001101111010", -- t[29562] = 13
      "001101" when "0111001101111011", -- t[29563] = 13
      "001101" when "0111001101111100", -- t[29564] = 13
      "001101" when "0111001101111101", -- t[29565] = 13
      "001101" when "0111001101111110", -- t[29566] = 13
      "001101" when "0111001101111111", -- t[29567] = 13
      "001101" when "0111001110000000", -- t[29568] = 13
      "001101" when "0111001110000001", -- t[29569] = 13
      "001101" when "0111001110000010", -- t[29570] = 13
      "001101" when "0111001110000011", -- t[29571] = 13
      "001101" when "0111001110000100", -- t[29572] = 13
      "001101" when "0111001110000101", -- t[29573] = 13
      "001101" when "0111001110000110", -- t[29574] = 13
      "001101" when "0111001110000111", -- t[29575] = 13
      "001101" when "0111001110001000", -- t[29576] = 13
      "001101" when "0111001110001001", -- t[29577] = 13
      "001101" when "0111001110001010", -- t[29578] = 13
      "001101" when "0111001110001011", -- t[29579] = 13
      "001101" when "0111001110001100", -- t[29580] = 13
      "001101" when "0111001110001101", -- t[29581] = 13
      "001101" when "0111001110001110", -- t[29582] = 13
      "001101" when "0111001110001111", -- t[29583] = 13
      "001101" when "0111001110010000", -- t[29584] = 13
      "001101" when "0111001110010001", -- t[29585] = 13
      "001101" when "0111001110010010", -- t[29586] = 13
      "001101" when "0111001110010011", -- t[29587] = 13
      "001101" when "0111001110010100", -- t[29588] = 13
      "001101" when "0111001110010101", -- t[29589] = 13
      "001101" when "0111001110010110", -- t[29590] = 13
      "001101" when "0111001110010111", -- t[29591] = 13
      "001110" when "0111001110011000", -- t[29592] = 14
      "001110" when "0111001110011001", -- t[29593] = 14
      "001110" when "0111001110011010", -- t[29594] = 14
      "001110" when "0111001110011011", -- t[29595] = 14
      "001110" when "0111001110011100", -- t[29596] = 14
      "001110" when "0111001110011101", -- t[29597] = 14
      "001110" when "0111001110011110", -- t[29598] = 14
      "001110" when "0111001110011111", -- t[29599] = 14
      "001110" when "0111001110100000", -- t[29600] = 14
      "001110" when "0111001110100001", -- t[29601] = 14
      "001110" when "0111001110100010", -- t[29602] = 14
      "001110" when "0111001110100011", -- t[29603] = 14
      "001110" when "0111001110100100", -- t[29604] = 14
      "001110" when "0111001110100101", -- t[29605] = 14
      "001110" when "0111001110100110", -- t[29606] = 14
      "001110" when "0111001110100111", -- t[29607] = 14
      "001110" when "0111001110101000", -- t[29608] = 14
      "001110" when "0111001110101001", -- t[29609] = 14
      "001110" when "0111001110101010", -- t[29610] = 14
      "001110" when "0111001110101011", -- t[29611] = 14
      "001110" when "0111001110101100", -- t[29612] = 14
      "001110" when "0111001110101101", -- t[29613] = 14
      "001110" when "0111001110101110", -- t[29614] = 14
      "001110" when "0111001110101111", -- t[29615] = 14
      "001110" when "0111001110110000", -- t[29616] = 14
      "001110" when "0111001110110001", -- t[29617] = 14
      "001110" when "0111001110110010", -- t[29618] = 14
      "001110" when "0111001110110011", -- t[29619] = 14
      "001110" when "0111001110110100", -- t[29620] = 14
      "001110" when "0111001110110101", -- t[29621] = 14
      "001110" when "0111001110110110", -- t[29622] = 14
      "001110" when "0111001110110111", -- t[29623] = 14
      "001110" when "0111001110111000", -- t[29624] = 14
      "001110" when "0111001110111001", -- t[29625] = 14
      "001110" when "0111001110111010", -- t[29626] = 14
      "001110" when "0111001110111011", -- t[29627] = 14
      "001110" when "0111001110111100", -- t[29628] = 14
      "001110" when "0111001110111101", -- t[29629] = 14
      "001110" when "0111001110111110", -- t[29630] = 14
      "001110" when "0111001110111111", -- t[29631] = 14
      "001110" when "0111001111000000", -- t[29632] = 14
      "001110" when "0111001111000001", -- t[29633] = 14
      "001110" when "0111001111000010", -- t[29634] = 14
      "001110" when "0111001111000011", -- t[29635] = 14
      "001110" when "0111001111000100", -- t[29636] = 14
      "001110" when "0111001111000101", -- t[29637] = 14
      "001110" when "0111001111000110", -- t[29638] = 14
      "001110" when "0111001111000111", -- t[29639] = 14
      "001110" when "0111001111001000", -- t[29640] = 14
      "001110" when "0111001111001001", -- t[29641] = 14
      "001110" when "0111001111001010", -- t[29642] = 14
      "001110" when "0111001111001011", -- t[29643] = 14
      "001110" when "0111001111001100", -- t[29644] = 14
      "001110" when "0111001111001101", -- t[29645] = 14
      "001110" when "0111001111001110", -- t[29646] = 14
      "001110" when "0111001111001111", -- t[29647] = 14
      "001110" when "0111001111010000", -- t[29648] = 14
      "001110" when "0111001111010001", -- t[29649] = 14
      "001110" when "0111001111010010", -- t[29650] = 14
      "001110" when "0111001111010011", -- t[29651] = 14
      "001110" when "0111001111010100", -- t[29652] = 14
      "001110" when "0111001111010101", -- t[29653] = 14
      "001110" when "0111001111010110", -- t[29654] = 14
      "001110" when "0111001111010111", -- t[29655] = 14
      "001110" when "0111001111011000", -- t[29656] = 14
      "001110" when "0111001111011001", -- t[29657] = 14
      "001110" when "0111001111011010", -- t[29658] = 14
      "001110" when "0111001111011011", -- t[29659] = 14
      "001110" when "0111001111011100", -- t[29660] = 14
      "001110" when "0111001111011101", -- t[29661] = 14
      "001110" when "0111001111011110", -- t[29662] = 14
      "001110" when "0111001111011111", -- t[29663] = 14
      "001110" when "0111001111100000", -- t[29664] = 14
      "001110" when "0111001111100001", -- t[29665] = 14
      "001110" when "0111001111100010", -- t[29666] = 14
      "001110" when "0111001111100011", -- t[29667] = 14
      "001110" when "0111001111100100", -- t[29668] = 14
      "001110" when "0111001111100101", -- t[29669] = 14
      "001110" when "0111001111100110", -- t[29670] = 14
      "001110" when "0111001111100111", -- t[29671] = 14
      "001110" when "0111001111101000", -- t[29672] = 14
      "001110" when "0111001111101001", -- t[29673] = 14
      "001110" when "0111001111101010", -- t[29674] = 14
      "001110" when "0111001111101011", -- t[29675] = 14
      "001110" when "0111001111101100", -- t[29676] = 14
      "001110" when "0111001111101101", -- t[29677] = 14
      "001110" when "0111001111101110", -- t[29678] = 14
      "001110" when "0111001111101111", -- t[29679] = 14
      "001110" when "0111001111110000", -- t[29680] = 14
      "001110" when "0111001111110001", -- t[29681] = 14
      "001110" when "0111001111110010", -- t[29682] = 14
      "001110" when "0111001111110011", -- t[29683] = 14
      "001110" when "0111001111110100", -- t[29684] = 14
      "001110" when "0111001111110101", -- t[29685] = 14
      "001110" when "0111001111110110", -- t[29686] = 14
      "001110" when "0111001111110111", -- t[29687] = 14
      "001110" when "0111001111111000", -- t[29688] = 14
      "001110" when "0111001111111001", -- t[29689] = 14
      "001110" when "0111001111111010", -- t[29690] = 14
      "001110" when "0111001111111011", -- t[29691] = 14
      "001110" when "0111001111111100", -- t[29692] = 14
      "001110" when "0111001111111101", -- t[29693] = 14
      "001110" when "0111001111111110", -- t[29694] = 14
      "001110" when "0111001111111111", -- t[29695] = 14
      "001110" when "0111010000000000", -- t[29696] = 14
      "001110" when "0111010000000001", -- t[29697] = 14
      "001110" when "0111010000000010", -- t[29698] = 14
      "001110" when "0111010000000011", -- t[29699] = 14
      "001110" when "0111010000000100", -- t[29700] = 14
      "001110" when "0111010000000101", -- t[29701] = 14
      "001110" when "0111010000000110", -- t[29702] = 14
      "001110" when "0111010000000111", -- t[29703] = 14
      "001110" when "0111010000001000", -- t[29704] = 14
      "001110" when "0111010000001001", -- t[29705] = 14
      "001110" when "0111010000001010", -- t[29706] = 14
      "001110" when "0111010000001011", -- t[29707] = 14
      "001110" when "0111010000001100", -- t[29708] = 14
      "001110" when "0111010000001101", -- t[29709] = 14
      "001110" when "0111010000001110", -- t[29710] = 14
      "001110" when "0111010000001111", -- t[29711] = 14
      "001110" when "0111010000010000", -- t[29712] = 14
      "001110" when "0111010000010001", -- t[29713] = 14
      "001110" when "0111010000010010", -- t[29714] = 14
      "001110" when "0111010000010011", -- t[29715] = 14
      "001110" when "0111010000010100", -- t[29716] = 14
      "001110" when "0111010000010101", -- t[29717] = 14
      "001110" when "0111010000010110", -- t[29718] = 14
      "001110" when "0111010000010111", -- t[29719] = 14
      "001110" when "0111010000011000", -- t[29720] = 14
      "001110" when "0111010000011001", -- t[29721] = 14
      "001110" when "0111010000011010", -- t[29722] = 14
      "001110" when "0111010000011011", -- t[29723] = 14
      "001110" when "0111010000011100", -- t[29724] = 14
      "001110" when "0111010000011101", -- t[29725] = 14
      "001110" when "0111010000011110", -- t[29726] = 14
      "001110" when "0111010000011111", -- t[29727] = 14
      "001110" when "0111010000100000", -- t[29728] = 14
      "001110" when "0111010000100001", -- t[29729] = 14
      "001110" when "0111010000100010", -- t[29730] = 14
      "001110" when "0111010000100011", -- t[29731] = 14
      "001110" when "0111010000100100", -- t[29732] = 14
      "001110" when "0111010000100101", -- t[29733] = 14
      "001110" when "0111010000100110", -- t[29734] = 14
      "001110" when "0111010000100111", -- t[29735] = 14
      "001110" when "0111010000101000", -- t[29736] = 14
      "001110" when "0111010000101001", -- t[29737] = 14
      "001110" when "0111010000101010", -- t[29738] = 14
      "001110" when "0111010000101011", -- t[29739] = 14
      "001110" when "0111010000101100", -- t[29740] = 14
      "001110" when "0111010000101101", -- t[29741] = 14
      "001110" when "0111010000101110", -- t[29742] = 14
      "001110" when "0111010000101111", -- t[29743] = 14
      "001110" when "0111010000110000", -- t[29744] = 14
      "001110" when "0111010000110001", -- t[29745] = 14
      "001110" when "0111010000110010", -- t[29746] = 14
      "001110" when "0111010000110011", -- t[29747] = 14
      "001110" when "0111010000110100", -- t[29748] = 14
      "001110" when "0111010000110101", -- t[29749] = 14
      "001110" when "0111010000110110", -- t[29750] = 14
      "001110" when "0111010000110111", -- t[29751] = 14
      "001110" when "0111010000111000", -- t[29752] = 14
      "001110" when "0111010000111001", -- t[29753] = 14
      "001110" when "0111010000111010", -- t[29754] = 14
      "001110" when "0111010000111011", -- t[29755] = 14
      "001110" when "0111010000111100", -- t[29756] = 14
      "001110" when "0111010000111101", -- t[29757] = 14
      "001110" when "0111010000111110", -- t[29758] = 14
      "001110" when "0111010000111111", -- t[29759] = 14
      "001110" when "0111010001000000", -- t[29760] = 14
      "001110" when "0111010001000001", -- t[29761] = 14
      "001110" when "0111010001000010", -- t[29762] = 14
      "001110" when "0111010001000011", -- t[29763] = 14
      "001110" when "0111010001000100", -- t[29764] = 14
      "001110" when "0111010001000101", -- t[29765] = 14
      "001110" when "0111010001000110", -- t[29766] = 14
      "001110" when "0111010001000111", -- t[29767] = 14
      "001110" when "0111010001001000", -- t[29768] = 14
      "001110" when "0111010001001001", -- t[29769] = 14
      "001110" when "0111010001001010", -- t[29770] = 14
      "001110" when "0111010001001011", -- t[29771] = 14
      "001110" when "0111010001001100", -- t[29772] = 14
      "001110" when "0111010001001101", -- t[29773] = 14
      "001110" when "0111010001001110", -- t[29774] = 14
      "001110" when "0111010001001111", -- t[29775] = 14
      "001110" when "0111010001010000", -- t[29776] = 14
      "001110" when "0111010001010001", -- t[29777] = 14
      "001110" when "0111010001010010", -- t[29778] = 14
      "001110" when "0111010001010011", -- t[29779] = 14
      "001110" when "0111010001010100", -- t[29780] = 14
      "001110" when "0111010001010101", -- t[29781] = 14
      "001110" when "0111010001010110", -- t[29782] = 14
      "001110" when "0111010001010111", -- t[29783] = 14
      "001110" when "0111010001011000", -- t[29784] = 14
      "001110" when "0111010001011001", -- t[29785] = 14
      "001110" when "0111010001011010", -- t[29786] = 14
      "001110" when "0111010001011011", -- t[29787] = 14
      "001110" when "0111010001011100", -- t[29788] = 14
      "001110" when "0111010001011101", -- t[29789] = 14
      "001110" when "0111010001011110", -- t[29790] = 14
      "001110" when "0111010001011111", -- t[29791] = 14
      "001110" when "0111010001100000", -- t[29792] = 14
      "001110" when "0111010001100001", -- t[29793] = 14
      "001110" when "0111010001100010", -- t[29794] = 14
      "001110" when "0111010001100011", -- t[29795] = 14
      "001110" when "0111010001100100", -- t[29796] = 14
      "001110" when "0111010001100101", -- t[29797] = 14
      "001110" when "0111010001100110", -- t[29798] = 14
      "001110" when "0111010001100111", -- t[29799] = 14
      "001110" when "0111010001101000", -- t[29800] = 14
      "001110" when "0111010001101001", -- t[29801] = 14
      "001110" when "0111010001101010", -- t[29802] = 14
      "001110" when "0111010001101011", -- t[29803] = 14
      "001110" when "0111010001101100", -- t[29804] = 14
      "001110" when "0111010001101101", -- t[29805] = 14
      "001110" when "0111010001101110", -- t[29806] = 14
      "001110" when "0111010001101111", -- t[29807] = 14
      "001110" when "0111010001110000", -- t[29808] = 14
      "001110" when "0111010001110001", -- t[29809] = 14
      "001110" when "0111010001110010", -- t[29810] = 14
      "001110" when "0111010001110011", -- t[29811] = 14
      "001110" when "0111010001110100", -- t[29812] = 14
      "001110" when "0111010001110101", -- t[29813] = 14
      "001110" when "0111010001110110", -- t[29814] = 14
      "001110" when "0111010001110111", -- t[29815] = 14
      "001110" when "0111010001111000", -- t[29816] = 14
      "001110" when "0111010001111001", -- t[29817] = 14
      "001110" when "0111010001111010", -- t[29818] = 14
      "001110" when "0111010001111011", -- t[29819] = 14
      "001110" when "0111010001111100", -- t[29820] = 14
      "001110" when "0111010001111101", -- t[29821] = 14
      "001110" when "0111010001111110", -- t[29822] = 14
      "001110" when "0111010001111111", -- t[29823] = 14
      "001110" when "0111010010000000", -- t[29824] = 14
      "001110" when "0111010010000001", -- t[29825] = 14
      "001110" when "0111010010000010", -- t[29826] = 14
      "001110" when "0111010010000011", -- t[29827] = 14
      "001110" when "0111010010000100", -- t[29828] = 14
      "001110" when "0111010010000101", -- t[29829] = 14
      "001110" when "0111010010000110", -- t[29830] = 14
      "001110" when "0111010010000111", -- t[29831] = 14
      "001110" when "0111010010001000", -- t[29832] = 14
      "001110" when "0111010010001001", -- t[29833] = 14
      "001110" when "0111010010001010", -- t[29834] = 14
      "001110" when "0111010010001011", -- t[29835] = 14
      "001110" when "0111010010001100", -- t[29836] = 14
      "001110" when "0111010010001101", -- t[29837] = 14
      "001110" when "0111010010001110", -- t[29838] = 14
      "001110" when "0111010010001111", -- t[29839] = 14
      "001110" when "0111010010010000", -- t[29840] = 14
      "001110" when "0111010010010001", -- t[29841] = 14
      "001110" when "0111010010010010", -- t[29842] = 14
      "001110" when "0111010010010011", -- t[29843] = 14
      "001110" when "0111010010010100", -- t[29844] = 14
      "001110" when "0111010010010101", -- t[29845] = 14
      "001110" when "0111010010010110", -- t[29846] = 14
      "001110" when "0111010010010111", -- t[29847] = 14
      "001110" when "0111010010011000", -- t[29848] = 14
      "001110" when "0111010010011001", -- t[29849] = 14
      "001110" when "0111010010011010", -- t[29850] = 14
      "001110" when "0111010010011011", -- t[29851] = 14
      "001110" when "0111010010011100", -- t[29852] = 14
      "001110" when "0111010010011101", -- t[29853] = 14
      "001110" when "0111010010011110", -- t[29854] = 14
      "001110" when "0111010010011111", -- t[29855] = 14
      "001110" when "0111010010100000", -- t[29856] = 14
      "001110" when "0111010010100001", -- t[29857] = 14
      "001110" when "0111010010100010", -- t[29858] = 14
      "001110" when "0111010010100011", -- t[29859] = 14
      "001110" when "0111010010100100", -- t[29860] = 14
      "001110" when "0111010010100101", -- t[29861] = 14
      "001110" when "0111010010100110", -- t[29862] = 14
      "001110" when "0111010010100111", -- t[29863] = 14
      "001110" when "0111010010101000", -- t[29864] = 14
      "001110" when "0111010010101001", -- t[29865] = 14
      "001110" when "0111010010101010", -- t[29866] = 14
      "001110" when "0111010010101011", -- t[29867] = 14
      "001110" when "0111010010101100", -- t[29868] = 14
      "001110" when "0111010010101101", -- t[29869] = 14
      "001110" when "0111010010101110", -- t[29870] = 14
      "001110" when "0111010010101111", -- t[29871] = 14
      "001110" when "0111010010110000", -- t[29872] = 14
      "001110" when "0111010010110001", -- t[29873] = 14
      "001110" when "0111010010110010", -- t[29874] = 14
      "001110" when "0111010010110011", -- t[29875] = 14
      "001110" when "0111010010110100", -- t[29876] = 14
      "001110" when "0111010010110101", -- t[29877] = 14
      "001110" when "0111010010110110", -- t[29878] = 14
      "001110" when "0111010010110111", -- t[29879] = 14
      "001110" when "0111010010111000", -- t[29880] = 14
      "001110" when "0111010010111001", -- t[29881] = 14
      "001110" when "0111010010111010", -- t[29882] = 14
      "001110" when "0111010010111011", -- t[29883] = 14
      "001110" when "0111010010111100", -- t[29884] = 14
      "001110" when "0111010010111101", -- t[29885] = 14
      "001110" when "0111010010111110", -- t[29886] = 14
      "001110" when "0111010010111111", -- t[29887] = 14
      "001110" when "0111010011000000", -- t[29888] = 14
      "001110" when "0111010011000001", -- t[29889] = 14
      "001110" when "0111010011000010", -- t[29890] = 14
      "001110" when "0111010011000011", -- t[29891] = 14
      "001110" when "0111010011000100", -- t[29892] = 14
      "001110" when "0111010011000101", -- t[29893] = 14
      "001110" when "0111010011000110", -- t[29894] = 14
      "001110" when "0111010011000111", -- t[29895] = 14
      "001110" when "0111010011001000", -- t[29896] = 14
      "001110" when "0111010011001001", -- t[29897] = 14
      "001110" when "0111010011001010", -- t[29898] = 14
      "001110" when "0111010011001011", -- t[29899] = 14
      "001110" when "0111010011001100", -- t[29900] = 14
      "001110" when "0111010011001101", -- t[29901] = 14
      "001110" when "0111010011001110", -- t[29902] = 14
      "001110" when "0111010011001111", -- t[29903] = 14
      "001110" when "0111010011010000", -- t[29904] = 14
      "001110" when "0111010011010001", -- t[29905] = 14
      "001110" when "0111010011010010", -- t[29906] = 14
      "001110" when "0111010011010011", -- t[29907] = 14
      "001110" when "0111010011010100", -- t[29908] = 14
      "001110" when "0111010011010101", -- t[29909] = 14
      "001110" when "0111010011010110", -- t[29910] = 14
      "001110" when "0111010011010111", -- t[29911] = 14
      "001110" when "0111010011011000", -- t[29912] = 14
      "001110" when "0111010011011001", -- t[29913] = 14
      "001110" when "0111010011011010", -- t[29914] = 14
      "001110" when "0111010011011011", -- t[29915] = 14
      "001110" when "0111010011011100", -- t[29916] = 14
      "001110" when "0111010011011101", -- t[29917] = 14
      "001110" when "0111010011011110", -- t[29918] = 14
      "001110" when "0111010011011111", -- t[29919] = 14
      "001110" when "0111010011100000", -- t[29920] = 14
      "001110" when "0111010011100001", -- t[29921] = 14
      "001110" when "0111010011100010", -- t[29922] = 14
      "001110" when "0111010011100011", -- t[29923] = 14
      "001110" when "0111010011100100", -- t[29924] = 14
      "001110" when "0111010011100101", -- t[29925] = 14
      "001110" when "0111010011100110", -- t[29926] = 14
      "001110" when "0111010011100111", -- t[29927] = 14
      "001110" when "0111010011101000", -- t[29928] = 14
      "001110" when "0111010011101001", -- t[29929] = 14
      "001110" when "0111010011101010", -- t[29930] = 14
      "001110" when "0111010011101011", -- t[29931] = 14
      "001110" when "0111010011101100", -- t[29932] = 14
      "001110" when "0111010011101101", -- t[29933] = 14
      "001110" when "0111010011101110", -- t[29934] = 14
      "001110" when "0111010011101111", -- t[29935] = 14
      "001110" when "0111010011110000", -- t[29936] = 14
      "001110" when "0111010011110001", -- t[29937] = 14
      "001110" when "0111010011110010", -- t[29938] = 14
      "001110" when "0111010011110011", -- t[29939] = 14
      "001110" when "0111010011110100", -- t[29940] = 14
      "001110" when "0111010011110101", -- t[29941] = 14
      "001110" when "0111010011110110", -- t[29942] = 14
      "001110" when "0111010011110111", -- t[29943] = 14
      "001110" when "0111010011111000", -- t[29944] = 14
      "001110" when "0111010011111001", -- t[29945] = 14
      "001110" when "0111010011111010", -- t[29946] = 14
      "001110" when "0111010011111011", -- t[29947] = 14
      "001110" when "0111010011111100", -- t[29948] = 14
      "001110" when "0111010011111101", -- t[29949] = 14
      "001110" when "0111010011111110", -- t[29950] = 14
      "001110" when "0111010011111111", -- t[29951] = 14
      "001110" when "0111010100000000", -- t[29952] = 14
      "001110" when "0111010100000001", -- t[29953] = 14
      "001110" when "0111010100000010", -- t[29954] = 14
      "001110" when "0111010100000011", -- t[29955] = 14
      "001110" when "0111010100000100", -- t[29956] = 14
      "001110" when "0111010100000101", -- t[29957] = 14
      "001110" when "0111010100000110", -- t[29958] = 14
      "001110" when "0111010100000111", -- t[29959] = 14
      "001110" when "0111010100001000", -- t[29960] = 14
      "001110" when "0111010100001001", -- t[29961] = 14
      "001110" when "0111010100001010", -- t[29962] = 14
      "001110" when "0111010100001011", -- t[29963] = 14
      "001110" when "0111010100001100", -- t[29964] = 14
      "001110" when "0111010100001101", -- t[29965] = 14
      "001110" when "0111010100001110", -- t[29966] = 14
      "001110" when "0111010100001111", -- t[29967] = 14
      "001110" when "0111010100010000", -- t[29968] = 14
      "001110" when "0111010100010001", -- t[29969] = 14
      "001110" when "0111010100010010", -- t[29970] = 14
      "001110" when "0111010100010011", -- t[29971] = 14
      "001110" when "0111010100010100", -- t[29972] = 14
      "001110" when "0111010100010101", -- t[29973] = 14
      "001110" when "0111010100010110", -- t[29974] = 14
      "001110" when "0111010100010111", -- t[29975] = 14
      "001110" when "0111010100011000", -- t[29976] = 14
      "001110" when "0111010100011001", -- t[29977] = 14
      "001110" when "0111010100011010", -- t[29978] = 14
      "001110" when "0111010100011011", -- t[29979] = 14
      "001110" when "0111010100011100", -- t[29980] = 14
      "001110" when "0111010100011101", -- t[29981] = 14
      "001110" when "0111010100011110", -- t[29982] = 14
      "001110" when "0111010100011111", -- t[29983] = 14
      "001110" when "0111010100100000", -- t[29984] = 14
      "001110" when "0111010100100001", -- t[29985] = 14
      "001110" when "0111010100100010", -- t[29986] = 14
      "001110" when "0111010100100011", -- t[29987] = 14
      "001110" when "0111010100100100", -- t[29988] = 14
      "001110" when "0111010100100101", -- t[29989] = 14
      "001110" when "0111010100100110", -- t[29990] = 14
      "001110" when "0111010100100111", -- t[29991] = 14
      "001110" when "0111010100101000", -- t[29992] = 14
      "001110" when "0111010100101001", -- t[29993] = 14
      "001110" when "0111010100101010", -- t[29994] = 14
      "001110" when "0111010100101011", -- t[29995] = 14
      "001110" when "0111010100101100", -- t[29996] = 14
      "001110" when "0111010100101101", -- t[29997] = 14
      "001110" when "0111010100101110", -- t[29998] = 14
      "001110" when "0111010100101111", -- t[29999] = 14
      "001110" when "0111010100110000", -- t[30000] = 14
      "001110" when "0111010100110001", -- t[30001] = 14
      "001110" when "0111010100110010", -- t[30002] = 14
      "001110" when "0111010100110011", -- t[30003] = 14
      "001110" when "0111010100110100", -- t[30004] = 14
      "001110" when "0111010100110101", -- t[30005] = 14
      "001110" when "0111010100110110", -- t[30006] = 14
      "001110" when "0111010100110111", -- t[30007] = 14
      "001110" when "0111010100111000", -- t[30008] = 14
      "001110" when "0111010100111001", -- t[30009] = 14
      "001110" when "0111010100111010", -- t[30010] = 14
      "001110" when "0111010100111011", -- t[30011] = 14
      "001110" when "0111010100111100", -- t[30012] = 14
      "001110" when "0111010100111101", -- t[30013] = 14
      "001111" when "0111010100111110", -- t[30014] = 15
      "001111" when "0111010100111111", -- t[30015] = 15
      "001111" when "0111010101000000", -- t[30016] = 15
      "001111" when "0111010101000001", -- t[30017] = 15
      "001111" when "0111010101000010", -- t[30018] = 15
      "001111" when "0111010101000011", -- t[30019] = 15
      "001111" when "0111010101000100", -- t[30020] = 15
      "001111" when "0111010101000101", -- t[30021] = 15
      "001111" when "0111010101000110", -- t[30022] = 15
      "001111" when "0111010101000111", -- t[30023] = 15
      "001111" when "0111010101001000", -- t[30024] = 15
      "001111" when "0111010101001001", -- t[30025] = 15
      "001111" when "0111010101001010", -- t[30026] = 15
      "001111" when "0111010101001011", -- t[30027] = 15
      "001111" when "0111010101001100", -- t[30028] = 15
      "001111" when "0111010101001101", -- t[30029] = 15
      "001111" when "0111010101001110", -- t[30030] = 15
      "001111" when "0111010101001111", -- t[30031] = 15
      "001111" when "0111010101010000", -- t[30032] = 15
      "001111" when "0111010101010001", -- t[30033] = 15
      "001111" when "0111010101010010", -- t[30034] = 15
      "001111" when "0111010101010011", -- t[30035] = 15
      "001111" when "0111010101010100", -- t[30036] = 15
      "001111" when "0111010101010101", -- t[30037] = 15
      "001111" when "0111010101010110", -- t[30038] = 15
      "001111" when "0111010101010111", -- t[30039] = 15
      "001111" when "0111010101011000", -- t[30040] = 15
      "001111" when "0111010101011001", -- t[30041] = 15
      "001111" when "0111010101011010", -- t[30042] = 15
      "001111" when "0111010101011011", -- t[30043] = 15
      "001111" when "0111010101011100", -- t[30044] = 15
      "001111" when "0111010101011101", -- t[30045] = 15
      "001111" when "0111010101011110", -- t[30046] = 15
      "001111" when "0111010101011111", -- t[30047] = 15
      "001111" when "0111010101100000", -- t[30048] = 15
      "001111" when "0111010101100001", -- t[30049] = 15
      "001111" when "0111010101100010", -- t[30050] = 15
      "001111" when "0111010101100011", -- t[30051] = 15
      "001111" when "0111010101100100", -- t[30052] = 15
      "001111" when "0111010101100101", -- t[30053] = 15
      "001111" when "0111010101100110", -- t[30054] = 15
      "001111" when "0111010101100111", -- t[30055] = 15
      "001111" when "0111010101101000", -- t[30056] = 15
      "001111" when "0111010101101001", -- t[30057] = 15
      "001111" when "0111010101101010", -- t[30058] = 15
      "001111" when "0111010101101011", -- t[30059] = 15
      "001111" when "0111010101101100", -- t[30060] = 15
      "001111" when "0111010101101101", -- t[30061] = 15
      "001111" when "0111010101101110", -- t[30062] = 15
      "001111" when "0111010101101111", -- t[30063] = 15
      "001111" when "0111010101110000", -- t[30064] = 15
      "001111" when "0111010101110001", -- t[30065] = 15
      "001111" when "0111010101110010", -- t[30066] = 15
      "001111" when "0111010101110011", -- t[30067] = 15
      "001111" when "0111010101110100", -- t[30068] = 15
      "001111" when "0111010101110101", -- t[30069] = 15
      "001111" when "0111010101110110", -- t[30070] = 15
      "001111" when "0111010101110111", -- t[30071] = 15
      "001111" when "0111010101111000", -- t[30072] = 15
      "001111" when "0111010101111001", -- t[30073] = 15
      "001111" when "0111010101111010", -- t[30074] = 15
      "001111" when "0111010101111011", -- t[30075] = 15
      "001111" when "0111010101111100", -- t[30076] = 15
      "001111" when "0111010101111101", -- t[30077] = 15
      "001111" when "0111010101111110", -- t[30078] = 15
      "001111" when "0111010101111111", -- t[30079] = 15
      "001111" when "0111010110000000", -- t[30080] = 15
      "001111" when "0111010110000001", -- t[30081] = 15
      "001111" when "0111010110000010", -- t[30082] = 15
      "001111" when "0111010110000011", -- t[30083] = 15
      "001111" when "0111010110000100", -- t[30084] = 15
      "001111" when "0111010110000101", -- t[30085] = 15
      "001111" when "0111010110000110", -- t[30086] = 15
      "001111" when "0111010110000111", -- t[30087] = 15
      "001111" when "0111010110001000", -- t[30088] = 15
      "001111" when "0111010110001001", -- t[30089] = 15
      "001111" when "0111010110001010", -- t[30090] = 15
      "001111" when "0111010110001011", -- t[30091] = 15
      "001111" when "0111010110001100", -- t[30092] = 15
      "001111" when "0111010110001101", -- t[30093] = 15
      "001111" when "0111010110001110", -- t[30094] = 15
      "001111" when "0111010110001111", -- t[30095] = 15
      "001111" when "0111010110010000", -- t[30096] = 15
      "001111" when "0111010110010001", -- t[30097] = 15
      "001111" when "0111010110010010", -- t[30098] = 15
      "001111" when "0111010110010011", -- t[30099] = 15
      "001111" when "0111010110010100", -- t[30100] = 15
      "001111" when "0111010110010101", -- t[30101] = 15
      "001111" when "0111010110010110", -- t[30102] = 15
      "001111" when "0111010110010111", -- t[30103] = 15
      "001111" when "0111010110011000", -- t[30104] = 15
      "001111" when "0111010110011001", -- t[30105] = 15
      "001111" when "0111010110011010", -- t[30106] = 15
      "001111" when "0111010110011011", -- t[30107] = 15
      "001111" when "0111010110011100", -- t[30108] = 15
      "001111" when "0111010110011101", -- t[30109] = 15
      "001111" when "0111010110011110", -- t[30110] = 15
      "001111" when "0111010110011111", -- t[30111] = 15
      "001111" when "0111010110100000", -- t[30112] = 15
      "001111" when "0111010110100001", -- t[30113] = 15
      "001111" when "0111010110100010", -- t[30114] = 15
      "001111" when "0111010110100011", -- t[30115] = 15
      "001111" when "0111010110100100", -- t[30116] = 15
      "001111" when "0111010110100101", -- t[30117] = 15
      "001111" when "0111010110100110", -- t[30118] = 15
      "001111" when "0111010110100111", -- t[30119] = 15
      "001111" when "0111010110101000", -- t[30120] = 15
      "001111" when "0111010110101001", -- t[30121] = 15
      "001111" when "0111010110101010", -- t[30122] = 15
      "001111" when "0111010110101011", -- t[30123] = 15
      "001111" when "0111010110101100", -- t[30124] = 15
      "001111" when "0111010110101101", -- t[30125] = 15
      "001111" when "0111010110101110", -- t[30126] = 15
      "001111" when "0111010110101111", -- t[30127] = 15
      "001111" when "0111010110110000", -- t[30128] = 15
      "001111" when "0111010110110001", -- t[30129] = 15
      "001111" when "0111010110110010", -- t[30130] = 15
      "001111" when "0111010110110011", -- t[30131] = 15
      "001111" when "0111010110110100", -- t[30132] = 15
      "001111" when "0111010110110101", -- t[30133] = 15
      "001111" when "0111010110110110", -- t[30134] = 15
      "001111" when "0111010110110111", -- t[30135] = 15
      "001111" when "0111010110111000", -- t[30136] = 15
      "001111" when "0111010110111001", -- t[30137] = 15
      "001111" when "0111010110111010", -- t[30138] = 15
      "001111" when "0111010110111011", -- t[30139] = 15
      "001111" when "0111010110111100", -- t[30140] = 15
      "001111" when "0111010110111101", -- t[30141] = 15
      "001111" when "0111010110111110", -- t[30142] = 15
      "001111" when "0111010110111111", -- t[30143] = 15
      "001111" when "0111010111000000", -- t[30144] = 15
      "001111" when "0111010111000001", -- t[30145] = 15
      "001111" when "0111010111000010", -- t[30146] = 15
      "001111" when "0111010111000011", -- t[30147] = 15
      "001111" when "0111010111000100", -- t[30148] = 15
      "001111" when "0111010111000101", -- t[30149] = 15
      "001111" when "0111010111000110", -- t[30150] = 15
      "001111" when "0111010111000111", -- t[30151] = 15
      "001111" when "0111010111001000", -- t[30152] = 15
      "001111" when "0111010111001001", -- t[30153] = 15
      "001111" when "0111010111001010", -- t[30154] = 15
      "001111" when "0111010111001011", -- t[30155] = 15
      "001111" when "0111010111001100", -- t[30156] = 15
      "001111" when "0111010111001101", -- t[30157] = 15
      "001111" when "0111010111001110", -- t[30158] = 15
      "001111" when "0111010111001111", -- t[30159] = 15
      "001111" when "0111010111010000", -- t[30160] = 15
      "001111" when "0111010111010001", -- t[30161] = 15
      "001111" when "0111010111010010", -- t[30162] = 15
      "001111" when "0111010111010011", -- t[30163] = 15
      "001111" when "0111010111010100", -- t[30164] = 15
      "001111" when "0111010111010101", -- t[30165] = 15
      "001111" when "0111010111010110", -- t[30166] = 15
      "001111" when "0111010111010111", -- t[30167] = 15
      "001111" when "0111010111011000", -- t[30168] = 15
      "001111" when "0111010111011001", -- t[30169] = 15
      "001111" when "0111010111011010", -- t[30170] = 15
      "001111" when "0111010111011011", -- t[30171] = 15
      "001111" when "0111010111011100", -- t[30172] = 15
      "001111" when "0111010111011101", -- t[30173] = 15
      "001111" when "0111010111011110", -- t[30174] = 15
      "001111" when "0111010111011111", -- t[30175] = 15
      "001111" when "0111010111100000", -- t[30176] = 15
      "001111" when "0111010111100001", -- t[30177] = 15
      "001111" when "0111010111100010", -- t[30178] = 15
      "001111" when "0111010111100011", -- t[30179] = 15
      "001111" when "0111010111100100", -- t[30180] = 15
      "001111" when "0111010111100101", -- t[30181] = 15
      "001111" when "0111010111100110", -- t[30182] = 15
      "001111" when "0111010111100111", -- t[30183] = 15
      "001111" when "0111010111101000", -- t[30184] = 15
      "001111" when "0111010111101001", -- t[30185] = 15
      "001111" when "0111010111101010", -- t[30186] = 15
      "001111" when "0111010111101011", -- t[30187] = 15
      "001111" when "0111010111101100", -- t[30188] = 15
      "001111" when "0111010111101101", -- t[30189] = 15
      "001111" when "0111010111101110", -- t[30190] = 15
      "001111" when "0111010111101111", -- t[30191] = 15
      "001111" when "0111010111110000", -- t[30192] = 15
      "001111" when "0111010111110001", -- t[30193] = 15
      "001111" when "0111010111110010", -- t[30194] = 15
      "001111" when "0111010111110011", -- t[30195] = 15
      "001111" when "0111010111110100", -- t[30196] = 15
      "001111" when "0111010111110101", -- t[30197] = 15
      "001111" when "0111010111110110", -- t[30198] = 15
      "001111" when "0111010111110111", -- t[30199] = 15
      "001111" when "0111010111111000", -- t[30200] = 15
      "001111" when "0111010111111001", -- t[30201] = 15
      "001111" when "0111010111111010", -- t[30202] = 15
      "001111" when "0111010111111011", -- t[30203] = 15
      "001111" when "0111010111111100", -- t[30204] = 15
      "001111" when "0111010111111101", -- t[30205] = 15
      "001111" when "0111010111111110", -- t[30206] = 15
      "001111" when "0111010111111111", -- t[30207] = 15
      "001111" when "0111011000000000", -- t[30208] = 15
      "001111" when "0111011000000001", -- t[30209] = 15
      "001111" when "0111011000000010", -- t[30210] = 15
      "001111" when "0111011000000011", -- t[30211] = 15
      "001111" when "0111011000000100", -- t[30212] = 15
      "001111" when "0111011000000101", -- t[30213] = 15
      "001111" when "0111011000000110", -- t[30214] = 15
      "001111" when "0111011000000111", -- t[30215] = 15
      "001111" when "0111011000001000", -- t[30216] = 15
      "001111" when "0111011000001001", -- t[30217] = 15
      "001111" when "0111011000001010", -- t[30218] = 15
      "001111" when "0111011000001011", -- t[30219] = 15
      "001111" when "0111011000001100", -- t[30220] = 15
      "001111" when "0111011000001101", -- t[30221] = 15
      "001111" when "0111011000001110", -- t[30222] = 15
      "001111" when "0111011000001111", -- t[30223] = 15
      "001111" when "0111011000010000", -- t[30224] = 15
      "001111" when "0111011000010001", -- t[30225] = 15
      "001111" when "0111011000010010", -- t[30226] = 15
      "001111" when "0111011000010011", -- t[30227] = 15
      "001111" when "0111011000010100", -- t[30228] = 15
      "001111" when "0111011000010101", -- t[30229] = 15
      "001111" when "0111011000010110", -- t[30230] = 15
      "001111" when "0111011000010111", -- t[30231] = 15
      "001111" when "0111011000011000", -- t[30232] = 15
      "001111" when "0111011000011001", -- t[30233] = 15
      "001111" when "0111011000011010", -- t[30234] = 15
      "001111" when "0111011000011011", -- t[30235] = 15
      "001111" when "0111011000011100", -- t[30236] = 15
      "001111" when "0111011000011101", -- t[30237] = 15
      "001111" when "0111011000011110", -- t[30238] = 15
      "001111" when "0111011000011111", -- t[30239] = 15
      "001111" when "0111011000100000", -- t[30240] = 15
      "001111" when "0111011000100001", -- t[30241] = 15
      "001111" when "0111011000100010", -- t[30242] = 15
      "001111" when "0111011000100011", -- t[30243] = 15
      "001111" when "0111011000100100", -- t[30244] = 15
      "001111" when "0111011000100101", -- t[30245] = 15
      "001111" when "0111011000100110", -- t[30246] = 15
      "001111" when "0111011000100111", -- t[30247] = 15
      "001111" when "0111011000101000", -- t[30248] = 15
      "001111" when "0111011000101001", -- t[30249] = 15
      "001111" when "0111011000101010", -- t[30250] = 15
      "001111" when "0111011000101011", -- t[30251] = 15
      "001111" when "0111011000101100", -- t[30252] = 15
      "001111" when "0111011000101101", -- t[30253] = 15
      "001111" when "0111011000101110", -- t[30254] = 15
      "001111" when "0111011000101111", -- t[30255] = 15
      "001111" when "0111011000110000", -- t[30256] = 15
      "001111" when "0111011000110001", -- t[30257] = 15
      "001111" when "0111011000110010", -- t[30258] = 15
      "001111" when "0111011000110011", -- t[30259] = 15
      "001111" when "0111011000110100", -- t[30260] = 15
      "001111" when "0111011000110101", -- t[30261] = 15
      "001111" when "0111011000110110", -- t[30262] = 15
      "001111" when "0111011000110111", -- t[30263] = 15
      "001111" when "0111011000111000", -- t[30264] = 15
      "001111" when "0111011000111001", -- t[30265] = 15
      "001111" when "0111011000111010", -- t[30266] = 15
      "001111" when "0111011000111011", -- t[30267] = 15
      "001111" when "0111011000111100", -- t[30268] = 15
      "001111" when "0111011000111101", -- t[30269] = 15
      "001111" when "0111011000111110", -- t[30270] = 15
      "001111" when "0111011000111111", -- t[30271] = 15
      "001111" when "0111011001000000", -- t[30272] = 15
      "001111" when "0111011001000001", -- t[30273] = 15
      "001111" when "0111011001000010", -- t[30274] = 15
      "001111" when "0111011001000011", -- t[30275] = 15
      "001111" when "0111011001000100", -- t[30276] = 15
      "001111" when "0111011001000101", -- t[30277] = 15
      "001111" when "0111011001000110", -- t[30278] = 15
      "001111" when "0111011001000111", -- t[30279] = 15
      "001111" when "0111011001001000", -- t[30280] = 15
      "001111" when "0111011001001001", -- t[30281] = 15
      "001111" when "0111011001001010", -- t[30282] = 15
      "001111" when "0111011001001011", -- t[30283] = 15
      "001111" when "0111011001001100", -- t[30284] = 15
      "001111" when "0111011001001101", -- t[30285] = 15
      "001111" when "0111011001001110", -- t[30286] = 15
      "001111" when "0111011001001111", -- t[30287] = 15
      "001111" when "0111011001010000", -- t[30288] = 15
      "001111" when "0111011001010001", -- t[30289] = 15
      "001111" when "0111011001010010", -- t[30290] = 15
      "001111" when "0111011001010011", -- t[30291] = 15
      "001111" when "0111011001010100", -- t[30292] = 15
      "001111" when "0111011001010101", -- t[30293] = 15
      "001111" when "0111011001010110", -- t[30294] = 15
      "001111" when "0111011001010111", -- t[30295] = 15
      "001111" when "0111011001011000", -- t[30296] = 15
      "001111" when "0111011001011001", -- t[30297] = 15
      "001111" when "0111011001011010", -- t[30298] = 15
      "001111" when "0111011001011011", -- t[30299] = 15
      "001111" when "0111011001011100", -- t[30300] = 15
      "001111" when "0111011001011101", -- t[30301] = 15
      "001111" when "0111011001011110", -- t[30302] = 15
      "001111" when "0111011001011111", -- t[30303] = 15
      "001111" when "0111011001100000", -- t[30304] = 15
      "001111" when "0111011001100001", -- t[30305] = 15
      "001111" when "0111011001100010", -- t[30306] = 15
      "001111" when "0111011001100011", -- t[30307] = 15
      "001111" when "0111011001100100", -- t[30308] = 15
      "001111" when "0111011001100101", -- t[30309] = 15
      "001111" when "0111011001100110", -- t[30310] = 15
      "001111" when "0111011001100111", -- t[30311] = 15
      "001111" when "0111011001101000", -- t[30312] = 15
      "001111" when "0111011001101001", -- t[30313] = 15
      "001111" when "0111011001101010", -- t[30314] = 15
      "001111" when "0111011001101011", -- t[30315] = 15
      "001111" when "0111011001101100", -- t[30316] = 15
      "001111" when "0111011001101101", -- t[30317] = 15
      "001111" when "0111011001101110", -- t[30318] = 15
      "001111" when "0111011001101111", -- t[30319] = 15
      "001111" when "0111011001110000", -- t[30320] = 15
      "001111" when "0111011001110001", -- t[30321] = 15
      "001111" when "0111011001110010", -- t[30322] = 15
      "001111" when "0111011001110011", -- t[30323] = 15
      "001111" when "0111011001110100", -- t[30324] = 15
      "001111" when "0111011001110101", -- t[30325] = 15
      "001111" when "0111011001110110", -- t[30326] = 15
      "001111" when "0111011001110111", -- t[30327] = 15
      "001111" when "0111011001111000", -- t[30328] = 15
      "001111" when "0111011001111001", -- t[30329] = 15
      "001111" when "0111011001111010", -- t[30330] = 15
      "001111" when "0111011001111011", -- t[30331] = 15
      "001111" when "0111011001111100", -- t[30332] = 15
      "001111" when "0111011001111101", -- t[30333] = 15
      "001111" when "0111011001111110", -- t[30334] = 15
      "001111" when "0111011001111111", -- t[30335] = 15
      "001111" when "0111011010000000", -- t[30336] = 15
      "001111" when "0111011010000001", -- t[30337] = 15
      "001111" when "0111011010000010", -- t[30338] = 15
      "001111" when "0111011010000011", -- t[30339] = 15
      "001111" when "0111011010000100", -- t[30340] = 15
      "001111" when "0111011010000101", -- t[30341] = 15
      "001111" when "0111011010000110", -- t[30342] = 15
      "001111" when "0111011010000111", -- t[30343] = 15
      "001111" when "0111011010001000", -- t[30344] = 15
      "001111" when "0111011010001001", -- t[30345] = 15
      "001111" when "0111011010001010", -- t[30346] = 15
      "001111" when "0111011010001011", -- t[30347] = 15
      "001111" when "0111011010001100", -- t[30348] = 15
      "001111" when "0111011010001101", -- t[30349] = 15
      "001111" when "0111011010001110", -- t[30350] = 15
      "001111" when "0111011010001111", -- t[30351] = 15
      "001111" when "0111011010010000", -- t[30352] = 15
      "001111" when "0111011010010001", -- t[30353] = 15
      "001111" when "0111011010010010", -- t[30354] = 15
      "001111" when "0111011010010011", -- t[30355] = 15
      "001111" when "0111011010010100", -- t[30356] = 15
      "001111" when "0111011010010101", -- t[30357] = 15
      "001111" when "0111011010010110", -- t[30358] = 15
      "001111" when "0111011010010111", -- t[30359] = 15
      "001111" when "0111011010011000", -- t[30360] = 15
      "001111" when "0111011010011001", -- t[30361] = 15
      "001111" when "0111011010011010", -- t[30362] = 15
      "001111" when "0111011010011011", -- t[30363] = 15
      "001111" when "0111011010011100", -- t[30364] = 15
      "001111" when "0111011010011101", -- t[30365] = 15
      "001111" when "0111011010011110", -- t[30366] = 15
      "001111" when "0111011010011111", -- t[30367] = 15
      "001111" when "0111011010100000", -- t[30368] = 15
      "001111" when "0111011010100001", -- t[30369] = 15
      "001111" when "0111011010100010", -- t[30370] = 15
      "001111" when "0111011010100011", -- t[30371] = 15
      "001111" when "0111011010100100", -- t[30372] = 15
      "001111" when "0111011010100101", -- t[30373] = 15
      "001111" when "0111011010100110", -- t[30374] = 15
      "001111" when "0111011010100111", -- t[30375] = 15
      "001111" when "0111011010101000", -- t[30376] = 15
      "001111" when "0111011010101001", -- t[30377] = 15
      "001111" when "0111011010101010", -- t[30378] = 15
      "001111" when "0111011010101011", -- t[30379] = 15
      "001111" when "0111011010101100", -- t[30380] = 15
      "001111" when "0111011010101101", -- t[30381] = 15
      "001111" when "0111011010101110", -- t[30382] = 15
      "001111" when "0111011010101111", -- t[30383] = 15
      "001111" when "0111011010110000", -- t[30384] = 15
      "001111" when "0111011010110001", -- t[30385] = 15
      "001111" when "0111011010110010", -- t[30386] = 15
      "001111" when "0111011010110011", -- t[30387] = 15
      "001111" when "0111011010110100", -- t[30388] = 15
      "001111" when "0111011010110101", -- t[30389] = 15
      "001111" when "0111011010110110", -- t[30390] = 15
      "001111" when "0111011010110111", -- t[30391] = 15
      "001111" when "0111011010111000", -- t[30392] = 15
      "001111" when "0111011010111001", -- t[30393] = 15
      "001111" when "0111011010111010", -- t[30394] = 15
      "001111" when "0111011010111011", -- t[30395] = 15
      "001111" when "0111011010111100", -- t[30396] = 15
      "001111" when "0111011010111101", -- t[30397] = 15
      "001111" when "0111011010111110", -- t[30398] = 15
      "001111" when "0111011010111111", -- t[30399] = 15
      "001111" when "0111011011000000", -- t[30400] = 15
      "001111" when "0111011011000001", -- t[30401] = 15
      "001111" when "0111011011000010", -- t[30402] = 15
      "001111" when "0111011011000011", -- t[30403] = 15
      "001111" when "0111011011000100", -- t[30404] = 15
      "001111" when "0111011011000101", -- t[30405] = 15
      "001111" when "0111011011000110", -- t[30406] = 15
      "010000" when "0111011011000111", -- t[30407] = 16
      "010000" when "0111011011001000", -- t[30408] = 16
      "010000" when "0111011011001001", -- t[30409] = 16
      "010000" when "0111011011001010", -- t[30410] = 16
      "010000" when "0111011011001011", -- t[30411] = 16
      "010000" when "0111011011001100", -- t[30412] = 16
      "010000" when "0111011011001101", -- t[30413] = 16
      "010000" when "0111011011001110", -- t[30414] = 16
      "010000" when "0111011011001111", -- t[30415] = 16
      "010000" when "0111011011010000", -- t[30416] = 16
      "010000" when "0111011011010001", -- t[30417] = 16
      "010000" when "0111011011010010", -- t[30418] = 16
      "010000" when "0111011011010011", -- t[30419] = 16
      "010000" when "0111011011010100", -- t[30420] = 16
      "010000" when "0111011011010101", -- t[30421] = 16
      "010000" when "0111011011010110", -- t[30422] = 16
      "010000" when "0111011011010111", -- t[30423] = 16
      "010000" when "0111011011011000", -- t[30424] = 16
      "010000" when "0111011011011001", -- t[30425] = 16
      "010000" when "0111011011011010", -- t[30426] = 16
      "010000" when "0111011011011011", -- t[30427] = 16
      "010000" when "0111011011011100", -- t[30428] = 16
      "010000" when "0111011011011101", -- t[30429] = 16
      "010000" when "0111011011011110", -- t[30430] = 16
      "010000" when "0111011011011111", -- t[30431] = 16
      "010000" when "0111011011100000", -- t[30432] = 16
      "010000" when "0111011011100001", -- t[30433] = 16
      "010000" when "0111011011100010", -- t[30434] = 16
      "010000" when "0111011011100011", -- t[30435] = 16
      "010000" when "0111011011100100", -- t[30436] = 16
      "010000" when "0111011011100101", -- t[30437] = 16
      "010000" when "0111011011100110", -- t[30438] = 16
      "010000" when "0111011011100111", -- t[30439] = 16
      "010000" when "0111011011101000", -- t[30440] = 16
      "010000" when "0111011011101001", -- t[30441] = 16
      "010000" when "0111011011101010", -- t[30442] = 16
      "010000" when "0111011011101011", -- t[30443] = 16
      "010000" when "0111011011101100", -- t[30444] = 16
      "010000" when "0111011011101101", -- t[30445] = 16
      "010000" when "0111011011101110", -- t[30446] = 16
      "010000" when "0111011011101111", -- t[30447] = 16
      "010000" when "0111011011110000", -- t[30448] = 16
      "010000" when "0111011011110001", -- t[30449] = 16
      "010000" when "0111011011110010", -- t[30450] = 16
      "010000" when "0111011011110011", -- t[30451] = 16
      "010000" when "0111011011110100", -- t[30452] = 16
      "010000" when "0111011011110101", -- t[30453] = 16
      "010000" when "0111011011110110", -- t[30454] = 16
      "010000" when "0111011011110111", -- t[30455] = 16
      "010000" when "0111011011111000", -- t[30456] = 16
      "010000" when "0111011011111001", -- t[30457] = 16
      "010000" when "0111011011111010", -- t[30458] = 16
      "010000" when "0111011011111011", -- t[30459] = 16
      "010000" when "0111011011111100", -- t[30460] = 16
      "010000" when "0111011011111101", -- t[30461] = 16
      "010000" when "0111011011111110", -- t[30462] = 16
      "010000" when "0111011011111111", -- t[30463] = 16
      "010000" when "0111011100000000", -- t[30464] = 16
      "010000" when "0111011100000001", -- t[30465] = 16
      "010000" when "0111011100000010", -- t[30466] = 16
      "010000" when "0111011100000011", -- t[30467] = 16
      "010000" when "0111011100000100", -- t[30468] = 16
      "010000" when "0111011100000101", -- t[30469] = 16
      "010000" when "0111011100000110", -- t[30470] = 16
      "010000" when "0111011100000111", -- t[30471] = 16
      "010000" when "0111011100001000", -- t[30472] = 16
      "010000" when "0111011100001001", -- t[30473] = 16
      "010000" when "0111011100001010", -- t[30474] = 16
      "010000" when "0111011100001011", -- t[30475] = 16
      "010000" when "0111011100001100", -- t[30476] = 16
      "010000" when "0111011100001101", -- t[30477] = 16
      "010000" when "0111011100001110", -- t[30478] = 16
      "010000" when "0111011100001111", -- t[30479] = 16
      "010000" when "0111011100010000", -- t[30480] = 16
      "010000" when "0111011100010001", -- t[30481] = 16
      "010000" when "0111011100010010", -- t[30482] = 16
      "010000" when "0111011100010011", -- t[30483] = 16
      "010000" when "0111011100010100", -- t[30484] = 16
      "010000" when "0111011100010101", -- t[30485] = 16
      "010000" when "0111011100010110", -- t[30486] = 16
      "010000" when "0111011100010111", -- t[30487] = 16
      "010000" when "0111011100011000", -- t[30488] = 16
      "010000" when "0111011100011001", -- t[30489] = 16
      "010000" when "0111011100011010", -- t[30490] = 16
      "010000" when "0111011100011011", -- t[30491] = 16
      "010000" when "0111011100011100", -- t[30492] = 16
      "010000" when "0111011100011101", -- t[30493] = 16
      "010000" when "0111011100011110", -- t[30494] = 16
      "010000" when "0111011100011111", -- t[30495] = 16
      "010000" when "0111011100100000", -- t[30496] = 16
      "010000" when "0111011100100001", -- t[30497] = 16
      "010000" when "0111011100100010", -- t[30498] = 16
      "010000" when "0111011100100011", -- t[30499] = 16
      "010000" when "0111011100100100", -- t[30500] = 16
      "010000" when "0111011100100101", -- t[30501] = 16
      "010000" when "0111011100100110", -- t[30502] = 16
      "010000" when "0111011100100111", -- t[30503] = 16
      "010000" when "0111011100101000", -- t[30504] = 16
      "010000" when "0111011100101001", -- t[30505] = 16
      "010000" when "0111011100101010", -- t[30506] = 16
      "010000" when "0111011100101011", -- t[30507] = 16
      "010000" when "0111011100101100", -- t[30508] = 16
      "010000" when "0111011100101101", -- t[30509] = 16
      "010000" when "0111011100101110", -- t[30510] = 16
      "010000" when "0111011100101111", -- t[30511] = 16
      "010000" when "0111011100110000", -- t[30512] = 16
      "010000" when "0111011100110001", -- t[30513] = 16
      "010000" when "0111011100110010", -- t[30514] = 16
      "010000" when "0111011100110011", -- t[30515] = 16
      "010000" when "0111011100110100", -- t[30516] = 16
      "010000" when "0111011100110101", -- t[30517] = 16
      "010000" when "0111011100110110", -- t[30518] = 16
      "010000" when "0111011100110111", -- t[30519] = 16
      "010000" when "0111011100111000", -- t[30520] = 16
      "010000" when "0111011100111001", -- t[30521] = 16
      "010000" when "0111011100111010", -- t[30522] = 16
      "010000" when "0111011100111011", -- t[30523] = 16
      "010000" when "0111011100111100", -- t[30524] = 16
      "010000" when "0111011100111101", -- t[30525] = 16
      "010000" when "0111011100111110", -- t[30526] = 16
      "010000" when "0111011100111111", -- t[30527] = 16
      "010000" when "0111011101000000", -- t[30528] = 16
      "010000" when "0111011101000001", -- t[30529] = 16
      "010000" when "0111011101000010", -- t[30530] = 16
      "010000" when "0111011101000011", -- t[30531] = 16
      "010000" when "0111011101000100", -- t[30532] = 16
      "010000" when "0111011101000101", -- t[30533] = 16
      "010000" when "0111011101000110", -- t[30534] = 16
      "010000" when "0111011101000111", -- t[30535] = 16
      "010000" when "0111011101001000", -- t[30536] = 16
      "010000" when "0111011101001001", -- t[30537] = 16
      "010000" when "0111011101001010", -- t[30538] = 16
      "010000" when "0111011101001011", -- t[30539] = 16
      "010000" when "0111011101001100", -- t[30540] = 16
      "010000" when "0111011101001101", -- t[30541] = 16
      "010000" when "0111011101001110", -- t[30542] = 16
      "010000" when "0111011101001111", -- t[30543] = 16
      "010000" when "0111011101010000", -- t[30544] = 16
      "010000" when "0111011101010001", -- t[30545] = 16
      "010000" when "0111011101010010", -- t[30546] = 16
      "010000" when "0111011101010011", -- t[30547] = 16
      "010000" when "0111011101010100", -- t[30548] = 16
      "010000" when "0111011101010101", -- t[30549] = 16
      "010000" when "0111011101010110", -- t[30550] = 16
      "010000" when "0111011101010111", -- t[30551] = 16
      "010000" when "0111011101011000", -- t[30552] = 16
      "010000" when "0111011101011001", -- t[30553] = 16
      "010000" when "0111011101011010", -- t[30554] = 16
      "010000" when "0111011101011011", -- t[30555] = 16
      "010000" when "0111011101011100", -- t[30556] = 16
      "010000" when "0111011101011101", -- t[30557] = 16
      "010000" when "0111011101011110", -- t[30558] = 16
      "010000" when "0111011101011111", -- t[30559] = 16
      "010000" when "0111011101100000", -- t[30560] = 16
      "010000" when "0111011101100001", -- t[30561] = 16
      "010000" when "0111011101100010", -- t[30562] = 16
      "010000" when "0111011101100011", -- t[30563] = 16
      "010000" when "0111011101100100", -- t[30564] = 16
      "010000" when "0111011101100101", -- t[30565] = 16
      "010000" when "0111011101100110", -- t[30566] = 16
      "010000" when "0111011101100111", -- t[30567] = 16
      "010000" when "0111011101101000", -- t[30568] = 16
      "010000" when "0111011101101001", -- t[30569] = 16
      "010000" when "0111011101101010", -- t[30570] = 16
      "010000" when "0111011101101011", -- t[30571] = 16
      "010000" when "0111011101101100", -- t[30572] = 16
      "010000" when "0111011101101101", -- t[30573] = 16
      "010000" when "0111011101101110", -- t[30574] = 16
      "010000" when "0111011101101111", -- t[30575] = 16
      "010000" when "0111011101110000", -- t[30576] = 16
      "010000" when "0111011101110001", -- t[30577] = 16
      "010000" when "0111011101110010", -- t[30578] = 16
      "010000" when "0111011101110011", -- t[30579] = 16
      "010000" when "0111011101110100", -- t[30580] = 16
      "010000" when "0111011101110101", -- t[30581] = 16
      "010000" when "0111011101110110", -- t[30582] = 16
      "010000" when "0111011101110111", -- t[30583] = 16
      "010000" when "0111011101111000", -- t[30584] = 16
      "010000" when "0111011101111001", -- t[30585] = 16
      "010000" when "0111011101111010", -- t[30586] = 16
      "010000" when "0111011101111011", -- t[30587] = 16
      "010000" when "0111011101111100", -- t[30588] = 16
      "010000" when "0111011101111101", -- t[30589] = 16
      "010000" when "0111011101111110", -- t[30590] = 16
      "010000" when "0111011101111111", -- t[30591] = 16
      "010000" when "0111011110000000", -- t[30592] = 16
      "010000" when "0111011110000001", -- t[30593] = 16
      "010000" when "0111011110000010", -- t[30594] = 16
      "010000" when "0111011110000011", -- t[30595] = 16
      "010000" when "0111011110000100", -- t[30596] = 16
      "010000" when "0111011110000101", -- t[30597] = 16
      "010000" when "0111011110000110", -- t[30598] = 16
      "010000" when "0111011110000111", -- t[30599] = 16
      "010000" when "0111011110001000", -- t[30600] = 16
      "010000" when "0111011110001001", -- t[30601] = 16
      "010000" when "0111011110001010", -- t[30602] = 16
      "010000" when "0111011110001011", -- t[30603] = 16
      "010000" when "0111011110001100", -- t[30604] = 16
      "010000" when "0111011110001101", -- t[30605] = 16
      "010000" when "0111011110001110", -- t[30606] = 16
      "010000" when "0111011110001111", -- t[30607] = 16
      "010000" when "0111011110010000", -- t[30608] = 16
      "010000" when "0111011110010001", -- t[30609] = 16
      "010000" when "0111011110010010", -- t[30610] = 16
      "010000" when "0111011110010011", -- t[30611] = 16
      "010000" when "0111011110010100", -- t[30612] = 16
      "010000" when "0111011110010101", -- t[30613] = 16
      "010000" when "0111011110010110", -- t[30614] = 16
      "010000" when "0111011110010111", -- t[30615] = 16
      "010000" when "0111011110011000", -- t[30616] = 16
      "010000" when "0111011110011001", -- t[30617] = 16
      "010000" when "0111011110011010", -- t[30618] = 16
      "010000" when "0111011110011011", -- t[30619] = 16
      "010000" when "0111011110011100", -- t[30620] = 16
      "010000" when "0111011110011101", -- t[30621] = 16
      "010000" when "0111011110011110", -- t[30622] = 16
      "010000" when "0111011110011111", -- t[30623] = 16
      "010000" when "0111011110100000", -- t[30624] = 16
      "010000" when "0111011110100001", -- t[30625] = 16
      "010000" when "0111011110100010", -- t[30626] = 16
      "010000" when "0111011110100011", -- t[30627] = 16
      "010000" when "0111011110100100", -- t[30628] = 16
      "010000" when "0111011110100101", -- t[30629] = 16
      "010000" when "0111011110100110", -- t[30630] = 16
      "010000" when "0111011110100111", -- t[30631] = 16
      "010000" when "0111011110101000", -- t[30632] = 16
      "010000" when "0111011110101001", -- t[30633] = 16
      "010000" when "0111011110101010", -- t[30634] = 16
      "010000" when "0111011110101011", -- t[30635] = 16
      "010000" when "0111011110101100", -- t[30636] = 16
      "010000" when "0111011110101101", -- t[30637] = 16
      "010000" when "0111011110101110", -- t[30638] = 16
      "010000" when "0111011110101111", -- t[30639] = 16
      "010000" when "0111011110110000", -- t[30640] = 16
      "010000" when "0111011110110001", -- t[30641] = 16
      "010000" when "0111011110110010", -- t[30642] = 16
      "010000" when "0111011110110011", -- t[30643] = 16
      "010000" when "0111011110110100", -- t[30644] = 16
      "010000" when "0111011110110101", -- t[30645] = 16
      "010000" when "0111011110110110", -- t[30646] = 16
      "010000" when "0111011110110111", -- t[30647] = 16
      "010000" when "0111011110111000", -- t[30648] = 16
      "010000" when "0111011110111001", -- t[30649] = 16
      "010000" when "0111011110111010", -- t[30650] = 16
      "010000" when "0111011110111011", -- t[30651] = 16
      "010000" when "0111011110111100", -- t[30652] = 16
      "010000" when "0111011110111101", -- t[30653] = 16
      "010000" when "0111011110111110", -- t[30654] = 16
      "010000" when "0111011110111111", -- t[30655] = 16
      "010000" when "0111011111000000", -- t[30656] = 16
      "010000" when "0111011111000001", -- t[30657] = 16
      "010000" when "0111011111000010", -- t[30658] = 16
      "010000" when "0111011111000011", -- t[30659] = 16
      "010000" when "0111011111000100", -- t[30660] = 16
      "010000" when "0111011111000101", -- t[30661] = 16
      "010000" when "0111011111000110", -- t[30662] = 16
      "010000" when "0111011111000111", -- t[30663] = 16
      "010000" when "0111011111001000", -- t[30664] = 16
      "010000" when "0111011111001001", -- t[30665] = 16
      "010000" when "0111011111001010", -- t[30666] = 16
      "010000" when "0111011111001011", -- t[30667] = 16
      "010000" when "0111011111001100", -- t[30668] = 16
      "010000" when "0111011111001101", -- t[30669] = 16
      "010000" when "0111011111001110", -- t[30670] = 16
      "010000" when "0111011111001111", -- t[30671] = 16
      "010000" when "0111011111010000", -- t[30672] = 16
      "010000" when "0111011111010001", -- t[30673] = 16
      "010000" when "0111011111010010", -- t[30674] = 16
      "010000" when "0111011111010011", -- t[30675] = 16
      "010000" when "0111011111010100", -- t[30676] = 16
      "010000" when "0111011111010101", -- t[30677] = 16
      "010000" when "0111011111010110", -- t[30678] = 16
      "010000" when "0111011111010111", -- t[30679] = 16
      "010000" when "0111011111011000", -- t[30680] = 16
      "010000" when "0111011111011001", -- t[30681] = 16
      "010000" when "0111011111011010", -- t[30682] = 16
      "010000" when "0111011111011011", -- t[30683] = 16
      "010000" when "0111011111011100", -- t[30684] = 16
      "010000" when "0111011111011101", -- t[30685] = 16
      "010000" when "0111011111011110", -- t[30686] = 16
      "010000" when "0111011111011111", -- t[30687] = 16
      "010000" when "0111011111100000", -- t[30688] = 16
      "010000" when "0111011111100001", -- t[30689] = 16
      "010000" when "0111011111100010", -- t[30690] = 16
      "010000" when "0111011111100011", -- t[30691] = 16
      "010000" when "0111011111100100", -- t[30692] = 16
      "010000" when "0111011111100101", -- t[30693] = 16
      "010000" when "0111011111100110", -- t[30694] = 16
      "010000" when "0111011111100111", -- t[30695] = 16
      "010000" when "0111011111101000", -- t[30696] = 16
      "010000" when "0111011111101001", -- t[30697] = 16
      "010000" when "0111011111101010", -- t[30698] = 16
      "010000" when "0111011111101011", -- t[30699] = 16
      "010000" when "0111011111101100", -- t[30700] = 16
      "010000" when "0111011111101101", -- t[30701] = 16
      "010000" when "0111011111101110", -- t[30702] = 16
      "010000" when "0111011111101111", -- t[30703] = 16
      "010000" when "0111011111110000", -- t[30704] = 16
      "010000" when "0111011111110001", -- t[30705] = 16
      "010000" when "0111011111110010", -- t[30706] = 16
      "010000" when "0111011111110011", -- t[30707] = 16
      "010000" when "0111011111110100", -- t[30708] = 16
      "010000" when "0111011111110101", -- t[30709] = 16
      "010000" when "0111011111110110", -- t[30710] = 16
      "010000" when "0111011111110111", -- t[30711] = 16
      "010000" when "0111011111111000", -- t[30712] = 16
      "010000" when "0111011111111001", -- t[30713] = 16
      "010000" when "0111011111111010", -- t[30714] = 16
      "010000" when "0111011111111011", -- t[30715] = 16
      "010000" when "0111011111111100", -- t[30716] = 16
      "010000" when "0111011111111101", -- t[30717] = 16
      "010000" when "0111011111111110", -- t[30718] = 16
      "010000" when "0111011111111111", -- t[30719] = 16
      "010000" when "0111100000000000", -- t[30720] = 16
      "010000" when "0111100000000001", -- t[30721] = 16
      "010000" when "0111100000000010", -- t[30722] = 16
      "010000" when "0111100000000011", -- t[30723] = 16
      "010000" when "0111100000000100", -- t[30724] = 16
      "010000" when "0111100000000101", -- t[30725] = 16
      "010000" when "0111100000000110", -- t[30726] = 16
      "010000" when "0111100000000111", -- t[30727] = 16
      "010000" when "0111100000001000", -- t[30728] = 16
      "010000" when "0111100000001001", -- t[30729] = 16
      "010000" when "0111100000001010", -- t[30730] = 16
      "010000" when "0111100000001011", -- t[30731] = 16
      "010000" when "0111100000001100", -- t[30732] = 16
      "010000" when "0111100000001101", -- t[30733] = 16
      "010000" when "0111100000001110", -- t[30734] = 16
      "010000" when "0111100000001111", -- t[30735] = 16
      "010000" when "0111100000010000", -- t[30736] = 16
      "010000" when "0111100000010001", -- t[30737] = 16
      "010000" when "0111100000010010", -- t[30738] = 16
      "010000" when "0111100000010011", -- t[30739] = 16
      "010000" when "0111100000010100", -- t[30740] = 16
      "010000" when "0111100000010101", -- t[30741] = 16
      "010000" when "0111100000010110", -- t[30742] = 16
      "010000" when "0111100000010111", -- t[30743] = 16
      "010000" when "0111100000011000", -- t[30744] = 16
      "010000" when "0111100000011001", -- t[30745] = 16
      "010000" when "0111100000011010", -- t[30746] = 16
      "010000" when "0111100000011011", -- t[30747] = 16
      "010000" when "0111100000011100", -- t[30748] = 16
      "010000" when "0111100000011101", -- t[30749] = 16
      "010000" when "0111100000011110", -- t[30750] = 16
      "010000" when "0111100000011111", -- t[30751] = 16
      "010000" when "0111100000100000", -- t[30752] = 16
      "010000" when "0111100000100001", -- t[30753] = 16
      "010000" when "0111100000100010", -- t[30754] = 16
      "010000" when "0111100000100011", -- t[30755] = 16
      "010000" when "0111100000100100", -- t[30756] = 16
      "010000" when "0111100000100101", -- t[30757] = 16
      "010000" when "0111100000100110", -- t[30758] = 16
      "010000" when "0111100000100111", -- t[30759] = 16
      "010000" when "0111100000101000", -- t[30760] = 16
      "010000" when "0111100000101001", -- t[30761] = 16
      "010000" when "0111100000101010", -- t[30762] = 16
      "010000" when "0111100000101011", -- t[30763] = 16
      "010000" when "0111100000101100", -- t[30764] = 16
      "010000" when "0111100000101101", -- t[30765] = 16
      "010000" when "0111100000101110", -- t[30766] = 16
      "010000" when "0111100000101111", -- t[30767] = 16
      "010000" when "0111100000110000", -- t[30768] = 16
      "010000" when "0111100000110001", -- t[30769] = 16
      "010000" when "0111100000110010", -- t[30770] = 16
      "010000" when "0111100000110011", -- t[30771] = 16
      "010000" when "0111100000110100", -- t[30772] = 16
      "010000" when "0111100000110101", -- t[30773] = 16
      "010000" when "0111100000110110", -- t[30774] = 16
      "010000" when "0111100000110111", -- t[30775] = 16
      "010001" when "0111100000111000", -- t[30776] = 17
      "010001" when "0111100000111001", -- t[30777] = 17
      "010001" when "0111100000111010", -- t[30778] = 17
      "010001" when "0111100000111011", -- t[30779] = 17
      "010001" when "0111100000111100", -- t[30780] = 17
      "010001" when "0111100000111101", -- t[30781] = 17
      "010001" when "0111100000111110", -- t[30782] = 17
      "010001" when "0111100000111111", -- t[30783] = 17
      "010001" when "0111100001000000", -- t[30784] = 17
      "010001" when "0111100001000001", -- t[30785] = 17
      "010001" when "0111100001000010", -- t[30786] = 17
      "010001" when "0111100001000011", -- t[30787] = 17
      "010001" when "0111100001000100", -- t[30788] = 17
      "010001" when "0111100001000101", -- t[30789] = 17
      "010001" when "0111100001000110", -- t[30790] = 17
      "010001" when "0111100001000111", -- t[30791] = 17
      "010001" when "0111100001001000", -- t[30792] = 17
      "010001" when "0111100001001001", -- t[30793] = 17
      "010001" when "0111100001001010", -- t[30794] = 17
      "010001" when "0111100001001011", -- t[30795] = 17
      "010001" when "0111100001001100", -- t[30796] = 17
      "010001" when "0111100001001101", -- t[30797] = 17
      "010001" when "0111100001001110", -- t[30798] = 17
      "010001" when "0111100001001111", -- t[30799] = 17
      "010001" when "0111100001010000", -- t[30800] = 17
      "010001" when "0111100001010001", -- t[30801] = 17
      "010001" when "0111100001010010", -- t[30802] = 17
      "010001" when "0111100001010011", -- t[30803] = 17
      "010001" when "0111100001010100", -- t[30804] = 17
      "010001" when "0111100001010101", -- t[30805] = 17
      "010001" when "0111100001010110", -- t[30806] = 17
      "010001" when "0111100001010111", -- t[30807] = 17
      "010001" when "0111100001011000", -- t[30808] = 17
      "010001" when "0111100001011001", -- t[30809] = 17
      "010001" when "0111100001011010", -- t[30810] = 17
      "010001" when "0111100001011011", -- t[30811] = 17
      "010001" when "0111100001011100", -- t[30812] = 17
      "010001" when "0111100001011101", -- t[30813] = 17
      "010001" when "0111100001011110", -- t[30814] = 17
      "010001" when "0111100001011111", -- t[30815] = 17
      "010001" when "0111100001100000", -- t[30816] = 17
      "010001" when "0111100001100001", -- t[30817] = 17
      "010001" when "0111100001100010", -- t[30818] = 17
      "010001" when "0111100001100011", -- t[30819] = 17
      "010001" when "0111100001100100", -- t[30820] = 17
      "010001" when "0111100001100101", -- t[30821] = 17
      "010001" when "0111100001100110", -- t[30822] = 17
      "010001" when "0111100001100111", -- t[30823] = 17
      "010001" when "0111100001101000", -- t[30824] = 17
      "010001" when "0111100001101001", -- t[30825] = 17
      "010001" when "0111100001101010", -- t[30826] = 17
      "010001" when "0111100001101011", -- t[30827] = 17
      "010001" when "0111100001101100", -- t[30828] = 17
      "010001" when "0111100001101101", -- t[30829] = 17
      "010001" when "0111100001101110", -- t[30830] = 17
      "010001" when "0111100001101111", -- t[30831] = 17
      "010001" when "0111100001110000", -- t[30832] = 17
      "010001" when "0111100001110001", -- t[30833] = 17
      "010001" when "0111100001110010", -- t[30834] = 17
      "010001" when "0111100001110011", -- t[30835] = 17
      "010001" when "0111100001110100", -- t[30836] = 17
      "010001" when "0111100001110101", -- t[30837] = 17
      "010001" when "0111100001110110", -- t[30838] = 17
      "010001" when "0111100001110111", -- t[30839] = 17
      "010001" when "0111100001111000", -- t[30840] = 17
      "010001" when "0111100001111001", -- t[30841] = 17
      "010001" when "0111100001111010", -- t[30842] = 17
      "010001" when "0111100001111011", -- t[30843] = 17
      "010001" when "0111100001111100", -- t[30844] = 17
      "010001" when "0111100001111101", -- t[30845] = 17
      "010001" when "0111100001111110", -- t[30846] = 17
      "010001" when "0111100001111111", -- t[30847] = 17
      "010001" when "0111100010000000", -- t[30848] = 17
      "010001" when "0111100010000001", -- t[30849] = 17
      "010001" when "0111100010000010", -- t[30850] = 17
      "010001" when "0111100010000011", -- t[30851] = 17
      "010001" when "0111100010000100", -- t[30852] = 17
      "010001" when "0111100010000101", -- t[30853] = 17
      "010001" when "0111100010000110", -- t[30854] = 17
      "010001" when "0111100010000111", -- t[30855] = 17
      "010001" when "0111100010001000", -- t[30856] = 17
      "010001" when "0111100010001001", -- t[30857] = 17
      "010001" when "0111100010001010", -- t[30858] = 17
      "010001" when "0111100010001011", -- t[30859] = 17
      "010001" when "0111100010001100", -- t[30860] = 17
      "010001" when "0111100010001101", -- t[30861] = 17
      "010001" when "0111100010001110", -- t[30862] = 17
      "010001" when "0111100010001111", -- t[30863] = 17
      "010001" when "0111100010010000", -- t[30864] = 17
      "010001" when "0111100010010001", -- t[30865] = 17
      "010001" when "0111100010010010", -- t[30866] = 17
      "010001" when "0111100010010011", -- t[30867] = 17
      "010001" when "0111100010010100", -- t[30868] = 17
      "010001" when "0111100010010101", -- t[30869] = 17
      "010001" when "0111100010010110", -- t[30870] = 17
      "010001" when "0111100010010111", -- t[30871] = 17
      "010001" when "0111100010011000", -- t[30872] = 17
      "010001" when "0111100010011001", -- t[30873] = 17
      "010001" when "0111100010011010", -- t[30874] = 17
      "010001" when "0111100010011011", -- t[30875] = 17
      "010001" when "0111100010011100", -- t[30876] = 17
      "010001" when "0111100010011101", -- t[30877] = 17
      "010001" when "0111100010011110", -- t[30878] = 17
      "010001" when "0111100010011111", -- t[30879] = 17
      "010001" when "0111100010100000", -- t[30880] = 17
      "010001" when "0111100010100001", -- t[30881] = 17
      "010001" when "0111100010100010", -- t[30882] = 17
      "010001" when "0111100010100011", -- t[30883] = 17
      "010001" when "0111100010100100", -- t[30884] = 17
      "010001" when "0111100010100101", -- t[30885] = 17
      "010001" when "0111100010100110", -- t[30886] = 17
      "010001" when "0111100010100111", -- t[30887] = 17
      "010001" when "0111100010101000", -- t[30888] = 17
      "010001" when "0111100010101001", -- t[30889] = 17
      "010001" when "0111100010101010", -- t[30890] = 17
      "010001" when "0111100010101011", -- t[30891] = 17
      "010001" when "0111100010101100", -- t[30892] = 17
      "010001" when "0111100010101101", -- t[30893] = 17
      "010001" when "0111100010101110", -- t[30894] = 17
      "010001" when "0111100010101111", -- t[30895] = 17
      "010001" when "0111100010110000", -- t[30896] = 17
      "010001" when "0111100010110001", -- t[30897] = 17
      "010001" when "0111100010110010", -- t[30898] = 17
      "010001" when "0111100010110011", -- t[30899] = 17
      "010001" when "0111100010110100", -- t[30900] = 17
      "010001" when "0111100010110101", -- t[30901] = 17
      "010001" when "0111100010110110", -- t[30902] = 17
      "010001" when "0111100010110111", -- t[30903] = 17
      "010001" when "0111100010111000", -- t[30904] = 17
      "010001" when "0111100010111001", -- t[30905] = 17
      "010001" when "0111100010111010", -- t[30906] = 17
      "010001" when "0111100010111011", -- t[30907] = 17
      "010001" when "0111100010111100", -- t[30908] = 17
      "010001" when "0111100010111101", -- t[30909] = 17
      "010001" when "0111100010111110", -- t[30910] = 17
      "010001" when "0111100010111111", -- t[30911] = 17
      "010001" when "0111100011000000", -- t[30912] = 17
      "010001" when "0111100011000001", -- t[30913] = 17
      "010001" when "0111100011000010", -- t[30914] = 17
      "010001" when "0111100011000011", -- t[30915] = 17
      "010001" when "0111100011000100", -- t[30916] = 17
      "010001" when "0111100011000101", -- t[30917] = 17
      "010001" when "0111100011000110", -- t[30918] = 17
      "010001" when "0111100011000111", -- t[30919] = 17
      "010001" when "0111100011001000", -- t[30920] = 17
      "010001" when "0111100011001001", -- t[30921] = 17
      "010001" when "0111100011001010", -- t[30922] = 17
      "010001" when "0111100011001011", -- t[30923] = 17
      "010001" when "0111100011001100", -- t[30924] = 17
      "010001" when "0111100011001101", -- t[30925] = 17
      "010001" when "0111100011001110", -- t[30926] = 17
      "010001" when "0111100011001111", -- t[30927] = 17
      "010001" when "0111100011010000", -- t[30928] = 17
      "010001" when "0111100011010001", -- t[30929] = 17
      "010001" when "0111100011010010", -- t[30930] = 17
      "010001" when "0111100011010011", -- t[30931] = 17
      "010001" when "0111100011010100", -- t[30932] = 17
      "010001" when "0111100011010101", -- t[30933] = 17
      "010001" when "0111100011010110", -- t[30934] = 17
      "010001" when "0111100011010111", -- t[30935] = 17
      "010001" when "0111100011011000", -- t[30936] = 17
      "010001" when "0111100011011001", -- t[30937] = 17
      "010001" when "0111100011011010", -- t[30938] = 17
      "010001" when "0111100011011011", -- t[30939] = 17
      "010001" when "0111100011011100", -- t[30940] = 17
      "010001" when "0111100011011101", -- t[30941] = 17
      "010001" when "0111100011011110", -- t[30942] = 17
      "010001" when "0111100011011111", -- t[30943] = 17
      "010001" when "0111100011100000", -- t[30944] = 17
      "010001" when "0111100011100001", -- t[30945] = 17
      "010001" when "0111100011100010", -- t[30946] = 17
      "010001" when "0111100011100011", -- t[30947] = 17
      "010001" when "0111100011100100", -- t[30948] = 17
      "010001" when "0111100011100101", -- t[30949] = 17
      "010001" when "0111100011100110", -- t[30950] = 17
      "010001" when "0111100011100111", -- t[30951] = 17
      "010001" when "0111100011101000", -- t[30952] = 17
      "010001" when "0111100011101001", -- t[30953] = 17
      "010001" when "0111100011101010", -- t[30954] = 17
      "010001" when "0111100011101011", -- t[30955] = 17
      "010001" when "0111100011101100", -- t[30956] = 17
      "010001" when "0111100011101101", -- t[30957] = 17
      "010001" when "0111100011101110", -- t[30958] = 17
      "010001" when "0111100011101111", -- t[30959] = 17
      "010001" when "0111100011110000", -- t[30960] = 17
      "010001" when "0111100011110001", -- t[30961] = 17
      "010001" when "0111100011110010", -- t[30962] = 17
      "010001" when "0111100011110011", -- t[30963] = 17
      "010001" when "0111100011110100", -- t[30964] = 17
      "010001" when "0111100011110101", -- t[30965] = 17
      "010001" when "0111100011110110", -- t[30966] = 17
      "010001" when "0111100011110111", -- t[30967] = 17
      "010001" when "0111100011111000", -- t[30968] = 17
      "010001" when "0111100011111001", -- t[30969] = 17
      "010001" when "0111100011111010", -- t[30970] = 17
      "010001" when "0111100011111011", -- t[30971] = 17
      "010001" when "0111100011111100", -- t[30972] = 17
      "010001" when "0111100011111101", -- t[30973] = 17
      "010001" when "0111100011111110", -- t[30974] = 17
      "010001" when "0111100011111111", -- t[30975] = 17
      "010001" when "0111100100000000", -- t[30976] = 17
      "010001" when "0111100100000001", -- t[30977] = 17
      "010001" when "0111100100000010", -- t[30978] = 17
      "010001" when "0111100100000011", -- t[30979] = 17
      "010001" when "0111100100000100", -- t[30980] = 17
      "010001" when "0111100100000101", -- t[30981] = 17
      "010001" when "0111100100000110", -- t[30982] = 17
      "010001" when "0111100100000111", -- t[30983] = 17
      "010001" when "0111100100001000", -- t[30984] = 17
      "010001" when "0111100100001001", -- t[30985] = 17
      "010001" when "0111100100001010", -- t[30986] = 17
      "010001" when "0111100100001011", -- t[30987] = 17
      "010001" when "0111100100001100", -- t[30988] = 17
      "010001" when "0111100100001101", -- t[30989] = 17
      "010001" when "0111100100001110", -- t[30990] = 17
      "010001" when "0111100100001111", -- t[30991] = 17
      "010001" when "0111100100010000", -- t[30992] = 17
      "010001" when "0111100100010001", -- t[30993] = 17
      "010001" when "0111100100010010", -- t[30994] = 17
      "010001" when "0111100100010011", -- t[30995] = 17
      "010001" when "0111100100010100", -- t[30996] = 17
      "010001" when "0111100100010101", -- t[30997] = 17
      "010001" when "0111100100010110", -- t[30998] = 17
      "010001" when "0111100100010111", -- t[30999] = 17
      "010001" when "0111100100011000", -- t[31000] = 17
      "010001" when "0111100100011001", -- t[31001] = 17
      "010001" when "0111100100011010", -- t[31002] = 17
      "010001" when "0111100100011011", -- t[31003] = 17
      "010001" when "0111100100011100", -- t[31004] = 17
      "010001" when "0111100100011101", -- t[31005] = 17
      "010001" when "0111100100011110", -- t[31006] = 17
      "010001" when "0111100100011111", -- t[31007] = 17
      "010001" when "0111100100100000", -- t[31008] = 17
      "010001" when "0111100100100001", -- t[31009] = 17
      "010001" when "0111100100100010", -- t[31010] = 17
      "010001" when "0111100100100011", -- t[31011] = 17
      "010001" when "0111100100100100", -- t[31012] = 17
      "010001" when "0111100100100101", -- t[31013] = 17
      "010001" when "0111100100100110", -- t[31014] = 17
      "010001" when "0111100100100111", -- t[31015] = 17
      "010001" when "0111100100101000", -- t[31016] = 17
      "010001" when "0111100100101001", -- t[31017] = 17
      "010001" when "0111100100101010", -- t[31018] = 17
      "010001" when "0111100100101011", -- t[31019] = 17
      "010001" when "0111100100101100", -- t[31020] = 17
      "010001" when "0111100100101101", -- t[31021] = 17
      "010001" when "0111100100101110", -- t[31022] = 17
      "010001" when "0111100100101111", -- t[31023] = 17
      "010001" when "0111100100110000", -- t[31024] = 17
      "010001" when "0111100100110001", -- t[31025] = 17
      "010001" when "0111100100110010", -- t[31026] = 17
      "010001" when "0111100100110011", -- t[31027] = 17
      "010001" when "0111100100110100", -- t[31028] = 17
      "010001" when "0111100100110101", -- t[31029] = 17
      "010001" when "0111100100110110", -- t[31030] = 17
      "010001" when "0111100100110111", -- t[31031] = 17
      "010001" when "0111100100111000", -- t[31032] = 17
      "010001" when "0111100100111001", -- t[31033] = 17
      "010001" when "0111100100111010", -- t[31034] = 17
      "010001" when "0111100100111011", -- t[31035] = 17
      "010001" when "0111100100111100", -- t[31036] = 17
      "010001" when "0111100100111101", -- t[31037] = 17
      "010001" when "0111100100111110", -- t[31038] = 17
      "010001" when "0111100100111111", -- t[31039] = 17
      "010001" when "0111100101000000", -- t[31040] = 17
      "010001" when "0111100101000001", -- t[31041] = 17
      "010001" when "0111100101000010", -- t[31042] = 17
      "010001" when "0111100101000011", -- t[31043] = 17
      "010001" when "0111100101000100", -- t[31044] = 17
      "010001" when "0111100101000101", -- t[31045] = 17
      "010001" when "0111100101000110", -- t[31046] = 17
      "010001" when "0111100101000111", -- t[31047] = 17
      "010001" when "0111100101001000", -- t[31048] = 17
      "010001" when "0111100101001001", -- t[31049] = 17
      "010001" when "0111100101001010", -- t[31050] = 17
      "010001" when "0111100101001011", -- t[31051] = 17
      "010001" when "0111100101001100", -- t[31052] = 17
      "010001" when "0111100101001101", -- t[31053] = 17
      "010001" when "0111100101001110", -- t[31054] = 17
      "010001" when "0111100101001111", -- t[31055] = 17
      "010001" when "0111100101010000", -- t[31056] = 17
      "010001" when "0111100101010001", -- t[31057] = 17
      "010001" when "0111100101010010", -- t[31058] = 17
      "010001" when "0111100101010011", -- t[31059] = 17
      "010001" when "0111100101010100", -- t[31060] = 17
      "010001" when "0111100101010101", -- t[31061] = 17
      "010001" when "0111100101010110", -- t[31062] = 17
      "010001" when "0111100101010111", -- t[31063] = 17
      "010001" when "0111100101011000", -- t[31064] = 17
      "010001" when "0111100101011001", -- t[31065] = 17
      "010001" when "0111100101011010", -- t[31066] = 17
      "010001" when "0111100101011011", -- t[31067] = 17
      "010001" when "0111100101011100", -- t[31068] = 17
      "010001" when "0111100101011101", -- t[31069] = 17
      "010001" when "0111100101011110", -- t[31070] = 17
      "010001" when "0111100101011111", -- t[31071] = 17
      "010001" when "0111100101100000", -- t[31072] = 17
      "010001" when "0111100101100001", -- t[31073] = 17
      "010001" when "0111100101100010", -- t[31074] = 17
      "010001" when "0111100101100011", -- t[31075] = 17
      "010001" when "0111100101100100", -- t[31076] = 17
      "010001" when "0111100101100101", -- t[31077] = 17
      "010001" when "0111100101100110", -- t[31078] = 17
      "010001" when "0111100101100111", -- t[31079] = 17
      "010001" when "0111100101101000", -- t[31080] = 17
      "010001" when "0111100101101001", -- t[31081] = 17
      "010001" when "0111100101101010", -- t[31082] = 17
      "010001" when "0111100101101011", -- t[31083] = 17
      "010001" when "0111100101101100", -- t[31084] = 17
      "010001" when "0111100101101101", -- t[31085] = 17
      "010001" when "0111100101101110", -- t[31086] = 17
      "010001" when "0111100101101111", -- t[31087] = 17
      "010001" when "0111100101110000", -- t[31088] = 17
      "010001" when "0111100101110001", -- t[31089] = 17
      "010001" when "0111100101110010", -- t[31090] = 17
      "010001" when "0111100101110011", -- t[31091] = 17
      "010001" when "0111100101110100", -- t[31092] = 17
      "010001" when "0111100101110101", -- t[31093] = 17
      "010001" when "0111100101110110", -- t[31094] = 17
      "010001" when "0111100101110111", -- t[31095] = 17
      "010001" when "0111100101111000", -- t[31096] = 17
      "010001" when "0111100101111001", -- t[31097] = 17
      "010001" when "0111100101111010", -- t[31098] = 17
      "010001" when "0111100101111011", -- t[31099] = 17
      "010001" when "0111100101111100", -- t[31100] = 17
      "010001" when "0111100101111101", -- t[31101] = 17
      "010001" when "0111100101111110", -- t[31102] = 17
      "010001" when "0111100101111111", -- t[31103] = 17
      "010001" when "0111100110000000", -- t[31104] = 17
      "010001" when "0111100110000001", -- t[31105] = 17
      "010001" when "0111100110000010", -- t[31106] = 17
      "010001" when "0111100110000011", -- t[31107] = 17
      "010001" when "0111100110000100", -- t[31108] = 17
      "010001" when "0111100110000101", -- t[31109] = 17
      "010001" when "0111100110000110", -- t[31110] = 17
      "010001" when "0111100110000111", -- t[31111] = 17
      "010001" when "0111100110001000", -- t[31112] = 17
      "010001" when "0111100110001001", -- t[31113] = 17
      "010001" when "0111100110001010", -- t[31114] = 17
      "010001" when "0111100110001011", -- t[31115] = 17
      "010001" when "0111100110001100", -- t[31116] = 17
      "010001" when "0111100110001101", -- t[31117] = 17
      "010001" when "0111100110001110", -- t[31118] = 17
      "010001" when "0111100110001111", -- t[31119] = 17
      "010001" when "0111100110010000", -- t[31120] = 17
      "010001" when "0111100110010001", -- t[31121] = 17
      "010001" when "0111100110010010", -- t[31122] = 17
      "010010" when "0111100110010011", -- t[31123] = 18
      "010010" when "0111100110010100", -- t[31124] = 18
      "010010" when "0111100110010101", -- t[31125] = 18
      "010010" when "0111100110010110", -- t[31126] = 18
      "010010" when "0111100110010111", -- t[31127] = 18
      "010010" when "0111100110011000", -- t[31128] = 18
      "010010" when "0111100110011001", -- t[31129] = 18
      "010010" when "0111100110011010", -- t[31130] = 18
      "010010" when "0111100110011011", -- t[31131] = 18
      "010010" when "0111100110011100", -- t[31132] = 18
      "010010" when "0111100110011101", -- t[31133] = 18
      "010010" when "0111100110011110", -- t[31134] = 18
      "010010" when "0111100110011111", -- t[31135] = 18
      "010010" when "0111100110100000", -- t[31136] = 18
      "010010" when "0111100110100001", -- t[31137] = 18
      "010010" when "0111100110100010", -- t[31138] = 18
      "010010" when "0111100110100011", -- t[31139] = 18
      "010010" when "0111100110100100", -- t[31140] = 18
      "010010" when "0111100110100101", -- t[31141] = 18
      "010010" when "0111100110100110", -- t[31142] = 18
      "010010" when "0111100110100111", -- t[31143] = 18
      "010010" when "0111100110101000", -- t[31144] = 18
      "010010" when "0111100110101001", -- t[31145] = 18
      "010010" when "0111100110101010", -- t[31146] = 18
      "010010" when "0111100110101011", -- t[31147] = 18
      "010010" when "0111100110101100", -- t[31148] = 18
      "010010" when "0111100110101101", -- t[31149] = 18
      "010010" when "0111100110101110", -- t[31150] = 18
      "010010" when "0111100110101111", -- t[31151] = 18
      "010010" when "0111100110110000", -- t[31152] = 18
      "010010" when "0111100110110001", -- t[31153] = 18
      "010010" when "0111100110110010", -- t[31154] = 18
      "010010" when "0111100110110011", -- t[31155] = 18
      "010010" when "0111100110110100", -- t[31156] = 18
      "010010" when "0111100110110101", -- t[31157] = 18
      "010010" when "0111100110110110", -- t[31158] = 18
      "010010" when "0111100110110111", -- t[31159] = 18
      "010010" when "0111100110111000", -- t[31160] = 18
      "010010" when "0111100110111001", -- t[31161] = 18
      "010010" when "0111100110111010", -- t[31162] = 18
      "010010" when "0111100110111011", -- t[31163] = 18
      "010010" when "0111100110111100", -- t[31164] = 18
      "010010" when "0111100110111101", -- t[31165] = 18
      "010010" when "0111100110111110", -- t[31166] = 18
      "010010" when "0111100110111111", -- t[31167] = 18
      "010010" when "0111100111000000", -- t[31168] = 18
      "010010" when "0111100111000001", -- t[31169] = 18
      "010010" when "0111100111000010", -- t[31170] = 18
      "010010" when "0111100111000011", -- t[31171] = 18
      "010010" when "0111100111000100", -- t[31172] = 18
      "010010" when "0111100111000101", -- t[31173] = 18
      "010010" when "0111100111000110", -- t[31174] = 18
      "010010" when "0111100111000111", -- t[31175] = 18
      "010010" when "0111100111001000", -- t[31176] = 18
      "010010" when "0111100111001001", -- t[31177] = 18
      "010010" when "0111100111001010", -- t[31178] = 18
      "010010" when "0111100111001011", -- t[31179] = 18
      "010010" when "0111100111001100", -- t[31180] = 18
      "010010" when "0111100111001101", -- t[31181] = 18
      "010010" when "0111100111001110", -- t[31182] = 18
      "010010" when "0111100111001111", -- t[31183] = 18
      "010010" when "0111100111010000", -- t[31184] = 18
      "010010" when "0111100111010001", -- t[31185] = 18
      "010010" when "0111100111010010", -- t[31186] = 18
      "010010" when "0111100111010011", -- t[31187] = 18
      "010010" when "0111100111010100", -- t[31188] = 18
      "010010" when "0111100111010101", -- t[31189] = 18
      "010010" when "0111100111010110", -- t[31190] = 18
      "010010" when "0111100111010111", -- t[31191] = 18
      "010010" when "0111100111011000", -- t[31192] = 18
      "010010" when "0111100111011001", -- t[31193] = 18
      "010010" when "0111100111011010", -- t[31194] = 18
      "010010" when "0111100111011011", -- t[31195] = 18
      "010010" when "0111100111011100", -- t[31196] = 18
      "010010" when "0111100111011101", -- t[31197] = 18
      "010010" when "0111100111011110", -- t[31198] = 18
      "010010" when "0111100111011111", -- t[31199] = 18
      "010010" when "0111100111100000", -- t[31200] = 18
      "010010" when "0111100111100001", -- t[31201] = 18
      "010010" when "0111100111100010", -- t[31202] = 18
      "010010" when "0111100111100011", -- t[31203] = 18
      "010010" when "0111100111100100", -- t[31204] = 18
      "010010" when "0111100111100101", -- t[31205] = 18
      "010010" when "0111100111100110", -- t[31206] = 18
      "010010" when "0111100111100111", -- t[31207] = 18
      "010010" when "0111100111101000", -- t[31208] = 18
      "010010" when "0111100111101001", -- t[31209] = 18
      "010010" when "0111100111101010", -- t[31210] = 18
      "010010" when "0111100111101011", -- t[31211] = 18
      "010010" when "0111100111101100", -- t[31212] = 18
      "010010" when "0111100111101101", -- t[31213] = 18
      "010010" when "0111100111101110", -- t[31214] = 18
      "010010" when "0111100111101111", -- t[31215] = 18
      "010010" when "0111100111110000", -- t[31216] = 18
      "010010" when "0111100111110001", -- t[31217] = 18
      "010010" when "0111100111110010", -- t[31218] = 18
      "010010" when "0111100111110011", -- t[31219] = 18
      "010010" when "0111100111110100", -- t[31220] = 18
      "010010" when "0111100111110101", -- t[31221] = 18
      "010010" when "0111100111110110", -- t[31222] = 18
      "010010" when "0111100111110111", -- t[31223] = 18
      "010010" when "0111100111111000", -- t[31224] = 18
      "010010" when "0111100111111001", -- t[31225] = 18
      "010010" when "0111100111111010", -- t[31226] = 18
      "010010" when "0111100111111011", -- t[31227] = 18
      "010010" when "0111100111111100", -- t[31228] = 18
      "010010" when "0111100111111101", -- t[31229] = 18
      "010010" when "0111100111111110", -- t[31230] = 18
      "010010" when "0111100111111111", -- t[31231] = 18
      "010010" when "0111101000000000", -- t[31232] = 18
      "010010" when "0111101000000001", -- t[31233] = 18
      "010010" when "0111101000000010", -- t[31234] = 18
      "010010" when "0111101000000011", -- t[31235] = 18
      "010010" when "0111101000000100", -- t[31236] = 18
      "010010" when "0111101000000101", -- t[31237] = 18
      "010010" when "0111101000000110", -- t[31238] = 18
      "010010" when "0111101000000111", -- t[31239] = 18
      "010010" when "0111101000001000", -- t[31240] = 18
      "010010" when "0111101000001001", -- t[31241] = 18
      "010010" when "0111101000001010", -- t[31242] = 18
      "010010" when "0111101000001011", -- t[31243] = 18
      "010010" when "0111101000001100", -- t[31244] = 18
      "010010" when "0111101000001101", -- t[31245] = 18
      "010010" when "0111101000001110", -- t[31246] = 18
      "010010" when "0111101000001111", -- t[31247] = 18
      "010010" when "0111101000010000", -- t[31248] = 18
      "010010" when "0111101000010001", -- t[31249] = 18
      "010010" when "0111101000010010", -- t[31250] = 18
      "010010" when "0111101000010011", -- t[31251] = 18
      "010010" when "0111101000010100", -- t[31252] = 18
      "010010" when "0111101000010101", -- t[31253] = 18
      "010010" when "0111101000010110", -- t[31254] = 18
      "010010" when "0111101000010111", -- t[31255] = 18
      "010010" when "0111101000011000", -- t[31256] = 18
      "010010" when "0111101000011001", -- t[31257] = 18
      "010010" when "0111101000011010", -- t[31258] = 18
      "010010" when "0111101000011011", -- t[31259] = 18
      "010010" when "0111101000011100", -- t[31260] = 18
      "010010" when "0111101000011101", -- t[31261] = 18
      "010010" when "0111101000011110", -- t[31262] = 18
      "010010" when "0111101000011111", -- t[31263] = 18
      "010010" when "0111101000100000", -- t[31264] = 18
      "010010" when "0111101000100001", -- t[31265] = 18
      "010010" when "0111101000100010", -- t[31266] = 18
      "010010" when "0111101000100011", -- t[31267] = 18
      "010010" when "0111101000100100", -- t[31268] = 18
      "010010" when "0111101000100101", -- t[31269] = 18
      "010010" when "0111101000100110", -- t[31270] = 18
      "010010" when "0111101000100111", -- t[31271] = 18
      "010010" when "0111101000101000", -- t[31272] = 18
      "010010" when "0111101000101001", -- t[31273] = 18
      "010010" when "0111101000101010", -- t[31274] = 18
      "010010" when "0111101000101011", -- t[31275] = 18
      "010010" when "0111101000101100", -- t[31276] = 18
      "010010" when "0111101000101101", -- t[31277] = 18
      "010010" when "0111101000101110", -- t[31278] = 18
      "010010" when "0111101000101111", -- t[31279] = 18
      "010010" when "0111101000110000", -- t[31280] = 18
      "010010" when "0111101000110001", -- t[31281] = 18
      "010010" when "0111101000110010", -- t[31282] = 18
      "010010" when "0111101000110011", -- t[31283] = 18
      "010010" when "0111101000110100", -- t[31284] = 18
      "010010" when "0111101000110101", -- t[31285] = 18
      "010010" when "0111101000110110", -- t[31286] = 18
      "010010" when "0111101000110111", -- t[31287] = 18
      "010010" when "0111101000111000", -- t[31288] = 18
      "010010" when "0111101000111001", -- t[31289] = 18
      "010010" when "0111101000111010", -- t[31290] = 18
      "010010" when "0111101000111011", -- t[31291] = 18
      "010010" when "0111101000111100", -- t[31292] = 18
      "010010" when "0111101000111101", -- t[31293] = 18
      "010010" when "0111101000111110", -- t[31294] = 18
      "010010" when "0111101000111111", -- t[31295] = 18
      "010010" when "0111101001000000", -- t[31296] = 18
      "010010" when "0111101001000001", -- t[31297] = 18
      "010010" when "0111101001000010", -- t[31298] = 18
      "010010" when "0111101001000011", -- t[31299] = 18
      "010010" when "0111101001000100", -- t[31300] = 18
      "010010" when "0111101001000101", -- t[31301] = 18
      "010010" when "0111101001000110", -- t[31302] = 18
      "010010" when "0111101001000111", -- t[31303] = 18
      "010010" when "0111101001001000", -- t[31304] = 18
      "010010" when "0111101001001001", -- t[31305] = 18
      "010010" when "0111101001001010", -- t[31306] = 18
      "010010" when "0111101001001011", -- t[31307] = 18
      "010010" when "0111101001001100", -- t[31308] = 18
      "010010" when "0111101001001101", -- t[31309] = 18
      "010010" when "0111101001001110", -- t[31310] = 18
      "010010" when "0111101001001111", -- t[31311] = 18
      "010010" when "0111101001010000", -- t[31312] = 18
      "010010" when "0111101001010001", -- t[31313] = 18
      "010010" when "0111101001010010", -- t[31314] = 18
      "010010" when "0111101001010011", -- t[31315] = 18
      "010010" when "0111101001010100", -- t[31316] = 18
      "010010" when "0111101001010101", -- t[31317] = 18
      "010010" when "0111101001010110", -- t[31318] = 18
      "010010" when "0111101001010111", -- t[31319] = 18
      "010010" when "0111101001011000", -- t[31320] = 18
      "010010" when "0111101001011001", -- t[31321] = 18
      "010010" when "0111101001011010", -- t[31322] = 18
      "010010" when "0111101001011011", -- t[31323] = 18
      "010010" when "0111101001011100", -- t[31324] = 18
      "010010" when "0111101001011101", -- t[31325] = 18
      "010010" when "0111101001011110", -- t[31326] = 18
      "010010" when "0111101001011111", -- t[31327] = 18
      "010010" when "0111101001100000", -- t[31328] = 18
      "010010" when "0111101001100001", -- t[31329] = 18
      "010010" when "0111101001100010", -- t[31330] = 18
      "010010" when "0111101001100011", -- t[31331] = 18
      "010010" when "0111101001100100", -- t[31332] = 18
      "010010" when "0111101001100101", -- t[31333] = 18
      "010010" when "0111101001100110", -- t[31334] = 18
      "010010" when "0111101001100111", -- t[31335] = 18
      "010010" when "0111101001101000", -- t[31336] = 18
      "010010" when "0111101001101001", -- t[31337] = 18
      "010010" when "0111101001101010", -- t[31338] = 18
      "010010" when "0111101001101011", -- t[31339] = 18
      "010010" when "0111101001101100", -- t[31340] = 18
      "010010" when "0111101001101101", -- t[31341] = 18
      "010010" when "0111101001101110", -- t[31342] = 18
      "010010" when "0111101001101111", -- t[31343] = 18
      "010010" when "0111101001110000", -- t[31344] = 18
      "010010" when "0111101001110001", -- t[31345] = 18
      "010010" when "0111101001110010", -- t[31346] = 18
      "010010" when "0111101001110011", -- t[31347] = 18
      "010010" when "0111101001110100", -- t[31348] = 18
      "010010" when "0111101001110101", -- t[31349] = 18
      "010010" when "0111101001110110", -- t[31350] = 18
      "010010" when "0111101001110111", -- t[31351] = 18
      "010010" when "0111101001111000", -- t[31352] = 18
      "010010" when "0111101001111001", -- t[31353] = 18
      "010010" when "0111101001111010", -- t[31354] = 18
      "010010" when "0111101001111011", -- t[31355] = 18
      "010010" when "0111101001111100", -- t[31356] = 18
      "010010" when "0111101001111101", -- t[31357] = 18
      "010010" when "0111101001111110", -- t[31358] = 18
      "010010" when "0111101001111111", -- t[31359] = 18
      "010010" when "0111101010000000", -- t[31360] = 18
      "010010" when "0111101010000001", -- t[31361] = 18
      "010010" when "0111101010000010", -- t[31362] = 18
      "010010" when "0111101010000011", -- t[31363] = 18
      "010010" when "0111101010000100", -- t[31364] = 18
      "010010" when "0111101010000101", -- t[31365] = 18
      "010010" when "0111101010000110", -- t[31366] = 18
      "010010" when "0111101010000111", -- t[31367] = 18
      "010010" when "0111101010001000", -- t[31368] = 18
      "010010" when "0111101010001001", -- t[31369] = 18
      "010010" when "0111101010001010", -- t[31370] = 18
      "010010" when "0111101010001011", -- t[31371] = 18
      "010010" when "0111101010001100", -- t[31372] = 18
      "010010" when "0111101010001101", -- t[31373] = 18
      "010010" when "0111101010001110", -- t[31374] = 18
      "010010" when "0111101010001111", -- t[31375] = 18
      "010010" when "0111101010010000", -- t[31376] = 18
      "010010" when "0111101010010001", -- t[31377] = 18
      "010010" when "0111101010010010", -- t[31378] = 18
      "010010" when "0111101010010011", -- t[31379] = 18
      "010010" when "0111101010010100", -- t[31380] = 18
      "010010" when "0111101010010101", -- t[31381] = 18
      "010010" when "0111101010010110", -- t[31382] = 18
      "010010" when "0111101010010111", -- t[31383] = 18
      "010010" when "0111101010011000", -- t[31384] = 18
      "010010" when "0111101010011001", -- t[31385] = 18
      "010010" when "0111101010011010", -- t[31386] = 18
      "010010" when "0111101010011011", -- t[31387] = 18
      "010010" when "0111101010011100", -- t[31388] = 18
      "010010" when "0111101010011101", -- t[31389] = 18
      "010010" when "0111101010011110", -- t[31390] = 18
      "010010" when "0111101010011111", -- t[31391] = 18
      "010010" when "0111101010100000", -- t[31392] = 18
      "010010" when "0111101010100001", -- t[31393] = 18
      "010010" when "0111101010100010", -- t[31394] = 18
      "010010" when "0111101010100011", -- t[31395] = 18
      "010010" when "0111101010100100", -- t[31396] = 18
      "010010" when "0111101010100101", -- t[31397] = 18
      "010010" when "0111101010100110", -- t[31398] = 18
      "010010" when "0111101010100111", -- t[31399] = 18
      "010010" when "0111101010101000", -- t[31400] = 18
      "010010" when "0111101010101001", -- t[31401] = 18
      "010010" when "0111101010101010", -- t[31402] = 18
      "010010" when "0111101010101011", -- t[31403] = 18
      "010010" when "0111101010101100", -- t[31404] = 18
      "010010" when "0111101010101101", -- t[31405] = 18
      "010010" when "0111101010101110", -- t[31406] = 18
      "010010" when "0111101010101111", -- t[31407] = 18
      "010010" when "0111101010110000", -- t[31408] = 18
      "010010" when "0111101010110001", -- t[31409] = 18
      "010010" when "0111101010110010", -- t[31410] = 18
      "010010" when "0111101010110011", -- t[31411] = 18
      "010010" when "0111101010110100", -- t[31412] = 18
      "010010" when "0111101010110101", -- t[31413] = 18
      "010010" when "0111101010110110", -- t[31414] = 18
      "010010" when "0111101010110111", -- t[31415] = 18
      "010010" when "0111101010111000", -- t[31416] = 18
      "010010" when "0111101010111001", -- t[31417] = 18
      "010010" when "0111101010111010", -- t[31418] = 18
      "010010" when "0111101010111011", -- t[31419] = 18
      "010010" when "0111101010111100", -- t[31420] = 18
      "010010" when "0111101010111101", -- t[31421] = 18
      "010010" when "0111101010111110", -- t[31422] = 18
      "010010" when "0111101010111111", -- t[31423] = 18
      "010010" when "0111101011000000", -- t[31424] = 18
      "010010" when "0111101011000001", -- t[31425] = 18
      "010010" when "0111101011000010", -- t[31426] = 18
      "010010" when "0111101011000011", -- t[31427] = 18
      "010010" when "0111101011000100", -- t[31428] = 18
      "010010" when "0111101011000101", -- t[31429] = 18
      "010010" when "0111101011000110", -- t[31430] = 18
      "010010" when "0111101011000111", -- t[31431] = 18
      "010010" when "0111101011001000", -- t[31432] = 18
      "010010" when "0111101011001001", -- t[31433] = 18
      "010010" when "0111101011001010", -- t[31434] = 18
      "010010" when "0111101011001011", -- t[31435] = 18
      "010010" when "0111101011001100", -- t[31436] = 18
      "010010" when "0111101011001101", -- t[31437] = 18
      "010010" when "0111101011001110", -- t[31438] = 18
      "010010" when "0111101011001111", -- t[31439] = 18
      "010010" when "0111101011010000", -- t[31440] = 18
      "010010" when "0111101011010001", -- t[31441] = 18
      "010010" when "0111101011010010", -- t[31442] = 18
      "010010" when "0111101011010011", -- t[31443] = 18
      "010010" when "0111101011010100", -- t[31444] = 18
      "010010" when "0111101011010101", -- t[31445] = 18
      "010010" when "0111101011010110", -- t[31446] = 18
      "010010" when "0111101011010111", -- t[31447] = 18
      "010010" when "0111101011011000", -- t[31448] = 18
      "010010" when "0111101011011001", -- t[31449] = 18
      "010010" when "0111101011011010", -- t[31450] = 18
      "010011" when "0111101011011011", -- t[31451] = 19
      "010011" when "0111101011011100", -- t[31452] = 19
      "010011" when "0111101011011101", -- t[31453] = 19
      "010011" when "0111101011011110", -- t[31454] = 19
      "010011" when "0111101011011111", -- t[31455] = 19
      "010011" when "0111101011100000", -- t[31456] = 19
      "010011" when "0111101011100001", -- t[31457] = 19
      "010011" when "0111101011100010", -- t[31458] = 19
      "010011" when "0111101011100011", -- t[31459] = 19
      "010011" when "0111101011100100", -- t[31460] = 19
      "010011" when "0111101011100101", -- t[31461] = 19
      "010011" when "0111101011100110", -- t[31462] = 19
      "010011" when "0111101011100111", -- t[31463] = 19
      "010011" when "0111101011101000", -- t[31464] = 19
      "010011" when "0111101011101001", -- t[31465] = 19
      "010011" when "0111101011101010", -- t[31466] = 19
      "010011" when "0111101011101011", -- t[31467] = 19
      "010011" when "0111101011101100", -- t[31468] = 19
      "010011" when "0111101011101101", -- t[31469] = 19
      "010011" when "0111101011101110", -- t[31470] = 19
      "010011" when "0111101011101111", -- t[31471] = 19
      "010011" when "0111101011110000", -- t[31472] = 19
      "010011" when "0111101011110001", -- t[31473] = 19
      "010011" when "0111101011110010", -- t[31474] = 19
      "010011" when "0111101011110011", -- t[31475] = 19
      "010011" when "0111101011110100", -- t[31476] = 19
      "010011" when "0111101011110101", -- t[31477] = 19
      "010011" when "0111101011110110", -- t[31478] = 19
      "010011" when "0111101011110111", -- t[31479] = 19
      "010011" when "0111101011111000", -- t[31480] = 19
      "010011" when "0111101011111001", -- t[31481] = 19
      "010011" when "0111101011111010", -- t[31482] = 19
      "010011" when "0111101011111011", -- t[31483] = 19
      "010011" when "0111101011111100", -- t[31484] = 19
      "010011" when "0111101011111101", -- t[31485] = 19
      "010011" when "0111101011111110", -- t[31486] = 19
      "010011" when "0111101011111111", -- t[31487] = 19
      "010011" when "0111101100000000", -- t[31488] = 19
      "010011" when "0111101100000001", -- t[31489] = 19
      "010011" when "0111101100000010", -- t[31490] = 19
      "010011" when "0111101100000011", -- t[31491] = 19
      "010011" when "0111101100000100", -- t[31492] = 19
      "010011" when "0111101100000101", -- t[31493] = 19
      "010011" when "0111101100000110", -- t[31494] = 19
      "010011" when "0111101100000111", -- t[31495] = 19
      "010011" when "0111101100001000", -- t[31496] = 19
      "010011" when "0111101100001001", -- t[31497] = 19
      "010011" when "0111101100001010", -- t[31498] = 19
      "010011" when "0111101100001011", -- t[31499] = 19
      "010011" when "0111101100001100", -- t[31500] = 19
      "010011" when "0111101100001101", -- t[31501] = 19
      "010011" when "0111101100001110", -- t[31502] = 19
      "010011" when "0111101100001111", -- t[31503] = 19
      "010011" when "0111101100010000", -- t[31504] = 19
      "010011" when "0111101100010001", -- t[31505] = 19
      "010011" when "0111101100010010", -- t[31506] = 19
      "010011" when "0111101100010011", -- t[31507] = 19
      "010011" when "0111101100010100", -- t[31508] = 19
      "010011" when "0111101100010101", -- t[31509] = 19
      "010011" when "0111101100010110", -- t[31510] = 19
      "010011" when "0111101100010111", -- t[31511] = 19
      "010011" when "0111101100011000", -- t[31512] = 19
      "010011" when "0111101100011001", -- t[31513] = 19
      "010011" when "0111101100011010", -- t[31514] = 19
      "010011" when "0111101100011011", -- t[31515] = 19
      "010011" when "0111101100011100", -- t[31516] = 19
      "010011" when "0111101100011101", -- t[31517] = 19
      "010011" when "0111101100011110", -- t[31518] = 19
      "010011" when "0111101100011111", -- t[31519] = 19
      "010011" when "0111101100100000", -- t[31520] = 19
      "010011" when "0111101100100001", -- t[31521] = 19
      "010011" when "0111101100100010", -- t[31522] = 19
      "010011" when "0111101100100011", -- t[31523] = 19
      "010011" when "0111101100100100", -- t[31524] = 19
      "010011" when "0111101100100101", -- t[31525] = 19
      "010011" when "0111101100100110", -- t[31526] = 19
      "010011" when "0111101100100111", -- t[31527] = 19
      "010011" when "0111101100101000", -- t[31528] = 19
      "010011" when "0111101100101001", -- t[31529] = 19
      "010011" when "0111101100101010", -- t[31530] = 19
      "010011" when "0111101100101011", -- t[31531] = 19
      "010011" when "0111101100101100", -- t[31532] = 19
      "010011" when "0111101100101101", -- t[31533] = 19
      "010011" when "0111101100101110", -- t[31534] = 19
      "010011" when "0111101100101111", -- t[31535] = 19
      "010011" when "0111101100110000", -- t[31536] = 19
      "010011" when "0111101100110001", -- t[31537] = 19
      "010011" when "0111101100110010", -- t[31538] = 19
      "010011" when "0111101100110011", -- t[31539] = 19
      "010011" when "0111101100110100", -- t[31540] = 19
      "010011" when "0111101100110101", -- t[31541] = 19
      "010011" when "0111101100110110", -- t[31542] = 19
      "010011" when "0111101100110111", -- t[31543] = 19
      "010011" when "0111101100111000", -- t[31544] = 19
      "010011" when "0111101100111001", -- t[31545] = 19
      "010011" when "0111101100111010", -- t[31546] = 19
      "010011" when "0111101100111011", -- t[31547] = 19
      "010011" when "0111101100111100", -- t[31548] = 19
      "010011" when "0111101100111101", -- t[31549] = 19
      "010011" when "0111101100111110", -- t[31550] = 19
      "010011" when "0111101100111111", -- t[31551] = 19
      "010011" when "0111101101000000", -- t[31552] = 19
      "010011" when "0111101101000001", -- t[31553] = 19
      "010011" when "0111101101000010", -- t[31554] = 19
      "010011" when "0111101101000011", -- t[31555] = 19
      "010011" when "0111101101000100", -- t[31556] = 19
      "010011" when "0111101101000101", -- t[31557] = 19
      "010011" when "0111101101000110", -- t[31558] = 19
      "010011" when "0111101101000111", -- t[31559] = 19
      "010011" when "0111101101001000", -- t[31560] = 19
      "010011" when "0111101101001001", -- t[31561] = 19
      "010011" when "0111101101001010", -- t[31562] = 19
      "010011" when "0111101101001011", -- t[31563] = 19
      "010011" when "0111101101001100", -- t[31564] = 19
      "010011" when "0111101101001101", -- t[31565] = 19
      "010011" when "0111101101001110", -- t[31566] = 19
      "010011" when "0111101101001111", -- t[31567] = 19
      "010011" when "0111101101010000", -- t[31568] = 19
      "010011" when "0111101101010001", -- t[31569] = 19
      "010011" when "0111101101010010", -- t[31570] = 19
      "010011" when "0111101101010011", -- t[31571] = 19
      "010011" when "0111101101010100", -- t[31572] = 19
      "010011" when "0111101101010101", -- t[31573] = 19
      "010011" when "0111101101010110", -- t[31574] = 19
      "010011" when "0111101101010111", -- t[31575] = 19
      "010011" when "0111101101011000", -- t[31576] = 19
      "010011" when "0111101101011001", -- t[31577] = 19
      "010011" when "0111101101011010", -- t[31578] = 19
      "010011" when "0111101101011011", -- t[31579] = 19
      "010011" when "0111101101011100", -- t[31580] = 19
      "010011" when "0111101101011101", -- t[31581] = 19
      "010011" when "0111101101011110", -- t[31582] = 19
      "010011" when "0111101101011111", -- t[31583] = 19
      "010011" when "0111101101100000", -- t[31584] = 19
      "010011" when "0111101101100001", -- t[31585] = 19
      "010011" when "0111101101100010", -- t[31586] = 19
      "010011" when "0111101101100011", -- t[31587] = 19
      "010011" when "0111101101100100", -- t[31588] = 19
      "010011" when "0111101101100101", -- t[31589] = 19
      "010011" when "0111101101100110", -- t[31590] = 19
      "010011" when "0111101101100111", -- t[31591] = 19
      "010011" when "0111101101101000", -- t[31592] = 19
      "010011" when "0111101101101001", -- t[31593] = 19
      "010011" when "0111101101101010", -- t[31594] = 19
      "010011" when "0111101101101011", -- t[31595] = 19
      "010011" when "0111101101101100", -- t[31596] = 19
      "010011" when "0111101101101101", -- t[31597] = 19
      "010011" when "0111101101101110", -- t[31598] = 19
      "010011" when "0111101101101111", -- t[31599] = 19
      "010011" when "0111101101110000", -- t[31600] = 19
      "010011" when "0111101101110001", -- t[31601] = 19
      "010011" when "0111101101110010", -- t[31602] = 19
      "010011" when "0111101101110011", -- t[31603] = 19
      "010011" when "0111101101110100", -- t[31604] = 19
      "010011" when "0111101101110101", -- t[31605] = 19
      "010011" when "0111101101110110", -- t[31606] = 19
      "010011" when "0111101101110111", -- t[31607] = 19
      "010011" when "0111101101111000", -- t[31608] = 19
      "010011" when "0111101101111001", -- t[31609] = 19
      "010011" when "0111101101111010", -- t[31610] = 19
      "010011" when "0111101101111011", -- t[31611] = 19
      "010011" when "0111101101111100", -- t[31612] = 19
      "010011" when "0111101101111101", -- t[31613] = 19
      "010011" when "0111101101111110", -- t[31614] = 19
      "010011" when "0111101101111111", -- t[31615] = 19
      "010011" when "0111101110000000", -- t[31616] = 19
      "010011" when "0111101110000001", -- t[31617] = 19
      "010011" when "0111101110000010", -- t[31618] = 19
      "010011" when "0111101110000011", -- t[31619] = 19
      "010011" when "0111101110000100", -- t[31620] = 19
      "010011" when "0111101110000101", -- t[31621] = 19
      "010011" when "0111101110000110", -- t[31622] = 19
      "010011" when "0111101110000111", -- t[31623] = 19
      "010011" when "0111101110001000", -- t[31624] = 19
      "010011" when "0111101110001001", -- t[31625] = 19
      "010011" when "0111101110001010", -- t[31626] = 19
      "010011" when "0111101110001011", -- t[31627] = 19
      "010011" when "0111101110001100", -- t[31628] = 19
      "010011" when "0111101110001101", -- t[31629] = 19
      "010011" when "0111101110001110", -- t[31630] = 19
      "010011" when "0111101110001111", -- t[31631] = 19
      "010011" when "0111101110010000", -- t[31632] = 19
      "010011" when "0111101110010001", -- t[31633] = 19
      "010011" when "0111101110010010", -- t[31634] = 19
      "010011" when "0111101110010011", -- t[31635] = 19
      "010011" when "0111101110010100", -- t[31636] = 19
      "010011" when "0111101110010101", -- t[31637] = 19
      "010011" when "0111101110010110", -- t[31638] = 19
      "010011" when "0111101110010111", -- t[31639] = 19
      "010011" when "0111101110011000", -- t[31640] = 19
      "010011" when "0111101110011001", -- t[31641] = 19
      "010011" when "0111101110011010", -- t[31642] = 19
      "010011" when "0111101110011011", -- t[31643] = 19
      "010011" when "0111101110011100", -- t[31644] = 19
      "010011" when "0111101110011101", -- t[31645] = 19
      "010011" when "0111101110011110", -- t[31646] = 19
      "010011" when "0111101110011111", -- t[31647] = 19
      "010011" when "0111101110100000", -- t[31648] = 19
      "010011" when "0111101110100001", -- t[31649] = 19
      "010011" when "0111101110100010", -- t[31650] = 19
      "010011" when "0111101110100011", -- t[31651] = 19
      "010011" when "0111101110100100", -- t[31652] = 19
      "010011" when "0111101110100101", -- t[31653] = 19
      "010011" when "0111101110100110", -- t[31654] = 19
      "010011" when "0111101110100111", -- t[31655] = 19
      "010011" when "0111101110101000", -- t[31656] = 19
      "010011" when "0111101110101001", -- t[31657] = 19
      "010011" when "0111101110101010", -- t[31658] = 19
      "010011" when "0111101110101011", -- t[31659] = 19
      "010011" when "0111101110101100", -- t[31660] = 19
      "010011" when "0111101110101101", -- t[31661] = 19
      "010011" when "0111101110101110", -- t[31662] = 19
      "010011" when "0111101110101111", -- t[31663] = 19
      "010011" when "0111101110110000", -- t[31664] = 19
      "010011" when "0111101110110001", -- t[31665] = 19
      "010011" when "0111101110110010", -- t[31666] = 19
      "010011" when "0111101110110011", -- t[31667] = 19
      "010011" when "0111101110110100", -- t[31668] = 19
      "010011" when "0111101110110101", -- t[31669] = 19
      "010011" when "0111101110110110", -- t[31670] = 19
      "010011" when "0111101110110111", -- t[31671] = 19
      "010011" when "0111101110111000", -- t[31672] = 19
      "010011" when "0111101110111001", -- t[31673] = 19
      "010011" when "0111101110111010", -- t[31674] = 19
      "010011" when "0111101110111011", -- t[31675] = 19
      "010011" when "0111101110111100", -- t[31676] = 19
      "010011" when "0111101110111101", -- t[31677] = 19
      "010011" when "0111101110111110", -- t[31678] = 19
      "010011" when "0111101110111111", -- t[31679] = 19
      "010011" when "0111101111000000", -- t[31680] = 19
      "010011" when "0111101111000001", -- t[31681] = 19
      "010011" when "0111101111000010", -- t[31682] = 19
      "010011" when "0111101111000011", -- t[31683] = 19
      "010011" when "0111101111000100", -- t[31684] = 19
      "010011" when "0111101111000101", -- t[31685] = 19
      "010011" when "0111101111000110", -- t[31686] = 19
      "010011" when "0111101111000111", -- t[31687] = 19
      "010011" when "0111101111001000", -- t[31688] = 19
      "010011" when "0111101111001001", -- t[31689] = 19
      "010011" when "0111101111001010", -- t[31690] = 19
      "010011" when "0111101111001011", -- t[31691] = 19
      "010011" when "0111101111001100", -- t[31692] = 19
      "010011" when "0111101111001101", -- t[31693] = 19
      "010011" when "0111101111001110", -- t[31694] = 19
      "010011" when "0111101111001111", -- t[31695] = 19
      "010011" when "0111101111010000", -- t[31696] = 19
      "010011" when "0111101111010001", -- t[31697] = 19
      "010011" when "0111101111010010", -- t[31698] = 19
      "010011" when "0111101111010011", -- t[31699] = 19
      "010011" when "0111101111010100", -- t[31700] = 19
      "010011" when "0111101111010101", -- t[31701] = 19
      "010011" when "0111101111010110", -- t[31702] = 19
      "010011" when "0111101111010111", -- t[31703] = 19
      "010011" when "0111101111011000", -- t[31704] = 19
      "010011" when "0111101111011001", -- t[31705] = 19
      "010011" when "0111101111011010", -- t[31706] = 19
      "010011" when "0111101111011011", -- t[31707] = 19
      "010011" when "0111101111011100", -- t[31708] = 19
      "010011" when "0111101111011101", -- t[31709] = 19
      "010011" when "0111101111011110", -- t[31710] = 19
      "010011" when "0111101111011111", -- t[31711] = 19
      "010011" when "0111101111100000", -- t[31712] = 19
      "010011" when "0111101111100001", -- t[31713] = 19
      "010011" when "0111101111100010", -- t[31714] = 19
      "010011" when "0111101111100011", -- t[31715] = 19
      "010011" when "0111101111100100", -- t[31716] = 19
      "010011" when "0111101111100101", -- t[31717] = 19
      "010011" when "0111101111100110", -- t[31718] = 19
      "010011" when "0111101111100111", -- t[31719] = 19
      "010011" when "0111101111101000", -- t[31720] = 19
      "010011" when "0111101111101001", -- t[31721] = 19
      "010011" when "0111101111101010", -- t[31722] = 19
      "010011" when "0111101111101011", -- t[31723] = 19
      "010011" when "0111101111101100", -- t[31724] = 19
      "010011" when "0111101111101101", -- t[31725] = 19
      "010011" when "0111101111101110", -- t[31726] = 19
      "010011" when "0111101111101111", -- t[31727] = 19
      "010011" when "0111101111110000", -- t[31728] = 19
      "010011" when "0111101111110001", -- t[31729] = 19
      "010011" when "0111101111110010", -- t[31730] = 19
      "010011" when "0111101111110011", -- t[31731] = 19
      "010011" when "0111101111110100", -- t[31732] = 19
      "010011" when "0111101111110101", -- t[31733] = 19
      "010011" when "0111101111110110", -- t[31734] = 19
      "010011" when "0111101111110111", -- t[31735] = 19
      "010011" when "0111101111111000", -- t[31736] = 19
      "010011" when "0111101111111001", -- t[31737] = 19
      "010011" when "0111101111111010", -- t[31738] = 19
      "010011" when "0111101111111011", -- t[31739] = 19
      "010011" when "0111101111111100", -- t[31740] = 19
      "010011" when "0111101111111101", -- t[31741] = 19
      "010011" when "0111101111111110", -- t[31742] = 19
      "010011" when "0111101111111111", -- t[31743] = 19
      "010011" when "0111110000000000", -- t[31744] = 19
      "010011" when "0111110000000001", -- t[31745] = 19
      "010011" when "0111110000000010", -- t[31746] = 19
      "010011" when "0111110000000011", -- t[31747] = 19
      "010011" when "0111110000000100", -- t[31748] = 19
      "010011" when "0111110000000101", -- t[31749] = 19
      "010011" when "0111110000000110", -- t[31750] = 19
      "010011" when "0111110000000111", -- t[31751] = 19
      "010011" when "0111110000001000", -- t[31752] = 19
      "010011" when "0111110000001001", -- t[31753] = 19
      "010011" when "0111110000001010", -- t[31754] = 19
      "010011" when "0111110000001011", -- t[31755] = 19
      "010011" when "0111110000001100", -- t[31756] = 19
      "010011" when "0111110000001101", -- t[31757] = 19
      "010011" when "0111110000001110", -- t[31758] = 19
      "010011" when "0111110000001111", -- t[31759] = 19
      "010011" when "0111110000010000", -- t[31760] = 19
      "010011" when "0111110000010001", -- t[31761] = 19
      "010100" when "0111110000010010", -- t[31762] = 20
      "010100" when "0111110000010011", -- t[31763] = 20
      "010100" when "0111110000010100", -- t[31764] = 20
      "010100" when "0111110000010101", -- t[31765] = 20
      "010100" when "0111110000010110", -- t[31766] = 20
      "010100" when "0111110000010111", -- t[31767] = 20
      "010100" when "0111110000011000", -- t[31768] = 20
      "010100" when "0111110000011001", -- t[31769] = 20
      "010100" when "0111110000011010", -- t[31770] = 20
      "010100" when "0111110000011011", -- t[31771] = 20
      "010100" when "0111110000011100", -- t[31772] = 20
      "010100" when "0111110000011101", -- t[31773] = 20
      "010100" when "0111110000011110", -- t[31774] = 20
      "010100" when "0111110000011111", -- t[31775] = 20
      "010100" when "0111110000100000", -- t[31776] = 20
      "010100" when "0111110000100001", -- t[31777] = 20
      "010100" when "0111110000100010", -- t[31778] = 20
      "010100" when "0111110000100011", -- t[31779] = 20
      "010100" when "0111110000100100", -- t[31780] = 20
      "010100" when "0111110000100101", -- t[31781] = 20
      "010100" when "0111110000100110", -- t[31782] = 20
      "010100" when "0111110000100111", -- t[31783] = 20
      "010100" when "0111110000101000", -- t[31784] = 20
      "010100" when "0111110000101001", -- t[31785] = 20
      "010100" when "0111110000101010", -- t[31786] = 20
      "010100" when "0111110000101011", -- t[31787] = 20
      "010100" when "0111110000101100", -- t[31788] = 20
      "010100" when "0111110000101101", -- t[31789] = 20
      "010100" when "0111110000101110", -- t[31790] = 20
      "010100" when "0111110000101111", -- t[31791] = 20
      "010100" when "0111110000110000", -- t[31792] = 20
      "010100" when "0111110000110001", -- t[31793] = 20
      "010100" when "0111110000110010", -- t[31794] = 20
      "010100" when "0111110000110011", -- t[31795] = 20
      "010100" when "0111110000110100", -- t[31796] = 20
      "010100" when "0111110000110101", -- t[31797] = 20
      "010100" when "0111110000110110", -- t[31798] = 20
      "010100" when "0111110000110111", -- t[31799] = 20
      "010100" when "0111110000111000", -- t[31800] = 20
      "010100" when "0111110000111001", -- t[31801] = 20
      "010100" when "0111110000111010", -- t[31802] = 20
      "010100" when "0111110000111011", -- t[31803] = 20
      "010100" when "0111110000111100", -- t[31804] = 20
      "010100" when "0111110000111101", -- t[31805] = 20
      "010100" when "0111110000111110", -- t[31806] = 20
      "010100" when "0111110000111111", -- t[31807] = 20
      "010100" when "0111110001000000", -- t[31808] = 20
      "010100" when "0111110001000001", -- t[31809] = 20
      "010100" when "0111110001000010", -- t[31810] = 20
      "010100" when "0111110001000011", -- t[31811] = 20
      "010100" when "0111110001000100", -- t[31812] = 20
      "010100" when "0111110001000101", -- t[31813] = 20
      "010100" when "0111110001000110", -- t[31814] = 20
      "010100" when "0111110001000111", -- t[31815] = 20
      "010100" when "0111110001001000", -- t[31816] = 20
      "010100" when "0111110001001001", -- t[31817] = 20
      "010100" when "0111110001001010", -- t[31818] = 20
      "010100" when "0111110001001011", -- t[31819] = 20
      "010100" when "0111110001001100", -- t[31820] = 20
      "010100" when "0111110001001101", -- t[31821] = 20
      "010100" when "0111110001001110", -- t[31822] = 20
      "010100" when "0111110001001111", -- t[31823] = 20
      "010100" when "0111110001010000", -- t[31824] = 20
      "010100" when "0111110001010001", -- t[31825] = 20
      "010100" when "0111110001010010", -- t[31826] = 20
      "010100" when "0111110001010011", -- t[31827] = 20
      "010100" when "0111110001010100", -- t[31828] = 20
      "010100" when "0111110001010101", -- t[31829] = 20
      "010100" when "0111110001010110", -- t[31830] = 20
      "010100" when "0111110001010111", -- t[31831] = 20
      "010100" when "0111110001011000", -- t[31832] = 20
      "010100" when "0111110001011001", -- t[31833] = 20
      "010100" when "0111110001011010", -- t[31834] = 20
      "010100" when "0111110001011011", -- t[31835] = 20
      "010100" when "0111110001011100", -- t[31836] = 20
      "010100" when "0111110001011101", -- t[31837] = 20
      "010100" when "0111110001011110", -- t[31838] = 20
      "010100" when "0111110001011111", -- t[31839] = 20
      "010100" when "0111110001100000", -- t[31840] = 20
      "010100" when "0111110001100001", -- t[31841] = 20
      "010100" when "0111110001100010", -- t[31842] = 20
      "010100" when "0111110001100011", -- t[31843] = 20
      "010100" when "0111110001100100", -- t[31844] = 20
      "010100" when "0111110001100101", -- t[31845] = 20
      "010100" when "0111110001100110", -- t[31846] = 20
      "010100" when "0111110001100111", -- t[31847] = 20
      "010100" when "0111110001101000", -- t[31848] = 20
      "010100" when "0111110001101001", -- t[31849] = 20
      "010100" when "0111110001101010", -- t[31850] = 20
      "010100" when "0111110001101011", -- t[31851] = 20
      "010100" when "0111110001101100", -- t[31852] = 20
      "010100" when "0111110001101101", -- t[31853] = 20
      "010100" when "0111110001101110", -- t[31854] = 20
      "010100" when "0111110001101111", -- t[31855] = 20
      "010100" when "0111110001110000", -- t[31856] = 20
      "010100" when "0111110001110001", -- t[31857] = 20
      "010100" when "0111110001110010", -- t[31858] = 20
      "010100" when "0111110001110011", -- t[31859] = 20
      "010100" when "0111110001110100", -- t[31860] = 20
      "010100" when "0111110001110101", -- t[31861] = 20
      "010100" when "0111110001110110", -- t[31862] = 20
      "010100" when "0111110001110111", -- t[31863] = 20
      "010100" when "0111110001111000", -- t[31864] = 20
      "010100" when "0111110001111001", -- t[31865] = 20
      "010100" when "0111110001111010", -- t[31866] = 20
      "010100" when "0111110001111011", -- t[31867] = 20
      "010100" when "0111110001111100", -- t[31868] = 20
      "010100" when "0111110001111101", -- t[31869] = 20
      "010100" when "0111110001111110", -- t[31870] = 20
      "010100" when "0111110001111111", -- t[31871] = 20
      "010100" when "0111110010000000", -- t[31872] = 20
      "010100" when "0111110010000001", -- t[31873] = 20
      "010100" when "0111110010000010", -- t[31874] = 20
      "010100" when "0111110010000011", -- t[31875] = 20
      "010100" when "0111110010000100", -- t[31876] = 20
      "010100" when "0111110010000101", -- t[31877] = 20
      "010100" when "0111110010000110", -- t[31878] = 20
      "010100" when "0111110010000111", -- t[31879] = 20
      "010100" when "0111110010001000", -- t[31880] = 20
      "010100" when "0111110010001001", -- t[31881] = 20
      "010100" when "0111110010001010", -- t[31882] = 20
      "010100" when "0111110010001011", -- t[31883] = 20
      "010100" when "0111110010001100", -- t[31884] = 20
      "010100" when "0111110010001101", -- t[31885] = 20
      "010100" when "0111110010001110", -- t[31886] = 20
      "010100" when "0111110010001111", -- t[31887] = 20
      "010100" when "0111110010010000", -- t[31888] = 20
      "010100" when "0111110010010001", -- t[31889] = 20
      "010100" when "0111110010010010", -- t[31890] = 20
      "010100" when "0111110010010011", -- t[31891] = 20
      "010100" when "0111110010010100", -- t[31892] = 20
      "010100" when "0111110010010101", -- t[31893] = 20
      "010100" when "0111110010010110", -- t[31894] = 20
      "010100" when "0111110010010111", -- t[31895] = 20
      "010100" when "0111110010011000", -- t[31896] = 20
      "010100" when "0111110010011001", -- t[31897] = 20
      "010100" when "0111110010011010", -- t[31898] = 20
      "010100" when "0111110010011011", -- t[31899] = 20
      "010100" when "0111110010011100", -- t[31900] = 20
      "010100" when "0111110010011101", -- t[31901] = 20
      "010100" when "0111110010011110", -- t[31902] = 20
      "010100" when "0111110010011111", -- t[31903] = 20
      "010100" when "0111110010100000", -- t[31904] = 20
      "010100" when "0111110010100001", -- t[31905] = 20
      "010100" when "0111110010100010", -- t[31906] = 20
      "010100" when "0111110010100011", -- t[31907] = 20
      "010100" when "0111110010100100", -- t[31908] = 20
      "010100" when "0111110010100101", -- t[31909] = 20
      "010100" when "0111110010100110", -- t[31910] = 20
      "010100" when "0111110010100111", -- t[31911] = 20
      "010100" when "0111110010101000", -- t[31912] = 20
      "010100" when "0111110010101001", -- t[31913] = 20
      "010100" when "0111110010101010", -- t[31914] = 20
      "010100" when "0111110010101011", -- t[31915] = 20
      "010100" when "0111110010101100", -- t[31916] = 20
      "010100" when "0111110010101101", -- t[31917] = 20
      "010100" when "0111110010101110", -- t[31918] = 20
      "010100" when "0111110010101111", -- t[31919] = 20
      "010100" when "0111110010110000", -- t[31920] = 20
      "010100" when "0111110010110001", -- t[31921] = 20
      "010100" when "0111110010110010", -- t[31922] = 20
      "010100" when "0111110010110011", -- t[31923] = 20
      "010100" when "0111110010110100", -- t[31924] = 20
      "010100" when "0111110010110101", -- t[31925] = 20
      "010100" when "0111110010110110", -- t[31926] = 20
      "010100" when "0111110010110111", -- t[31927] = 20
      "010100" when "0111110010111000", -- t[31928] = 20
      "010100" when "0111110010111001", -- t[31929] = 20
      "010100" when "0111110010111010", -- t[31930] = 20
      "010100" when "0111110010111011", -- t[31931] = 20
      "010100" when "0111110010111100", -- t[31932] = 20
      "010100" when "0111110010111101", -- t[31933] = 20
      "010100" when "0111110010111110", -- t[31934] = 20
      "010100" when "0111110010111111", -- t[31935] = 20
      "010100" when "0111110011000000", -- t[31936] = 20
      "010100" when "0111110011000001", -- t[31937] = 20
      "010100" when "0111110011000010", -- t[31938] = 20
      "010100" when "0111110011000011", -- t[31939] = 20
      "010100" when "0111110011000100", -- t[31940] = 20
      "010100" when "0111110011000101", -- t[31941] = 20
      "010100" when "0111110011000110", -- t[31942] = 20
      "010100" when "0111110011000111", -- t[31943] = 20
      "010100" when "0111110011001000", -- t[31944] = 20
      "010100" when "0111110011001001", -- t[31945] = 20
      "010100" when "0111110011001010", -- t[31946] = 20
      "010100" when "0111110011001011", -- t[31947] = 20
      "010100" when "0111110011001100", -- t[31948] = 20
      "010100" when "0111110011001101", -- t[31949] = 20
      "010100" when "0111110011001110", -- t[31950] = 20
      "010100" when "0111110011001111", -- t[31951] = 20
      "010100" when "0111110011010000", -- t[31952] = 20
      "010100" when "0111110011010001", -- t[31953] = 20
      "010100" when "0111110011010010", -- t[31954] = 20
      "010100" when "0111110011010011", -- t[31955] = 20
      "010100" when "0111110011010100", -- t[31956] = 20
      "010100" when "0111110011010101", -- t[31957] = 20
      "010100" when "0111110011010110", -- t[31958] = 20
      "010100" when "0111110011010111", -- t[31959] = 20
      "010100" when "0111110011011000", -- t[31960] = 20
      "010100" when "0111110011011001", -- t[31961] = 20
      "010100" when "0111110011011010", -- t[31962] = 20
      "010100" when "0111110011011011", -- t[31963] = 20
      "010100" when "0111110011011100", -- t[31964] = 20
      "010100" when "0111110011011101", -- t[31965] = 20
      "010100" when "0111110011011110", -- t[31966] = 20
      "010100" when "0111110011011111", -- t[31967] = 20
      "010100" when "0111110011100000", -- t[31968] = 20
      "010100" when "0111110011100001", -- t[31969] = 20
      "010100" when "0111110011100010", -- t[31970] = 20
      "010100" when "0111110011100011", -- t[31971] = 20
      "010100" when "0111110011100100", -- t[31972] = 20
      "010100" when "0111110011100101", -- t[31973] = 20
      "010100" when "0111110011100110", -- t[31974] = 20
      "010100" when "0111110011100111", -- t[31975] = 20
      "010100" when "0111110011101000", -- t[31976] = 20
      "010100" when "0111110011101001", -- t[31977] = 20
      "010100" when "0111110011101010", -- t[31978] = 20
      "010100" when "0111110011101011", -- t[31979] = 20
      "010100" when "0111110011101100", -- t[31980] = 20
      "010100" when "0111110011101101", -- t[31981] = 20
      "010100" when "0111110011101110", -- t[31982] = 20
      "010100" when "0111110011101111", -- t[31983] = 20
      "010100" when "0111110011110000", -- t[31984] = 20
      "010100" when "0111110011110001", -- t[31985] = 20
      "010100" when "0111110011110010", -- t[31986] = 20
      "010100" when "0111110011110011", -- t[31987] = 20
      "010100" when "0111110011110100", -- t[31988] = 20
      "010100" when "0111110011110101", -- t[31989] = 20
      "010100" when "0111110011110110", -- t[31990] = 20
      "010100" when "0111110011110111", -- t[31991] = 20
      "010100" when "0111110011111000", -- t[31992] = 20
      "010100" when "0111110011111001", -- t[31993] = 20
      "010100" when "0111110011111010", -- t[31994] = 20
      "010100" when "0111110011111011", -- t[31995] = 20
      "010100" when "0111110011111100", -- t[31996] = 20
      "010100" when "0111110011111101", -- t[31997] = 20
      "010100" when "0111110011111110", -- t[31998] = 20
      "010100" when "0111110011111111", -- t[31999] = 20
      "010100" when "0111110100000000", -- t[32000] = 20
      "010100" when "0111110100000001", -- t[32001] = 20
      "010100" when "0111110100000010", -- t[32002] = 20
      "010100" when "0111110100000011", -- t[32003] = 20
      "010100" when "0111110100000100", -- t[32004] = 20
      "010100" when "0111110100000101", -- t[32005] = 20
      "010100" when "0111110100000110", -- t[32006] = 20
      "010100" when "0111110100000111", -- t[32007] = 20
      "010100" when "0111110100001000", -- t[32008] = 20
      "010100" when "0111110100001001", -- t[32009] = 20
      "010100" when "0111110100001010", -- t[32010] = 20
      "010100" when "0111110100001011", -- t[32011] = 20
      "010100" when "0111110100001100", -- t[32012] = 20
      "010100" when "0111110100001101", -- t[32013] = 20
      "010100" when "0111110100001110", -- t[32014] = 20
      "010100" when "0111110100001111", -- t[32015] = 20
      "010100" when "0111110100010000", -- t[32016] = 20
      "010100" when "0111110100010001", -- t[32017] = 20
      "010100" when "0111110100010010", -- t[32018] = 20
      "010100" when "0111110100010011", -- t[32019] = 20
      "010100" when "0111110100010100", -- t[32020] = 20
      "010100" when "0111110100010101", -- t[32021] = 20
      "010100" when "0111110100010110", -- t[32022] = 20
      "010100" when "0111110100010111", -- t[32023] = 20
      "010100" when "0111110100011000", -- t[32024] = 20
      "010100" when "0111110100011001", -- t[32025] = 20
      "010100" when "0111110100011010", -- t[32026] = 20
      "010100" when "0111110100011011", -- t[32027] = 20
      "010100" when "0111110100011100", -- t[32028] = 20
      "010100" when "0111110100011101", -- t[32029] = 20
      "010100" when "0111110100011110", -- t[32030] = 20
      "010100" when "0111110100011111", -- t[32031] = 20
      "010100" when "0111110100100000", -- t[32032] = 20
      "010100" when "0111110100100001", -- t[32033] = 20
      "010100" when "0111110100100010", -- t[32034] = 20
      "010100" when "0111110100100011", -- t[32035] = 20
      "010100" when "0111110100100100", -- t[32036] = 20
      "010100" when "0111110100100101", -- t[32037] = 20
      "010100" when "0111110100100110", -- t[32038] = 20
      "010100" when "0111110100100111", -- t[32039] = 20
      "010100" when "0111110100101000", -- t[32040] = 20
      "010100" when "0111110100101001", -- t[32041] = 20
      "010100" when "0111110100101010", -- t[32042] = 20
      "010100" when "0111110100101011", -- t[32043] = 20
      "010100" when "0111110100101100", -- t[32044] = 20
      "010100" when "0111110100101101", -- t[32045] = 20
      "010100" when "0111110100101110", -- t[32046] = 20
      "010100" when "0111110100101111", -- t[32047] = 20
      "010100" when "0111110100110000", -- t[32048] = 20
      "010100" when "0111110100110001", -- t[32049] = 20
      "010100" when "0111110100110010", -- t[32050] = 20
      "010100" when "0111110100110011", -- t[32051] = 20
      "010100" when "0111110100110100", -- t[32052] = 20
      "010100" when "0111110100110101", -- t[32053] = 20
      "010100" when "0111110100110110", -- t[32054] = 20
      "010100" when "0111110100110111", -- t[32055] = 20
      "010100" when "0111110100111000", -- t[32056] = 20
      "010101" when "0111110100111001", -- t[32057] = 21
      "010101" when "0111110100111010", -- t[32058] = 21
      "010101" when "0111110100111011", -- t[32059] = 21
      "010101" when "0111110100111100", -- t[32060] = 21
      "010101" when "0111110100111101", -- t[32061] = 21
      "010101" when "0111110100111110", -- t[32062] = 21
      "010101" when "0111110100111111", -- t[32063] = 21
      "010101" when "0111110101000000", -- t[32064] = 21
      "010101" when "0111110101000001", -- t[32065] = 21
      "010101" when "0111110101000010", -- t[32066] = 21
      "010101" when "0111110101000011", -- t[32067] = 21
      "010101" when "0111110101000100", -- t[32068] = 21
      "010101" when "0111110101000101", -- t[32069] = 21
      "010101" when "0111110101000110", -- t[32070] = 21
      "010101" when "0111110101000111", -- t[32071] = 21
      "010101" when "0111110101001000", -- t[32072] = 21
      "010101" when "0111110101001001", -- t[32073] = 21
      "010101" when "0111110101001010", -- t[32074] = 21
      "010101" when "0111110101001011", -- t[32075] = 21
      "010101" when "0111110101001100", -- t[32076] = 21
      "010101" when "0111110101001101", -- t[32077] = 21
      "010101" when "0111110101001110", -- t[32078] = 21
      "010101" when "0111110101001111", -- t[32079] = 21
      "010101" when "0111110101010000", -- t[32080] = 21
      "010101" when "0111110101010001", -- t[32081] = 21
      "010101" when "0111110101010010", -- t[32082] = 21
      "010101" when "0111110101010011", -- t[32083] = 21
      "010101" when "0111110101010100", -- t[32084] = 21
      "010101" when "0111110101010101", -- t[32085] = 21
      "010101" when "0111110101010110", -- t[32086] = 21
      "010101" when "0111110101010111", -- t[32087] = 21
      "010101" when "0111110101011000", -- t[32088] = 21
      "010101" when "0111110101011001", -- t[32089] = 21
      "010101" when "0111110101011010", -- t[32090] = 21
      "010101" when "0111110101011011", -- t[32091] = 21
      "010101" when "0111110101011100", -- t[32092] = 21
      "010101" when "0111110101011101", -- t[32093] = 21
      "010101" when "0111110101011110", -- t[32094] = 21
      "010101" when "0111110101011111", -- t[32095] = 21
      "010101" when "0111110101100000", -- t[32096] = 21
      "010101" when "0111110101100001", -- t[32097] = 21
      "010101" when "0111110101100010", -- t[32098] = 21
      "010101" when "0111110101100011", -- t[32099] = 21
      "010101" when "0111110101100100", -- t[32100] = 21
      "010101" when "0111110101100101", -- t[32101] = 21
      "010101" when "0111110101100110", -- t[32102] = 21
      "010101" when "0111110101100111", -- t[32103] = 21
      "010101" when "0111110101101000", -- t[32104] = 21
      "010101" when "0111110101101001", -- t[32105] = 21
      "010101" when "0111110101101010", -- t[32106] = 21
      "010101" when "0111110101101011", -- t[32107] = 21
      "010101" when "0111110101101100", -- t[32108] = 21
      "010101" when "0111110101101101", -- t[32109] = 21
      "010101" when "0111110101101110", -- t[32110] = 21
      "010101" when "0111110101101111", -- t[32111] = 21
      "010101" when "0111110101110000", -- t[32112] = 21
      "010101" when "0111110101110001", -- t[32113] = 21
      "010101" when "0111110101110010", -- t[32114] = 21
      "010101" when "0111110101110011", -- t[32115] = 21
      "010101" when "0111110101110100", -- t[32116] = 21
      "010101" when "0111110101110101", -- t[32117] = 21
      "010101" when "0111110101110110", -- t[32118] = 21
      "010101" when "0111110101110111", -- t[32119] = 21
      "010101" when "0111110101111000", -- t[32120] = 21
      "010101" when "0111110101111001", -- t[32121] = 21
      "010101" when "0111110101111010", -- t[32122] = 21
      "010101" when "0111110101111011", -- t[32123] = 21
      "010101" when "0111110101111100", -- t[32124] = 21
      "010101" when "0111110101111101", -- t[32125] = 21
      "010101" when "0111110101111110", -- t[32126] = 21
      "010101" when "0111110101111111", -- t[32127] = 21
      "010101" when "0111110110000000", -- t[32128] = 21
      "010101" when "0111110110000001", -- t[32129] = 21
      "010101" when "0111110110000010", -- t[32130] = 21
      "010101" when "0111110110000011", -- t[32131] = 21
      "010101" when "0111110110000100", -- t[32132] = 21
      "010101" when "0111110110000101", -- t[32133] = 21
      "010101" when "0111110110000110", -- t[32134] = 21
      "010101" when "0111110110000111", -- t[32135] = 21
      "010101" when "0111110110001000", -- t[32136] = 21
      "010101" when "0111110110001001", -- t[32137] = 21
      "010101" when "0111110110001010", -- t[32138] = 21
      "010101" when "0111110110001011", -- t[32139] = 21
      "010101" when "0111110110001100", -- t[32140] = 21
      "010101" when "0111110110001101", -- t[32141] = 21
      "010101" when "0111110110001110", -- t[32142] = 21
      "010101" when "0111110110001111", -- t[32143] = 21
      "010101" when "0111110110010000", -- t[32144] = 21
      "010101" when "0111110110010001", -- t[32145] = 21
      "010101" when "0111110110010010", -- t[32146] = 21
      "010101" when "0111110110010011", -- t[32147] = 21
      "010101" when "0111110110010100", -- t[32148] = 21
      "010101" when "0111110110010101", -- t[32149] = 21
      "010101" when "0111110110010110", -- t[32150] = 21
      "010101" when "0111110110010111", -- t[32151] = 21
      "010101" when "0111110110011000", -- t[32152] = 21
      "010101" when "0111110110011001", -- t[32153] = 21
      "010101" when "0111110110011010", -- t[32154] = 21
      "010101" when "0111110110011011", -- t[32155] = 21
      "010101" when "0111110110011100", -- t[32156] = 21
      "010101" when "0111110110011101", -- t[32157] = 21
      "010101" when "0111110110011110", -- t[32158] = 21
      "010101" when "0111110110011111", -- t[32159] = 21
      "010101" when "0111110110100000", -- t[32160] = 21
      "010101" when "0111110110100001", -- t[32161] = 21
      "010101" when "0111110110100010", -- t[32162] = 21
      "010101" when "0111110110100011", -- t[32163] = 21
      "010101" when "0111110110100100", -- t[32164] = 21
      "010101" when "0111110110100101", -- t[32165] = 21
      "010101" when "0111110110100110", -- t[32166] = 21
      "010101" when "0111110110100111", -- t[32167] = 21
      "010101" when "0111110110101000", -- t[32168] = 21
      "010101" when "0111110110101001", -- t[32169] = 21
      "010101" when "0111110110101010", -- t[32170] = 21
      "010101" when "0111110110101011", -- t[32171] = 21
      "010101" when "0111110110101100", -- t[32172] = 21
      "010101" when "0111110110101101", -- t[32173] = 21
      "010101" when "0111110110101110", -- t[32174] = 21
      "010101" when "0111110110101111", -- t[32175] = 21
      "010101" when "0111110110110000", -- t[32176] = 21
      "010101" when "0111110110110001", -- t[32177] = 21
      "010101" when "0111110110110010", -- t[32178] = 21
      "010101" when "0111110110110011", -- t[32179] = 21
      "010101" when "0111110110110100", -- t[32180] = 21
      "010101" when "0111110110110101", -- t[32181] = 21
      "010101" when "0111110110110110", -- t[32182] = 21
      "010101" when "0111110110110111", -- t[32183] = 21
      "010101" when "0111110110111000", -- t[32184] = 21
      "010101" when "0111110110111001", -- t[32185] = 21
      "010101" when "0111110110111010", -- t[32186] = 21
      "010101" when "0111110110111011", -- t[32187] = 21
      "010101" when "0111110110111100", -- t[32188] = 21
      "010101" when "0111110110111101", -- t[32189] = 21
      "010101" when "0111110110111110", -- t[32190] = 21
      "010101" when "0111110110111111", -- t[32191] = 21
      "010101" when "0111110111000000", -- t[32192] = 21
      "010101" when "0111110111000001", -- t[32193] = 21
      "010101" when "0111110111000010", -- t[32194] = 21
      "010101" when "0111110111000011", -- t[32195] = 21
      "010101" when "0111110111000100", -- t[32196] = 21
      "010101" when "0111110111000101", -- t[32197] = 21
      "010101" when "0111110111000110", -- t[32198] = 21
      "010101" when "0111110111000111", -- t[32199] = 21
      "010101" when "0111110111001000", -- t[32200] = 21
      "010101" when "0111110111001001", -- t[32201] = 21
      "010101" when "0111110111001010", -- t[32202] = 21
      "010101" when "0111110111001011", -- t[32203] = 21
      "010101" when "0111110111001100", -- t[32204] = 21
      "010101" when "0111110111001101", -- t[32205] = 21
      "010101" when "0111110111001110", -- t[32206] = 21
      "010101" when "0111110111001111", -- t[32207] = 21
      "010101" when "0111110111010000", -- t[32208] = 21
      "010101" when "0111110111010001", -- t[32209] = 21
      "010101" when "0111110111010010", -- t[32210] = 21
      "010101" when "0111110111010011", -- t[32211] = 21
      "010101" when "0111110111010100", -- t[32212] = 21
      "010101" when "0111110111010101", -- t[32213] = 21
      "010101" when "0111110111010110", -- t[32214] = 21
      "010101" when "0111110111010111", -- t[32215] = 21
      "010101" when "0111110111011000", -- t[32216] = 21
      "010101" when "0111110111011001", -- t[32217] = 21
      "010101" when "0111110111011010", -- t[32218] = 21
      "010101" when "0111110111011011", -- t[32219] = 21
      "010101" when "0111110111011100", -- t[32220] = 21
      "010101" when "0111110111011101", -- t[32221] = 21
      "010101" when "0111110111011110", -- t[32222] = 21
      "010101" when "0111110111011111", -- t[32223] = 21
      "010101" when "0111110111100000", -- t[32224] = 21
      "010101" when "0111110111100001", -- t[32225] = 21
      "010101" when "0111110111100010", -- t[32226] = 21
      "010101" when "0111110111100011", -- t[32227] = 21
      "010101" when "0111110111100100", -- t[32228] = 21
      "010101" when "0111110111100101", -- t[32229] = 21
      "010101" when "0111110111100110", -- t[32230] = 21
      "010101" when "0111110111100111", -- t[32231] = 21
      "010101" when "0111110111101000", -- t[32232] = 21
      "010101" when "0111110111101001", -- t[32233] = 21
      "010101" when "0111110111101010", -- t[32234] = 21
      "010101" when "0111110111101011", -- t[32235] = 21
      "010101" when "0111110111101100", -- t[32236] = 21
      "010101" when "0111110111101101", -- t[32237] = 21
      "010101" when "0111110111101110", -- t[32238] = 21
      "010101" when "0111110111101111", -- t[32239] = 21
      "010101" when "0111110111110000", -- t[32240] = 21
      "010101" when "0111110111110001", -- t[32241] = 21
      "010101" when "0111110111110010", -- t[32242] = 21
      "010101" when "0111110111110011", -- t[32243] = 21
      "010101" when "0111110111110100", -- t[32244] = 21
      "010101" when "0111110111110101", -- t[32245] = 21
      "010101" when "0111110111110110", -- t[32246] = 21
      "010101" when "0111110111110111", -- t[32247] = 21
      "010101" when "0111110111111000", -- t[32248] = 21
      "010101" when "0111110111111001", -- t[32249] = 21
      "010101" when "0111110111111010", -- t[32250] = 21
      "010101" when "0111110111111011", -- t[32251] = 21
      "010101" when "0111110111111100", -- t[32252] = 21
      "010101" when "0111110111111101", -- t[32253] = 21
      "010101" when "0111110111111110", -- t[32254] = 21
      "010101" when "0111110111111111", -- t[32255] = 21
      "010101" when "0111111000000000", -- t[32256] = 21
      "010101" when "0111111000000001", -- t[32257] = 21
      "010101" when "0111111000000010", -- t[32258] = 21
      "010101" when "0111111000000011", -- t[32259] = 21
      "010101" when "0111111000000100", -- t[32260] = 21
      "010101" when "0111111000000101", -- t[32261] = 21
      "010101" when "0111111000000110", -- t[32262] = 21
      "010101" when "0111111000000111", -- t[32263] = 21
      "010101" when "0111111000001000", -- t[32264] = 21
      "010101" when "0111111000001001", -- t[32265] = 21
      "010101" when "0111111000001010", -- t[32266] = 21
      "010101" when "0111111000001011", -- t[32267] = 21
      "010101" when "0111111000001100", -- t[32268] = 21
      "010101" when "0111111000001101", -- t[32269] = 21
      "010101" when "0111111000001110", -- t[32270] = 21
      "010101" when "0111111000001111", -- t[32271] = 21
      "010101" when "0111111000010000", -- t[32272] = 21
      "010101" when "0111111000010001", -- t[32273] = 21
      "010101" when "0111111000010010", -- t[32274] = 21
      "010101" when "0111111000010011", -- t[32275] = 21
      "010101" when "0111111000010100", -- t[32276] = 21
      "010101" when "0111111000010101", -- t[32277] = 21
      "010101" when "0111111000010110", -- t[32278] = 21
      "010101" when "0111111000010111", -- t[32279] = 21
      "010101" when "0111111000011000", -- t[32280] = 21
      "010101" when "0111111000011001", -- t[32281] = 21
      "010101" when "0111111000011010", -- t[32282] = 21
      "010101" when "0111111000011011", -- t[32283] = 21
      "010101" when "0111111000011100", -- t[32284] = 21
      "010101" when "0111111000011101", -- t[32285] = 21
      "010101" when "0111111000011110", -- t[32286] = 21
      "010101" when "0111111000011111", -- t[32287] = 21
      "010101" when "0111111000100000", -- t[32288] = 21
      "010101" when "0111111000100001", -- t[32289] = 21
      "010101" when "0111111000100010", -- t[32290] = 21
      "010101" when "0111111000100011", -- t[32291] = 21
      "010101" when "0111111000100100", -- t[32292] = 21
      "010101" when "0111111000100101", -- t[32293] = 21
      "010101" when "0111111000100110", -- t[32294] = 21
      "010101" when "0111111000100111", -- t[32295] = 21
      "010101" when "0111111000101000", -- t[32296] = 21
      "010101" when "0111111000101001", -- t[32297] = 21
      "010101" when "0111111000101010", -- t[32298] = 21
      "010101" when "0111111000101011", -- t[32299] = 21
      "010101" when "0111111000101100", -- t[32300] = 21
      "010101" when "0111111000101101", -- t[32301] = 21
      "010101" when "0111111000101110", -- t[32302] = 21
      "010101" when "0111111000101111", -- t[32303] = 21
      "010101" when "0111111000110000", -- t[32304] = 21
      "010101" when "0111111000110001", -- t[32305] = 21
      "010101" when "0111111000110010", -- t[32306] = 21
      "010101" when "0111111000110011", -- t[32307] = 21
      "010101" when "0111111000110100", -- t[32308] = 21
      "010101" when "0111111000110101", -- t[32309] = 21
      "010101" when "0111111000110110", -- t[32310] = 21
      "010101" when "0111111000110111", -- t[32311] = 21
      "010101" when "0111111000111000", -- t[32312] = 21
      "010101" when "0111111000111001", -- t[32313] = 21
      "010101" when "0111111000111010", -- t[32314] = 21
      "010101" when "0111111000111011", -- t[32315] = 21
      "010101" when "0111111000111100", -- t[32316] = 21
      "010101" when "0111111000111101", -- t[32317] = 21
      "010101" when "0111111000111110", -- t[32318] = 21
      "010101" when "0111111000111111", -- t[32319] = 21
      "010101" when "0111111001000000", -- t[32320] = 21
      "010101" when "0111111001000001", -- t[32321] = 21
      "010101" when "0111111001000010", -- t[32322] = 21
      "010101" when "0111111001000011", -- t[32323] = 21
      "010101" when "0111111001000100", -- t[32324] = 21
      "010101" when "0111111001000101", -- t[32325] = 21
      "010101" when "0111111001000110", -- t[32326] = 21
      "010101" when "0111111001000111", -- t[32327] = 21
      "010101" when "0111111001001000", -- t[32328] = 21
      "010101" when "0111111001001001", -- t[32329] = 21
      "010101" when "0111111001001010", -- t[32330] = 21
      "010101" when "0111111001001011", -- t[32331] = 21
      "010101" when "0111111001001100", -- t[32332] = 21
      "010101" when "0111111001001101", -- t[32333] = 21
      "010101" when "0111111001001110", -- t[32334] = 21
      "010101" when "0111111001001111", -- t[32335] = 21
      "010101" when "0111111001010000", -- t[32336] = 21
      "010101" when "0111111001010001", -- t[32337] = 21
      "010110" when "0111111001010010", -- t[32338] = 22
      "010110" when "0111111001010011", -- t[32339] = 22
      "010110" when "0111111001010100", -- t[32340] = 22
      "010110" when "0111111001010101", -- t[32341] = 22
      "010110" when "0111111001010110", -- t[32342] = 22
      "010110" when "0111111001010111", -- t[32343] = 22
      "010110" when "0111111001011000", -- t[32344] = 22
      "010110" when "0111111001011001", -- t[32345] = 22
      "010110" when "0111111001011010", -- t[32346] = 22
      "010110" when "0111111001011011", -- t[32347] = 22
      "010110" when "0111111001011100", -- t[32348] = 22
      "010110" when "0111111001011101", -- t[32349] = 22
      "010110" when "0111111001011110", -- t[32350] = 22
      "010110" when "0111111001011111", -- t[32351] = 22
      "010110" when "0111111001100000", -- t[32352] = 22
      "010110" when "0111111001100001", -- t[32353] = 22
      "010110" when "0111111001100010", -- t[32354] = 22
      "010110" when "0111111001100011", -- t[32355] = 22
      "010110" when "0111111001100100", -- t[32356] = 22
      "010110" when "0111111001100101", -- t[32357] = 22
      "010110" when "0111111001100110", -- t[32358] = 22
      "010110" when "0111111001100111", -- t[32359] = 22
      "010110" when "0111111001101000", -- t[32360] = 22
      "010110" when "0111111001101001", -- t[32361] = 22
      "010110" when "0111111001101010", -- t[32362] = 22
      "010110" when "0111111001101011", -- t[32363] = 22
      "010110" when "0111111001101100", -- t[32364] = 22
      "010110" when "0111111001101101", -- t[32365] = 22
      "010110" when "0111111001101110", -- t[32366] = 22
      "010110" when "0111111001101111", -- t[32367] = 22
      "010110" when "0111111001110000", -- t[32368] = 22
      "010110" when "0111111001110001", -- t[32369] = 22
      "010110" when "0111111001110010", -- t[32370] = 22
      "010110" when "0111111001110011", -- t[32371] = 22
      "010110" when "0111111001110100", -- t[32372] = 22
      "010110" when "0111111001110101", -- t[32373] = 22
      "010110" when "0111111001110110", -- t[32374] = 22
      "010110" when "0111111001110111", -- t[32375] = 22
      "010110" when "0111111001111000", -- t[32376] = 22
      "010110" when "0111111001111001", -- t[32377] = 22
      "010110" when "0111111001111010", -- t[32378] = 22
      "010110" when "0111111001111011", -- t[32379] = 22
      "010110" when "0111111001111100", -- t[32380] = 22
      "010110" when "0111111001111101", -- t[32381] = 22
      "010110" when "0111111001111110", -- t[32382] = 22
      "010110" when "0111111001111111", -- t[32383] = 22
      "010110" when "0111111010000000", -- t[32384] = 22
      "010110" when "0111111010000001", -- t[32385] = 22
      "010110" when "0111111010000010", -- t[32386] = 22
      "010110" when "0111111010000011", -- t[32387] = 22
      "010110" when "0111111010000100", -- t[32388] = 22
      "010110" when "0111111010000101", -- t[32389] = 22
      "010110" when "0111111010000110", -- t[32390] = 22
      "010110" when "0111111010000111", -- t[32391] = 22
      "010110" when "0111111010001000", -- t[32392] = 22
      "010110" when "0111111010001001", -- t[32393] = 22
      "010110" when "0111111010001010", -- t[32394] = 22
      "010110" when "0111111010001011", -- t[32395] = 22
      "010110" when "0111111010001100", -- t[32396] = 22
      "010110" when "0111111010001101", -- t[32397] = 22
      "010110" when "0111111010001110", -- t[32398] = 22
      "010110" when "0111111010001111", -- t[32399] = 22
      "010110" when "0111111010010000", -- t[32400] = 22
      "010110" when "0111111010010001", -- t[32401] = 22
      "010110" when "0111111010010010", -- t[32402] = 22
      "010110" when "0111111010010011", -- t[32403] = 22
      "010110" when "0111111010010100", -- t[32404] = 22
      "010110" when "0111111010010101", -- t[32405] = 22
      "010110" when "0111111010010110", -- t[32406] = 22
      "010110" when "0111111010010111", -- t[32407] = 22
      "010110" when "0111111010011000", -- t[32408] = 22
      "010110" when "0111111010011001", -- t[32409] = 22
      "010110" when "0111111010011010", -- t[32410] = 22
      "010110" when "0111111010011011", -- t[32411] = 22
      "010110" when "0111111010011100", -- t[32412] = 22
      "010110" when "0111111010011101", -- t[32413] = 22
      "010110" when "0111111010011110", -- t[32414] = 22
      "010110" when "0111111010011111", -- t[32415] = 22
      "010110" when "0111111010100000", -- t[32416] = 22
      "010110" when "0111111010100001", -- t[32417] = 22
      "010110" when "0111111010100010", -- t[32418] = 22
      "010110" when "0111111010100011", -- t[32419] = 22
      "010110" when "0111111010100100", -- t[32420] = 22
      "010110" when "0111111010100101", -- t[32421] = 22
      "010110" when "0111111010100110", -- t[32422] = 22
      "010110" when "0111111010100111", -- t[32423] = 22
      "010110" when "0111111010101000", -- t[32424] = 22
      "010110" when "0111111010101001", -- t[32425] = 22
      "010110" when "0111111010101010", -- t[32426] = 22
      "010110" when "0111111010101011", -- t[32427] = 22
      "010110" when "0111111010101100", -- t[32428] = 22
      "010110" when "0111111010101101", -- t[32429] = 22
      "010110" when "0111111010101110", -- t[32430] = 22
      "010110" when "0111111010101111", -- t[32431] = 22
      "010110" when "0111111010110000", -- t[32432] = 22
      "010110" when "0111111010110001", -- t[32433] = 22
      "010110" when "0111111010110010", -- t[32434] = 22
      "010110" when "0111111010110011", -- t[32435] = 22
      "010110" when "0111111010110100", -- t[32436] = 22
      "010110" when "0111111010110101", -- t[32437] = 22
      "010110" when "0111111010110110", -- t[32438] = 22
      "010110" when "0111111010110111", -- t[32439] = 22
      "010110" when "0111111010111000", -- t[32440] = 22
      "010110" when "0111111010111001", -- t[32441] = 22
      "010110" when "0111111010111010", -- t[32442] = 22
      "010110" when "0111111010111011", -- t[32443] = 22
      "010110" when "0111111010111100", -- t[32444] = 22
      "010110" when "0111111010111101", -- t[32445] = 22
      "010110" when "0111111010111110", -- t[32446] = 22
      "010110" when "0111111010111111", -- t[32447] = 22
      "010110" when "0111111011000000", -- t[32448] = 22
      "010110" when "0111111011000001", -- t[32449] = 22
      "010110" when "0111111011000010", -- t[32450] = 22
      "010110" when "0111111011000011", -- t[32451] = 22
      "010110" when "0111111011000100", -- t[32452] = 22
      "010110" when "0111111011000101", -- t[32453] = 22
      "010110" when "0111111011000110", -- t[32454] = 22
      "010110" when "0111111011000111", -- t[32455] = 22
      "010110" when "0111111011001000", -- t[32456] = 22
      "010110" when "0111111011001001", -- t[32457] = 22
      "010110" when "0111111011001010", -- t[32458] = 22
      "010110" when "0111111011001011", -- t[32459] = 22
      "010110" when "0111111011001100", -- t[32460] = 22
      "010110" when "0111111011001101", -- t[32461] = 22
      "010110" when "0111111011001110", -- t[32462] = 22
      "010110" when "0111111011001111", -- t[32463] = 22
      "010110" when "0111111011010000", -- t[32464] = 22
      "010110" when "0111111011010001", -- t[32465] = 22
      "010110" when "0111111011010010", -- t[32466] = 22
      "010110" when "0111111011010011", -- t[32467] = 22
      "010110" when "0111111011010100", -- t[32468] = 22
      "010110" when "0111111011010101", -- t[32469] = 22
      "010110" when "0111111011010110", -- t[32470] = 22
      "010110" when "0111111011010111", -- t[32471] = 22
      "010110" when "0111111011011000", -- t[32472] = 22
      "010110" when "0111111011011001", -- t[32473] = 22
      "010110" when "0111111011011010", -- t[32474] = 22
      "010110" when "0111111011011011", -- t[32475] = 22
      "010110" when "0111111011011100", -- t[32476] = 22
      "010110" when "0111111011011101", -- t[32477] = 22
      "010110" when "0111111011011110", -- t[32478] = 22
      "010110" when "0111111011011111", -- t[32479] = 22
      "010110" when "0111111011100000", -- t[32480] = 22
      "010110" when "0111111011100001", -- t[32481] = 22
      "010110" when "0111111011100010", -- t[32482] = 22
      "010110" when "0111111011100011", -- t[32483] = 22
      "010110" when "0111111011100100", -- t[32484] = 22
      "010110" when "0111111011100101", -- t[32485] = 22
      "010110" when "0111111011100110", -- t[32486] = 22
      "010110" when "0111111011100111", -- t[32487] = 22
      "010110" when "0111111011101000", -- t[32488] = 22
      "010110" when "0111111011101001", -- t[32489] = 22
      "010110" when "0111111011101010", -- t[32490] = 22
      "010110" when "0111111011101011", -- t[32491] = 22
      "010110" when "0111111011101100", -- t[32492] = 22
      "010110" when "0111111011101101", -- t[32493] = 22
      "010110" when "0111111011101110", -- t[32494] = 22
      "010110" when "0111111011101111", -- t[32495] = 22
      "010110" when "0111111011110000", -- t[32496] = 22
      "010110" when "0111111011110001", -- t[32497] = 22
      "010110" when "0111111011110010", -- t[32498] = 22
      "010110" when "0111111011110011", -- t[32499] = 22
      "010110" when "0111111011110100", -- t[32500] = 22
      "010110" when "0111111011110101", -- t[32501] = 22
      "010110" when "0111111011110110", -- t[32502] = 22
      "010110" when "0111111011110111", -- t[32503] = 22
      "010110" when "0111111011111000", -- t[32504] = 22
      "010110" when "0111111011111001", -- t[32505] = 22
      "010110" when "0111111011111010", -- t[32506] = 22
      "010110" when "0111111011111011", -- t[32507] = 22
      "010110" when "0111111011111100", -- t[32508] = 22
      "010110" when "0111111011111101", -- t[32509] = 22
      "010110" when "0111111011111110", -- t[32510] = 22
      "010110" when "0111111011111111", -- t[32511] = 22
      "010110" when "0111111100000000", -- t[32512] = 22
      "010110" when "0111111100000001", -- t[32513] = 22
      "010110" when "0111111100000010", -- t[32514] = 22
      "010110" when "0111111100000011", -- t[32515] = 22
      "010110" when "0111111100000100", -- t[32516] = 22
      "010110" when "0111111100000101", -- t[32517] = 22
      "010110" when "0111111100000110", -- t[32518] = 22
      "010110" when "0111111100000111", -- t[32519] = 22
      "010110" when "0111111100001000", -- t[32520] = 22
      "010110" when "0111111100001001", -- t[32521] = 22
      "010110" when "0111111100001010", -- t[32522] = 22
      "010110" when "0111111100001011", -- t[32523] = 22
      "010110" when "0111111100001100", -- t[32524] = 22
      "010110" when "0111111100001101", -- t[32525] = 22
      "010110" when "0111111100001110", -- t[32526] = 22
      "010110" when "0111111100001111", -- t[32527] = 22
      "010110" when "0111111100010000", -- t[32528] = 22
      "010110" when "0111111100010001", -- t[32529] = 22
      "010110" when "0111111100010010", -- t[32530] = 22
      "010110" when "0111111100010011", -- t[32531] = 22
      "010110" when "0111111100010100", -- t[32532] = 22
      "010110" when "0111111100010101", -- t[32533] = 22
      "010110" when "0111111100010110", -- t[32534] = 22
      "010110" when "0111111100010111", -- t[32535] = 22
      "010110" when "0111111100011000", -- t[32536] = 22
      "010110" when "0111111100011001", -- t[32537] = 22
      "010110" when "0111111100011010", -- t[32538] = 22
      "010110" when "0111111100011011", -- t[32539] = 22
      "010110" when "0111111100011100", -- t[32540] = 22
      "010110" when "0111111100011101", -- t[32541] = 22
      "010110" when "0111111100011110", -- t[32542] = 22
      "010110" when "0111111100011111", -- t[32543] = 22
      "010110" when "0111111100100000", -- t[32544] = 22
      "010110" when "0111111100100001", -- t[32545] = 22
      "010110" when "0111111100100010", -- t[32546] = 22
      "010110" when "0111111100100011", -- t[32547] = 22
      "010110" when "0111111100100100", -- t[32548] = 22
      "010110" when "0111111100100101", -- t[32549] = 22
      "010110" when "0111111100100110", -- t[32550] = 22
      "010110" when "0111111100100111", -- t[32551] = 22
      "010110" when "0111111100101000", -- t[32552] = 22
      "010110" when "0111111100101001", -- t[32553] = 22
      "010110" when "0111111100101010", -- t[32554] = 22
      "010110" when "0111111100101011", -- t[32555] = 22
      "010110" when "0111111100101100", -- t[32556] = 22
      "010110" when "0111111100101101", -- t[32557] = 22
      "010110" when "0111111100101110", -- t[32558] = 22
      "010110" when "0111111100101111", -- t[32559] = 22
      "010110" when "0111111100110000", -- t[32560] = 22
      "010110" when "0111111100110001", -- t[32561] = 22
      "010110" when "0111111100110010", -- t[32562] = 22
      "010110" when "0111111100110011", -- t[32563] = 22
      "010110" when "0111111100110100", -- t[32564] = 22
      "010110" when "0111111100110101", -- t[32565] = 22
      "010110" when "0111111100110110", -- t[32566] = 22
      "010110" when "0111111100110111", -- t[32567] = 22
      "010110" when "0111111100111000", -- t[32568] = 22
      "010110" when "0111111100111001", -- t[32569] = 22
      "010110" when "0111111100111010", -- t[32570] = 22
      "010110" when "0111111100111011", -- t[32571] = 22
      "010110" when "0111111100111100", -- t[32572] = 22
      "010110" when "0111111100111101", -- t[32573] = 22
      "010110" when "0111111100111110", -- t[32574] = 22
      "010110" when "0111111100111111", -- t[32575] = 22
      "010110" when "0111111101000000", -- t[32576] = 22
      "010110" when "0111111101000001", -- t[32577] = 22
      "010110" when "0111111101000010", -- t[32578] = 22
      "010110" when "0111111101000011", -- t[32579] = 22
      "010110" when "0111111101000100", -- t[32580] = 22
      "010110" when "0111111101000101", -- t[32581] = 22
      "010110" when "0111111101000110", -- t[32582] = 22
      "010110" when "0111111101000111", -- t[32583] = 22
      "010110" when "0111111101001000", -- t[32584] = 22
      "010110" when "0111111101001001", -- t[32585] = 22
      "010110" when "0111111101001010", -- t[32586] = 22
      "010110" when "0111111101001011", -- t[32587] = 22
      "010110" when "0111111101001100", -- t[32588] = 22
      "010110" when "0111111101001101", -- t[32589] = 22
      "010110" when "0111111101001110", -- t[32590] = 22
      "010110" when "0111111101001111", -- t[32591] = 22
      "010110" when "0111111101010000", -- t[32592] = 22
      "010110" when "0111111101010001", -- t[32593] = 22
      "010110" when "0111111101010010", -- t[32594] = 22
      "010110" when "0111111101010011", -- t[32595] = 22
      "010110" when "0111111101010100", -- t[32596] = 22
      "010110" when "0111111101010101", -- t[32597] = 22
      "010110" when "0111111101010110", -- t[32598] = 22
      "010110" when "0111111101010111", -- t[32599] = 22
      "010110" when "0111111101011000", -- t[32600] = 22
      "010110" when "0111111101011001", -- t[32601] = 22
      "010110" when "0111111101011010", -- t[32602] = 22
      "010110" when "0111111101011011", -- t[32603] = 22
      "010110" when "0111111101011100", -- t[32604] = 22
      "010110" when "0111111101011101", -- t[32605] = 22
      "010111" when "0111111101011110", -- t[32606] = 23
      "010111" when "0111111101011111", -- t[32607] = 23
      "010111" when "0111111101100000", -- t[32608] = 23
      "010111" when "0111111101100001", -- t[32609] = 23
      "010111" when "0111111101100010", -- t[32610] = 23
      "010111" when "0111111101100011", -- t[32611] = 23
      "010111" when "0111111101100100", -- t[32612] = 23
      "010111" when "0111111101100101", -- t[32613] = 23
      "010111" when "0111111101100110", -- t[32614] = 23
      "010111" when "0111111101100111", -- t[32615] = 23
      "010111" when "0111111101101000", -- t[32616] = 23
      "010111" when "0111111101101001", -- t[32617] = 23
      "010111" when "0111111101101010", -- t[32618] = 23
      "010111" when "0111111101101011", -- t[32619] = 23
      "010111" when "0111111101101100", -- t[32620] = 23
      "010111" when "0111111101101101", -- t[32621] = 23
      "010111" when "0111111101101110", -- t[32622] = 23
      "010111" when "0111111101101111", -- t[32623] = 23
      "010111" when "0111111101110000", -- t[32624] = 23
      "010111" when "0111111101110001", -- t[32625] = 23
      "010111" when "0111111101110010", -- t[32626] = 23
      "010111" when "0111111101110011", -- t[32627] = 23
      "010111" when "0111111101110100", -- t[32628] = 23
      "010111" when "0111111101110101", -- t[32629] = 23
      "010111" when "0111111101110110", -- t[32630] = 23
      "010111" when "0111111101110111", -- t[32631] = 23
      "010111" when "0111111101111000", -- t[32632] = 23
      "010111" when "0111111101111001", -- t[32633] = 23
      "010111" when "0111111101111010", -- t[32634] = 23
      "010111" when "0111111101111011", -- t[32635] = 23
      "010111" when "0111111101111100", -- t[32636] = 23
      "010111" when "0111111101111101", -- t[32637] = 23
      "010111" when "0111111101111110", -- t[32638] = 23
      "010111" when "0111111101111111", -- t[32639] = 23
      "010111" when "0111111110000000", -- t[32640] = 23
      "010111" when "0111111110000001", -- t[32641] = 23
      "010111" when "0111111110000010", -- t[32642] = 23
      "010111" when "0111111110000011", -- t[32643] = 23
      "010111" when "0111111110000100", -- t[32644] = 23
      "010111" when "0111111110000101", -- t[32645] = 23
      "010111" when "0111111110000110", -- t[32646] = 23
      "010111" when "0111111110000111", -- t[32647] = 23
      "010111" when "0111111110001000", -- t[32648] = 23
      "010111" when "0111111110001001", -- t[32649] = 23
      "010111" when "0111111110001010", -- t[32650] = 23
      "010111" when "0111111110001011", -- t[32651] = 23
      "010111" when "0111111110001100", -- t[32652] = 23
      "010111" when "0111111110001101", -- t[32653] = 23
      "010111" when "0111111110001110", -- t[32654] = 23
      "010111" when "0111111110001111", -- t[32655] = 23
      "010111" when "0111111110010000", -- t[32656] = 23
      "010111" when "0111111110010001", -- t[32657] = 23
      "010111" when "0111111110010010", -- t[32658] = 23
      "010111" when "0111111110010011", -- t[32659] = 23
      "010111" when "0111111110010100", -- t[32660] = 23
      "010111" when "0111111110010101", -- t[32661] = 23
      "010111" when "0111111110010110", -- t[32662] = 23
      "010111" when "0111111110010111", -- t[32663] = 23
      "010111" when "0111111110011000", -- t[32664] = 23
      "010111" when "0111111110011001", -- t[32665] = 23
      "010111" when "0111111110011010", -- t[32666] = 23
      "010111" when "0111111110011011", -- t[32667] = 23
      "010111" when "0111111110011100", -- t[32668] = 23
      "010111" when "0111111110011101", -- t[32669] = 23
      "010111" when "0111111110011110", -- t[32670] = 23
      "010111" when "0111111110011111", -- t[32671] = 23
      "010111" when "0111111110100000", -- t[32672] = 23
      "010111" when "0111111110100001", -- t[32673] = 23
      "010111" when "0111111110100010", -- t[32674] = 23
      "010111" when "0111111110100011", -- t[32675] = 23
      "010111" when "0111111110100100", -- t[32676] = 23
      "010111" when "0111111110100101", -- t[32677] = 23
      "010111" when "0111111110100110", -- t[32678] = 23
      "010111" when "0111111110100111", -- t[32679] = 23
      "010111" when "0111111110101000", -- t[32680] = 23
      "010111" when "0111111110101001", -- t[32681] = 23
      "010111" when "0111111110101010", -- t[32682] = 23
      "010111" when "0111111110101011", -- t[32683] = 23
      "010111" when "0111111110101100", -- t[32684] = 23
      "010111" when "0111111110101101", -- t[32685] = 23
      "010111" when "0111111110101110", -- t[32686] = 23
      "010111" when "0111111110101111", -- t[32687] = 23
      "010111" when "0111111110110000", -- t[32688] = 23
      "010111" when "0111111110110001", -- t[32689] = 23
      "010111" when "0111111110110010", -- t[32690] = 23
      "010111" when "0111111110110011", -- t[32691] = 23
      "010111" when "0111111110110100", -- t[32692] = 23
      "010111" when "0111111110110101", -- t[32693] = 23
      "010111" when "0111111110110110", -- t[32694] = 23
      "010111" when "0111111110110111", -- t[32695] = 23
      "010111" when "0111111110111000", -- t[32696] = 23
      "010111" when "0111111110111001", -- t[32697] = 23
      "010111" when "0111111110111010", -- t[32698] = 23
      "010111" when "0111111110111011", -- t[32699] = 23
      "010111" when "0111111110111100", -- t[32700] = 23
      "010111" when "0111111110111101", -- t[32701] = 23
      "010111" when "0111111110111110", -- t[32702] = 23
      "010111" when "0111111110111111", -- t[32703] = 23
      "010111" when "0111111111000000", -- t[32704] = 23
      "010111" when "0111111111000001", -- t[32705] = 23
      "010111" when "0111111111000010", -- t[32706] = 23
      "010111" when "0111111111000011", -- t[32707] = 23
      "010111" when "0111111111000100", -- t[32708] = 23
      "010111" when "0111111111000101", -- t[32709] = 23
      "010111" when "0111111111000110", -- t[32710] = 23
      "010111" when "0111111111000111", -- t[32711] = 23
      "010111" when "0111111111001000", -- t[32712] = 23
      "010111" when "0111111111001001", -- t[32713] = 23
      "010111" when "0111111111001010", -- t[32714] = 23
      "010111" when "0111111111001011", -- t[32715] = 23
      "010111" when "0111111111001100", -- t[32716] = 23
      "010111" when "0111111111001101", -- t[32717] = 23
      "010111" when "0111111111001110", -- t[32718] = 23
      "010111" when "0111111111001111", -- t[32719] = 23
      "010111" when "0111111111010000", -- t[32720] = 23
      "010111" when "0111111111010001", -- t[32721] = 23
      "010111" when "0111111111010010", -- t[32722] = 23
      "010111" when "0111111111010011", -- t[32723] = 23
      "010111" when "0111111111010100", -- t[32724] = 23
      "010111" when "0111111111010101", -- t[32725] = 23
      "010111" when "0111111111010110", -- t[32726] = 23
      "010111" when "0111111111010111", -- t[32727] = 23
      "010111" when "0111111111011000", -- t[32728] = 23
      "010111" when "0111111111011001", -- t[32729] = 23
      "010111" when "0111111111011010", -- t[32730] = 23
      "010111" when "0111111111011011", -- t[32731] = 23
      "010111" when "0111111111011100", -- t[32732] = 23
      "010111" when "0111111111011101", -- t[32733] = 23
      "010111" when "0111111111011110", -- t[32734] = 23
      "010111" when "0111111111011111", -- t[32735] = 23
      "010111" when "0111111111100000", -- t[32736] = 23
      "010111" when "0111111111100001", -- t[32737] = 23
      "010111" when "0111111111100010", -- t[32738] = 23
      "010111" when "0111111111100011", -- t[32739] = 23
      "010111" when "0111111111100100", -- t[32740] = 23
      "010111" when "0111111111100101", -- t[32741] = 23
      "010111" when "0111111111100110", -- t[32742] = 23
      "010111" when "0111111111100111", -- t[32743] = 23
      "010111" when "0111111111101000", -- t[32744] = 23
      "010111" when "0111111111101001", -- t[32745] = 23
      "010111" when "0111111111101010", -- t[32746] = 23
      "010111" when "0111111111101011", -- t[32747] = 23
      "010111" when "0111111111101100", -- t[32748] = 23
      "010111" when "0111111111101101", -- t[32749] = 23
      "010111" when "0111111111101110", -- t[32750] = 23
      "010111" when "0111111111101111", -- t[32751] = 23
      "010111" when "0111111111110000", -- t[32752] = 23
      "010111" when "0111111111110001", -- t[32753] = 23
      "010111" when "0111111111110010", -- t[32754] = 23
      "010111" when "0111111111110011", -- t[32755] = 23
      "010111" when "0111111111110100", -- t[32756] = 23
      "010111" when "0111111111110101", -- t[32757] = 23
      "010111" when "0111111111110110", -- t[32758] = 23
      "010111" when "0111111111110111", -- t[32759] = 23
      "010111" when "0111111111111000", -- t[32760] = 23
      "010111" when "0111111111111001", -- t[32761] = 23
      "010111" when "0111111111111010", -- t[32762] = 23
      "010111" when "0111111111111011", -- t[32763] = 23
      "010111" when "0111111111111100", -- t[32764] = 23
      "010111" when "0111111111111101", -- t[32765] = 23
      "010111" when "0111111111111110", -- t[32766] = 23
      "010111" when "0111111111111111", -- t[32767] = 23
      "------" when others;
end architecture;


-- MultiPartite: LNS subtraction function: [-7.999999999999998 -4.0[ -> [0.0 0.12500000000000003[
-- wI = 14 bits
-- wO = 9 bits
-- Decomposition: 8, 6 / 7, 3 / 2, 4
-- Guard bits: 3
-- Size: 4224 = 12.2^8 + 4.2^8 + 2.2^6

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T1_12 is
  component LNSSub_MPT_T1_12_tiv is
    port( x : in  std_logic_vector(7 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T1_12_to1 is
    port( x : in  std_logic_vector(7 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T1_12_to0 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(1 downto 0) );
  end component;

  component LNSSub_MPT_T1_12_to1_xor is
    port( a : in  std_logic_vector(6 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T1_12_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_12_tiv is
  port( x : in  std_logic_vector(7 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12_tiv is
begin
  with x select
    r <=
      "000010111111" when "00000000", -- t[0] = 191
      "000011000001" when "00000001", -- t[1] = 193
      "000011000011" when "00000010", -- t[2] = 195
      "000011000101" when "00000011", -- t[3] = 197
      "000011000111" when "00000100", -- t[4] = 199
      "000011001001" when "00000101", -- t[5] = 201
      "000011001011" when "00000110", -- t[6] = 203
      "000011001101" when "00000111", -- t[7] = 205
      "000011001111" when "00001000", -- t[8] = 207
      "000011010010" when "00001001", -- t[9] = 210
      "000011010100" when "00001010", -- t[10] = 212
      "000011010110" when "00001011", -- t[11] = 214
      "000011011000" when "00001100", -- t[12] = 216
      "000011011011" when "00001101", -- t[13] = 219
      "000011011101" when "00001110", -- t[14] = 221
      "000011011111" when "00001111", -- t[15] = 223
      "000011100010" when "00010000", -- t[16] = 226
      "000011100100" when "00010001", -- t[17] = 228
      "000011100111" when "00010010", -- t[18] = 231
      "000011101001" when "00010011", -- t[19] = 233
      "000011101100" when "00010100", -- t[20] = 236
      "000011101110" when "00010101", -- t[21] = 238
      "000011110001" when "00010110", -- t[22] = 241
      "000011110011" when "00010111", -- t[23] = 243
      "000011110110" when "00011000", -- t[24] = 246
      "000011111001" when "00011001", -- t[25] = 249
      "000011111011" when "00011010", -- t[26] = 251
      "000011111110" when "00011011", -- t[27] = 254
      "000100000001" when "00011100", -- t[28] = 257
      "000100000011" when "00011101", -- t[29] = 259
      "000100000110" when "00011110", -- t[30] = 262
      "000100001001" when "00011111", -- t[31] = 265
      "000100001100" when "00100000", -- t[32] = 268
      "000100001111" when "00100001", -- t[33] = 271
      "000100010010" when "00100010", -- t[34] = 274
      "000100010101" when "00100011", -- t[35] = 277
      "000100010111" when "00100100", -- t[36] = 279
      "000100011010" when "00100101", -- t[37] = 282
      "000100011110" when "00100110", -- t[38] = 286
      "000100100001" when "00100111", -- t[39] = 289
      "000100100100" when "00101000", -- t[40] = 292
      "000100100111" when "00101001", -- t[41] = 295
      "000100101010" when "00101010", -- t[42] = 298
      "000100101101" when "00101011", -- t[43] = 301
      "000100110000" when "00101100", -- t[44] = 304
      "000100110100" when "00101101", -- t[45] = 308
      "000100110111" when "00101110", -- t[46] = 311
      "000100111010" when "00101111", -- t[47] = 314
      "000100111110" when "00110000", -- t[48] = 318
      "000101000001" when "00110001", -- t[49] = 321
      "000101000101" when "00110010", -- t[50] = 325
      "000101001000" when "00110011", -- t[51] = 328
      "000101001100" when "00110100", -- t[52] = 332
      "000101001111" when "00110101", -- t[53] = 335
      "000101010011" when "00110110", -- t[54] = 339
      "000101010111" when "00110111", -- t[55] = 343
      "000101011010" when "00111000", -- t[56] = 346
      "000101011110" when "00111001", -- t[57] = 350
      "000101100010" when "00111010", -- t[58] = 354
      "000101100110" when "00111011", -- t[59] = 358
      "000101101001" when "00111100", -- t[60] = 361
      "000101101101" when "00111101", -- t[61] = 365
      "000101110001" when "00111110", -- t[62] = 369
      "000101110101" when "00111111", -- t[63] = 373
      "000101111001" when "01000000", -- t[64] = 377
      "000101111101" when "01000001", -- t[65] = 381
      "000110000001" when "01000010", -- t[66] = 385
      "000110000110" when "01000011", -- t[67] = 390
      "000110001010" when "01000100", -- t[68] = 394
      "000110001110" when "01000101", -- t[69] = 398
      "000110010010" when "01000110", -- t[70] = 402
      "000110010111" when "01000111", -- t[71] = 407
      "000110011011" when "01001000", -- t[72] = 411
      "000110100000" when "01001001", -- t[73] = 416
      "000110100100" when "01001010", -- t[74] = 420
      "000110101001" when "01001011", -- t[75] = 425
      "000110101101" when "01001100", -- t[76] = 429
      "000110110010" when "01001101", -- t[77] = 434
      "000110110111" when "01001110", -- t[78] = 439
      "000110111011" when "01001111", -- t[79] = 443
      "000111000000" when "01010000", -- t[80] = 448
      "000111000101" when "01010001", -- t[81] = 453
      "000111001010" when "01010010", -- t[82] = 458
      "000111001111" when "01010011", -- t[83] = 463
      "000111010100" when "01010100", -- t[84] = 468
      "000111011001" when "01010101", -- t[85] = 473
      "000111011110" when "01010110", -- t[86] = 478
      "000111100011" when "01010111", -- t[87] = 483
      "000111101000" when "01011000", -- t[88] = 488
      "000111101110" when "01011001", -- t[89] = 494
      "000111110011" when "01011010", -- t[90] = 499
      "000111111001" when "01011011", -- t[91] = 505
      "000111111110" when "01011100", -- t[92] = 510
      "001000000100" when "01011101", -- t[93] = 516
      "001000001001" when "01011110", -- t[94] = 521
      "001000001111" when "01011111", -- t[95] = 527
      "001000010101" when "01100000", -- t[96] = 533
      "001000011010" when "01100001", -- t[97] = 538
      "001000100000" when "01100010", -- t[98] = 544
      "001000100110" when "01100011", -- t[99] = 550
      "001000101100" when "01100100", -- t[100] = 556
      "001000110010" when "01100101", -- t[101] = 562
      "001000111000" when "01100110", -- t[102] = 568
      "001000111110" when "01100111", -- t[103] = 574
      "001001000101" when "01101000", -- t[104] = 581
      "001001001011" when "01101001", -- t[105] = 587
      "001001010001" when "01101010", -- t[106] = 593
      "001001011000" when "01101011", -- t[107] = 600
      "001001011110" when "01101100", -- t[108] = 606
      "001001100101" when "01101101", -- t[109] = 613
      "001001101100" when "01101110", -- t[110] = 620
      "001001110010" when "01101111", -- t[111] = 626
      "001001111001" when "01110000", -- t[112] = 633
      "001010000000" when "01110001", -- t[113] = 640
      "001010000111" when "01110010", -- t[114] = 647
      "001010001110" when "01110011", -- t[115] = 654
      "001010010101" when "01110100", -- t[116] = 661
      "001010011100" when "01110101", -- t[117] = 668
      "001010100100" when "01110110", -- t[118] = 676
      "001010101011" when "01110111", -- t[119] = 683
      "001010110010" when "01111000", -- t[120] = 690
      "001010111010" when "01111001", -- t[121] = 698
      "001011000010" when "01111010", -- t[122] = 706
      "001011001001" when "01111011", -- t[123] = 713
      "001011010001" when "01111100", -- t[124] = 721
      "001011011001" when "01111101", -- t[125] = 729
      "001011100001" when "01111110", -- t[126] = 737
      "001011101001" when "01111111", -- t[127] = 745
      "001011110001" when "10000000", -- t[128] = 753
      "001011111001" when "10000001", -- t[129] = 761
      "001100000010" when "10000010", -- t[130] = 770
      "001100001010" when "10000011", -- t[131] = 778
      "001100010010" when "10000100", -- t[132] = 786
      "001100011011" when "10000101", -- t[133] = 795
      "001100100100" when "10000110", -- t[134] = 804
      "001100101100" when "10000111", -- t[135] = 812
      "001100110101" when "10001000", -- t[136] = 821
      "001100111110" when "10001001", -- t[137] = 830
      "001101000111" when "10001010", -- t[138] = 839
      "001101010001" when "10001011", -- t[139] = 849
      "001101011010" when "10001100", -- t[140] = 858
      "001101100011" when "10001101", -- t[141] = 867
      "001101101101" when "10001110", -- t[142] = 877
      "001101110110" when "10001111", -- t[143] = 886
      "001110000000" when "10010000", -- t[144] = 896
      "001110001010" when "10010001", -- t[145] = 906
      "001110010100" when "10010010", -- t[146] = 916
      "001110011110" when "10010011", -- t[147] = 926
      "001110101000" when "10010100", -- t[148] = 936
      "001110110010" when "10010101", -- t[149] = 946
      "001110111100" when "10010110", -- t[150] = 956
      "001111000111" when "10010111", -- t[151] = 967
      "001111010010" when "10011000", -- t[152] = 978
      "001111011100" when "10011001", -- t[153] = 988
      "001111100111" when "10011010", -- t[154] = 999
      "001111110010" when "10011011", -- t[155] = 1010
      "001111111101" when "10011100", -- t[156] = 1021
      "010000001000" when "10011101", -- t[157] = 1032
      "010000010100" when "10011110", -- t[158] = 1044
      "010000011111" when "10011111", -- t[159] = 1055
      "010000101011" when "10100000", -- t[160] = 1067
      "010000110110" when "10100001", -- t[161] = 1078
      "010001000010" when "10100010", -- t[162] = 1090
      "010001001110" when "10100011", -- t[163] = 1102
      "010001011010" when "10100100", -- t[164] = 1114
      "010001100110" when "10100101", -- t[165] = 1126
      "010001110011" when "10100110", -- t[166] = 1139
      "010001111111" when "10100111", -- t[167] = 1151
      "010010001100" when "10101000", -- t[168] = 1164
      "010010011001" when "10101001", -- t[169] = 1177
      "010010100110" when "10101010", -- t[170] = 1190
      "010010110011" when "10101011", -- t[171] = 1203
      "010011000000" when "10101100", -- t[172] = 1216
      "010011001101" when "10101101", -- t[173] = 1229
      "010011011011" when "10101110", -- t[174] = 1243
      "010011101000" when "10101111", -- t[175] = 1256
      "010011110110" when "10110000", -- t[176] = 1270
      "010100000100" when "10110001", -- t[177] = 1284
      "010100010010" when "10110010", -- t[178] = 1298
      "010100100001" when "10110011", -- t[179] = 1313
      "010100101111" when "10110100", -- t[180] = 1327
      "010100111110" when "10110101", -- t[181] = 1342
      "010101001100" when "10110110", -- t[182] = 1356
      "010101011011" when "10110111", -- t[183] = 1371
      "010101101010" when "10111000", -- t[184] = 1386
      "010101111010" when "10111001", -- t[185] = 1402
      "010110001001" when "10111010", -- t[186] = 1417
      "010110011001" when "10111011", -- t[187] = 1433
      "010110101001" when "10111100", -- t[188] = 1449
      "010110111001" when "10111101", -- t[189] = 1465
      "010111001001" when "10111110", -- t[190] = 1481
      "010111011001" when "10111111", -- t[191] = 1497
      "010111101010" when "11000000", -- t[192] = 1514
      "010111111010" when "11000001", -- t[193] = 1530
      "011000001011" when "11000010", -- t[194] = 1547
      "011000011100" when "11000011", -- t[195] = 1564
      "011000101110" when "11000100", -- t[196] = 1582
      "011000111111" when "11000101", -- t[197] = 1599
      "011001010001" when "11000110", -- t[198] = 1617
      "011001100010" when "11000111", -- t[199] = 1634
      "011001110101" when "11001000", -- t[200] = 1653
      "011010000111" when "11001001", -- t[201] = 1671
      "011010011001" when "11001010", -- t[202] = 1689
      "011010101100" when "11001011", -- t[203] = 1708
      "011010111111" when "11001100", -- t[204] = 1727
      "011011010010" when "11001101", -- t[205] = 1746
      "011011100101" when "11001110", -- t[206] = 1765
      "011011111001" when "11001111", -- t[207] = 1785
      "011100001101" when "11010000", -- t[208] = 1805
      "011100100001" when "11010001", -- t[209] = 1825
      "011100110101" when "11010010", -- t[210] = 1845
      "011101001001" when "11010011", -- t[211] = 1865
      "011101011110" when "11010100", -- t[212] = 1886
      "011101110011" when "11010101", -- t[213] = 1907
      "011110001000" when "11010110", -- t[214] = 1928
      "011110011101" when "11010111", -- t[215] = 1949
      "011110110011" when "11011000", -- t[216] = 1971
      "011111001001" when "11011001", -- t[217] = 1993
      "011111011111" when "11011010", -- t[218] = 2015
      "011111110101" when "11011011", -- t[219] = 2037
      "100000001100" when "11011100", -- t[220] = 2060
      "100000100011" when "11011101", -- t[221] = 2083
      "100000111010" when "11011110", -- t[222] = 2106
      "100001010001" when "11011111", -- t[223] = 2129
      "100001101001" when "11100000", -- t[224] = 2153
      "100010000001" when "11100001", -- t[225] = 2177
      "100010011001" when "11100010", -- t[226] = 2201
      "100010110010" when "11100011", -- t[227] = 2226
      "100011001010" when "11100100", -- t[228] = 2250
      "100011100100" when "11100101", -- t[229] = 2276
      "100011111101" when "11100110", -- t[230] = 2301
      "100100010110" when "11100111", -- t[231] = 2326
      "100100110000" when "11101000", -- t[232] = 2352
      "100101001011" when "11101001", -- t[233] = 2379
      "100101100101" when "11101010", -- t[234] = 2405
      "100110000000" when "11101011", -- t[235] = 2432
      "100110011011" when "11101100", -- t[236] = 2459
      "100110110111" when "11101101", -- t[237] = 2487
      "100111010010" when "11101110", -- t[238] = 2514
      "100111101110" when "11101111", -- t[239] = 2542
      "101000001011" when "11110000", -- t[240] = 2571
      "101000101000" when "11110001", -- t[241] = 2600
      "101001000101" when "11110010", -- t[242] = 2629
      "101001100010" when "11110011", -- t[243] = 2658
      "101010000000" when "11110100", -- t[244] = 2688
      "101010011110" when "11110101", -- t[245] = 2718
      "101010111100" when "11110110", -- t[246] = 2748
      "101011011011" when "11110111", -- t[247] = 2779
      "101011111010" when "11111000", -- t[248] = 2810
      "101100011010" when "11111001", -- t[249] = 2842
      "101100111001" when "11111010", -- t[250] = 2873
      "101101011010" when "11111011", -- t[251] = 2906
      "101101111010" when "11111100", -- t[252] = 2938
      "101110011011" when "11111101", -- t[253] = 2971
      "101110111101" when "11111110", -- t[254] = 3005
      "101111011110" when "11111111", -- t[255] = 3038
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_12_to1 is
  port( x : in  std_logic_vector(7 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12_to1 is
begin
  with x select
    r <=
      "0000" when "00000000", -- t[0] = 0
      "0000" when "00000001", -- t[1] = 0
      "0000" when "00000010", -- t[2] = 0
      "0000" when "00000011", -- t[3] = 0
      "0000" when "00000100", -- t[4] = 0
      "0000" when "00000101", -- t[5] = 0
      "0000" when "00000110", -- t[6] = 0
      "0000" when "00000111", -- t[7] = 0
      "0000" when "00001000", -- t[8] = 0
      "0000" when "00001001", -- t[9] = 0
      "0000" when "00001010", -- t[10] = 0
      "0000" when "00001011", -- t[11] = 0
      "0000" when "00001100", -- t[12] = 0
      "0000" when "00001101", -- t[13] = 0
      "0000" when "00001110", -- t[14] = 0
      "0000" when "00001111", -- t[15] = 0
      "0000" when "00010000", -- t[16] = 0
      "0000" when "00010001", -- t[17] = 0
      "0000" when "00010010", -- t[18] = 0
      "0000" when "00010011", -- t[19] = 0
      "0000" when "00010100", -- t[20] = 0
      "0000" when "00010101", -- t[21] = 0
      "0000" when "00010110", -- t[22] = 0
      "0000" when "00010111", -- t[23] = 0
      "0000" when "00011000", -- t[24] = 0
      "0000" when "00011001", -- t[25] = 0
      "0000" when "00011010", -- t[26] = 0
      "0001" when "00011011", -- t[27] = 1
      "0000" when "00011100", -- t[28] = 0
      "0001" when "00011101", -- t[29] = 1
      "0000" when "00011110", -- t[30] = 0
      "0001" when "00011111", -- t[31] = 1
      "0000" when "00100000", -- t[32] = 0
      "0001" when "00100001", -- t[33] = 1
      "0000" when "00100010", -- t[34] = 0
      "0001" when "00100011", -- t[35] = 1
      "0000" when "00100100", -- t[36] = 0
      "0001" when "00100101", -- t[37] = 1
      "0000" when "00100110", -- t[38] = 0
      "0001" when "00100111", -- t[39] = 1
      "0000" when "00101000", -- t[40] = 0
      "0001" when "00101001", -- t[41] = 1
      "0000" when "00101010", -- t[42] = 0
      "0001" when "00101011", -- t[43] = 1
      "0000" when "00101100", -- t[44] = 0
      "0001" when "00101101", -- t[45] = 1
      "0000" when "00101110", -- t[46] = 0
      "0001" when "00101111", -- t[47] = 1
      "0000" when "00110000", -- t[48] = 0
      "0001" when "00110001", -- t[49] = 1
      "0000" when "00110010", -- t[50] = 0
      "0001" when "00110011", -- t[51] = 1
      "0000" when "00110100", -- t[52] = 0
      "0001" when "00110101", -- t[53] = 1
      "0000" when "00110110", -- t[54] = 0
      "0001" when "00110111", -- t[55] = 1
      "0000" when "00111000", -- t[56] = 0
      "0001" when "00111001", -- t[57] = 1
      "0000" when "00111010", -- t[58] = 0
      "0001" when "00111011", -- t[59] = 1
      "0000" when "00111100", -- t[60] = 0
      "0001" when "00111101", -- t[61] = 1
      "0000" when "00111110", -- t[62] = 0
      "0001" when "00111111", -- t[63] = 1
      "0000" when "01000000", -- t[64] = 0
      "0001" when "01000001", -- t[65] = 1
      "0000" when "01000010", -- t[66] = 0
      "0001" when "01000011", -- t[67] = 1
      "0000" when "01000100", -- t[68] = 0
      "0001" when "01000101", -- t[69] = 1
      "0000" when "01000110", -- t[70] = 0
      "0001" when "01000111", -- t[71] = 1
      "0000" when "01001000", -- t[72] = 0
      "0001" when "01001001", -- t[73] = 1
      "0000" when "01001010", -- t[74] = 0
      "0001" when "01001011", -- t[75] = 1
      "0000" when "01001100", -- t[76] = 0
      "0001" when "01001101", -- t[77] = 1
      "0000" when "01001110", -- t[78] = 0
      "0001" when "01001111", -- t[79] = 1
      "0000" when "01010000", -- t[80] = 0
      "0001" when "01010001", -- t[81] = 1
      "0000" when "01010010", -- t[82] = 0
      "0001" when "01010011", -- t[83] = 1
      "0000" when "01010100", -- t[84] = 0
      "0001" when "01010101", -- t[85] = 1
      "0000" when "01010110", -- t[86] = 0
      "0001" when "01010111", -- t[87] = 1
      "0000" when "01011000", -- t[88] = 0
      "0001" when "01011001", -- t[89] = 1
      "0000" when "01011010", -- t[90] = 0
      "0010" when "01011011", -- t[91] = 2
      "0000" when "01011100", -- t[92] = 0
      "0010" when "01011101", -- t[93] = 2
      "0000" when "01011110", -- t[94] = 0
      "0010" when "01011111", -- t[95] = 2
      "0000" when "01100000", -- t[96] = 0
      "0010" when "01100001", -- t[97] = 2
      "0000" when "01100010", -- t[98] = 0
      "0010" when "01100011", -- t[99] = 2
      "0000" when "01100100", -- t[100] = 0
      "0010" when "01100101", -- t[101] = 2
      "0000" when "01100110", -- t[102] = 0
      "0010" when "01100111", -- t[103] = 2
      "0000" when "01101000", -- t[104] = 0
      "0010" when "01101001", -- t[105] = 2
      "0000" when "01101010", -- t[106] = 0
      "0010" when "01101011", -- t[107] = 2
      "0000" when "01101100", -- t[108] = 0
      "0010" when "01101101", -- t[109] = 2
      "0000" when "01101110", -- t[110] = 0
      "0010" when "01101111", -- t[111] = 2
      "0000" when "01110000", -- t[112] = 0
      "0010" when "01110001", -- t[113] = 2
      "0000" when "01110010", -- t[114] = 0
      "0010" when "01110011", -- t[115] = 2
      "0000" when "01110100", -- t[116] = 0
      "0010" when "01110101", -- t[117] = 2
      "0000" when "01110110", -- t[118] = 0
      "0010" when "01110111", -- t[119] = 2
      "0000" when "01111000", -- t[120] = 0
      "0010" when "01111001", -- t[121] = 2
      "0000" when "01111010", -- t[122] = 0
      "0010" when "01111011", -- t[123] = 2
      "0000" when "01111100", -- t[124] = 0
      "0010" when "01111101", -- t[125] = 2
      "0001" when "01111110", -- t[126] = 1
      "0011" when "01111111", -- t[127] = 3
      "0001" when "10000000", -- t[128] = 1
      "0011" when "10000001", -- t[129] = 3
      "0001" when "10000010", -- t[130] = 1
      "0011" when "10000011", -- t[131] = 3
      "0001" when "10000100", -- t[132] = 1
      "0011" when "10000101", -- t[133] = 3
      "0001" when "10000110", -- t[134] = 1
      "0011" when "10000111", -- t[135] = 3
      "0001" when "10001000", -- t[136] = 1
      "0011" when "10001001", -- t[137] = 3
      "0001" when "10001010", -- t[138] = 1
      "0011" when "10001011", -- t[139] = 3
      "0001" when "10001100", -- t[140] = 1
      "0011" when "10001101", -- t[141] = 3
      "0001" when "10001110", -- t[142] = 1
      "0011" when "10001111", -- t[143] = 3
      "0001" when "10010000", -- t[144] = 1
      "0011" when "10010001", -- t[145] = 3
      "0001" when "10010010", -- t[146] = 1
      "0011" when "10010011", -- t[147] = 3
      "0001" when "10010100", -- t[148] = 1
      "0011" when "10010101", -- t[149] = 3
      "0001" when "10010110", -- t[150] = 1
      "0011" when "10010111", -- t[151] = 3
      "0001" when "10011000", -- t[152] = 1
      "0100" when "10011001", -- t[153] = 4
      "0001" when "10011010", -- t[154] = 1
      "0100" when "10011011", -- t[155] = 4
      "0001" when "10011100", -- t[156] = 1
      "0100" when "10011101", -- t[157] = 4
      "0001" when "10011110", -- t[158] = 1
      "0100" when "10011111", -- t[159] = 4
      "0001" when "10100000", -- t[160] = 1
      "0100" when "10100001", -- t[161] = 4
      "0001" when "10100010", -- t[162] = 1
      "0100" when "10100011", -- t[163] = 4
      "0001" when "10100100", -- t[164] = 1
      "0100" when "10100101", -- t[165] = 4
      "0001" when "10100110", -- t[166] = 1
      "0100" when "10100111", -- t[167] = 4
      "0001" when "10101000", -- t[168] = 1
      "0100" when "10101001", -- t[169] = 4
      "0001" when "10101010", -- t[170] = 1
      "0100" when "10101011", -- t[171] = 4
      "0001" when "10101100", -- t[172] = 1
      "0101" when "10101101", -- t[173] = 5
      "0001" when "10101110", -- t[174] = 1
      "0101" when "10101111", -- t[175] = 5
      "0001" when "10110000", -- t[176] = 1
      "0101" when "10110001", -- t[177] = 5
      "0001" when "10110010", -- t[178] = 1
      "0101" when "10110011", -- t[179] = 5
      "0001" when "10110100", -- t[180] = 1
      "0101" when "10110101", -- t[181] = 5
      "0001" when "10110110", -- t[182] = 1
      "0101" when "10110111", -- t[183] = 5
      "0001" when "10111000", -- t[184] = 1
      "0101" when "10111001", -- t[185] = 5
      "0001" when "10111010", -- t[186] = 1
      "0101" when "10111011", -- t[187] = 5
      "0001" when "10111100", -- t[188] = 1
      "0101" when "10111101", -- t[189] = 5
      "0010" when "10111110", -- t[190] = 2
      "0110" when "10111111", -- t[191] = 6
      "0010" when "11000000", -- t[192] = 2
      "0110" when "11000001", -- t[193] = 6
      "0010" when "11000010", -- t[194] = 2
      "0110" when "11000011", -- t[195] = 6
      "0010" when "11000100", -- t[196] = 2
      "0110" when "11000101", -- t[197] = 6
      "0010" when "11000110", -- t[198] = 2
      "0110" when "11000111", -- t[199] = 6
      "0010" when "11001000", -- t[200] = 2
      "0110" when "11001001", -- t[201] = 6
      "0010" when "11001010", -- t[202] = 2
      "0110" when "11001011", -- t[203] = 6
      "0010" when "11001100", -- t[204] = 2
      "0111" when "11001101", -- t[205] = 7
      "0010" when "11001110", -- t[206] = 2
      "0111" when "11001111", -- t[207] = 7
      "0010" when "11010000", -- t[208] = 2
      "0111" when "11010001", -- t[209] = 7
      "0010" when "11010010", -- t[210] = 2
      "0111" when "11010011", -- t[211] = 7
      "0010" when "11010100", -- t[212] = 2
      "0111" when "11010101", -- t[213] = 7
      "0010" when "11010110", -- t[214] = 2
      "1000" when "11010111", -- t[215] = 8
      "0010" when "11011000", -- t[216] = 2
      "1000" when "11011001", -- t[217] = 8
      "0010" when "11011010", -- t[218] = 2
      "1000" when "11011011", -- t[219] = 8
      "0010" when "11011100", -- t[220] = 2
      "1000" when "11011101", -- t[221] = 8
      "0010" when "11011110", -- t[222] = 2
      "1000" when "11011111", -- t[223] = 8
      "0010" when "11100000", -- t[224] = 2
      "1000" when "11100001", -- t[225] = 8
      "0011" when "11100010", -- t[226] = 3
      "1001" when "11100011", -- t[227] = 9
      "0011" when "11100100", -- t[228] = 3
      "1001" when "11100101", -- t[229] = 9
      "0011" when "11100110", -- t[230] = 3
      "1001" when "11100111", -- t[231] = 9
      "0011" when "11101000", -- t[232] = 3
      "1001" when "11101001", -- t[233] = 9
      "0011" when "11101010", -- t[234] = 3
      "1010" when "11101011", -- t[235] = 10
      "0011" when "11101100", -- t[236] = 3
      "1010" when "11101101", -- t[237] = 10
      "0011" when "11101110", -- t[238] = 3
      "1010" when "11101111", -- t[239] = 10
      "0011" when "11110000", -- t[240] = 3
      "1010" when "11110001", -- t[241] = 10
      "0011" when "11110010", -- t[242] = 3
      "1011" when "11110011", -- t[243] = 11
      "0011" when "11110100", -- t[244] = 3
      "1011" when "11110101", -- t[245] = 11
      "0011" when "11110110", -- t[246] = 3
      "1011" when "11110111", -- t[247] = 11
      "0011" when "11111000", -- t[248] = 3
      "1011" when "11111001", -- t[249] = 11
      "0100" when "11111010", -- t[250] = 4
      "1100" when "11111011", -- t[251] = 12
      "0100" when "11111100", -- t[252] = 4
      "1100" when "11111101", -- t[253] = 12
      "0100" when "11111110", -- t[254] = 4
      "1100" when "11111111", -- t[255] = 12
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T1_12_to0 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(1 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12_to0 is
begin
  with x select
    r <=
      "00" when "000000", -- t[0] = 0
      "00" when "000001", -- t[1] = 0
      "00" when "000010", -- t[2] = 0
      "00" when "000011", -- t[3] = 0
      "00" when "000100", -- t[4] = 0
      "00" when "000101", -- t[5] = 0
      "00" when "000110", -- t[6] = 0
      "00" when "000111", -- t[7] = 0
      "00" when "001000", -- t[8] = 0
      "00" when "001001", -- t[9] = 0
      "00" when "001010", -- t[10] = 0
      "00" when "001011", -- t[11] = 0
      "00" when "001100", -- t[12] = 0
      "00" when "001101", -- t[13] = 0
      "00" when "001110", -- t[14] = 0
      "00" when "001111", -- t[15] = 0
      "00" when "010000", -- t[16] = 0
      "00" when "010001", -- t[17] = 0
      "00" when "010010", -- t[18] = 0
      "00" when "010011", -- t[19] = 0
      "00" when "010100", -- t[20] = 0
      "00" when "010101", -- t[21] = 0
      "00" when "010110", -- t[22] = 0
      "00" when "010111", -- t[23] = 0
      "00" when "011000", -- t[24] = 0
      "00" when "011001", -- t[25] = 0
      "00" when "011010", -- t[26] = 0
      "00" when "011011", -- t[27] = 0
      "00" when "011100", -- t[28] = 0
      "00" when "011101", -- t[29] = 0
      "00" when "011110", -- t[30] = 0
      "00" when "011111", -- t[31] = 0
      "00" when "100000", -- t[32] = 0
      "00" when "100001", -- t[33] = 0
      "00" when "100010", -- t[34] = 0
      "00" when "100011", -- t[35] = 0
      "00" when "100100", -- t[36] = 0
      "00" when "100101", -- t[37] = 0
      "00" when "100110", -- t[38] = 0
      "01" when "100111", -- t[39] = 1
      "00" when "101000", -- t[40] = 0
      "00" when "101001", -- t[41] = 0
      "00" when "101010", -- t[42] = 0
      "00" when "101011", -- t[43] = 0
      "00" when "101100", -- t[44] = 0
      "01" when "101101", -- t[45] = 1
      "01" when "101110", -- t[46] = 1
      "01" when "101111", -- t[47] = 1
      "00" when "110000", -- t[48] = 0
      "00" when "110001", -- t[49] = 0
      "00" when "110010", -- t[50] = 0
      "01" when "110011", -- t[51] = 1
      "01" when "110100", -- t[52] = 1
      "01" when "110101", -- t[53] = 1
      "10" when "110110", -- t[54] = 2
      "10" when "110111", -- t[55] = 2
      "00" when "111000", -- t[56] = 0
      "00" when "111001", -- t[57] = 0
      "01" when "111010", -- t[58] = 1
      "01" when "111011", -- t[59] = 1
      "10" when "111100", -- t[60] = 2
      "10" when "111101", -- t[61] = 2
      "10" when "111110", -- t[62] = 2
      "11" when "111111", -- t[63] = 3
      "--" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_12.all;

entity LNSSub_MPT_T1_12_to1_xor is
  port( a : in  std_logic_vector(6 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(7 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(7 downto 1) <= a(6 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T1_12_to1
    port map( x => in_t,
              r => out_t );

  r(11 downto 4) <= (11 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_12.all;

entity LNSSub_MPT_T1_12_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(1 downto 0);
begin
  sign <= not b(3);
  in_t(5 downto 3) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;
  in_t(2) <= b(2) xor sign;

  inst_to0 : LNSSub_MPT_T1_12_to0
    port map( x => in_t,
              r => out_t );

  r(11 downto 2) <= (11 downto 2 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_12.all;

entity LNSSub_MPT_T1_12 is
  port( x : in  std_logic_vector(13 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T1_12 is
  signal in_tiv  : std_logic_vector(7 downto 0);
  signal out_tiv : std_logic_vector(11 downto 0);
  signal a1      : std_logic_vector(6 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(11 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(3 downto 0);
  signal out0    : std_logic_vector(11 downto 0);
  signal sum     : std_logic_vector(11 downto 0);
begin
  in_tiv <= x(13 downto 6);
  inst_tiv : LNSSub_MPT_T1_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(13 downto 7);
  b1 <= x(5 downto 4);
  inst_to1_xor : LNSSub_MPT_T1_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(13 downto 11);
  b0 <= x(3 downto 0);
  inst_to0_xor : LNSSub_MPT_T1_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(11 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T1_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T1_12_Clk is
  port( x   : in  std_logic_vector(13 downto 0);
        r   : out std_logic_vector(8 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T1_12_Clk is
  signal in_tiv_1  : std_logic_vector(7 downto 0);
  signal out_tiv_1 : std_logic_vector(11 downto 0);
  signal out_tiv_2 : std_logic_vector(11 downto 0);
  signal a1_1      : std_logic_vector(6 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(11 downto 0);
  signal out1_2    : std_logic_vector(11 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(3 downto 0);
  signal out0_1    : std_logic_vector(11 downto 0);
  signal out0_2    : std_logic_vector(11 downto 0);
  signal psum1_2     : std_logic_vector(11 downto 0);
  signal psum1_3     : std_logic_vector(11 downto 0);
  signal psum2_2     : std_logic_vector(11 downto 0);
  signal psum2_3     : std_logic_vector(11 downto 0);
  signal sum_3     : std_logic_vector(11 downto 0);
begin
  in_tiv_1 <= x(13 downto 6);
  inst_tiv : LNSSub_MPT_T1_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(13 downto 7);
  b1_1 <= x(5 downto 4);
  inst_to1_xor : LNSSub_MPT_T1_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(13 downto 11);
  b0_1 <= x(3 downto 0);
  inst_to0_xor : LNSSub_MPT_T1_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(11 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-4.0 -2.0[ -> [0.0 0.5[
-- wI = 13 bits
-- wO = 11 bits
-- Decomposition: 7, 6 / 6, 4, 2 / 2, 2, 2
-- Guard bits: 2
-- Size: 2408 = 13.2^7 + 5.2^7 + 3.2^5 + 1.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T2_12 is
  component LNSSub_MPT_T2_12_tiv is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to2 is
    port( x : in  std_logic_vector(6 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to2_xor is
    port( a : in  std_logic_vector(5 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T2_12_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_12_tiv is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_tiv is
begin
  with x select
    r <=
      "0011000000001" when "0000000", -- t[0] = 1537
      "0011000010010" when "0000001", -- t[1] = 1554
      "0011000100100" when "0000010", -- t[2] = 1572
      "0011000110101" when "0000011", -- t[3] = 1589
      "0011001000111" when "0000100", -- t[4] = 1607
      "0011001011001" when "0000101", -- t[5] = 1625
      "0011001101100" when "0000110", -- t[6] = 1644
      "0011001111110" when "0000111", -- t[7] = 1662
      "0011010010001" when "0001000", -- t[8] = 1681
      "0011010100100" when "0001001", -- t[9] = 1700
      "0011010110111" when "0001010", -- t[10] = 1719
      "0011011001010" when "0001011", -- t[11] = 1738
      "0011011011110" when "0001100", -- t[12] = 1758
      "0011011110010" when "0001101", -- t[13] = 1778
      "0011100000110" when "0001110", -- t[14] = 1798
      "0011100011010" when "0001111", -- t[15] = 1818
      "0011100101111" when "0010000", -- t[16] = 1839
      "0011101000100" when "0010001", -- t[17] = 1860
      "0011101011001" when "0010010", -- t[18] = 1881
      "0011101101110" when "0010011", -- t[19] = 1902
      "0011110000011" when "0010100", -- t[20] = 1923
      "0011110011001" when "0010101", -- t[21] = 1945
      "0011110101111" when "0010110", -- t[22] = 1967
      "0011111000110" when "0010111", -- t[23] = 1990
      "0011111011100" when "0011000", -- t[24] = 2012
      "0011111110011" when "0011001", -- t[25] = 2035
      "0100000001010" when "0011010", -- t[26] = 2058
      "0100000100001" when "0011011", -- t[27] = 2081
      "0100000111001" when "0011100", -- t[28] = 2105
      "0100001010001" when "0011101", -- t[29] = 2129
      "0100001101001" when "0011110", -- t[30] = 2153
      "0100010000010" when "0011111", -- t[31] = 2178
      "0100010011011" when "0100000", -- t[32] = 2203
      "0100010110100" when "0100001", -- t[33] = 2228
      "0100011001101" when "0100010", -- t[34] = 2253
      "0100011100111" when "0100011", -- t[35] = 2279
      "0100100000001" when "0100100", -- t[36] = 2305
      "0100100011011" when "0100101", -- t[37] = 2331
      "0100100110110" when "0100110", -- t[38] = 2358
      "0100101010001" when "0100111", -- t[39] = 2385
      "0100101101100" when "0101000", -- t[40] = 2412
      "0100110001000" when "0101001", -- t[41] = 2440
      "0100110100100" when "0101010", -- t[42] = 2468
      "0100111000000" when "0101011", -- t[43] = 2496
      "0100111011101" when "0101100", -- t[44] = 2525
      "0100111111010" when "0101101", -- t[45] = 2554
      "0101000010111" when "0101110", -- t[46] = 2583
      "0101000110101" when "0101111", -- t[47] = 2613
      "0101001010011" when "0110000", -- t[48] = 2643
      "0101001110001" when "0110001", -- t[49] = 2673
      "0101010010000" when "0110010", -- t[50] = 2704
      "0101010101111" when "0110011", -- t[51] = 2735
      "0101011001111" when "0110100", -- t[52] = 2767
      "0101011101111" when "0110101", -- t[53] = 2799
      "0101100001111" when "0110110", -- t[54] = 2831
      "0101100110000" when "0110111", -- t[55] = 2864
      "0101101010001" when "0111000", -- t[56] = 2897
      "0101101110011" when "0111001", -- t[57] = 2931
      "0101110010101" when "0111010", -- t[58] = 2965
      "0101110110111" when "0111011", -- t[59] = 2999
      "0101111011010" when "0111100", -- t[60] = 3034
      "0101111111101" when "0111101", -- t[61] = 3069
      "0110000100001" when "0111110", -- t[62] = 3105
      "0110001000101" when "0111111", -- t[63] = 3141
      "0110001101001" when "1000000", -- t[64] = 3177
      "0110010001110" when "1000001", -- t[65] = 3214
      "0110010110100" when "1000010", -- t[66] = 3252
      "0110011011010" when "1000011", -- t[67] = 3290
      "0110100000000" when "1000100", -- t[68] = 3328
      "0110100100111" when "1000101", -- t[69] = 3367
      "0110101001111" when "1000110", -- t[70] = 3407
      "0110101110111" when "1000111", -- t[71] = 3447
      "0110110011111" when "1001000", -- t[72] = 3487
      "0110111001000" when "1001001", -- t[73] = 3528
      "0110111110001" when "1001010", -- t[74] = 3569
      "0111000011011" when "1001011", -- t[75] = 3611
      "0111001000110" when "1001100", -- t[76] = 3654
      "0111001110001" when "1001101", -- t[77] = 3697
      "0111010011100" when "1001110", -- t[78] = 3740
      "0111011001000" when "1001111", -- t[79] = 3784
      "0111011110101" when "1010000", -- t[80] = 3829
      "0111100100010" when "1010001", -- t[81] = 3874
      "0111101010000" when "1010010", -- t[82] = 3920
      "0111101111111" when "1010011", -- t[83] = 3967
      "0111110101110" when "1010100", -- t[84] = 4014
      "0111111011101" when "1010101", -- t[85] = 4061
      "1000000001110" when "1010110", -- t[86] = 4110
      "1000000111111" when "1010111", -- t[87] = 4159
      "1000001110000" when "1011000", -- t[88] = 4208
      "1000010100010" when "1011001", -- t[89] = 4258
      "1000011010101" when "1011010", -- t[90] = 4309
      "1000100001001" when "1011011", -- t[91] = 4361
      "1000100111101" when "1011100", -- t[92] = 4413
      "1000101110010" when "1011101", -- t[93] = 4466
      "1000110100111" when "1011110", -- t[94] = 4519
      "1000111011101" when "1011111", -- t[95] = 4573
      "1001000010100" when "1100000", -- t[96] = 4628
      "1001001001100" when "1100001", -- t[97] = 4684
      "1001010000100" when "1100010", -- t[98] = 4740
      "1001010111110" when "1100011", -- t[99] = 4798
      "1001011111000" when "1100100", -- t[100] = 4856
      "1001100110010" when "1100101", -- t[101] = 4914
      "1001101101110" when "1100110", -- t[102] = 4974
      "1001110101010" when "1100111", -- t[103] = 5034
      "1001111100111" when "1101000", -- t[104] = 5095
      "1010000100101" when "1101001", -- t[105] = 5157
      "1010001100100" when "1101010", -- t[106] = 5220
      "1010010100100" when "1101011", -- t[107] = 5284
      "1010011100100" when "1101100", -- t[108] = 5348
      "1010100100110" when "1101101", -- t[109] = 5414
      "1010101101000" when "1101110", -- t[110] = 5480
      "1010110101011" when "1101111", -- t[111] = 5547
      "1010111101111" when "1110000", -- t[112] = 5615
      "1011000110100" when "1110001", -- t[113] = 5684
      "1011001111010" when "1110010", -- t[114] = 5754
      "1011011000001" when "1110011", -- t[115] = 5825
      "1011100001001" when "1110100", -- t[116] = 5897
      "1011101010010" when "1110101", -- t[117] = 5970
      "1011110011100" when "1110110", -- t[118] = 6044
      "1011111101000" when "1110111", -- t[119] = 6120
      "1100000110100" when "1111000", -- t[120] = 6196
      "1100010000001" when "1111001", -- t[121] = 6273
      "1100011001111" when "1111010", -- t[122] = 6351
      "1100100011111" when "1111011", -- t[123] = 6431
      "1100101101111" when "1111100", -- t[124] = 6511
      "1100111000001" when "1111101", -- t[125] = 6593
      "1101000010100" when "1111110", -- t[126] = 6676
      "1101001101000" when "1111111", -- t[127] = 6760
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_12_to2 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to2 is
begin
  with x select
    r <=
      "00010" when "0000000", -- t[0] = 2
      "00110" when "0000001", -- t[1] = 6
      "00010" when "0000010", -- t[2] = 2
      "00110" when "0000011", -- t[3] = 6
      "00010" when "0000100", -- t[4] = 2
      "00110" when "0000101", -- t[5] = 6
      "00010" when "0000110", -- t[6] = 2
      "00110" when "0000111", -- t[7] = 6
      "00010" when "0001000", -- t[8] = 2
      "00111" when "0001001", -- t[9] = 7
      "00010" when "0001010", -- t[10] = 2
      "00111" when "0001011", -- t[11] = 7
      "00010" when "0001100", -- t[12] = 2
      "00111" when "0001101", -- t[13] = 7
      "00010" when "0001110", -- t[14] = 2
      "00111" when "0001111", -- t[15] = 7
      "00010" when "0010000", -- t[16] = 2
      "00111" when "0010001", -- t[17] = 7
      "00010" when "0010010", -- t[18] = 2
      "00111" when "0010011", -- t[19] = 7
      "00010" when "0010100", -- t[20] = 2
      "01000" when "0010101", -- t[21] = 8
      "00010" when "0010110", -- t[22] = 2
      "01000" when "0010111", -- t[23] = 8
      "00010" when "0011000", -- t[24] = 2
      "01000" when "0011001", -- t[25] = 8
      "00010" when "0011010", -- t[26] = 2
      "01000" when "0011011", -- t[27] = 8
      "00010" when "0011100", -- t[28] = 2
      "01000" when "0011101", -- t[29] = 8
      "00011" when "0011110", -- t[30] = 3
      "01001" when "0011111", -- t[31] = 9
      "00011" when "0100000", -- t[32] = 3
      "01001" when "0100001", -- t[33] = 9
      "00011" when "0100010", -- t[34] = 3
      "01001" when "0100011", -- t[35] = 9
      "00011" when "0100100", -- t[36] = 3
      "01001" when "0100101", -- t[37] = 9
      "00011" when "0100110", -- t[38] = 3
      "01010" when "0100111", -- t[39] = 10
      "00011" when "0101000", -- t[40] = 3
      "01010" when "0101001", -- t[41] = 10
      "00011" when "0101010", -- t[42] = 3
      "01010" when "0101011", -- t[43] = 10
      "00011" when "0101100", -- t[44] = 3
      "01010" when "0101101", -- t[45] = 10
      "00011" when "0101110", -- t[46] = 3
      "01011" when "0101111", -- t[47] = 11
      "00011" when "0110000", -- t[48] = 3
      "01011" when "0110001", -- t[49] = 11
      "00011" when "0110010", -- t[50] = 3
      "01011" when "0110011", -- t[51] = 11
      "00011" when "0110100", -- t[52] = 3
      "01011" when "0110101", -- t[53] = 11
      "00100" when "0110110", -- t[54] = 4
      "01100" when "0110111", -- t[55] = 12
      "00100" when "0111000", -- t[56] = 4
      "01100" when "0111001", -- t[57] = 12
      "00100" when "0111010", -- t[58] = 4
      "01100" when "0111011", -- t[59] = 12
      "00100" when "0111100", -- t[60] = 4
      "01101" when "0111101", -- t[61] = 13
      "00100" when "0111110", -- t[62] = 4
      "01101" when "0111111", -- t[63] = 13
      "00100" when "1000000", -- t[64] = 4
      "01101" when "1000001", -- t[65] = 13
      "00100" when "1000010", -- t[66] = 4
      "01110" when "1000011", -- t[67] = 14
      "00100" when "1000100", -- t[68] = 4
      "01110" when "1000101", -- t[69] = 14
      "00100" when "1000110", -- t[70] = 4
      "01110" when "1000111", -- t[71] = 14
      "00101" when "1001000", -- t[72] = 5
      "01111" when "1001001", -- t[73] = 15
      "00101" when "1001010", -- t[74] = 5
      "01111" when "1001011", -- t[75] = 15
      "00101" when "1001100", -- t[76] = 5
      "10000" when "1001101", -- t[77] = 16
      "00101" when "1001110", -- t[78] = 5
      "10000" when "1001111", -- t[79] = 16
      "00101" when "1010000", -- t[80] = 5
      "10000" when "1010001", -- t[81] = 16
      "00101" when "1010010", -- t[82] = 5
      "10001" when "1010011", -- t[83] = 17
      "00101" when "1010100", -- t[84] = 5
      "10001" when "1010101", -- t[85] = 17
      "00110" when "1010110", -- t[86] = 6
      "10010" when "1010111", -- t[87] = 18
      "00110" when "1011000", -- t[88] = 6
      "10010" when "1011001", -- t[89] = 18
      "00110" when "1011010", -- t[90] = 6
      "10011" when "1011011", -- t[91] = 19
      "00110" when "1011100", -- t[92] = 6
      "10011" when "1011101", -- t[93] = 19
      "00110" when "1011110", -- t[94] = 6
      "10100" when "1011111", -- t[95] = 20
      "00110" when "1100000", -- t[96] = 6
      "10100" when "1100001", -- t[97] = 20
      "00111" when "1100010", -- t[98] = 7
      "10101" when "1100011", -- t[99] = 21
      "00111" when "1100100", -- t[100] = 7
      "10101" when "1100101", -- t[101] = 21
      "00111" when "1100110", -- t[102] = 7
      "10110" when "1100111", -- t[103] = 22
      "00111" when "1101000", -- t[104] = 7
      "10111" when "1101001", -- t[105] = 23
      "00111" when "1101010", -- t[106] = 7
      "10111" when "1101011", -- t[107] = 23
      "01000" when "1101100", -- t[108] = 8
      "11000" when "1101101", -- t[109] = 24
      "01000" when "1101110", -- t[110] = 8
      "11001" when "1101111", -- t[111] = 25
      "01000" when "1110000", -- t[112] = 8
      "11001" when "1110001", -- t[113] = 25
      "01000" when "1110010", -- t[114] = 8
      "11010" when "1110011", -- t[115] = 26
      "01001" when "1110100", -- t[116] = 9
      "11011" when "1110101", -- t[117] = 27
      "01001" when "1110110", -- t[118] = 9
      "11100" when "1110111", -- t[119] = 28
      "01001" when "1111000", -- t[120] = 9
      "11100" when "1111001", -- t[121] = 28
      "01001" when "1111010", -- t[122] = 9
      "11101" when "1111011", -- t[123] = 29
      "01010" when "1111100", -- t[124] = 10
      "11110" when "1111101", -- t[125] = 30
      "01010" when "1111110", -- t[126] = 10
      "11111" when "1111111", -- t[127] = 31
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_12_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to1 is
begin
  with x select
    r <=
      "000" when "00000", -- t[0] = 0
      "001" when "00001", -- t[1] = 1
      "000" when "00010", -- t[2] = 0
      "001" when "00011", -- t[3] = 1
      "000" when "00100", -- t[4] = 0
      "010" when "00101", -- t[5] = 2
      "000" when "00110", -- t[6] = 0
      "010" when "00111", -- t[7] = 2
      "000" when "01000", -- t[8] = 0
      "010" when "01001", -- t[9] = 2
      "000" when "01010", -- t[10] = 0
      "010" when "01011", -- t[11] = 2
      "000" when "01100", -- t[12] = 0
      "010" when "01101", -- t[13] = 2
      "001" when "01110", -- t[14] = 1
      "011" when "01111", -- t[15] = 3
      "001" when "10000", -- t[16] = 1
      "011" when "10001", -- t[17] = 3
      "001" when "10010", -- t[18] = 1
      "011" when "10011", -- t[19] = 3
      "001" when "10100", -- t[20] = 1
      "100" when "10101", -- t[21] = 4
      "001" when "10110", -- t[22] = 1
      "100" when "10111", -- t[23] = 4
      "001" when "11000", -- t[24] = 1
      "101" when "11001", -- t[25] = 5
      "010" when "11010", -- t[26] = 2
      "110" when "11011", -- t[27] = 6
      "010" when "11100", -- t[28] = 2
      "110" when "11101", -- t[29] = 6
      "010" when "11110", -- t[30] = 2
      "111" when "11111", -- t[31] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T2_12_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to0 is
begin
  with x select
    r <=
      "0" when "000", -- t[0] = 0
      "0" when "001", -- t[1] = 0
      "0" when "010", -- t[2] = 0
      "0" when "011", -- t[3] = 0
      "0" when "100", -- t[4] = 0
      "1" when "101", -- t[5] = 1
      "0" when "110", -- t[6] = 0
      "1" when "111", -- t[7] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_12.all;

entity LNSSub_MPT_T2_12_to2_xor is
  port( a : in  std_logic_vector(5 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(6 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(6 downto 1) <= a(5 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T2_12_to2
    port map( x => in_t,
              r => out_t );

  r(12 downto 5) <= (12 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_12.all;

entity LNSSub_MPT_T2_12_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T2_12_to1
    port map( x => in_t,
              r => out_t );

  r(12 downto 3) <= (12 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_12.all;

entity LNSSub_MPT_T2_12_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T2_12_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 1) <= (12 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_12.all;

entity LNSSub_MPT_T2_12 is
  port( x : in  std_logic_vector(12 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T2_12 is
  signal in_tiv  : std_logic_vector(6 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a2      : std_logic_vector(5 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(12 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(12 downto 6);
  inst_tiv : LNSSub_MPT_T2_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(12 downto 7);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T2_12_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(12 downto 9);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T2_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(12 downto 11);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T2_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(12 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T2_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T2_12_Clk is
  port( x   : in  std_logic_vector(12 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T2_12_Clk is
  signal in_tiv_1  : std_logic_vector(6 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a2_1      : std_logic_vector(5 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(12 downto 0);
  signal out2_2    : std_logic_vector(12 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(12 downto 0);
  signal out1_2    : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(12 downto 6);
  inst_tiv : LNSSub_MPT_T2_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(12 downto 7);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T2_12_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(12 downto 9);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T2_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(12 downto 11);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T2_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 2);
end architecture;


-- MultiPartite: LNS subtraction function: [-2.0 -1.0[ -> [0.0 1.0[
-- wI = 12 bits
-- wO = 11 bits
-- Decomposition: 6, 6 / 5, 3, 2 / 2, 2, 2
-- Guard bits: 4
-- Size: 1600 = 15.2^6 + 8.2^6 + 6.2^4 + 4.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T3_12 is
  component LNSSub_MPT_T3_12_tiv is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to2 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(7 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to1 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(3 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to2_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to1_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T3_12_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_12_tiv is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_tiv is
begin
  with x select
    r <=
      "011010101111110" when "000000", -- t[0] = 13694
      "011011000101011" when "000001", -- t[1] = 13867
      "011011011011010" when "000010", -- t[2] = 14042
      "011011110001101" when "000011", -- t[3] = 14221
      "011100001000001" when "000100", -- t[4] = 14401
      "011100011111001" when "000101", -- t[5] = 14585
      "011100110110011" when "000110", -- t[6] = 14771
      "011101001110000" when "000111", -- t[7] = 14960
      "011101100110000" when "001000", -- t[8] = 15152
      "011101111110011" when "001001", -- t[9] = 15347
      "011110010111001" when "001010", -- t[10] = 15545
      "011110110000001" when "001011", -- t[11] = 15745
      "011111001001101" when "001100", -- t[12] = 15949
      "011111100011100" when "001101", -- t[13] = 16156
      "011111111101110" when "001110", -- t[14] = 16366
      "100000011000011" when "001111", -- t[15] = 16579
      "100000110011100" when "010000", -- t[16] = 16796
      "100001001111000" when "010001", -- t[17] = 17016
      "100001101010111" when "010010", -- t[18] = 17239
      "100010000111010" when "010011", -- t[19] = 17466
      "100010100100001" when "010100", -- t[20] = 17697
      "100011000001011" when "010101", -- t[21] = 17931
      "100011011111001" when "010110", -- t[22] = 18169
      "100011111101011" when "010111", -- t[23] = 18411
      "100100011100000" when "011000", -- t[24] = 18656
      "100100111011010" when "011001", -- t[25] = 18906
      "100101011011000" when "011010", -- t[26] = 19160
      "100101111011001" when "011011", -- t[27] = 19417
      "100110011011111" when "011100", -- t[28] = 19679
      "100110111101010" when "011101", -- t[29] = 19946
      "100111011111001" when "011110", -- t[30] = 20217
      "101000000001100" when "011111", -- t[31] = 20492
      "101000100100100" when "100000", -- t[32] = 20772
      "101001001000001" when "100001", -- t[33] = 21057
      "101001101100010" when "100010", -- t[34] = 21346
      "101010010001001" when "100011", -- t[35] = 21641
      "101010110110101" when "100100", -- t[36] = 21941
      "101011011100101" when "100101", -- t[37] = 22245
      "101100000011100" when "100110", -- t[38] = 22556
      "101100101010111" when "100111", -- t[39] = 22871
      "101101010011001" when "101000", -- t[40] = 23193
      "101101111100000" when "101001", -- t[41] = 23520
      "101110100101100" when "101010", -- t[42] = 23852
      "101111001111111" when "101011", -- t[43] = 24191
      "101111111011000" when "101100", -- t[44] = 24536
      "110000100111000" when "101101", -- t[45] = 24888
      "110001010011110" when "101110", -- t[46] = 25246
      "110010000001010" when "101111", -- t[47] = 25610
      "110010101111110" when "110000", -- t[48] = 25982
      "110011011111000" when "110001", -- t[49] = 26360
      "110100001111010" when "110010", -- t[50] = 26746
      "110101000000011" when "110011", -- t[51] = 27139
      "110101110010100" when "110100", -- t[52] = 27540
      "110110100101100" when "110101", -- t[53] = 27948
      "110111011001101" when "110110", -- t[54] = 28365
      "111000001110110" when "110111", -- t[55] = 28790
      "111001000100111" when "111000", -- t[56] = 29223
      "111001111100010" when "111001", -- t[57] = 29666
      "111010110100101" when "111010", -- t[58] = 30117
      "111011101110010" when "111011", -- t[59] = 30578
      "111100101001000" when "111100", -- t[60] = 31048
      "111101100101000" when "111101", -- t[61] = 31528
      "111110100010011" when "111110", -- t[62] = 32019
      "111111100001000" when "111111", -- t[63] = 32520
      "---------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_12_to2 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to2 is
begin
  with x select
    r <=
      "00010101" when "000000", -- t[0] = 21
      "01000000" when "000001", -- t[1] = 64
      "00010110" when "000010", -- t[2] = 22
      "01000010" when "000011", -- t[3] = 66
      "00010110" when "000100", -- t[4] = 22
      "01000100" when "000101", -- t[5] = 68
      "00010111" when "000110", -- t[6] = 23
      "01000110" when "000111", -- t[7] = 70
      "00011000" when "001000", -- t[8] = 24
      "01001000" when "001001", -- t[9] = 72
      "00011001" when "001010", -- t[10] = 25
      "01001011" when "001011", -- t[11] = 75
      "00011001" when "001100", -- t[12] = 25
      "01001101" when "001101", -- t[13] = 77
      "00011010" when "001110", -- t[14] = 26
      "01001111" when "001111", -- t[15] = 79
      "00011011" when "010000", -- t[16] = 27
      "01010010" when "010001", -- t[17] = 82
      "00011100" when "010010", -- t[18] = 28
      "01010100" when "010011", -- t[19] = 84
      "00011101" when "010100", -- t[20] = 29
      "01010111" when "010101", -- t[21] = 87
      "00011110" when "010110", -- t[22] = 30
      "01011010" when "010111", -- t[23] = 90
      "00011111" when "011000", -- t[24] = 31
      "01011101" when "011001", -- t[25] = 93
      "00100000" when "011010", -- t[26] = 32
      "01100000" when "011011", -- t[27] = 96
      "00100001" when "011100", -- t[28] = 33
      "01100011" when "011101", -- t[29] = 99
      "00100010" when "011110", -- t[30] = 34
      "01100111" when "011111", -- t[31] = 103
      "00100011" when "100000", -- t[32] = 35
      "01101010" when "100001", -- t[33] = 106
      "00100100" when "100010", -- t[34] = 36
      "01101110" when "100011", -- t[35] = 110
      "00100110" when "100100", -- t[36] = 38
      "01110010" when "100101", -- t[37] = 114
      "00100111" when "100110", -- t[38] = 39
      "01110110" when "100111", -- t[39] = 118
      "00101000" when "101000", -- t[40] = 40
      "01111010" when "101001", -- t[41] = 122
      "00101010" when "101010", -- t[42] = 42
      "01111110" when "101011", -- t[43] = 126
      "00101011" when "101100", -- t[44] = 43
      "10000011" when "101101", -- t[45] = 131
      "00101101" when "101110", -- t[46] = 45
      "10001000" when "101111", -- t[47] = 136
      "00101111" when "110000", -- t[48] = 47
      "10001101" when "110001", -- t[49] = 141
      "00110001" when "110010", -- t[50] = 49
      "10010011" when "110011", -- t[51] = 147
      "00110010" when "110100", -- t[52] = 50
      "10011000" when "110101", -- t[53] = 152
      "00110100" when "110110", -- t[54] = 52
      "10011110" when "110111", -- t[55] = 158
      "00110111" when "111000", -- t[56] = 55
      "10100101" when "111001", -- t[57] = 165
      "00111001" when "111010", -- t[58] = 57
      "10101100" when "111011", -- t[59] = 172
      "00111011" when "111100", -- t[60] = 59
      "10110011" when "111101", -- t[61] = 179
      "00111110" when "111110", -- t[62] = 62
      "10111011" when "111111", -- t[63] = 187
      "--------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_12_to1 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to1 is
begin
  with x select
    r <=
      "000101" when "0000", -- t[0] = 5
      "010000" when "0001", -- t[1] = 16
      "000110" when "0010", -- t[2] = 6
      "010011" when "0011", -- t[3] = 19
      "000111" when "0100", -- t[4] = 7
      "010101" when "0101", -- t[5] = 21
      "001000" when "0110", -- t[6] = 8
      "011000" when "0111", -- t[7] = 24
      "001001" when "1000", -- t[8] = 9
      "011100" when "1001", -- t[9] = 28
      "001010" when "1010", -- t[10] = 10
      "100000" when "1011", -- t[11] = 32
      "001100" when "1100", -- t[12] = 12
      "100101" when "1101", -- t[13] = 37
      "001110" when "1110", -- t[14] = 14
      "101100" when "1111", -- t[15] = 44
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T3_12_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(3 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to0 is
begin
  with x select
    r <=
      "0001" when "000", -- t[0] = 1
      "0100" when "001", -- t[1] = 4
      "0001" when "010", -- t[2] = 1
      "0101" when "011", -- t[3] = 5
      "0010" when "100", -- t[4] = 2
      "0111" when "101", -- t[5] = 7
      "0011" when "110", -- t[6] = 3
      "1010" when "111", -- t[7] = 10
      "----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_12.all;

entity LNSSub_MPT_T3_12_to2_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(7 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T3_12_to2
    port map( x => in_t,
              r => out_t );

  r(14 downto 8) <= (14 downto 8 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_12.all;

entity LNSSub_MPT_T3_12_to1_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(5 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T3_12_to1
    port map( x => in_t,
              r => out_t );

  r(14 downto 6) <= (14 downto 6 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_12.all;

entity LNSSub_MPT_T3_12_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(3 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T3_12_to0
    port map( x => in_t,
              r => out_t );

  r(14 downto 4) <= (14 downto 4 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_12.all;

entity LNSSub_MPT_T3_12 is
  port( x : in  std_logic_vector(11 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T3_12 is
  signal in_tiv  : std_logic_vector(5 downto 0);
  signal out_tiv : std_logic_vector(14 downto 0);
  signal a2      : std_logic_vector(4 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(14 downto 0);
  signal a1      : std_logic_vector(2 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(14 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(14 downto 0);
  signal sum     : std_logic_vector(14 downto 0);
begin
  in_tiv <= x(11 downto 6);
  inst_tiv : LNSSub_MPT_T3_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(11 downto 7);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T3_12_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(11 downto 9);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T3_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(11 downto 10);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T3_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(14 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T3_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T3_12_Clk is
  port( x   : in  std_logic_vector(11 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T3_12_Clk is
  signal in_tiv_1  : std_logic_vector(5 downto 0);
  signal out_tiv_1 : std_logic_vector(14 downto 0);
  signal out_tiv_2 : std_logic_vector(14 downto 0);
  signal a2_1      : std_logic_vector(4 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(14 downto 0);
  signal out2_2    : std_logic_vector(14 downto 0);
  signal a1_1      : std_logic_vector(2 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(14 downto 0);
  signal out1_2    : std_logic_vector(14 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(14 downto 0);
  signal out0_2    : std_logic_vector(14 downto 0);
  signal psum1_2     : std_logic_vector(14 downto 0);
  signal psum1_3     : std_logic_vector(14 downto 0);
  signal psum2_2     : std_logic_vector(14 downto 0);
  signal psum2_3     : std_logic_vector(14 downto 0);
  signal sum_3     : std_logic_vector(14 downto 0);
begin
  in_tiv_1 <= x(11 downto 6);
  inst_tiv : LNSSub_MPT_T3_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(11 downto 7);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T3_12_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(11 downto 9);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T3_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(11 downto 10);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T3_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(14 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-1.0 -0.5[ -> [0.0 2.0[
-- wI = 11 bits
-- wO = 11 bits
-- Decomposition: 5, 6 / 5, 4, 2 / 2, 2, 2
-- Guard bits: 5
-- Size: 1352 = 16.2^5 + 9.2^6 + 7.2^5 + 5.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T4_12 is
  component LNSSub_MPT_T4_12_tiv is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to2 is
    port( x : in  std_logic_vector(5 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to2_xor is
    port( a : in  std_logic_vector(4 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;

  component LNSSub_MPT_T4_12_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(15 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_12_tiv is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_tiv is
begin
  with x select
    r <=
      "1000000100010000" when "00000", -- t[0] = 33040
      "1000001100011011" when "00001", -- t[1] = 33563
      "1000010100110010" when "00010", -- t[2] = 34098
      "1000011101010101" when "00011", -- t[3] = 34645
      "1000100110000100" when "00100", -- t[4] = 35204
      "1000101111000001" when "00101", -- t[5] = 35777
      "1000111000001010" when "00110", -- t[6] = 36362
      "1001000001100010" when "00111", -- t[7] = 36962
      "1001001011001000" when "01000", -- t[8] = 37576
      "1001010100111100" when "01001", -- t[9] = 38204
      "1001011111000001" when "01010", -- t[10] = 38849
      "1001101001010101" when "01011", -- t[11] = 39509
      "1001110011111010" when "01100", -- t[12] = 40186
      "1001111110110000" when "01101", -- t[13] = 40880
      "1010001001111001" when "01110", -- t[14] = 41593
      "1010010101010100" when "01111", -- t[15] = 42324
      "1010100001000011" when "10000", -- t[16] = 43075
      "1010101101000110" when "10001", -- t[17] = 43846
      "1010111001011111" when "10010", -- t[18] = 44639
      "1011000110001111" when "10011", -- t[19] = 45455
      "1011010011010101" when "10100", -- t[20] = 46293
      "1011100000110100" when "10101", -- t[21] = 47156
      "1011101110101101" when "10110", -- t[22] = 48045
      "1011111101000001" when "10111", -- t[23] = 48961
      "1100001011110010" when "11000", -- t[24] = 49906
      "1100011011000000" when "11001", -- t[25] = 50880
      "1100101010101101" when "11010", -- t[26] = 51885
      "1100111010111100" when "11011", -- t[27] = 52924
      "1101001011101110" when "11100", -- t[28] = 53998
      "1101011101000101" when "11101", -- t[29] = 55109
      "1101101111000011" when "11110", -- t[30] = 56259
      "1110000001101011" when "11111", -- t[31] = 57451
      "----------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_12_to2 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to2 is
begin
  with x select
    r <=
      "001000000" when "000000", -- t[0] = 64
      "011000001" when "000001", -- t[1] = 193
      "001000001" when "000010", -- t[2] = 65
      "011000101" when "000011", -- t[3] = 197
      "001000011" when "000100", -- t[4] = 67
      "011001010" when "000101", -- t[5] = 202
      "001000100" when "000110", -- t[6] = 68
      "011001110" when "000111", -- t[7] = 206
      "001000110" when "001000", -- t[8] = 70
      "011010011" when "001001", -- t[9] = 211
      "001001000" when "001010", -- t[10] = 72
      "011011000" when "001011", -- t[11] = 216
      "001001001" when "001100", -- t[12] = 73
      "011011101" when "001101", -- t[13] = 221
      "001001011" when "001110", -- t[14] = 75
      "011100010" when "001111", -- t[15] = 226
      "001001101" when "010000", -- t[16] = 77
      "011101000" when "010001", -- t[17] = 232
      "001001111" when "010010", -- t[18] = 79
      "011101101" when "010011", -- t[19] = 237
      "001010001" when "010100", -- t[20] = 81
      "011110011" when "010101", -- t[21] = 243
      "001010011" when "010110", -- t[22] = 83
      "011111001" when "010111", -- t[23] = 249
      "001010101" when "011000", -- t[24] = 85
      "100000000" when "011001", -- t[25] = 256
      "001010111" when "011010", -- t[26] = 87
      "100000110" when "011011", -- t[27] = 262
      "001011001" when "011100", -- t[28] = 89
      "100001101" when "011101", -- t[29] = 269
      "001011100" when "011110", -- t[30] = 92
      "100010100" when "011111", -- t[31] = 276
      "001011110" when "100000", -- t[32] = 94
      "100011100" when "100001", -- t[33] = 284
      "001100001" when "100010", -- t[34] = 97
      "100100100" when "100011", -- t[35] = 292
      "001100100" when "100100", -- t[36] = 100
      "100101100" when "100101", -- t[37] = 300
      "001100110" when "100110", -- t[38] = 102
      "100110100" when "100111", -- t[39] = 308
      "001101001" when "101000", -- t[40] = 105
      "100111101" when "101001", -- t[41] = 317
      "001101101" when "101010", -- t[42] = 109
      "101000111" when "101011", -- t[43] = 327
      "001110000" when "101100", -- t[44] = 112
      "101010001" when "101101", -- t[45] = 337
      "001110011" when "101110", -- t[46] = 115
      "101011011" when "101111", -- t[47] = 347
      "001110111" when "110000", -- t[48] = 119
      "101100110" when "110001", -- t[49] = 358
      "001111011" when "110010", -- t[50] = 123
      "101110001" when "110011", -- t[51] = 369
      "001111111" when "110100", -- t[52] = 127
      "101111101" when "110101", -- t[53] = 381
      "010000011" when "110110", -- t[54] = 131
      "110001010" when "110111", -- t[55] = 394
      "010000111" when "111000", -- t[56] = 135
      "110010111" when "111001", -- t[57] = 407
      "010001100" when "111010", -- t[58] = 140
      "110100110" when "111011", -- t[59] = 422
      "010010001" when "111100", -- t[60] = 145
      "110110101" when "111101", -- t[61] = 437
      "010010111" when "111110", -- t[62] = 151
      "111000101" when "111111", -- t[63] = 453
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_12_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to1 is
begin
  with x select
    r <=
      "0010000" when "00000", -- t[0] = 16
      "0110001" when "00001", -- t[1] = 49
      "0010001" when "00010", -- t[2] = 17
      "0110011" when "00011", -- t[3] = 51
      "0010001" when "00100", -- t[4] = 17
      "0110101" when "00101", -- t[5] = 53
      "0010010" when "00110", -- t[6] = 18
      "0111000" when "00111", -- t[7] = 56
      "0010011" when "01000", -- t[8] = 19
      "0111010" when "01001", -- t[9] = 58
      "0010100" when "01010", -- t[10] = 20
      "0111101" when "01011", -- t[11] = 61
      "0010101" when "01100", -- t[12] = 21
      "1000001" when "01101", -- t[13] = 65
      "0010110" when "01110", -- t[14] = 22
      "1000100" when "01111", -- t[15] = 68
      "0011000" when "10000", -- t[16] = 24
      "1001000" when "10001", -- t[17] = 72
      "0011001" when "10010", -- t[18] = 25
      "1001100" when "10011", -- t[19] = 76
      "0011010" when "10100", -- t[20] = 26
      "1010000" when "10101", -- t[21] = 80
      "0011100" when "10110", -- t[22] = 28
      "1010101" when "10111", -- t[23] = 85
      "0011110" when "11000", -- t[24] = 30
      "1011011" when "11001", -- t[25] = 91
      "0100000" when "11010", -- t[26] = 32
      "1100001" when "11011", -- t[27] = 97
      "0100010" when "11100", -- t[28] = 34
      "1101000" when "11101", -- t[29] = 104
      "0100101" when "11110", -- t[30] = 37
      "1101111" when "11111", -- t[31] = 111
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T4_12_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to0 is
begin
  with x select
    r <=
      "00100" when "000", -- t[0] = 4
      "01101" when "001", -- t[1] = 13
      "00101" when "010", -- t[2] = 5
      "01111" when "011", -- t[3] = 15
      "00110" when "100", -- t[4] = 6
      "10011" when "101", -- t[5] = 19
      "01000" when "110", -- t[6] = 8
      "11001" when "111", -- t[7] = 25
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_12.all;

entity LNSSub_MPT_T4_12_to2_xor is
  port( a : in  std_logic_vector(4 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to2_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(5 downto 0);
  signal out_t : std_logic_vector(8 downto 0);
begin
  sign <= not b(1);
  in_t(5 downto 1) <= a(4 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to2 : LNSSub_MPT_T4_12_to2
    port map( x => in_t,
              r => out_t );

  r(15 downto 9) <= (15 downto 9 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
  r(7) <= out_t(7) xor sign;
  r(8) <= out_t(8) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_12.all;

entity LNSSub_MPT_T4_12_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(6 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T4_12_to1
    port map( x => in_t,
              r => out_t );

  r(15 downto 7) <= (15 downto 7 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_12.all;

entity LNSSub_MPT_T4_12_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T4_12_to0
    port map( x => in_t,
              r => out_t );

  r(15 downto 5) <= (15 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_12.all;

entity LNSSub_MPT_T4_12 is
  port( x : in  std_logic_vector(10 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T4_12 is
  signal in_tiv  : std_logic_vector(4 downto 0);
  signal out_tiv : std_logic_vector(15 downto 0);
  signal a2      : std_logic_vector(4 downto 0);
  signal b2      : std_logic_vector(1 downto 0);
  signal out2    : std_logic_vector(15 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(15 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(15 downto 0);
  signal sum     : std_logic_vector(15 downto 0);
begin
  in_tiv <= x(10 downto 6);
  inst_tiv : LNSSub_MPT_T4_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a2 <= x(10 downto 6);
  b2 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T4_12_to2_xor
    port map( a => a2,
              b => b2,
              r => out2 );

  a1 <= x(10 downto 7);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T4_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(10 downto 9);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T4_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out2 + out1 + out0;
  r <= sum(15 downto 5);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T4_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T4_12_Clk is
  port( x   : in  std_logic_vector(10 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T4_12_Clk is
  signal in_tiv_1  : std_logic_vector(4 downto 0);
  signal out_tiv_1 : std_logic_vector(15 downto 0);
  signal out_tiv_2 : std_logic_vector(15 downto 0);
  signal a2_1      : std_logic_vector(4 downto 0);
  signal b2_1      : std_logic_vector(1 downto 0);
  signal out2_1    : std_logic_vector(15 downto 0);
  signal out2_2    : std_logic_vector(15 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(15 downto 0);
  signal out1_2    : std_logic_vector(15 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(15 downto 0);
  signal out0_2    : std_logic_vector(15 downto 0);
  signal psum1_2     : std_logic_vector(15 downto 0);
  signal psum1_3     : std_logic_vector(15 downto 0);
  signal psum2_2     : std_logic_vector(15 downto 0);
  signal psum2_3     : std_logic_vector(15 downto 0);
  signal sum_3     : std_logic_vector(15 downto 0);
begin
  in_tiv_1 <= x(10 downto 6);
  inst_tiv : LNSSub_MPT_T4_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a2_1 <= x(10 downto 6);
  b2_1 <= x(5 downto 4);
  inst_to2_xor : LNSSub_MPT_T4_12_to2_xor
    port map( a => a2_1,
              b => b2_1,
              r => out2_1 );

  a1_1 <= x(10 downto 7);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T4_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(10 downto 9);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T4_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out2_2    <= out2_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out2_2;
  psum2_2 <= out1_2 + out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(15 downto 5);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.5 -0.25[ -> [0.0 4.0[
-- wI = 10 bits
-- wO = 11 bits
-- Decomposition: 5, 5 / 4, 3 / 2, 3
-- Guard bits: 4
-- Size: 896 = 15.2^5 + 7.2^5 + 6.2^5

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T5_12 is
  component LNSSub_MPT_T5_12_tiv is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T5_12_to1 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T5_12_to0 is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(5 downto 0) );
  end component;

  component LNSSub_MPT_T5_12_to1_xor is
    port( a : in  std_logic_vector(3 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;

  component LNSSub_MPT_T5_12_to0_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(14 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_12_tiv is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12_tiv is
begin
  with x select
    r <=
      "011100100000101" when "00000", -- t[0] = 14597
      "011100110100010" when "00001", -- t[1] = 14754
      "011101001000010" when "00010", -- t[2] = 14914
      "011101011100110" when "00011", -- t[3] = 15078
      "011101110001100" when "00100", -- t[4] = 15244
      "011110000110110" when "00101", -- t[5] = 15414
      "011110011100100" when "00110", -- t[6] = 15588
      "011110110010101" when "00111", -- t[7] = 15765
      "011111001001001" when "01000", -- t[8] = 15945
      "011111100000010" when "01001", -- t[9] = 16130
      "011111110111110" when "01010", -- t[10] = 16318
      "100000001111111" when "01011", -- t[11] = 16511
      "100000101000011" when "01100", -- t[12] = 16707
      "100001000001101" when "01101", -- t[13] = 16909
      "100001011011010" when "01110", -- t[14] = 17114
      "100001110101101" when "01111", -- t[15] = 17325
      "100010010000101" when "10000", -- t[16] = 17541
      "100010101100001" when "10001", -- t[17] = 17761
      "100011001000100" when "10010", -- t[18] = 17988
      "100011100101011" when "10011", -- t[19] = 18219
      "100100000011001" when "10100", -- t[20] = 18457
      "100100100001101" when "10101", -- t[21] = 18701
      "100101000001000" when "10110", -- t[22] = 18952
      "100101100001001" when "10111", -- t[23] = 19209
      "100110000010010" when "11000", -- t[24] = 19474
      "100110100100010" when "11001", -- t[25] = 19746
      "100111000111010" when "11010", -- t[26] = 20026
      "100111101011010" when "11011", -- t[27] = 20314
      "101000010000100" when "11100", -- t[28] = 20612
      "101000110110110" when "11101", -- t[29] = 20918
      "101001011110011" when "11110", -- t[30] = 21235
      "101010000111010" when "11111", -- t[31] = 21562
      "---------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_12_to1 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12_to1 is
begin
  with x select
    r <=
      "0010011" when "00000", -- t[0] = 19
      "0111010" when "00001", -- t[1] = 58
      "0010100" when "00010", -- t[2] = 20
      "0111101" when "00011", -- t[3] = 61
      "0010101" when "00100", -- t[4] = 21
      "0111111" when "00101", -- t[5] = 63
      "0010110" when "00110", -- t[6] = 22
      "1000010" when "00111", -- t[7] = 66
      "0010110" when "01000", -- t[8] = 22
      "1000100" when "01001", -- t[9] = 68
      "0011000" when "01010", -- t[10] = 24
      "1001000" when "01011", -- t[11] = 72
      "0011001" when "01100", -- t[12] = 25
      "1001011" when "01101", -- t[13] = 75
      "0011010" when "01110", -- t[14] = 26
      "1001110" when "01111", -- t[15] = 78
      "0011011" when "10000", -- t[16] = 27
      "1010010" when "10001", -- t[17] = 82
      "0011100" when "10010", -- t[18] = 28
      "1010110" when "10011", -- t[19] = 86
      "0011110" when "10100", -- t[20] = 30
      "1011011" when "10101", -- t[21] = 91
      "0100000" when "10110", -- t[22] = 32
      "1100000" when "10111", -- t[23] = 96
      "0100001" when "11000", -- t[24] = 33
      "1100101" when "11001", -- t[25] = 101
      "0100011" when "11010", -- t[26] = 35
      "1101011" when "11011", -- t[27] = 107
      "0100110" when "11100", -- t[28] = 38
      "1110010" when "11101", -- t[29] = 114
      "0101000" when "11110", -- t[30] = 40
      "1111010" when "11111", -- t[31] = 122
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T5_12_to0 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(5 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12_to0 is
begin
  with x select
    r <=
      "000010" when "00000", -- t[0] = 2
      "000111" when "00001", -- t[1] = 7
      "001100" when "00010", -- t[2] = 12
      "010001" when "00011", -- t[3] = 17
      "000010" when "00100", -- t[4] = 2
      "001000" when "00101", -- t[5] = 8
      "001101" when "00110", -- t[6] = 13
      "010010" when "00111", -- t[7] = 18
      "000010" when "01000", -- t[8] = 2
      "001000" when "01001", -- t[9] = 8
      "001110" when "01010", -- t[10] = 14
      "010100" when "01011", -- t[11] = 20
      "000011" when "01100", -- t[12] = 3
      "001001" when "01101", -- t[13] = 9
      "010000" when "01110", -- t[14] = 16
      "010110" when "01111", -- t[15] = 22
      "000011" when "10000", -- t[16] = 3
      "001010" when "10001", -- t[17] = 10
      "010001" when "10010", -- t[18] = 17
      "011000" when "10011", -- t[19] = 24
      "000011" when "10100", -- t[20] = 3
      "001011" when "10101", -- t[21] = 11
      "010011" when "10110", -- t[22] = 19
      "011011" when "10111", -- t[23] = 27
      "000100" when "11000", -- t[24] = 4
      "001101" when "11001", -- t[25] = 13
      "010101" when "11010", -- t[26] = 21
      "011110" when "11011", -- t[27] = 30
      "000100" when "11100", -- t[28] = 4
      "001110" when "11101", -- t[29] = 14
      "011000" when "11110", -- t[30] = 24
      "100010" when "11111", -- t[31] = 34
      "------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_12.all;

entity LNSSub_MPT_T5_12_to1_xor is
  port( a : in  std_logic_vector(3 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(6 downto 0);
begin
  sign <= not b(1);
  in_t(4 downto 1) <= a(3 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T5_12_to1
    port map( x => in_t,
              r => out_t );

  r(14 downto 7) <= (14 downto 7 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
  r(6) <= out_t(6) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_12.all;

entity LNSSub_MPT_T5_12_to0_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(14 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(4 downto 0);
  signal out_t : std_logic_vector(5 downto 0);
begin
  sign <= not b(2);
  in_t(4 downto 2) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T5_12_to0
    port map( x => in_t,
              r => out_t );

  r(14 downto 6) <= (14 downto 6 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
  r(5) <= out_t(5) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_12.all;

entity LNSSub_MPT_T5_12 is
  port( x : in  std_logic_vector(9 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T5_12 is
  signal in_tiv  : std_logic_vector(4 downto 0);
  signal out_tiv : std_logic_vector(14 downto 0);
  signal a1      : std_logic_vector(3 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(14 downto 0);
  signal a0      : std_logic_vector(2 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(14 downto 0);
  signal sum     : std_logic_vector(14 downto 0);
begin
  in_tiv <= x(9 downto 5);
  inst_tiv : LNSSub_MPT_T5_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(9 downto 6);
  b1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T5_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(9 downto 7);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T5_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(14 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T5_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T5_12_Clk is
  port( x   : in  std_logic_vector(9 downto 0);
        r   : out std_logic_vector(10 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T5_12_Clk is
  signal in_tiv_1  : std_logic_vector(4 downto 0);
  signal out_tiv_1 : std_logic_vector(14 downto 0);
  signal out_tiv_2 : std_logic_vector(14 downto 0);
  signal a1_1      : std_logic_vector(3 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(14 downto 0);
  signal out1_2    : std_logic_vector(14 downto 0);
  signal a0_1      : std_logic_vector(2 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(14 downto 0);
  signal out0_2    : std_logic_vector(14 downto 0);
  signal psum1_2     : std_logic_vector(14 downto 0);
  signal psum1_3     : std_logic_vector(14 downto 0);
  signal psum2_2     : std_logic_vector(14 downto 0);
  signal psum2_3     : std_logic_vector(14 downto 0);
  signal sum_3     : std_logic_vector(14 downto 0);
begin
  in_tiv_1 <= x(9 downto 5);
  inst_tiv : LNSSub_MPT_T5_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(9 downto 6);
  b1_1 <= x(4 downto 3);
  inst_to1_xor : LNSSub_MPT_T5_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(9 downto 7);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T5_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(14 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.25 -0.12500000000000003[ -> [0.0 4.0[
-- wI = 9 bits
-- wO = 10 bits
-- Decomposition: 5, 4 / 3, 1 / 2, 2
-- Guard bits: 3
-- Size: 508 = 13.2^5 + 5.2^4 + 3.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T6_12 is
  component LNSSub_MPT_T6_12_tiv is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T6_12_to1 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T6_12_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T6_12_to1_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T6_12_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_12_tiv is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12_tiv is
begin
  with x select
    r <=
      "1010101010000" when "00000", -- t[0] = 5456
      "1010101111011" when "00001", -- t[1] = 5499
      "1010110100110" when "00010", -- t[2] = 5542
      "1010111010011" when "00011", -- t[3] = 5587
      "1011000000000" when "00100", -- t[4] = 5632
      "1011000101110" when "00101", -- t[5] = 5678
      "1011001011101" when "00110", -- t[6] = 5725
      "1011010001101" when "00111", -- t[7] = 5773
      "1011010111110" when "01000", -- t[8] = 5822
      "1011011110000" when "01001", -- t[9] = 5872
      "1011100100011" when "01010", -- t[10] = 5923
      "1011101010111" when "01011", -- t[11] = 5975
      "1011110001100" when "01100", -- t[12] = 6028
      "1011111000010" when "01101", -- t[13] = 6082
      "1011111111001" when "01110", -- t[14] = 6137
      "1100000110001" when "01111", -- t[15] = 6193
      "1100001101011" when "10000", -- t[16] = 6251
      "1100010100110" when "10001", -- t[17] = 6310
      "1100011100010" when "10010", -- t[18] = 6370
      "1100100100000" when "10011", -- t[19] = 6432
      "1100101011111" when "10100", -- t[20] = 6495
      "1100110011111" when "10101", -- t[21] = 6559
      "1100111100010" when "10110", -- t[22] = 6626
      "1101000100110" when "10111", -- t[23] = 6694
      "1101001101100" when "11000", -- t[24] = 6764
      "1101010110100" when "11001", -- t[25] = 6836
      "1101011111101" when "11010", -- t[26] = 6909
      "1101101001001" when "11011", -- t[27] = 6985
      "1101110010111" when "11100", -- t[28] = 7063
      "1101111101000" when "11101", -- t[29] = 7144
      "1110000111011" when "11110", -- t[30] = 7227
      "1110010010000" when "11111", -- t[31] = 7312
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_12_to1 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12_to1 is
begin
  with x select
    r <=
      "00101" when "0000", -- t[0] = 5
      "10000" when "0001", -- t[1] = 16
      "00101" when "0010", -- t[2] = 5
      "10001" when "0011", -- t[3] = 17
      "00110" when "0100", -- t[4] = 6
      "10011" when "0101", -- t[5] = 19
      "00110" when "0110", -- t[6] = 6
      "10100" when "0111", -- t[7] = 20
      "00111" when "1000", -- t[8] = 7
      "10110" when "1001", -- t[9] = 22
      "01000" when "1010", -- t[10] = 8
      "11000" when "1011", -- t[11] = 24
      "01001" when "1100", -- t[12] = 9
      "11011" when "1101", -- t[13] = 27
      "01010" when "1110", -- t[14] = 10
      "11110" when "1111", -- t[15] = 30
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T6_12_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12_to0 is
begin
  with x select
    r <=
      "001" when "00", -- t[0] = 1
      "100" when "01", -- t[1] = 4
      "010" when "10", -- t[2] = 2
      "110" when "11", -- t[3] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_12.all;

entity LNSSub_MPT_T6_12_to1_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T6_12_to1
    port map( x => in_t,
              r => out_t );

  r(12 downto 5) <= (12 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_12.all;

entity LNSSub_MPT_T6_12_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T6_12_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 3) <= (12 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_12.all;

entity LNSSub_MPT_T6_12 is
  port( x : in  std_logic_vector(8 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T6_12 is
  signal in_tiv  : std_logic_vector(4 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a1      : std_logic_vector(2 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(8 downto 4);
  inst_tiv : LNSSub_MPT_T6_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(8 downto 6);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T6_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(8 downto 8);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T6_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(12 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T6_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T6_12_Clk is
  port( x   : in  std_logic_vector(8 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T6_12_Clk is
  signal in_tiv_1  : std_logic_vector(4 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a1_1      : std_logic_vector(2 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(12 downto 0);
  signal out1_2    : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(8 downto 4);
  inst_tiv : LNSSub_MPT_T6_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(8 downto 6);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T6_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(8 downto 8);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T6_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.12500000000000003 -0.0625[ -> [0.0 7.999999999999998[
-- wI = 8 bits
-- wO = 10 bits
-- Decomposition: 5, 3 / 2 / 3
-- Guard bits: 3
-- Size: 496 = 13.2^5 + 5.2^4

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T7_12 is
  component LNSSub_MPT_T7_12_tiv is
    port( x : in  std_logic_vector(4 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;

  component LNSSub_MPT_T7_12_to0 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T7_12_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(12 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T7_12_tiv is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_12_tiv is
begin
  with x select
    r <=
      "0111001101011" when "00000", -- t[0] = 3691
      "0111010000001" when "00001", -- t[1] = 3713
      "0111010011000" when "00010", -- t[2] = 3736
      "0111010101111" when "00011", -- t[3] = 3759
      "0111011000111" when "00100", -- t[4] = 3783
      "0111011011111" when "00101", -- t[5] = 3807
      "0111011110111" when "00110", -- t[6] = 3831
      "0111100010000" when "00111", -- t[7] = 3856
      "0111100101010" when "01000", -- t[8] = 3882
      "0111101000011" when "01001", -- t[9] = 3907
      "0111101011110" when "01010", -- t[10] = 3934
      "0111101111001" when "01011", -- t[11] = 3961
      "0111110010100" when "01100", -- t[12] = 3988
      "0111110110000" when "01101", -- t[13] = 4016
      "0111111001100" when "01110", -- t[14] = 4044
      "0111111101010" when "01111", -- t[15] = 4074
      "1000000000111" when "10000", -- t[16] = 4103
      "1000000100110" when "10001", -- t[17] = 4134
      "1000001000101" when "10010", -- t[18] = 4165
      "1000001100101" when "10011", -- t[19] = 4197
      "1000010000101" when "10100", -- t[20] = 4229
      "1000010100111" when "10101", -- t[21] = 4263
      "1000011001001" when "10110", -- t[22] = 4297
      "1000011101100" when "10111", -- t[23] = 4332
      "1000100010000" when "11000", -- t[24] = 4368
      "1000100110100" when "11001", -- t[25] = 4404
      "1000101011010" when "11010", -- t[26] = 4442
      "1000110000001" when "11011", -- t[27] = 4481
      "1000110101001" when "11100", -- t[28] = 4521
      "1000111010010" when "11101", -- t[29] = 4562
      "1000111111101" when "11110", -- t[30] = 4605
      "1001000101000" when "11111", -- t[31] = 4648
      "-------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T7_12_to0 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_12_to0 is
begin
  with x select
    r <=
      "00001" when "0000", -- t[0] = 1
      "00100" when "0001", -- t[1] = 4
      "00111" when "0010", -- t[2] = 7
      "01010" when "0011", -- t[3] = 10
      "00001" when "0100", -- t[4] = 1
      "00101" when "0101", -- t[5] = 5
      "01000" when "0110", -- t[6] = 8
      "01011" when "0111", -- t[7] = 11
      "00010" when "1000", -- t[8] = 2
      "00110" when "1001", -- t[9] = 6
      "01010" when "1010", -- t[10] = 10
      "01110" when "1011", -- t[11] = 14
      "00010" when "1100", -- t[12] = 2
      "00111" when "1101", -- t[13] = 7
      "01100" when "1110", -- t[14] = 12
      "10001" when "1111", -- t[15] = 17
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_12.all;

entity LNSSub_MPT_T7_12_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(12 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(2);
  in_t(3 downto 2) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T7_12_to0
    port map( x => in_t,
              r => out_t );

  r(12 downto 5) <= (12 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_12.all;

entity LNSSub_MPT_T7_12 is
  port( x : in  std_logic_vector(7 downto 0);
        r : out std_logic_vector(9 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T7_12 is
  signal in_tiv  : std_logic_vector(4 downto 0);
  signal out_tiv : std_logic_vector(12 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(12 downto 0);
  signal sum     : std_logic_vector(12 downto 0);
begin
  in_tiv <= x(7 downto 3);
  inst_tiv : LNSSub_MPT_T7_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a0 <= x(7 downto 6);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T7_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(12 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T7_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T7_12_Clk is
  port( x   : in  std_logic_vector(7 downto 0);
        r   : out std_logic_vector(9 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T7_12_Clk is
  signal in_tiv_1  : std_logic_vector(4 downto 0);
  signal out_tiv_1 : std_logic_vector(12 downto 0);
  signal out_tiv_2 : std_logic_vector(12 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(12 downto 0);
  signal out0_2    : std_logic_vector(12 downto 0);
  signal psum1_2     : std_logic_vector(12 downto 0);
  signal psum1_3     : std_logic_vector(12 downto 0);
  signal psum2_2     : std_logic_vector(12 downto 0);
  signal psum2_3     : std_logic_vector(12 downto 0);
  signal sum_3     : std_logic_vector(12 downto 0);
begin
  in_tiv_1 <= x(7 downto 3);
  inst_tiv : LNSSub_MPT_T7_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a0_1 <= x(7 downto 6);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T7_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(12 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.0625 -0.03125[ -> [0.0 7.999999999999998[
-- wI = 7 bits
-- wO = 9 bits
-- Decomposition: 3, 4 / 3, 1 / 2, 2
-- Guard bits: 3
-- Size: 188 = 12.2^3 + 5.2^4 + 3.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T8_12 is
  component LNSSub_MPT_T8_12_tiv is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T8_12_to1 is
    port( x : in  std_logic_vector(3 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T8_12_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T8_12_to1_xor is
    port( a : in  std_logic_vector(2 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;

  component LNSSub_MPT_T8_12_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(11 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_12_tiv is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12_tiv is
begin
  with x select
    r <=
      "100100111001" when "000", -- t[0] = 2361
      "100101101001" when "001", -- t[1] = 2409
      "100110011101" when "010", -- t[2] = 2461
      "100111010101" when "011", -- t[3] = 2517
      "101000010001" when "100", -- t[4] = 2577
      "101001010011" when "101", -- t[5] = 2643
      "101010011100" when "110", -- t[6] = 2716
      "101011101101" when "111", -- t[7] = 2797
      "------------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_12_to1 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12_to1 is
begin
  with x select
    r <=
      "00101" when "0000", -- t[0] = 5
      "10001" when "0001", -- t[1] = 17
      "00110" when "0010", -- t[2] = 6
      "10010" when "0011", -- t[3] = 18
      "00110" when "0100", -- t[4] = 6
      "10011" when "0101", -- t[5] = 19
      "00111" when "0110", -- t[6] = 7
      "10101" when "0111", -- t[7] = 21
      "00111" when "1000", -- t[8] = 7
      "10111" when "1001", -- t[9] = 23
      "01000" when "1010", -- t[10] = 8
      "11001" when "1011", -- t[11] = 25
      "01001" when "1100", -- t[12] = 9
      "11100" when "1101", -- t[13] = 28
      "01010" when "1110", -- t[14] = 10
      "11111" when "1111", -- t[15] = 31
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T8_12_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12_to0 is
begin
  with x select
    r <=
      "001" when "00", -- t[0] = 1
      "100" when "01", -- t[1] = 4
      "010" when "10", -- t[2] = 2
      "110" when "11", -- t[3] = 6
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_12.all;

entity LNSSub_MPT_T8_12_to1_xor is
  port( a : in  std_logic_vector(2 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(3 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(1);
  in_t(3 downto 1) <= a(2 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T8_12_to1
    port map( x => in_t,
              r => out_t );

  r(11 downto 5) <= (11 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_12.all;

entity LNSSub_MPT_T8_12_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(11 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T8_12_to0
    port map( x => in_t,
              r => out_t );

  r(11 downto 3) <= (11 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_12.all;

entity LNSSub_MPT_T8_12 is
  port( x : in  std_logic_vector(6 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T8_12 is
  signal in_tiv  : std_logic_vector(2 downto 0);
  signal out_tiv : std_logic_vector(11 downto 0);
  signal a1      : std_logic_vector(2 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(11 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(11 downto 0);
  signal sum     : std_logic_vector(11 downto 0);
begin
  in_tiv <= x(6 downto 4);
  inst_tiv : LNSSub_MPT_T8_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(6 downto 4);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T8_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(6 downto 6);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T8_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(11 downto 3);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T8_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T8_12_Clk is
  port( x   : in  std_logic_vector(6 downto 0);
        r   : out std_logic_vector(8 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T8_12_Clk is
  signal in_tiv_1  : std_logic_vector(2 downto 0);
  signal out_tiv_1 : std_logic_vector(11 downto 0);
  signal out_tiv_2 : std_logic_vector(11 downto 0);
  signal a1_1      : std_logic_vector(2 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(11 downto 0);
  signal out1_2    : std_logic_vector(11 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(11 downto 0);
  signal out0_2    : std_logic_vector(11 downto 0);
  signal psum1_2     : std_logic_vector(11 downto 0);
  signal psum1_3     : std_logic_vector(11 downto 0);
  signal psum2_2     : std_logic_vector(11 downto 0);
  signal psum2_3     : std_logic_vector(11 downto 0);
  signal sum_3     : std_logic_vector(11 downto 0);
begin
  in_tiv_1 <= x(6 downto 4);
  inst_tiv : LNSSub_MPT_T8_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(6 downto 4);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T8_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(6 downto 6);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T8_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(11 downto 3);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.03125 -0.015625000000000007[ -> [0.0 7.999999999999998[
-- wI = 6 bits
-- wO = 8 bits
-- Decomposition: 2, 4 / 2, 1 / 2, 2
-- Guard bits: 1
-- Size: 64 = 9.2^2 + 3.2^3 + 1.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T9_12 is
  component LNSSub_MPT_T9_12_tiv is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T9_12_to1 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T9_12_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(0 downto 0) );
  end component;

  component LNSSub_MPT_T9_12_to1_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T9_12_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_12_tiv is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12_tiv is
begin
  with x select
    r <=
      "101101010" when "00", -- t[0] = 362
      "101110111" when "01", -- t[1] = 375
      "110000110" when "10", -- t[2] = 390
      "110011001" when "11", -- t[3] = 409
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_12_to1 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12_to1 is
begin
  with x select
    r <=
      "001" when "000", -- t[0] = 1
      "100" when "001", -- t[1] = 4
      "001" when "010", -- t[2] = 1
      "101" when "011", -- t[3] = 5
      "010" when "100", -- t[4] = 2
      "110" when "101", -- t[5] = 6
      "010" when "110", -- t[6] = 2
      "111" when "111", -- t[7] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T9_12_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(0 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12_to0 is
begin
  with x select
    r <=
      "0" when "00", -- t[0] = 0
      "1" when "01", -- t[1] = 1
      "0" when "10", -- t[2] = 0
      "1" when "11", -- t[3] = 1
      "-" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_12.all;

entity LNSSub_MPT_T9_12_to1_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12_to1_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to1 : LNSSub_MPT_T9_12_to1
    port map( x => in_t,
              r => out_t );

  r(8 downto 3) <= (8 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_12.all;

entity LNSSub_MPT_T9_12_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(0 downto 0);
begin
  sign <= not b(1);
  in_t(1 downto 1) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T9_12_to0
    port map( x => in_t,
              r => out_t );

  r(8 downto 1) <= (8 downto 1 => sign);
  r(0) <= out_t(0) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_12.all;

entity LNSSub_MPT_T9_12 is
  port( x : in  std_logic_vector(5 downto 0);
        r : out std_logic_vector(7 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T9_12 is
  signal in_tiv  : std_logic_vector(1 downto 0);
  signal out_tiv : std_logic_vector(8 downto 0);
  signal a1      : std_logic_vector(1 downto 0);
  signal b1      : std_logic_vector(1 downto 0);
  signal out1    : std_logic_vector(8 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(8 downto 0);
  signal sum     : std_logic_vector(8 downto 0);
begin
  in_tiv <= x(5 downto 4);
  inst_tiv : LNSSub_MPT_T9_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a1 <= x(5 downto 4);
  b1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T9_12_to1_xor
    port map( a => a1,
              b => b1,
              r => out1 );

  a0 <= x(5 downto 5);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T9_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out1 + out0;
  r <= sum(8 downto 1);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T9_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T9_12_Clk is
  port( x   : in  std_logic_vector(5 downto 0);
        r   : out std_logic_vector(7 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T9_12_Clk is
  signal in_tiv_1  : std_logic_vector(1 downto 0);
  signal out_tiv_1 : std_logic_vector(8 downto 0);
  signal out_tiv_2 : std_logic_vector(8 downto 0);
  signal a1_1      : std_logic_vector(1 downto 0);
  signal b1_1      : std_logic_vector(1 downto 0);
  signal out1_1    : std_logic_vector(8 downto 0);
  signal out1_2    : std_logic_vector(8 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(8 downto 0);
  signal out0_2    : std_logic_vector(8 downto 0);
  signal psum1_2     : std_logic_vector(8 downto 0);
  signal psum1_3     : std_logic_vector(8 downto 0);
  signal psum2_2     : std_logic_vector(8 downto 0);
  signal psum2_3     : std_logic_vector(8 downto 0);
  signal sum_3     : std_logic_vector(8 downto 0);
begin
  in_tiv_1 <= x(5 downto 4);
  inst_tiv : LNSSub_MPT_T9_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a1_1 <= x(5 downto 4);
  b1_1 <= x(3 downto 2);
  inst_to1_xor : LNSSub_MPT_T9_12_to1_xor
    port map( a => a1_1,
              b => b1_1,
              r => out1_1 );

  a0_1 <= x(5 downto 5);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T9_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out1_2    <= out1_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2 + out1_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(8 downto 1);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.015625000000000007 -0.007812500000000002[ -> [0.0 7.999999999999998[
-- wI = 5 bits
-- wO = 7 bits
-- Decomposition: 2, 3 / 1 / 3
-- Guard bits: 2
-- Size: 60 = 9.2^2 + 3.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T10_12 is
  component LNSSub_MPT_T10_12_tiv is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;

  component LNSSub_MPT_T10_12_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T10_12_to0_xor is
    port( a : in  std_logic_vector(0 downto 0);
          b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(8 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T10_12_tiv is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_12_tiv is
begin
  with x select
    r <=
      "110101010" when "00", -- t[0] = 426
      "110110111" when "01", -- t[1] = 439
      "111000110" when "10", -- t[2] = 454
      "111011000" when "11", -- t[3] = 472
      "---------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T10_12_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_12_to0 is
begin
  with x select
    r <=
      "000" when "000", -- t[0] = 0
      "010" when "001", -- t[1] = 2
      "100" when "010", -- t[2] = 4
      "101" when "011", -- t[3] = 5
      "001" when "100", -- t[4] = 1
      "011" when "101", -- t[5] = 3
      "101" when "110", -- t[6] = 5
      "111" when "111", -- t[7] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_12.all;

entity LNSSub_MPT_T10_12_to0_xor is
  port( a : in  std_logic_vector(0 downto 0);
        b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(8 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(2);
  in_t(2 downto 2) <= a(0 downto 0);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T10_12_to0
    port map( x => in_t,
              r => out_t );

  r(8 downto 3) <= (8 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_12.all;

entity LNSSub_MPT_T10_12 is
  port( x : in  std_logic_vector(4 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T10_12 is
  signal in_tiv  : std_logic_vector(1 downto 0);
  signal out_tiv : std_logic_vector(8 downto 0);
  signal a0      : std_logic_vector(0 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(8 downto 0);
  signal sum     : std_logic_vector(8 downto 0);
begin
  in_tiv <= x(4 downto 3);
  inst_tiv : LNSSub_MPT_T10_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a0 <= x(4 downto 4);
  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T10_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(8 downto 2);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T10_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T10_12_Clk is
  port( x   : in  std_logic_vector(4 downto 0);
        r   : out std_logic_vector(6 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T10_12_Clk is
  signal in_tiv_1  : std_logic_vector(1 downto 0);
  signal out_tiv_1 : std_logic_vector(8 downto 0);
  signal out_tiv_2 : std_logic_vector(8 downto 0);
  signal a0_1      : std_logic_vector(0 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(8 downto 0);
  signal out0_2    : std_logic_vector(8 downto 0);
  signal psum1_2     : std_logic_vector(8 downto 0);
  signal psum1_3     : std_logic_vector(8 downto 0);
  signal psum2_2     : std_logic_vector(8 downto 0);
  signal psum2_3     : std_logic_vector(8 downto 0);
  signal sum_3     : std_logic_vector(8 downto 0);
begin
  in_tiv_1 <= x(4 downto 3);
  inst_tiv : LNSSub_MPT_T10_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a0_1 <= x(4 downto 4);
  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T10_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(8 downto 2);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.007812500000000002 -0.003906250000000001[ -> [0.0 15.999999999999998[
-- wI = 4 bits
-- wO = 7 bits
-- Decomposition: 1, 3 / 0 / 3
-- Guard bits: 4
-- Size: 42 = 11.2^1 + 5.2^2

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T11_12 is
  component LNSSub_MPT_T11_12_tiv is
    port( x : in  std_logic_vector(0 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;

  component LNSSub_MPT_T11_12_to0 is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(4 downto 0) );
  end component;

  component LNSSub_MPT_T11_12_to0_xor is
    port( b : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(10 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T11_12_tiv is
  port( x : in  std_logic_vector(0 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_12_tiv is
begin
  with x select
    r <=
      "01111100011" when "0", -- t[0] = 995
      "10000100001" when "1", -- t[1] = 1057
      "-----------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T11_12_to0 is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(4 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_12_to0 is
begin
  with x select
    r <=
      "00011" when "00", -- t[0] = 3
      "01011" when "01", -- t[1] = 11
      "10010" when "10", -- t[2] = 18
      "11010" when "11", -- t[3] = 26
      "-----" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_12.all;

entity LNSSub_MPT_T11_12_to0_xor is
  port( b : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(10 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(1 downto 0);
  signal out_t : std_logic_vector(4 downto 0);
begin
  sign <= not b(2);
  in_t(0) <= b(0) xor sign;
  in_t(1) <= b(1) xor sign;

  inst_to0 : LNSSub_MPT_T11_12_to0
    port map( x => in_t,
              r => out_t );

  r(10 downto 5) <= (10 downto 5 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
  r(3) <= out_t(3) xor sign;
  r(4) <= out_t(4) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_12.all;

entity LNSSub_MPT_T11_12 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T11_12 is
  signal in_tiv  : std_logic_vector(0 downto 0);
  signal out_tiv : std_logic_vector(10 downto 0);
  signal b0      : std_logic_vector(2 downto 0);
  signal out0    : std_logic_vector(10 downto 0);
  signal sum     : std_logic_vector(10 downto 0);
begin
  in_tiv <= x(3 downto 3);
  inst_tiv : LNSSub_MPT_T11_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  b0 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T11_12_to0_xor
    port map( b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(10 downto 4);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T11_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T11_12_Clk is
  port( x   : in  std_logic_vector(3 downto 0);
        r   : out std_logic_vector(6 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T11_12_Clk is
  signal in_tiv_1  : std_logic_vector(0 downto 0);
  signal out_tiv_1 : std_logic_vector(10 downto 0);
  signal out_tiv_2 : std_logic_vector(10 downto 0);
  signal b0_1      : std_logic_vector(2 downto 0);
  signal out0_1    : std_logic_vector(10 downto 0);
  signal out0_2    : std_logic_vector(10 downto 0);
  signal psum1_2     : std_logic_vector(10 downto 0);
  signal psum1_3     : std_logic_vector(10 downto 0);
  signal psum2_2     : std_logic_vector(10 downto 0);
  signal psum2_3     : std_logic_vector(10 downto 0);
  signal sum_3     : std_logic_vector(10 downto 0);
begin
  in_tiv_1 <= x(3 downto 3);
  inst_tiv : LNSSub_MPT_T11_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  b0_1 <= x(2 downto 0);
  inst_to0_xor : LNSSub_MPT_T11_12_to0_xor
    port map( b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(10 downto 4);
end architecture;


-- MultiPartite: LNS subtraction function: [-0.003906250000000001 0.0[ -> [0.0 15.999999999999998[
-- wI = 4 bits
-- wO = 7 bits
-- Decomposition: 2, 2 / 2 / 2
-- Guard bits: 0
-- Size: 52 = 7.2^2 + 3.2^3

library ieee;
use ieee.std_logic_1164.all;

package pkg_LNSSub_MPT_T12_12 is
  component LNSSub_MPT_T12_12_tiv is
    port( x : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;

  component LNSSub_MPT_T12_12_to0 is
    port( x : in  std_logic_vector(2 downto 0);
          r : out std_logic_vector(2 downto 0) );
  end component;

  component LNSSub_MPT_T12_12_to0_xor is
    port( a : in  std_logic_vector(1 downto 0);
          b : in  std_logic_vector(1 downto 0);
          r : out std_logic_vector(6 downto 0) );
  end component;
end package;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T12_12_tiv is
  port( x : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_12_tiv is
begin
  with x select
    r <=
      "1000110" when "00", -- t[0] = 70
      "1001010" when "01", -- t[1] = 74
      "1001111" when "10", -- t[2] = 79
      "1011101" when "11", -- t[3] = 93
      "-------" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;

entity LNSSub_MPT_T12_12_to0 is
  port( x : in  std_logic_vector(2 downto 0);
        r : out std_logic_vector(2 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_12_to0 is
begin
  with x select
    r <=
      "000" when "000", -- t[0] = 0
      "001" when "001", -- t[1] = 1
      "000" when "010", -- t[2] = 0
      "001" when "011", -- t[3] = 1
      "000" when "100", -- t[4] = 0
      "010" when "101", -- t[5] = 2
      "010" when "110", -- t[6] = 2
      "111" when "111", -- t[7] = 7
      "---" when others;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_12.all;

entity LNSSub_MPT_T12_12_to0_xor is
  port( a : in  std_logic_vector(1 downto 0);
        b : in  std_logic_vector(1 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_12_to0_xor is
  signal sign  : std_logic;
  signal in_t  : std_logic_vector(2 downto 0);
  signal out_t : std_logic_vector(2 downto 0);
begin
  sign <= not b(1);
  in_t(2 downto 1) <= a(1 downto 0);
  in_t(0) <= b(0) xor sign;

  inst_to0 : LNSSub_MPT_T12_12_to0
    port map( x => in_t,
              r => out_t );

  r(6 downto 3) <= (6 downto 3 => sign);
  r(0) <= out_t(0) xor sign;
  r(1) <= out_t(1) xor sign;
  r(2) <= out_t(2) xor sign;
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_12.all;

entity LNSSub_MPT_T12_12 is
  port( x : in  std_logic_vector(3 downto 0);
        r : out std_logic_vector(6 downto 0) );
end entity;

architecture arch of LNSSub_MPT_T12_12 is
  signal in_tiv  : std_logic_vector(1 downto 0);
  signal out_tiv : std_logic_vector(6 downto 0);
  signal a0      : std_logic_vector(1 downto 0);
  signal b0      : std_logic_vector(1 downto 0);
  signal out0    : std_logic_vector(6 downto 0);
  signal sum     : std_logic_vector(6 downto 0);
begin
  in_tiv <= x(3 downto 2);
  inst_tiv : LNSSub_MPT_T12_12_tiv
    port map( x => in_tiv,
              r => out_tiv );

  a0 <= x(3 downto 2);
  b0 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T12_12_to0_xor
    port map( a => a0,
              b => b0,
              r => out0 );


  sum <= out_tiv + out0;
  r <= sum(6 downto 0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_LNSSub_MPT_T12_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_T12_12_Clk is
  port( x   : in  std_logic_vector(3 downto 0);
        r   : out std_logic_vector(6 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_T12_12_Clk is
  signal in_tiv_1  : std_logic_vector(1 downto 0);
  signal out_tiv_1 : std_logic_vector(6 downto 0);
  signal out_tiv_2 : std_logic_vector(6 downto 0);
  signal a0_1      : std_logic_vector(1 downto 0);
  signal b0_1      : std_logic_vector(1 downto 0);
  signal out0_1    : std_logic_vector(6 downto 0);
  signal out0_2    : std_logic_vector(6 downto 0);
  signal psum1_2     : std_logic_vector(6 downto 0);
  signal psum1_3     : std_logic_vector(6 downto 0);
  signal psum2_2     : std_logic_vector(6 downto 0);
  signal psum2_3     : std_logic_vector(6 downto 0);
  signal sum_3     : std_logic_vector(6 downto 0);
begin
  in_tiv_1 <= x(3 downto 2);
  inst_tiv : LNSSub_MPT_T12_12_tiv
    port map( x => in_tiv_1,
              r => out_tiv_1 );

  a0_1 <= x(3 downto 2);
  b0_1 <= x(1 downto 0);
  inst_to0_xor : LNSSub_MPT_T12_12_to0_xor
    port map( a => a0_1,
              b => b0_1,
              r => out0_1 );

      out_tiv_2 <= out_tiv_1;
      out0_2    <= out0_1;

  psum1_2 <= out_tiv_2;
  psum2_2 <= out0_2;
  process(clk)
  begin
    if clk'event and clk='1' then
      psum1_3 <= psum1_2;
      psum2_3 <= psum2_2;
    end if;
  end process;
  sum_3 <= psum1_3 + psum2_3;
  r <= sum_3(6 downto 0);
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnssub_mpt_12.all;

entity LNSSub_MPT_12 is
  port( x : in  std_logic_vector(15 downto 0);
        r : out std_logic_vector(15 downto 0) );
end entity;

architecture arch of LNSSub_MPT_12 is

  signal out_t0 : std_logic_vector(5 downto 0);
  signal out_t1 : std_logic_vector(8 downto 0);
  signal out_t2 : std_logic_vector(10 downto 0);
  signal out_t3 : std_logic_vector(10 downto 0);
  signal out_t4 : std_logic_vector(10 downto 0);
  signal out_t5 : std_logic_vector(10 downto 0);
  signal out_t6 : std_logic_vector(9 downto 0);
  signal out_t7 : std_logic_vector(9 downto 0);
  signal out_t8 : std_logic_vector(8 downto 0);
  signal out_t9 : std_logic_vector(7 downto 0);
  signal out_t10 : std_logic_vector(6 downto 0);
  signal out_t11 : std_logic_vector(6 downto 0);
  signal out_t12 : std_logic_vector(6 downto 0);
begin
  inst_t0 : LNSSub_MPT_T0_12
    port map( x => x,
              r => out_t0 );

  inst_t1 : LNSSub_MPT_T1_12
    port map( x => x(13 downto 0),
              r => out_t1 );

  inst_t2 : LNSSub_MPT_T2_12
    port map( x => x(12 downto 0),
              r => out_t2 );

  inst_t3 : LNSSub_MPT_T3_12
    port map( x => x(11 downto 0),
              r => out_t3 );

  inst_t4 : LNSSub_MPT_T4_12
    port map( x => x(10 downto 0),
              r => out_t4 );

  inst_t5 : LNSSub_MPT_T5_12
    port map( x => x(9 downto 0),
              r => out_t5 );

  inst_t6 : LNSSub_MPT_T6_12
    port map( x => x(8 downto 0),
              r => out_t6 );

  inst_t7 : LNSSub_MPT_T7_12
    port map( x => x(7 downto 0),
              r => out_t7 );

  inst_t8 : LNSSub_MPT_T8_12
    port map( x => x(6 downto 0),
              r => out_t8 );

  inst_t9 : LNSSub_MPT_T9_12
    port map( x => x(5 downto 0),
              r => out_t9 );

  inst_t10 : LNSSub_MPT_T10_12
    port map( x => x(4 downto 0),
              r => out_t10 );

  inst_t11 : LNSSub_MPT_T11_12
    port map( x => x(3 downto 0),
              r => out_t11 );

  inst_t12 : LNSSub_MPT_T12_12
    port map( x => x(3 downto 0),
              r => out_t12 );

  r <= (15 downto 6 => '0') & out_t0
         when x(15 downto 15) /= (15 downto 15 => '1') else
       (15 downto 9 => '0') & out_t1
         when x(14) /= '1' else
       (15 downto 11 => '0') & out_t2
         when x(13) /= '1' else
       (15 downto 12 => '0') & out_t3 & (0 downto 0 => '0')
         when x(12) /= '1' else
       (15 downto 13 => '0') & out_t4 & (1 downto 0 => '0')
         when x(11) /= '1' else
       (15 downto 14 => '0') & out_t5 & (2 downto 0 => '0')
         when x(10) /= '1' else
       (15 downto 14 => '0') & out_t6 & (3 downto 0 => '0')
         when x(9) /= '1' else
       (15 downto 15 => '0') & out_t7 & (4 downto 0 => '0')
         when x(8) /= '1' else
       (15 downto 15 => '0') & out_t8 & (5 downto 0 => '0')
         when x(7) /= '1' else
       (15 downto 15 => '0') & out_t9 & (6 downto 0 => '0')
         when x(6) /= '1' else
       (15 downto 15 => '0') & out_t10 & (7 downto 0 => '0')
         when x(5) /= '1' else
       out_t11 & (8 downto 0 => '0')
         when x(4) /= '1' else
       out_t12 & (8 downto 0 => '0');
end architecture;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library fplib;
use fplib.pkg_lnssub_mpt_12.all;
use fplib.pkg_misc.all;

entity LNSSub_MPT_12_Clk is
  port( x   : in  std_logic_vector(15 downto 0);
        r   : out std_logic_vector(15 downto 0);
        clk : in  std_logic );
end entity;

architecture arch of LNSSub_MPT_12_Clk is
  signal x_1  : std_logic_vector(15 downto 0);
  signal x_10 : std_logic_vector(15 downto 0);

  signal out_t0_1  : std_logic_vector(5 downto 0);
  signal out_t0_10 : std_logic_vector(5 downto 0);
  signal out_t1_10 : std_logic_vector(8 downto 0);
  signal out_t2_10 : std_logic_vector(10 downto 0);
  signal out_t3_10 : std_logic_vector(10 downto 0);
  signal out_t4_10 : std_logic_vector(10 downto 0);
  signal out_t5_10 : std_logic_vector(10 downto 0);
  signal out_t6_10 : std_logic_vector(9 downto 0);
  signal out_t7_10 : std_logic_vector(9 downto 0);
  signal out_t8_10 : std_logic_vector(8 downto 0);
  signal out_t9_10 : std_logic_vector(7 downto 0);
  signal out_t10_10 : std_logic_vector(6 downto 0);
  signal out_t11_10 : std_logic_vector(6 downto 0);
  signal out_t12_10 : std_logic_vector(6 downto 0);
begin
  x_1 <= x;

  inst_t0 : LNSSub_MPT_T0_12
    port map( x   => x_1,
              r   => out_t0_1 );

  out_t0_delay : Delay
    generic map ( w => 6,
                  n => 1 )
    port map ( input  => out_t0_1,
               output => out_t0_10,
               clk    => clk );

  inst_t1 : LNSSub_MPT_T1_12_Clk
    port map( x   => x_1(13 downto 0),
              r   => out_t1_10,
              clk => clk );

  inst_t2 : LNSSub_MPT_T2_12_Clk
    port map( x   => x_1(12 downto 0),
              r   => out_t2_10,
              clk => clk );

  inst_t3 : LNSSub_MPT_T3_12_Clk
    port map( x   => x_1(11 downto 0),
              r   => out_t3_10,
              clk => clk );

  inst_t4 : LNSSub_MPT_T4_12_Clk
    port map( x   => x_1(10 downto 0),
              r   => out_t4_10,
              clk => clk );

  inst_t5 : LNSSub_MPT_T5_12_Clk
    port map( x   => x_1(9 downto 0),
              r   => out_t5_10,
              clk => clk );

  inst_t6 : LNSSub_MPT_T6_12_Clk
    port map( x   => x_1(8 downto 0),
              r   => out_t6_10,
              clk => clk );

  inst_t7 : LNSSub_MPT_T7_12_Clk
    port map( x   => x_1(7 downto 0),
              r   => out_t7_10,
              clk => clk );

  inst_t8 : LNSSub_MPT_T8_12_Clk
    port map( x   => x_1(6 downto 0),
              r   => out_t8_10,
              clk => clk );

  inst_t9 : LNSSub_MPT_T9_12_Clk
    port map( x   => x_1(5 downto 0),
              r   => out_t9_10,
              clk => clk );

  inst_t10 : LNSSub_MPT_T10_12_Clk
    port map( x   => x_1(4 downto 0),
              r   => out_t10_10,
              clk => clk );

  inst_t11 : LNSSub_MPT_T11_12_Clk
    port map( x   => x_1(3 downto 0),
              r   => out_t11_10,
              clk => clk );

  inst_t12 : LNSSub_MPT_T12_12_Clk
    port map( x   => x_1(3 downto 0),
              r   => out_t12_10,
              clk => clk );

  x_delay : Delay
    generic map ( w => 16,
                  n => 1 )
    port map ( input  => x_1,
               output => x_10,
               clk    => clk );

  r <= (15 downto 6 => '0') & out_t0_10
         when x_10(15 downto 15) /= (15 downto 15 => '1') else
       (15 downto 9 => '0') & out_t1_10
         when x_10(14) /= '1' else
       (15 downto 11 => '0') & out_t2_10
         when x_10(13) /= '1' else
       (15 downto 12 => '0') & out_t3_10 & (0 downto 0 => '0')
         when x_10(12) /= '1' else
       (15 downto 13 => '0') & out_t4_10 & (1 downto 0 => '0')
         when x_10(11) /= '1' else
       (15 downto 14 => '0') & out_t5_10 & (2 downto 0 => '0')
         when x_10(10) /= '1' else
       (15 downto 14 => '0') & out_t6_10 & (3 downto 0 => '0')
         when x_10(9) /= '1' else
       (15 downto 15 => '0') & out_t7_10 & (4 downto 0 => '0')
         when x_10(8) /= '1' else
       (15 downto 15 => '0') & out_t8_10 & (5 downto 0 => '0')
         when x_10(7) /= '1' else
       (15 downto 15 => '0') & out_t9_10 & (6 downto 0 => '0')
         when x_10(6) /= '1' else
       (15 downto 15 => '0') & out_t10_10 & (7 downto 0 => '0')
         when x_10(5) /= '1' else
       out_t11_10 & (8 downto 0 => '0')
         when x_10(4) /= '1' else
       out_t12_10 & (8 downto 0 => '0');
end architecture;
