-- Copyright 2003-2004 J�r�mie Detrey, Florent de Dinechin
--
-- This file is part of FPLibrary
--
-- FPLibrary is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- FPLibrary is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with FPLibrary; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA


library ieee;
use ieee.std_logic_1164.all;

-- ROM file for LNSAdd with wE = 8, wF = 23
entity Test_ROM is
  port ( addr   : in  std_logic_vector(9 downto 0);
         inVal  : out std_logic_vector(67 downto 0);
         outVal : out std_logic_vector(67 downto 0) );
end entity;

architecture arch of Test_ROM is
begin
with addr(9 downto 0) select
  inVal(67 downto 0) <=
    "00100000000000000000000000000000001001111111111111111111111111111111" when "0000000000",
    "00000000000000000000000000000000000110111101001100001011010111101100" when "0000000001",
    "01010110011110000111100001001000100101101011000110001001011001011110" when "0000000010",
    "11011111111111111111111111111111111111111111111111111111111111111111" when "0000000011",
    "00000000000000000000000000000000000101011101010011010000100101100100" when "0000000100",
    "10011111111111111111111111111111110101010100100111101101101110010100" when "0000000101",
    "00000000000000000000000000000000000110000101110010101000010101001111" when "0000000110",
    "00000000000000000000000000000000000100101101111001110011001111010101" when "0000000111",
    "01011100101110001110110110100011010110111001010011011100100011100010" when "0000001000",
    "11011111111111111111111111111111110100010110100010000101100101011101" when "0000001001",
    "00000000000000000000000000000000000101111000011100010000101110110100" when "0000001010",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "0000001011",
    "01001110110110010000010100011001110000000000000000000000000000000000" when "0000001100",
    "01100111000000100111011101101011100110011001010100010100011010001110" when "0000001101",
    "01000110111100101111010110001110110000000000000000000000000000000000" when "0000001110",
    "01001001110000111110010101011111000111100101100011100110111111000100" when "0000001111",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0000010000",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "0000010001",
    "01010010010111010101111101001110111101111111111111111111111111111111" when "0000010010",
    "00000000000000000000000000000000000111110010111100010000111010010001" when "0000010011",
    "01110000100001111100010011000110100110101000000110011000100111101111" when "0000010100",
    "01010000110100111001000000000010010101100011000100111000011001100000" when "0000010101",
    "10111111111111111111111111111111110110110101000110110100001110010101" when "0000010110",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "0000010111",
    "01110011100100111110110010111000101111111111111111111111111111111111" when "0000011000",
    "01101011100010110100011110010010100110011100000010011100011001000110" when "0000011001",
    "01000101011111101101101010000011110010000000000000000000000000000000" when "0000011010",
    "00100000000000000000000000000000000100101100000110000010110110010000" when "0000011011",
    "11111111111111111111111111111111110100010011101111000010000010001111" when "0000011100",
    "11111111111111111111111111111111110100011001011001101000101010010001" when "0000011101",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0000011110",
    "01111010110100101101111100001001100000000000000000000000000000000000" when "0000011111",
    "01010000001110100111101100011110001011111111111111111111111111111111" when "0000100000",
    "10011111111111111111111111111111110101101010100000100100001010100011" when "0000100001",
    "01000011111111000101011001111001110100001110110001101000100001111101" when "0000100010",
    "01010110011101001110111000110110111111111111111111111111111111111111" when "0000100011",
    "01010001010111011100010001100101110101100011111001110100010101001111" when "0000100100",
    "00000000000000000000000000000000000100100100111111000111110100001111" when "0000100101",
    "01100000011000101100110000000100010101110110101010011100010111100001" when "0000100110",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "0000100111",
    "01010001110001001000110010100111110111100111100011100100010101111101" when "0000101000",
    "00000000000000000000000000000000000110010010011101111110000000000000" when "0000101001",
    "01010000010011000000110100010100100110000101010101011101000110001000" when "0000101010",
    "11111111111111111111111111111111110101000110000001001010100010000110" when "0000101011",
    "11011111111111111111111111111111110111111011010010011001000000011011" when "0000101100",
    "01110011010100110111110010010110101011111111111111111111111111111111" when "0000101101",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0000101110",
    "01000101011110000001111011101011101001111111111111111111111111111111" when "0000101111",
    "11011111111111111111111111111111110101010010110010000111010010111111" when "0000110000",
    "11011111111111111111111111111111110101000111110110010000110110000101" when "0000110001",
    "01011111000101111000011011110101100010000000000000000000000000000000" when "0000110010",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0000110011",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0000110100",
    "01101010100100000000000000111001110010000000000000000000000000000000" when "0000110101",
    "01011111111101001000010001101001000000000000000000000000000000000000" when "0000110110",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0000110111",
    "11011111111111111111111111111111110100100111010011111010100001101011" when "0000111000",
    "01011110010100010000000111010010000110001010010111011100111101110000" when "0000111001",
    "11011111111111111111111111111111110110101011000001010101000000011000" when "0000111010",
    "01101001000111111100011011000111110000000000000000000000000000000000" when "0000111011",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "0000111100",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0000111101",
    "01110111000101000011010001011100101001111111111111111111111111111111" when "0000111110",
    "01011011100011110110100100001111010010000000000000000000000000000000" when "0000111111",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0001000000",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "0001000001",
    "10011111111111111111111111111111110111011101100011110001000100100100" when "0001000010",
    "01010110110010001111001001111111100100111010111010010001011001110111" when "0001000011",
    "00000000000000000000000000000000000100111110111100010101010111011100" when "0001000100",
    "01010010101001001100101101101111010010000000000000000000000000000000" when "0001000101",
    "11111111111111111111111111111111110100100001011111000010101011110110" when "0001000110",
    "01110011101111101010000101101111010000000000000000000000000000000000" when "0001000111",
    "10111111111111111111111111111111110100100111000000101001111010100110" when "0001001000",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0001001001",
    "01011111001100100000100111101111111111111111111111111111111111111111" when "0001001010",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "0001001011",
    "01110111010011011101110101110100100110011010101011101110011000111000" when "0001001100",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "0001001101",
    "01001100110010000000110111100001011101111111111111111111111111111111" when "0001001110",
    "01100001001010001100001010110011010100001111100011101101100001100010" when "0001001111",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "0001010000",
    "01001100010101000100000010110001000000000000000000000000000000000000" when "0001010001",
    "01101010110011010000011011101110100000000000000000000000000000000000" when "0001010010",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "0001010011",
    "01111010110000000000011000000110110101101011110111000001100110010001" when "0001010100",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0001010101",
    "01100011100110000011111011001101000000000000000000000000000000000000" when "0001010110",
    "01001010101011001000010000001010111001111111111111111111111111111111" when "0001010111",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0001011000",
    "01000000010001100101010110100110101011111111111111111111111111111111" when "0001011001",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "0001011010",
    "10111111111111111111111111111111110101110110001001110100100000100100" when "0001011011",
    "11011111111111111111111111111111110100100110010100001001010111111010" when "0001011100",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "0001011101",
    "01100000001011110001101110101001101001111111111111111111111111111111" when "0001011110",
    "00000000000000000000000000000000000101101000011100101011100001000011" when "0001011111",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0001100000",
    "01010100111000110010111010001100100110000100100100000110101100110111" when "0001100001",
    "01011010111101011101001100000010110000000000000000000000000000000000" when "0001100010",
    "01111101000100111011101010100011000100000100011000110001010101110010" when "0001100011",
    "00100000000000000000000000000000000110001001100111010000110000000100" when "0001100100",
    "01010000011001011000111011101011010000000000000000000000000000000000" when "0001100101",
    "00100000000000000000000000000000001001111111111111111111111111111111" when "0001100110",
    "01100011000111110011101111001001010000000000000000000000000000000000" when "0001100111",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "0001101000",
    "01010111010101000001101101000011100100111010011101100101001001100011" when "0001101001",
    "00000000000000000000000000000000000111010100011111000001101010111101" when "0001101010",
    "01110001101100111001111010101001100101000101111011110010111111001110" when "0001101011",
    "00000000000000000000000000000000000110100101011100101011001101010010" when "0001101100",
    "00000000000000000000000000000000000110101000111111011101110011100100" when "0001101101",
    "01000100100110010100001000111110010000000000000000000000000000000000" when "0001101110",
    "01100000100101100011001011111111110110111011001000010100000000110110" when "0001101111",
    "01001100000101010101101111110001000100001000011110110101110001001001" when "0001110000",
    "00000000000000000000000000000000000110111000110110110110110011100011" when "0001110001",
    "01001110100111100101111101000000101011111111111111111111111111111111" when "0001110010",
    "10111111111111111111111111111111111101111111111111111111111111111111" when "0001110011",
    "01011010101100011111111001001111110000000000000000000000000000000000" when "0001110100",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0001110101",
    "01000110111111110110111011110101100000000000000000000000000000000000" when "0001110110",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "0001110111",
    "10111111111111111111111111111111110100001111000011011010100000000001" when "0001111000",
    "01011001010100000101011001001001010110110000100110100110010100101000" when "0001111001",
    "11011111111111111111111111111111110111110000111100111101110011101010" when "0001111010",
    "01111110001000001000010010101111111001111111111111111111111111111111" when "0001111011",
    "01000110001111001101011111001111100100111110011110001000010010011010" when "0001111100",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "0001111101",
    "01111100111010010011101101011010010000000000000000000000000000000000" when "0001111110",
    "01110001100110011111111101000011110100100100010011100101101110011111" when "0001111111",
    "01111011011001011001011100100010011111111111111111111111111111111111" when "0010000000",
    "00000000000000000000000000000000000111110000000110010110100000100110" when "0010000001",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "0010000010",
    "00000000000000000000000000000000000101100101111000111111110110100001" when "0010000011",
    "01111100101010100100010100011001100111100011101011111111000001010011" when "0010000100",
    "01001100001110111111100100110111100110011011111100010011100010011110" when "0010000101",
    "00100000000000000000000000000000000100101110101110110101111111110100" when "0010000110",
    "00100000000000000000000000000000000110100000011101000100110111101011" when "0010000111",
    "01101000110010100000110101001011010101000010111000111011010010011101" when "0010001000",
    "01111110011010010001101000111001100000000000000000000000000000000000" when "0010001001",
    "01100010100101010101000010001011000000000000000000000000000000000000" when "0010001010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0010001011",
    "01110101101010010100100000011010010100011100110011011001011001010110" when "0010001100",
    "01011011011111111010000000000100111011111111111111111111111111111111" when "0010001101",
    "00000000000000000000000000000000000111110101100111001011100101011010" when "0010001110",
    "10011111111111111111111111111111110110100011011000011011011111010100" when "0010001111",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0010010000",
    "01100011011010110101010110000111100111011011110101010001000011110110" when "0010010001",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "0010010010",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "0010010011",
    "01110000101111000100100111000100000110110100010000000001110010010001" when "0010010100",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0010010101",
    "01000110101100110000000000111010100101110110100100010111000111000011" when "0010010110",
    "10011111111111111111111111111111110101100010000100110011111101110011" when "0010010111",
    "01110101001000000101011000011001001011111111111111111111111111111111" when "0010011000",
    "01001101010101111111101110000100110010000000000000000000000000000000" when "0010011001",
    "01011010000010001010010101011010110101011101100010000111011011001001" when "0010011010",
    "01101001110100010110110010100001000111011010111110000010010000111001" when "0010011011",
    "01111001100010100111000111110101110101011100000010100101000011100111" when "0010011100",
    "00000000000000000000000000000000000100110011111111100111001101110111" when "0010011101",
    "10011111111111111111111111111111110100100011001111001010010011011000" when "0010011110",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0010011111",
    "01010111111011110101011000100101010111010111100101000010101111010010" when "0010100000",
    "11111111111111111111111111111111110110011110011001110001000110010100" when "0010100001",
    "01100010000111001101010100101100111001111111111111111111111111111111" when "0010100010",
    "01011011011001011000000100111000100000000000000000000000000000000000" when "0010100011",
    "01111100100110100101011001011100000101111100110111111101000100011100" when "0010100100",
    "01100011111000000101001001101011010000000000000000000000000000000000" when "0010100101",
    "01100100001111110111011011110100110000000000000000000000000000000000" when "0010100110",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0010100111",
    "01110011001010100001111101011100110101111111010010000000011001000010" when "0010101000",
    "01011001100100110100010001001100001011111111111111111111111111111111" when "0010101001",
    "11111111111111111111111111111111110101000111101100100101001010011010" when "0010101010",
    "10011111111111111111111111111111110101100110010101011011011111111101" when "0010101011",
    "00000000000000000000000000000000000101010100011100110101100100100100" when "0010101100",
    "11111111111111111111111111111111111101111111111111111111111111111111" when "0010101101",
    "01110110010010000001110010011011000010000000000000000000000000000000" when "0010101110",
    "11011111111111111111111111111111110101010100111001100000001010110010" when "0010101111",
    "11111111111111111111111111111111110110101110000011111110111111000110" when "0010110000",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "0010110001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0010110010",
    "01000000100001010110011101110010110000000000000000000000000000000000" when "0010110011",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0010110100",
    "11111111111111111111111111111111110100100000100100000001110011011000" when "0010110101",
    "01011100011000000101100100000010111101111111111111111111111111111111" when "0010110110",
    "01010101110010110010100001011000011001111111111111111111111111111111" when "0010110111",
    "00000000000000000000000000000000000111101010011110101001100110010010" when "0010111000",
    "00000000000000000000000000000000000111101010100010010000011001010111" when "0010111001",
    "00100000000000000000000000000000000101110101010111010010011111000100" when "0010111010",
    "01110010001101111001000100011001010111001100110001000101111100010010" when "0010111011",
    "11111111111111111111111111111111110111000010001101001100000111010110" when "0010111100",
    "00100000000000000000000000000000000111011000111110010001100110000000" when "0010111101",
    "01111000000001000011111101101111110000000000000000000000000000000000" when "0010111110",
    "01010100001110100111110110100001010110101101111100010010111010000000" when "0010111111",
    "01111010011010101110110110100000010100100101010111110001110010011100" when "0011000000",
    "01101101111001010101011010110110010111011011101101101000100111011111" when "0011000001",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0011000010",
    "01110101000101011000000111110111000100001100111000110011111110011000" when "0011000011",
    "11011111111111111111111111111111110111110100001110101011011101010111" when "0011000100",
    "01100111010010110111001110000110000111010110001110100011000010001001" when "0011000101",
    "00100000000000000000000000000000000100110011010110001011010011110010" when "0011000110",
    "01100110010100000100010101110000000010000000000000000000000000000000" when "0011000111",
    "01110000010011001111100101110111110101110111001100111111110011011110" when "0011001000",
    "01001011000111010001010010111010110111100101001010101010010101110011" when "0011001001",
    "01100011010011110101100100101001010000000000000000000000000000000000" when "0011001010",
    "01110011111110010001100101111010110110011010100001110101010010101111" when "0011001011",
    "00000000000000000000000000000000000111100011100001110001001011010100" when "0011001100",
    "10111111111111111111111111111111111101111111111111111111111111111111" when "0011001101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011001110",
    "10011111111111111111111111111111110101000101111010000010110011001000" when "0011001111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011010000",
    "01001110010101110111100000101001010111100001001001011000000011110010" when "0011010001",
    "00100000000000000000000000000000000101001100110101010111100011010100" when "0011010010",
    "01101110000100100011100110101111111001111111111111111111111111111111" when "0011010011",
    "01000000111111011111001001011101001011111111111111111111111111111111" when "0011010100",
    "01110011101001001011110111100101000111000010001001010110101111101000" when "0011010101",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0011010110",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0011010111",
    "01011110100111100100100001010011010000000000000000000000000000000000" when "0011011000",
    "01010000101110011010100110101110000101100111101100101010101000000001" when "0011011001",
    "01001110101000111001111001011101100010000000000000000000000000000000" when "0011011010",
    "01110101001010111000001101111101110100110010011110000111010100101100" when "0011011011",
    "01100100110011100001101011010111000100011101100100011000110101110000" when "0011011100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011011101",
    "01001000011011010100100000000000101001111111111111111111111111111111" when "0011011110",
    "01010010100010101011100110110110010100110100000111011100000100010101" when "0011011111",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0011100000",
    "11011111111111111111111111111111110110000110000010011101000011101000" when "0011100001",
    "01101101110000010101011111110111110110101010101100111000000101101011" when "0011100010",
    "00000000000000000000000000000000000111111100110000110110111110110000" when "0011100011",
    "11011111111111111111111111111111110101101100110111001110101011100100" when "0011100100",
    "01110000111001001101110001110101010000000000000000000000000000000000" when "0011100101",
    "11111111111111111111111111111111110101110111111000011001111000001011" when "0011100110",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0011100111",
    "01110001010101011011100010110101010110110010110111101101000101011000" when "0011101000",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0011101001",
    "01111000000000000110011000110011011001111111111111111111111111111111" when "0011101010",
    "01000101001110010111001110011010000101110101101001011001011001001001" when "0011101011",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0011101100",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0011101101",
    "01000101000001010010111000110001110101001011001011110001110000010110" when "0011101110",
    "11111111111111111111111111111111111001111111111111111111111111111111" when "0011101111",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0011110000",
    "11111111111111111111111111111111110111010011000000001111001001001010" when "0011110001",
    "01011100011011110111011001001100100111110001110000001011000110101101" when "0011110010",
    "01001001011111111111000010100011100110011110001101111101111110001011" when "0011110011",
    "01110000101100010101111100110010000010000000000000000000000000000000" when "0011110100",
    "01000101110000000010000100100000111101111111111111111111111111111111" when "0011110101",
    "01111110001111101011101101001001001001111111111111111111111111111111" when "0011110110",
    "01110100000001101100100000100011000000000000000000000000000000000000" when "0011110111",
    "00100000000000000000000000000000000110011010011010111010110100100000" when "0011111000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011111001",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "0011111010",
    "01001100111000100001110111001101110010000000000000000000000000000000" when "0011111011",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0011111100",
    "00000000000000000000000000000000000110010011010100100011101101010110" when "0011111101",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0011111110",
    "10111111111111111111111111111111111111111111111111111111111111111111" when "0011111111",
    "11111111111111111111111111111111111001111111111111111111111111111111" when "0100000000",
    "01101011011101011000000011000100011001111111111111111111111111111111" when "0100000001",
    "00100000000000000000000000000000000111010000010010101000100000001011" when "0100000010",
    "10011111111111111111111111111111110100010101111000101101001001010101" when "0100000011",
    "01000111111111111000111000000100100100001110010110111110010000110100" when "0100000100",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "0100000101",
    "01011101111111100111001011011000010110010100001110011110001000001110" when "0100000110",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "0100000111",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "0100001000",
    "01100110000001010010111011000001010101110000010110000011010100011110" when "0100001001",
    "01001010001010100011100100010011110000000000000000000000000000000000" when "0100001010",
    "01010111100100110101100101000110010111011101101000110011010001111100" when "0100001011",
    "01110101010001011101101000001011010000000000000000000000000000000000" when "0100001100",
    "10111111111111111111111111111111110101011000010100111100101100110010" when "0100001101",
    "10011111111111111111111111111111110111001100010110100110100100001010" when "0100001110",
    "00000000000000000000000000000000000111001010101011111111000001111101" when "0100001111",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "0100010000",
    "00000000000000000000000000000000000100001010010101000001110000100101" when "0100010001",
    "01000101000111001000001000100100000110010100110000101011000111000000" when "0100010010",
    "01101101001101011010110000101111110010000000000000000000000000000000" when "0100010011",
    "01111111101001111000101001110110001111111111111111111111111111111111" when "0100010100",
    "01001010011110111010000000010001010010000000000000000000000000000000" when "0100010101",
    "01011010010111000100101000100000110111000100000100111010011010111011" when "0100010110",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0100010111",
    "00100000000000000000000000000000000110111010010101001110011001011111" when "0100011000",
    "01011100000001010010110101011101100110000101010100110010101100011111" when "0100011001",
    "01001011010100001011100101001100110101101110111100010100011000001010" when "0100011010",
    "01110010101001101110101001010010010101001110101011100101101110111010" when "0100011011",
    "01001101011111011111111001011101000010000000000000000000000000000000" when "0100011100",
    "10011111111111111111111111111111110110000101000100000001011001010011" when "0100011101",
    "00100000000000000000000000000000000111010010100111010111101010101111" when "0100011110",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0100011111",
    "11111111111111111111111111111111111111111111111111111111111111111111" when "0100100000",
    "11111111111111111111111111111111111001111111111111111111111111111111" when "0100100001",
    "11011111111111111111111111111111110101000000101110101001101011001000" when "0100100010",
    "01110000011011110010011001011100000110100000000100011101001001110100" when "0100100011",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "0100100100",
    "01011010101100101101001001111111110000000000000000000000000000000000" when "0100100101",
    "01011110011011011000000100111001010101011110100111000001011000000110" when "0100100110",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "0100100111",
    "00100000000000000000000000000000000111010000111111101011110000010111" when "0100101000",
    "01001111011101100000101011001001100101011100010111111011011011001000" when "0100101001",
    "01011111111001110001010001101010100110100001001011110110010110111001" when "0100101010",
    "01101000100101011011010100001010110100111011011100111011101101100000" when "0100101011",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0100101100",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0100101101",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "0100101110",
    "01011011110010011001100001101000101111111111111111111111111111111111" when "0100101111",
    "01101001001010010011100111111111100010000000000000000000000000000000" when "0100110000",
    "11111111111111111111111111111111110110101111111101110001100101011001" when "0100110001",
    "10111111111111111111111111111111110101110000000101011110011011100100" when "0100110010",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0100110011",
    "01110100100100011110101000001000000110110011111000011010111101111001" when "0100110100",
    "01000011000010010010100100111010100000000000000000000000000000000000" when "0100110101",
    "11111111111111111111111111111111110101111110011011100111010110001000" when "0100110110",
    "01010101010101101010010011010001010101000011000011010010011111010110" when "0100110111",
    "01000110011100001010100011101001010101110010100100001000100000100001" when "0100111000",
    "01011111010011000010111110010011011001111111111111111111111111111111" when "0100111001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0100111010",
    "01011101110101101001010001111111010010000000000000000000000000000000" when "0100111011",
    "10111111111111111111111111111111110100000001011110110100001000011010" when "0100111100",
    "01000111000011111101001101010110010111111010010011101000010111101001" when "0100111101",
    "01001011010101010010010000011110010111011011110111101101011101101010" when "0100111110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0100111111",
    "10011111111111111111111111111111110111110100010011001001110010010110" when "0101000000",
    "01000010101101010001011111100011101111111111111111111111111111111111" when "0101000001",
    "01001010100011111110100000101000100100011110100001111100000001110000" when "0101000010",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0101000011",
    "10111111111111111111111111111111110100011101010000110101100101000001" when "0101000100",
    "10011111111111111111111111111111111101111111111111111111111111111111" when "0101000101",
    "01111100100011011110101010110101010100111000110111100101110010000001" when "0101000110",
    "01000101000100101111111000110010010110111100000010010010111010111101" when "0101000111",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0101001000",
    "11011111111111111111111111111111110101111000110101000110010100010001" when "0101001001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0101001010",
    "01100100001001001000101110011111100110101100010111111111001101100001" when "0101001011",
    "01101011000011001100000000101000010000000000000000000000000000000000" when "0101001100",
    "01000111101101101111001100011110110000000000000000000000000000000000" when "0101001101",
    "01001100010110101100100110010001000000000000000000000000000000000000" when "0101001110",
    "10011111111111111111111111111111110111111011001101010000000001111111" when "0101001111",
    "01111000000011111011010011100010100101001101100010111111110001100101" when "0101010000",
    "01101100101110011011110111000000010000000000000000000000000000000000" when "0101010001",
    "00000000000000000000000000000000000101000011110000101001000010101000" when "0101010010",
    "01000000110001110011010100100011011011111111111111111111111111111111" when "0101010011",
    "01100111101111101011111111000011100100110111100100011100110100011111" when "0101010100",
    "01001001011000101110001011001100101111111111111111111111111111111111" when "0101010101",
    "10011111111111111111111111111111110101110101111100011010000111101111" when "0101010110",
    "01010111010000011100010111000001000100001101011001000110010000011001" when "0101010111",
    "11111111111111111111111111111111110100110111010011110010011111000000" when "0101011000",
    "01100000000001010001110011011011000110000001011011101001001001111111" when "0101011001",
    "00000000000000000000000000000000000100101000110010110001011111000010" when "0101011010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0101011011",
    "01011010011010100111011010110101010100001100011010110001100001000111" when "0101011100",
    "00000000000000000000000000000000000110101111111101101101010010001000" when "0101011101",
    "01001011110111110101100100001110110000000000000000000000000000000000" when "0101011110",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "0101011111",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "0101100000",
    "00100000000000000000000000000000000101101100011001010000000101001000" when "0101100001",
    "01100100110101101100000111000010000010000000000000000000000000000000" when "0101100010",
    "00000000000000000000000000000000000110101100010000011001010111011101" when "0101100011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101100100",
    "01110111001001110100100010011110010101010110101101100001111100101011" when "0101100101",
    "10111111111111111111111111111111110101111010110011001100101010100100" when "0101100110",
    "10111111111111111111111111111111110110100001010101010011100000010001" when "0101100111",
    "01110100000100010100111110100000000000000000000000000000000000000000" when "0101101000",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "0101101001",
    "10111111111111111111111111111111111111111111111111111111111111111111" when "0101101010",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0101101011",
    "01010000110001111001001010100001111001111111111111111111111111111111" when "0101101100",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0101101101",
    "01011000011011000000011001101001000110000100000001100001111000101000" when "0101101110",
    "01110111101010100100001110111011000110000000001111001000010100101100" when "0101101111",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0101110000",
    "01101011001100101000111111010111101101111111111111111111111111111111" when "0101110001",
    "01100111110101111110000000100110100010000000000000000000000000000000" when "0101110010",
    "11111111111111111111111111111111111111111111111111111111111111111111" when "0101110011",
    "01010010010010100101101110000101100010000000000000000000000000000000" when "0101110100",
    "01101001111011010010011101001011111101111111111111111111111111111111" when "0101110101",
    "01100101011000001111110011111111110111011010110000100000101110111011" when "0101110110",
    "11011111111111111111111111111111110100110101101000101001010100100011" when "0101110111",
    "00100000000000000000000000000000000110111110000100000001111110010101" when "0101111000",
    "10111111111111111111111111111111110100100000111100100100010100001100" when "0101111001",
    "01010110100010100100000000101000101111111111111111111111111111111111" when "0101111010",
    "01101011011110110001101001011000100000000000000000000000000000000000" when "0101111011",
    "11011111111111111111111111111111110101101110011110011101110101000011" when "0101111100",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0101111101",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "0101111110",
    "00000000000000000000000000000000000101011100001000010111100000101111" when "0101111111",
    "01111000001111100110010001111100100101001000001101100100010011001100" when "0110000000",
    "01000100101110100100100110000110111011111111111111111111111111111111" when "0110000001",
    "00100000000000000000000000000000001001111111111111111111111111111111" when "0110000010",
    "00000000000000000000000000000000000111111100101101111100001000101111" when "0110000011",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "0110000100",
    "11111111111111111111111111111111111101111111111111111111111111111111" when "0110000101",
    "10011111111111111111111111111111110110000001101011000001000000001101" when "0110000110",
    "01101011010101100001000001111110001111111111111111111111111111111111" when "0110000111",
    "11111111111111111111111111111111110110000000100010001100111001001100" when "0110001000",
    "01001001110000011000100101111111011011111111111111111111111111111111" when "0110001001",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "0110001010",
    "01001011010111000101111111001010101111111111111111111111111111111111" when "0110001011",
    "00100000000000000000000000000000000101001100011001111010000111000101" when "0110001100",
    "01101000001011111000111101111000100101010110100101010011111100101111" when "0110001101",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "0110001110",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "0110001111",
    "01010001110000100001001000110000011011111111111111111111111111111111" when "0110010000",
    "00100000000000000000000000000000000111100010110100110101011000011111" when "0110010001",
    "01010111011011101100011010000111100101101101101111011100110000111000" when "0110010010",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0110010011",
    "10111111111111111111111111111111110111110101010011001110111000001010" when "0110010100",
    "01000001010100010101110110111101010100011011101111100011111000101010" when "0110010101",
    "11111111111111111111111111111111111111111111111111111111111111111111" when "0110010110",
    "01101010010011010101111111101001110010000000000000000000000000000000" when "0110010111",
    "01111000010100011011010000101100001011111111111111111111111111111111" when "0110011000",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0110011001",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "0110011010",
    "10111111111111111111111111111111110111011110000001001001001110110100" when "0110011011",
    "01101011111011111111101110000010110010000000000000000000000000000000" when "0110011100",
    "01101110101011011010001111010110100010000000000000000000000000000000" when "0110011101",
    "01100000010110110110011000001001000101010000000011001101101011001001" when "0110011110",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0110011111",
    "01001111010110001001101101010010000111111001001110010101010000001111" when "0110100000",
    "01110010110100010000001100101011000101010100100010011100111001000111" when "0110100001",
    "00000000000000000000000000000000000101001111100011100101101110100101" when "0110100010",
    "11111111111111111111111111111111110110101111001110011100011010011011" when "0110100011",
    "11011111111111111111111111111111110101111111000011000000111001011100" when "0110100100",
    "01100111011010100000001111111100111011111111111111111111111111111111" when "0110100101",
    "01000110100001001001011000010111100100110000100111110110110000001100" when "0110100110",
    "00000000000000000000000000000000000110110111111000000110010101001011" when "0110100111",
    "01001111011101000101010000110011010000000000000000000000000000000000" when "0110101000",
    "01001000100111110110100111101111010000000000000000000000000000000000" when "0110101001",
    "10111111111111111111111111111111110111110000001000101111000111000100" when "0110101010",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "0110101011",
    "01011110010011111010011010111111100101110010111101011110110110011000" when "0110101100",
    "01101010110011100111001100111010100100101000110001001010000011111010" when "0110101101",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "0110101110",
    "01111110010100011101011010101110000010000000000000000000000000000000" when "0110101111",
    "00100000000000000000000000000000000110111110000111010001101110011100" when "0110110000",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "0110110001",
    "01101011101100111110011101111110010111011110101110011110100101000000" when "0110110010",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "0110110011",
    "01010101010011111010011010100100100111111100100110110010010111011111" when "0110110100",
    "11111111111111111111111111111111111101111111111111111111111111111111" when "0110110101",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "0110110110",
    "01001011011110011100110011000001110000000000000000000000000000000000" when "0110110111",
    "01011000111011111010110101110110000110011000000101110000010001010101" when "0110111000",
    "00100000000000000000000000000000000101110011100010110101010010001100" when "0110111001",
    "01111100101000010001001011011100000000000000000000000000000000000000" when "0110111010",
    "01000100101010011001110100111011100100001001111111110111100100110000" when "0110111011",
    "01010110010001100010110010110100010010000000000000000000000000000000" when "0110111100",
    "00100000000000000000000000000000000111011110101100000001101111001000" when "0110111101",
    "01110100111010101101001100011000000010000000000000000000000000000000" when "0110111110",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "0110111111",
    "10011111111111111111111111111111110100110111100011011110110011011000" when "0111000000",
    "01001111111000101111010110111110010110000001111000001010011010101000" when "0111000001",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "0111000010",
    "01100001110011010111101000011001000111110010011110111001101010100000" when "0111000011",
    "01011100010000100110111010010011100101001010010100111001001110101011" when "0111000100",
    "01000010101000000001010100001011100000000000000000000000000000000000" when "0111000101",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0111000110",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0111000111",
    "01010001110111111000100011001100101101111111111111111111111111111111" when "0111001000",
    "01001001110000101110000110000010110100111010000111010000100011001011" when "0111001001",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0111001010",
    "00100000000000000000000000000000000111001111011100010011011100101001" when "0111001011",
    "01100011101111111101001111000000100101000010001110110001000000101100" when "0111001100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111001101",
    "01110010000010111111101100100110010111000111110101110011110111010101" when "0111001110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111001111",
    "01000001011001101101101101011110000010000000000000000000000000000000" when "0111010000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111010001",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0111010010",
    "01000110100111110111101011000010101011111111111111111111111111111111" when "0111010011",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "0111010100",
    "01101011001111010110100101000110010000000000000000000000000000000000" when "0111010101",
    "01001010110011011101111110001100010101001000010101010100000110011110" when "0111010110",
    "01010011101100101100100100111100010101110100101000101001110101000001" when "0111010111",
    "00000000000000000000000000000000000110010011110110000110010111011101" when "0111011000",
    "00100000000000000000000000000000000110100100001001110111101001010101" when "0111011001",
    "01000111000101110101100011011110110100110001100000011010010000100111" when "0111011010",
    "01000000111001011101011011110101001011111111111111111111111111111111" when "0111011011",
    "00000000000000000000000000000000000100110110110101100100110001111001" when "0111011100",
    "01001100001100100011010110000001010100110011000101100001111100000010" when "0111011101",
    "10011111111111111111111111111111110110010111010001110101011001011011" when "0111011110",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "0111011111",
    "01111000101001110111001101100110100010000000000000000000000000000000" when "0111100000",
    "01000110000010001000011110111000001111111111111111111111111111111111" when "0111100001",
    "01100110010010101010001101001001000100101011100010110101001011011011" when "0111100010",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "0111100011",
    "00100000000000000000000000000000000111001111011110001010110100111111" when "0111100100",
    "11111111111111111111111111111111110111010011111111000110011011100001" when "0111100101",
    "00100000000000000000000000000000001001111111111111111111111111111111" when "0111100110",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "0111100111",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "0111101000",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "0111101001",
    "01010010100111010001101110001000010100010101011100101010101011010111" when "0111101010",
    "01001111110100010011100001000110000000000000000000000000000000000000" when "0111101011",
    "10011111111111111111111111111111110101001001111010111000000010111000" when "0111101100",
    "01001001001110000101100010000101011111111111111111111111111111111111" when "0111101101",
    "01010100111101110000101101010111010000000000000000000000000000000000" when "0111101110",
    "01010100101010110001000110000101100100000010001111010010111000001110" when "0111101111",
    "11111111111111111111111111111111110100111100010111110001111000100111" when "0111110000",
    "01001011100111000001000011100000010101001001111000111100011000100100" when "0111110001",
    "01011110110101001001101010110101010100101100111111011110110101011001" when "0111110010",
    "11111111111111111111111111111111111011111111111111111111111111111111" when "0111110011",
    "01011100111011010101100011100000101111111111111111111111111111111111" when "0111110100",
    "10011111111111111111111111111111111101111111111111111111111111111111" when "0111110101",
    "00000000000000000000000000000000000101011111001110100000111101110001" when "0111110110",
    "00000000000000000000000000000000000100101100001100010000011000101110" when "0111110111",
    "10111111111111111111111111111111110101000101100001110110100000010101" when "0111111000",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "0111111001",
    "01000010000101110010100001111101000100100100000111100110110101011010" when "0111111010",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "0111111011",
    "01000011011110000100100001101111110010000000000000000000000000000000" when "0111111100",
    "01001100101100111010101011000100101001111111111111111111111111111111" when "0111111101",
    "01011010111000010110011000001011100010000000000000000000000000000000" when "0111111110",
    "01100000001010111100100110111101100111111100011101110100001100011101" when "0111111111",
    "01011111100011010110010001000010011011111111111111111111111111111111" when "1000000000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1000000001",
    "01001010000110100111000101111001100000000000000000000000000000000000" when "1000000010",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "1000000011",
    "01100101110001010010011010110110010110110010010111001001100000101100" when "1000000100",
    "01011101001110111100011100010000001101111111111111111111111111111111" when "1000000101",
    "01010110100010001111010110001100100101100100111100100110111001001101" when "1000000110",
    "10011111111111111111111111111111110100000110000100011001001010010001" when "1000000111",
    "11011111111111111111111111111111110101101010111000011010001010111000" when "1000001000",
    "00100000000000000000000000000000000100001101010001110010101101110011" when "1000001001",
    "01101000001011001111010101000110000101010010011110000101110011110011" when "1000001010",
    "01100001100101011111000000110110110010000000000000000000000000000000" when "1000001011",
    "01000000000001010000110000110110100100110010100101100101101011001010" when "1000001100",
    "01111111101100011100111010101011110000000000000000000000000000000000" when "1000001101",
    "00000000000000000000000000000000000101100001111000111001110010000111" when "1000001110",
    "10111111111111111111111111111111110110011000001001101011001111000001" when "1000001111",
    "01110011010111011110111000010010110101010101001001001101100111000000" when "1000010000",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1000010001",
    "11111111111111111111111111111111110100100110101011010111110110001111" when "1000010010",
    "01101011100011111010100111011011000110000100001100111011110110110110" when "1000010011",
    "00000000000000000000000000000000000110000001111011101000110101000100" when "1000010100",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1000010101",
    "01110001111111101111001011100011001111111111111111111111111111111111" when "1000010110",
    "01110101010101101011000011101111010000000000000000000000000000000000" when "1000010111",
    "10111111111111111111111111111111111111111111111111111111111111111111" when "1000011000",
    "01011101011100001000011000101010100100001010001000010001001000001111" when "1000011001",
    "01011100001000000110101111110010100111000110110101011001101101101110" when "1000011010",
    "01010001101011001000101111101111000111011001110110110100100000001001" when "1000011011",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1000011100",
    "01000101000111000111011110010111101001111111111111111111111111111111" when "1000011101",
    "00100000000000000000000000000000000101010110111010011010001010110001" when "1000011110",
    "00100000000000000000000000000000000111111010000100100100011111010011" when "1000011111",
    "01100100000001110000101000111110110111010110010011111010100111010111" when "1000100000",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "1000100001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1000100010",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1000100011",
    "01110110100101110100100110001101110110010010001000100111010100110011" when "1000100100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000100101",
    "01011111101101011110111101100000000000000000000000000000000000000000" when "1000100110",
    "01001000111000011001001011111101011011111111111111111111111111111111" when "1000100111",
    "00000000000000000000000000000000000110110100011110100010011011111011" when "1000101000",
    "01110001011110101111100110111100011011111111111111111111111111111111" when "1000101001",
    "11111111111111111111111111111111110111100000100000110001110000100011" when "1000101010",
    "00100000000000000000000000000000000100100110100011101001000010100010" when "1000101011",
    "01100011010110011110001000000000111111111111111111111111111111111111" when "1000101100",
    "01101100010000001000000000010110010110000001010001111010001000011011" when "1000101101",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "1000101110",
    "01110100001111110101000111101110001011111111111111111111111111111111" when "1000101111",
    "11111111111111111111111111111111110111000101010110111001001111100011" when "1000110000",
    "00000000000000000000000000000000000110011111001011000111000100100011" when "1000110001",
    "01011110100011011001000001101001100101000101110110100001101100110110" when "1000110010",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "1000110011",
    "01110011110001010100111111011001110000000000000000000000000000000000" when "1000110100",
    "01000010001011010111100101001111110110110010011010101100101101100110" when "1000110101",
    "11111111111111111111111111111111110101001101100010111110000010100001" when "1000110110",
    "01011110000101110010001101111000110111011101000000010010010000101111" when "1000110111",
    "00100000000000000000000000000000000101111010011000011001100110101101" when "1000111000",
    "11111111111111111111111111111111110100011111010101010010011001000001" when "1000111001",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1000111010",
    "01000110011101010001111101000111110110010011111000001110010101000010" when "1000111011",
    "11011111111111111111111111111111110100101000100111011111101001100001" when "1000111100",
    "01111000011011100101001110111011100111010001001001101101110100010101" when "1000111101",
    "01100010100000110100101111010100000000000000000000000000000000000000" when "1000111110",
    "01010001111111011011101001110000101101111111111111111111111111111111" when "1000111111",
    "00100000000000000000000000000000000111100101110000011111100000011011" when "1001000000",
    "01101111111110100010100000110000111101111111111111111111111111111111" when "1001000001",
    "01010011101110001111111100101010100101101011101101100111100010110101" when "1001000010",
    "11111111111111111111111111111111111111111111111111111111111111111111" when "1001000011",
    "00100000000000000000000000000000000101110111100110101010100110110010" when "1001000100",
    "01001011101001111100111000100011100100101110011110101111010001101101" when "1001000101",
    "10111111111111111111111111111111110100101010000101100010111011100010" when "1001000110",
    "00000000000000000000000000000000000100000011001011000110011110100110" when "1001000111",
    "11011111111111111111111111111111111111111111111111111111111111111111" when "1001001000",
    "01100101010100011110010011110111101001111111111111111111111111111111" when "1001001001",
    "11011111111111111111111111111111110110000011010111010111110000101001" when "1001001010",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1001001011",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1001001100",
    "00000000000000000000000000000000000110001000100011000001000000100000" when "1001001101",
    "01101101001001011001001011111100010010000000000000000000000000000000" when "1001001110",
    "01101011100111001001011100100000010111010110110011000100011101111101" when "1001001111",
    "10011111111111111111111111111111110101100111000011010001011100101000" when "1001010000",
    "10011111111111111111111111111111111101111111111111111111111111111111" when "1001010001",
    "01110010000101010010000010101110100111000110001111100110111010111101" when "1001010010",
    "11011111111111111111111111111111110100011111000111011110100001111111" when "1001010011",
    "01000110100010110000101100001001001101111111111111111111111111111111" when "1001010100",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1001010101",
    "01010111110010110100110100001001010100110000101011101001100100000111" when "1001010110",
    "00100000000000000000000000000000000111000001011001101011001000011010" when "1001010111",
    "00000000000000000000000000000000000110111001010111001011001100011000" when "1001011000",
    "00100000000000000000000000000000000100111011000101111001001101110110" when "1001011001",
    "01110100010110000011101100111010010000000000000000000000000000000000" when "1001011010",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "1001011011",
    "01000010001111011000001010101101100100110011000000101000011000001100" when "1001011100",
    "01000111111110110011010101110001010000000000000000000000000000000000" when "1001011101",
    "10011111111111111111111111111111110101011001111000101110001110010011" when "1001011110",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1001011111",
    "11011111111111111111111111111111110110111111001111110101001001010111" when "1001100000",
    "01011110100001101001000100110010000000000000000000000000000000000000" when "1001100001",
    "00100000000000000000000000000000000101111111100100000011001011101110" when "1001100010",
    "01010110010110111011111010101001110100010000101111111100000111100010" when "1001100011",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "1001100100",
    "10011111111111111111111111111111110110001111101101010101001110000011" when "1001100101",
    "01011010011010110010011001001101111111111111111111111111111111111111" when "1001100110",
    "01001110100111011001101001111101110101111010111101010111010001011100" when "1001100111",
    "01111011001100110000111101011011100010000000000000000000000000000000" when "1001101000",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1001101001",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1001101010",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1001101011",
    "10011111111111111111111111111111110101111001011101010010101011111110" when "1001101100",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1001101101",
    "00000000000000000000000000000000000101011100011010111001000110010110" when "1001101110",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1001101111",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1001110000",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1001110001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1001110010",
    "01001101000111000111000111001011010000000000000000000000000000000000" when "1001110011",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "1001110100",
    "01010110000001111011111001110011110100101011111100010000110000001011" when "1001110101",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1001110110",
    "01000011111001111101111010011011110000000000000000000000000000000000" when "1001110111",
    "00100000000000000000000000000000000101000010110111100111001100010001" when "1001111000",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1001111001",
    "00000000000000000000000000000000001001111111111111111111111111111111" when "1001111010",
    "11111111111111111111111111111111110110100100100110111100101110100000" when "1001111011",
    "01101101110100110111000111001100010010000000000000000000000000000000" when "1001111100",
    "00100000000000000000000000000000000101001010001100100110110010010010" when "1001111101",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "1001111110",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "1001111111",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "1010000000",
    "01100101001101001100000000010001110101110111000000110110110011101010" when "1010000001",
    "00100000000000000000000000000000000111110110101010001010100101110001" when "1010000010",
    "01100011000100110011110100000100010000000000000000000000000000000000" when "1010000011",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1010000100",
    "01101001110000000011100011010000110110100110000010001111100000011111" when "1010000101",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "1010000110",
    "01000101011011110101110010101001001001111111111111111111111111111111" when "1010000111",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1010001000",
    "01011100110000000011000000000011111011111111111111111111111111111111" when "1010001001",
    "01100001110000011110111100111110111111111111111111111111111111111111" when "1010001010",
    "10111111111111111111111111111111110110001000100101100101011000100010" when "1010001011",
    "00100000000000000000000000000000000100000000100100000000011000010000" when "1010001100",
    "01100000100101011000000111010101000111001101010011100011000111011000" when "1010001101",
    "01100000001011100000011011110110011011111111111111111111111111111111" when "1010001110",
    "01110010000100110111011110101001010000000000000000000000000000000000" when "1010001111",
    "11011111111111111111111111111111110111111010000011110000110010111010" when "1010010000",
    "01011111100011111110100011010000110100011011010110100011111101011111" when "1010010001",
    "01001111001110010111110101010011011101111111111111111111111111111111" when "1010010010",
    "11011111111111111111111111111111110110100110000011110000011000000000" when "1010010011",
    "01001001001000010000110010111111000111110111011111010000101101100011" when "1010010100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010010101",
    "01001000011111011110111100001011110110000001100100000101100000000100" when "1010010110",
    "11111111111111111111111111111111110110011010100101011000111100100010" when "1010010111",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1010011000",
    "01011101101011100000110100001011111011111111111111111111111111111111" when "1010011001",
    "10111111111111111111111111111111110100100000111110100110011011001101" when "1010011010",
    "01110000101110111011001110101000111011111111111111111111111111111111" when "1010011011",
    "01100011100100010001001001111100000111000110110101111111111011101010" when "1010011100",
    "10011111111111111111111111111111110010000000000000000000000000000000" when "1010011101",
    "11011111111111111111111111111111110100010000101000110101101000100100" when "1010011110",
    "01111111101011111111011111010110101111111111111111111111111111111111" when "1010011111",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "1010100000",
    "01100111001110011100101100100010100010000000000000000000000000000000" when "1010100001",
    "01000110100001010010101110111011100111111110000101100100000011010000" when "1010100010",
    "01100000010000101001010011011100100100001111101000010101111000000001" when "1010100011",
    "01101100110101010100010111001001110111010001110110000111000000011111" when "1010100100",
    "01101010001000010010101010011100010000000000000000000000000000000000" when "1010100101",
    "01010001110110100001000100101001010100100000111101110111110110110110" when "1010100110",
    "01010001111011011010101000001001010000000000000000000000000000000000" when "1010100111",
    "00000000000000000000000000000000000100000100101001011010101110001001" when "1010101000",
    "01111001110111010010110111001101010010000000000000000000000000000000" when "1010101001",
    "00000000000000000000000000000000000110010111101111001001010100111111" when "1010101010",
    "00000000000000000000000000000000000100111001110010011011001000100100" when "1010101011",
    "01110100010110011110110001110010100100110001011011010011011111010000" when "1010101100",
    "00100000000000000000000000000000000111001011110110001000101101111001" when "1010101101",
    "00100000000000000000000000000000000111100101000111110000011101011110" when "1010101110",
    "00100000000000000000000000000000000101100001100100101111000111111100" when "1010101111",
    "00000000000000000000000000000000000100101000111000000000110101111100" when "1010110000",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1010110001",
    "01010010000100000110101011000000000100011011100110111001101010101000" when "1010110010",
    "01010001101100000100110101110111100100010010011011110100010100011011" when "1010110011",
    "00100000000000000000000000000000000110100110000100011011000001110100" when "1010110100",
    "01101011010010010001111000111100100000000000000000000000000000000000" when "1010110101",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "1010110110",
    "10011111111111111111111111111111110111110100011111111011011100110000" when "1010110111",
    "00100000000000000000000000000000000101100111101100001010101001110111" when "1010111000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1010111001",
    "01111001010110110101101010101010110010000000000000000000000000000000" when "1010111010",
    "01010000101110101000001100100000100110100001111110111101010111111011" when "1010111011",
    "01111111010001000010011101110111010010000000000000000000000000000000" when "1010111100",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "1010111101",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "1010111110",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1010111111",
    "01000101111001001111010010111000010000000000000000000000000000000000" when "1011000000",
    "01101111010110010001010001101100011111111111111111111111111111111111" when "1011000001",
    "01111001000000111001011110000110000111010100110101100101111111000011" when "1011000010",
    "11111111111111111111111111111111110100010001111110110100111110101010" when "1011000011",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "1011000100",
    "01000110110101100101101000001101110101010010001000000001000110010000" when "1011000101",
    "01101001110100101011101000101111000111110011101010000010101001101110" when "1011000110",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "1011000111",
    "01001110110011000110010010001101000100010011000000100110010110010110" when "1011001000",
    "00100000000000000000000000000000001001111111111111111111111111111111" when "1011001001",
    "01000110010111011000011100010111100111100101000101111110000111010100" when "1011001010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011001011",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1011001100",
    "01001111100011111010101000010011010110101101010010011100100110000100" when "1011001101",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011001110",
    "00100000000000000000000000000000000110010111011011010001000000110001" when "1011001111",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "1011010000",
    "00000000000000000000000000000000000111011101001111100001010111101010" when "1011010001",
    "01111010110110001101100101010101011101111111111111111111111111111111" when "1011010010",
    "11111111111111111111111111111111110110110100011111101110101100000110" when "1011010011",
    "00100000000000000000000000000000000101001101001110011001010010101110" when "1011010100",
    "01100001010100100000000110110110010100010110010100010110101100000111" when "1011010101",
    "01111000101101001111100101010001010111101111101000000010111010110010" when "1011010110",
    "01011110011101111001001011111010110101010000010110010111000001101000" when "1011010111",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1011011000",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1011011001",
    "10011111111111111111111111111111110101010011001110000011001001110001" when "1011011010",
    "00000000000000000000000000000000000110000010110000011011010100110011" when "1011011011",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1011011100",
    "01100000111100011001010001011001101101111111111111111111111111111111" when "1011011101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011011110",
    "01010100000000111111010100011111010000000000000000000000000000000000" when "1011011111",
    "00000000000000000000000000000000000111100001001000100100001110101011" when "1011100000",
    "01011111111010010011110101110010000000000000000000000000000000000000" when "1011100001",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1011100010",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011100011",
    "01110111100111001000110000100101010010000000000000000000000000000000" when "1011100100",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011100101",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1011100110",
    "01011000101010001000100000000111001001111111111111111111111111111111" when "1011100111",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1011101000",
    "10011111111111111111111111111111110111010011010110110010111100110000" when "1011101001",
    "00000000000000000000000000000000000110011100101000010011100110101100" when "1011101010",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1011101011",
    "00000000000000000000000000000000000111111111111110100001010100100011" when "1011101100",
    "00000000000000000000000000000000000101011111101011101101101001111101" when "1011101101",
    "00000000000000000000000000000000000100010110011101111000010101010100" when "1011101110",
    "01011101110100111001101110101011100010000000000000000000000000000000" when "1011101111",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1011110000",
    "01110111000010101011001110010000000110111100100100001001010011011001" when "1011110001",
    "11111111111111111111111111111111110100101001110001100001101001100110" when "1011110010",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "1011110011",
    "01011111100101010011000010100011000000000000000000000000000000000000" when "1011110100",
    "10111111111111111111111111111111110101110111010000111011010101001111" when "1011110101",
    "01011000101000011010010101101001001101111111111111111111111111111111" when "1011110110",
    "01111000110011110001011011101101010000000000000000000000000000000000" when "1011110111",
    "01101010100100100100110001011001000111011000001111100010011110100011" when "1011111000",
    "00100000000000000000000000000000000111100000000100010110011111111101" when "1011111001",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "1011111010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011111011",
    "01000111101110100001110010101101010010000000000000000000000000000000" when "1011111100",
    "00100000000000000000000000000000000110110100000101011101111001000000" when "1011111101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1011111110",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1011111111",
    "01000000101111111110101000111011010000000000000000000000000000000000" when "1100000000",
    "00100000000000000000000000000000000100101110011011010011100010011011" when "1100000001",
    "01011011010000011101111010100101110100110110001110011111101010100110" when "1100000010",
    "01111110100100101111101011110011100000000000000000000000000000000000" when "1100000011",
    "01101100111100001101101000011001011111111111111111111111111111111111" when "1100000100",
    "10011111111111111111111111111111110101001000001111001011100010001101" when "1100000101",
    "01100111010001011111010000000101110110101101101101000000111110111000" when "1100000110",
    "01010000101101101001011011111111000000000000000000000000000000000000" when "1100000111",
    "01101100001000101110110111111100000010000000000000000000000000000000" when "1100001000",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1100001001",
    "01111011100101011010011000001011000110110001010111001110110100011010" when "1100001010",
    "00100000000000000000000000000000000111111101111100010101101011000101" when "1100001011",
    "01111110111101010100110000001111000100111011010010101010111010001111" when "1100001100",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1100001101",
    "01111110111101001000010100111101000101110111100011000110011111011001" when "1100001110",
    "11011111111111111111111111111111110101010010100000011001001110101100" when "1100001111",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "1100010000",
    "01111000110010000100110100110000110100101010010111000001011001010000" when "1100010001",
    "10011111111111111111111111111111110000000000000000000000000000000000" when "1100010010",
    "01100101011101101110100110101110010100000000111100100100110000001001" when "1100010011",
    "01000000101001110010111111001100000000000000000000000000000000000000" when "1100010100",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1100010101",
    "00000000000000000000000000000000000110010001001010110011100111011111" when "1100010110",
    "01001000110010100110010111010110100100011111000101001100011001101101" when "1100010111",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "1100011000",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1100011001",
    "11011111111111111111111111111111111111111111111111111111111111111111" when "1100011010",
    "01010110011011100101110100101101010111111000111111100101000000110011" when "1100011011",
    "10111111111111111111111111111111110111111011010011100011011111000110" when "1100011100",
    "00000000000000000000000000000000001011111111111111111111111111111111" when "1100011101",
    "01110100111100000010100011001110010010000000000000000000000000000000" when "1100011110",
    "01110001011110111101100101001100111111111111111111111111111111111111" when "1100011111",
    "10011111111111111111111111111111110101000011101000101010110110011011" when "1100100000",
    "01100110110000000110101111011110000101011011010100001001000001011011" when "1100100001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1100100010",
    "01111100001000011010010111001111110000000000000000000000000000000000" when "1100100011",
    "01101100101100100000101001001011100010000000000000000000000000000000" when "1100100100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100100101",
    "01100000010000010000101100111110010010000000000000000000000000000000" when "1100100110",
    "01100010111101000100101101010010001011111111111111111111111111111111" when "1100100111",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "1100101000",
    "11011111111111111111111111111111110100001101110011011100001111100110" when "1100101001",
    "00100000000000000000000000000000000101101110100101111000100101110011" when "1100101010",
    "11111111111111111111111111111111110110101010001110111101000111010110" when "1100101011",
    "01001110010110001001110101100010000010000000000000000000000000000000" when "1100101100",
    "01110101110000000010010110000011110000000000000000000000000000000000" when "1100101101",
    "01101011100100110010000001011011100101101110001010100001111111101001" when "1100101110",
    "01111110110100011001111000010010100100110101000000001101010000011011" when "1100101111",
    "01101100111110100110110100011010010101111100110101110001100000000101" when "1100110000",
    "11011111111111111111111111111111111001111111111111111111111111111111" when "1100110001",
    "00100000000000000000000000000000000110010101110000110001000000110100" when "1100110010",
    "00100000000000000000000000000000000111111011000011010011100000000000" when "1100110011",
    "01101000111000101100101100000001001101111111111111111111111111111111" when "1100110100",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "1100110101",
    "01111001010010000100111010001101000101000101110101110010110011111011" when "1100110110",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "1100110111",
    "01111111010111110100001001001100110010000000000000000000000000000000" when "1100111000",
    "01110101110101101000000000000011110000000000000000000000000000000000" when "1100111001",
    "01001110101011110010101110010001110110101111011011101001100110001000" when "1100111010",
    "01110010111101010101001000111010110100011000111101011010001011100111" when "1100111011",
    "00000000000000000000000000000000000111111000101000011100100110011101" when "1100111100",
    "01111000001100101000000111000001111001111111111111111111111111111111" when "1100111101",
    "10011111111111111111111111111111110101110111110000010001001111011011" when "1100111110",
    "10111111111111111111111111111111110100000000111110000110010011111000" when "1100111111",
    "11111111111111111111111111111111111101111111111111111111111111111111" when "1101000000",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "1101000001",
    "11011111111111111111111111111111111011111111111111111111111111111111" when "1101000010",
    "01100001011110110101110000111101011101111111111111111111111111111111" when "1101000011",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1101000100",
    "10111111111111111111111111111111110111110101101001111011101010111001" when "1101000101",
    "01001110000011110111010101101101110010000000000000000000000000000000" when "1101000110",
    "00100000000000000000000000000000000101110000001000001101001001000001" when "1101000111",
    "01000100001001111010001101001100010101000110111101101010110111001011" when "1101001000",
    "01110000111010011010100011001011110000000000000000000000000000000000" when "1101001001",
    "01111011011010101111011100011001010010000000000000000000000000000000" when "1101001010",
    "10011111111111111111111111111111111111111111111111111111111111111111" when "1101001011",
    "01011100100110111011011111110100010111100101110101111101011011000000" when "1101001100",
    "00000000000000000000000000000000000101101000110011100010101110101001" when "1101001101",
    "01000001000110110100011100001000110010000000000000000000000000000000" when "1101001110",
    "01010000010011101111100111111010110111000001100100110110111010010000" when "1101001111",
    "01111011100010101000001110101101010111110011111000000011101111000101" when "1101010000",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "1101010001",
    "01001000111100001101111100110110110111000100001001001001111110010100" when "1101010010",
    "11011111111111111111111111111111110110001111100110010001110010010010" when "1101010011",
    "01100000010110000010111110100100100100001110110011011011111111110000" when "1101010100",
    "11111111111111111111111111111111111001111111111111111111111111111111" when "1101010101",
    "01111000000111111111011000010100110000000000000000000000000000000000" when "1101010110",
    "11011111111111111111111111111111110010000000000000000000000000000000" when "1101010111",
    "10111111111111111111111111111111110111001000000111111011100010000110" when "1101011000",
    "01001001100110001100110110111101010000000000000000000000000000000000" when "1101011001",
    "01110101101111010010001000011000000101100011000100110010001011100100" when "1101011010",
    "01111100000110010101010110110000000010000000000000000000000000000000" when "1101011011",
    "01111111001001000001101001011001011101111111111111111111111111111111" when "1101011100",
    "01111100111010011001001100001000000110110011010011100101110101001010" when "1101011101",
    "10111111111111111111111111111111110111001011111000100100011011101100" when "1101011110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1101011111",
    "01101100111000010101011010101001110010000000000000000000000000000000" when "1101100000",
    "01010010001110100100001111110001000111010001100010000101100111111111" when "1101100001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1101100010",
    "10111111111111111111111111111111111101111111111111111111111111111111" when "1101100011",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1101100100",
    "11111111111111111111111111111111110111100000100111010100110000011000" when "1101100101",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1101100110",
    "01011011011001010111001111011100010111111010110110101100100010110000" when "1101100111",
    "11011111111111111111111111111111110100101011000100001101111111111111" when "1101101000",
    "01101110111010010110010110000101110100100010100100101010010110010110" when "1101101001",
    "11011111111111111111111111111111110110101011110100001110101100011110" when "1101101010",
    "00100000000000000000000000000000000100000101101000010100011001101111" when "1101101011",
    "11111111111111111111111111111111110101001100010000101011111000011111" when "1101101100",
    "01111110100101111000010101111110001111111111111111111111111111111111" when "1101101101",
    "01100110000001111011001101000111110100111001100000111111001001000110" when "1101101110",
    "01010001111101011110101011111101110111110100111101010011000010000101" when "1101101111",
    "01111001000111100010110011010111110010000000000000000000000000000000" when "1101110000",
    "01111001010101010001001110110010000100001000010110101110110000001010" when "1101110001",
    "01100000000110100110001011111110011001111111111111111111111111111111" when "1101110010",
    "01101110001010100011001011101010111011111111111111111111111111111111" when "1101110011",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1101110100",
    "01010010000100010100111011110100111101111111111111111111111111111111" when "1101110101",
    "10011111111111111111111111111111110110100000000100100001010101110000" when "1101110110",
    "01000100010110010001010000100111001101111111111111111111111111111111" when "1101110111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101111000",
    "01011100111010111101010100111101010111100110000011011000010100100111" when "1101111001",
    "11011111111111111111111111111111110111100001011001010100101111000011" when "1101111010",
    "01011101110000110101010001000000000111101101111101111011111001111000" when "1101111011",
    "01111110101011101010001100010001101001111111111111111111111111111111" when "1101111100",
    "10011111111111111111111111111111110101100000010001101010011110011100" when "1101111101",
    "01111001010111100100100001001011000000000000000000000000000000000000" when "1101111110",
    "01101101110001010011011011010010010110111111111101001001101100110010" when "1101111111",
    "10111111111111111111111111111111111001111111111111111111111111111111" when "1110000000",
    "00000000000000000000000000000000000101000101001111010101010110010100" when "1110000001",
    "01010010010100101110000111010000110000000000000000000000000000000000" when "1110000010",
    "10111111111111111111111111111111111001111111111111111111111111111111" when "1110000011",
    "01101111100011001010010111100010000111011000101011101001011011011110" when "1110000100",
    "01100101110011001000100000100000001011111111111111111111111111111111" when "1110000101",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1110000110",
    "01111111000000010000010010101111100110101010001101100111011000100110" when "1110000111",
    "01101101110001101011111110110010101101111111111111111111111111111111" when "1110001000",
    "10011111111111111111111111111111110101011001001110001111111101001010" when "1110001001",
    "01110101001011101011000000001100110010000000000000000000000000000000" when "1110001010",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "1110001011",
    "01101000101100010100111011101000100010000000000000000000000000000000" when "1110001100",
    "01111000001110100101100000001011001111111111111111111111111111111111" when "1110001101",
    "00100000000000000000000000000000001111111111111111111111111111111111" when "1110001110",
    "01100010010010001001011000011111101111111111111111111111111111111111" when "1110001111",
    "11011111111111111111111111111111110101111011010110011010100011011110" when "1110010000",
    "01011011111111000001001000110101010010000000000000000000000000000000" when "1110010001",
    "01010101111011000111010001000000001011111111111111111111111111111111" when "1110010010",
    "01010010100001001100100110111110100010000000000000000000000000000000" when "1110010011",
    "10111111111111111111111111111111110110111001110000111100010000000110" when "1110010100",
    "01110100100110010110100111011010010101110110111011010000011101001111" when "1110010101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1110010110",
    "01110000011101000010111111001101010100010011100001100110110000100110" when "1110010111",
    "01111000010010000010110001101110111101111111111111111111111111111111" when "1110011000",
    "01101101000101010010011010101001000010000000000000000000000000000000" when "1110011001",
    "00000000000000000000000000000000000111001000100001010110010111011001" when "1110011010",
    "01001001111001011111001011010100111011111111111111111111111111111111" when "1110011011",
    "00000000000000000000000000000000000110111100001010111111010110110001" when "1110011100",
    "01100010100011100010000001110010010101111110110100111000101010111100" when "1110011101",
    "01001011011100111000001001000011011011111111111111111111111111111111" when "1110011110",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "1110011111",
    "01101010001001101100111110010000110101111000011110011100010011110111" when "1110100000",
    "11011111111111111111111111111111110111000110000000100010110110010111" when "1110100001",
    "01101001000011010000010110010101011101111111111111111111111111111111" when "1110100010",
    "01010100111010011001100111100011000010000000000000000000000000000000" when "1110100011",
    "01011101010110000101000001111000101101111111111111111111111111111111" when "1110100100",
    "10111111111111111111111111111111110100011000111101001010001100000110" when "1110100101",
    "01100100100010111110001111101011100000000000000000000000000000000000" when "1110100110",
    "01100011011101110110111101110101011011111111111111111111111111111111" when "1110100111",
    "10111111111111111111111111111111110101001111101111110100111000010001" when "1110101000",
    "00100000000000000000000000000000001011111111111111111111111111111111" when "1110101001",
    "01100001101011000011111110011100011111111111111111111111111111111111" when "1110101010",
    "10011111111111111111111111111111110101100110010011001100100011011011" when "1110101011",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "1110101100",
    "01101101100100010000010101000011001001111111111111111111111111111111" when "1110101101",
    "01000110111101110110010110001010110101001011000100011111011110001011" when "1110101110",
    "01001110000000010110100100001110100101010101111010010110011000111100" when "1110101111",
    "10011111111111111111111111111111111011111111111111111111111111111111" when "1110110000",
    "01010000000100010100100101111001011011111111111111111111111111111111" when "1110110001",
    "01100110001000010011100000110100101111111111111111111111111111111111" when "1110110010",
    "01101100110010110011000100100111000110001001011011011111111111110101" when "1110110011",
    "01000010011000011110111001010001000110001100111111111000011111011011" when "1110110100",
    "01000001011011011010111001100001001101111111111111111111111111111111" when "1110110101",
    "11111111111111111111111111111111110000000000000000000000000000000000" when "1110110110",
    "01011111100111100010100010110010100100110011110010001011011101000100" when "1110110111",
    "01011000100010110110110101110000000100011111000101001100011111101000" when "1110111000",
    "01001111010001111000011000010000011111111111111111111111111111111111" when "1110111001",
    "00000000000000000000000000000000001111111111111111111111111111111111" when "1110111010",
    "01000001011011101110000110100101010110000100000111001100010011010111" when "1110111011",
    "10111111111111111111111111111111110100100001011100101010100011110001" when "1110111100",
    "01101100011000001011111010110101111001111111111111111111111111111111" when "1110111101",
    "01110110101110101001000010111001100000000000000000000000000000000000" when "1110111110",
    "01010111010001001001111001111100010010000000000000000000000000000000" when "1110111111",
    "01001100010100001101001011010111111001111111111111111111111111111111" when "1111000000",
    "11011111111111111111111111111111110101110000100110000111010001111101" when "1111000001",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1111000010",
    "10111111111111111111111111111111111001111111111111111111111111111111" when "1111000011",
    "10111111111111111111111111111111111101111111111111111111111111111111" when "1111000100",
    "01100100001001010000010001011011111101111111111111111111111111111111" when "1111000101",
    "00000000000000000000000000000000000010000000000000000000000000000000" when "1111000110",
    "11111111111111111111111111111111110010000000000000000000000000000000" when "1111000111",
    "10111111111111111111111111111111110010000000000000000000000000000000" when "1111001000",
    "11111111111111111111111111111111110101010001111111100110000101100101" when "1111001001",
    "01100101000111010011011010000000010110010101110101110111001111001111" when "1111001010",
    "10011111111111111111111111111111110111101111001001110100100001110001" when "1111001011",
    "01111011101100101001100011111001011001111111111111111111111111111111" when "1111001100",
    "01000010101000110110000100110000110101010101110010101000100110010100" when "1111001101",
    "00100000000000000000000000000000001001111111111111111111111111111111" when "1111001110",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1111001111",
    "00100000000000000000000000000000001101111111111111111111111111111111" when "1111010000",
    "01000110110010010110011000101011110101110110001000110110100101011010" when "1111010001",
    "01101101101111001010000010111001000010000000000000000000000000000000" when "1111010010",
    "10111111111111111111111111111111110101101110110011111101011111000110" when "1111010011",
    "11011111111111111111111111111111110000000000000000000000000000000000" when "1111010100",
    "01010011001011011111010001100100100101011011010011101101100100000011" when "1111010101",
    "01110000100101101100010001010111011001111111111111111111111111111111" when "1111010110",
    "01001101101110101101100010000011111101111111111111111111111111111111" when "1111010111",
    "01000110010110000101111110100111100101001011000010101010110101011000" when "1111011000",
    "01100111111001100110001101111001010111110010111111011100110101011111" when "1111011001",
    "01110101111101001000011000111001101101111111111111111111111111111111" when "1111011010",
    "01001000010101111100110110100111100110101010110111010110111001110010" when "1111011011",
    "01111110100000111000110110110111110101111101000011101111100001010000" when "1111011100",
    "10111111111111111111111111111111110110110010101010100101111100100010" when "1111011101",
    "01111100010001100000001110111110100101100111110000001011110000100000" when "1111011110",
    "01010100111111000000011110101010010110000110101001100111101111000010" when "1111011111",
    "01110011110010110000000000010010010000000000000000000000000000000000" when "1111100000",
    "01010111001000100001100000101111110100111001001011111000010110010010" when "1111100001",
    "00100000000000000000000000000000000000000000000000000000000000000000" when "1111100010",
    "01011001000110111101110010011010100000000000000000000000000000000000" when "1111100011",
    "01101001001101001111010010110011010111000101001100010111011010101011" when "1111100100",
    "01110010001100100110001010101000100111010010001111011011100001110001" when "1111100101",
    "01111110110111110100101011011110111101111111111111111111111111111111" when "1111100110",
    "01001101001001000111000010101000110111001011110101011000110110011011" when "1111100111",
    "01110111000101111001111100010101110101010010110110010100111101011010" when "1111101000",
    "00000000000000000000000000000000000100111110001011001000010010011000" when "1111101001",
    "01101110110100110100001011100101101101111111111111111111111111111111" when "1111101010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111101011",
    "01111100111101111000010110010011001001111111111111111111111111111111" when "1111101100",
    "11011111111111111111111111111111110100111110001010010111100101001011" when "1111101101",
    "01101110001111110011100110011101110110000110000111111110001111100011" when "1111101110",
    "01011110000110001101111011000011111011111111111111111111111111111111" when "1111101111",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1111110000",
    "10111111111111111111111111111111110000000000000000000000000000000000" when "1111110001",
    "00100000000000000000000000000000000111000110000000001100000011111111" when "1111110010",
    "01110001011011000110000011010010011001111111111111111111111111111111" when "1111110011",
    "01011111001001110011010001010010010100100000111110000110000111000101" when "1111110100",
    "10111111111111111111111111111111111001111111111111111111111111111111" when "1111110101",
    "00000000000000000000000000000000001101111111111111111111111111111111" when "1111110110",
    "01101011101101011010000110101110001111111111111111111111111111111111" when "1111110111",
    "01001000011101101000000000001111010100100011110011100101100011011011" when "1111111000",
    "01100110111101001111101000101000100101001111110010000001010000100101" when "1111111001",
    "00000000000000000000000000000000000100011110101011011111111111110110" when "1111111010",
    "01110111110010111010111110111100101101111111111111111111111111111111" when "1111111011",
    "11111111111111111111111111111111110100000111111100110010111110111101" when "1111111100",
    "01001001011101011010100001000011001101111111111111111111111111111111" when "1111111101",
    "01010110101101110011001001101011000010000000000000000000000000000000" when "1111111110",
    "01110011000000011001111000101001110110010111010111111100100011010111" when "1111111111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when others;

with addr(9 downto 0) select
  outVal(67 downto 0) <=
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000000000",
    "01101111010011000010110101111011000110111101001100001011010111101100" when "0000000001",
    "01011010110001100010010110010111100101101011000110001001011001011110" when "0000000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000000011",
    "01010111010100110100001001011001000101011101010011010000100101100100" when "0000000100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000000101",
    "01100001011100101010000101010011110110000101110010101000010101001111" when "0000000110",
    "01001011011110011100110011110101010100101101111001110011001111010101" when "0000000111",
    "01101110010100110111001000111000100110111001010011011100100011100010" when "0000001000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000001001",
    "01011110000111000100001011101101000101111000011100010000101110110100" when "0000001010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000001011",
    "01001110110110010000010100011001110100111011011001000001010001100111" when "0000001100",
    "01100111000000111000010000110000000110011100000011100001000011000001" when "0000001101",
    "01000110111100101111010110001110110100011011110010111101011000111011" when "0000001110",
    "01001001110000111110010101011111000100100111000011111001010101111100" when "0000001111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0000010000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000010001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000010010",
    "01111100101111000100001110100100010111110010111100010000111010010001" when "0000010011",
    "01101010000001100110001001111011110110101000000110011000100111101111" when "0000010100",
    "01011000110001001110000110011000000101100011000100111000011001100000" when "0000010101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000010110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000010111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000011000",
    "01101011100010110100011110010010100110101110001011010001111001001010" when "0000011001",
    "01000101011111101101101010000011110100010101111110110110101000001111" when "0000011010",
    "01001011000001100000101101100100000100101100000110000010110110010000" when "0000011011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000011100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000011101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000011110",
    "01111010110100101101111100001001100111101011010010110111110000100110" when "0000011111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000100000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000100001",
    "01000100000001001011000000100001000100010000000100101100000010000101" when "0000100010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000100011",
    "01011000111110011101000101010011110101100011111001110100010101001111" when "0000100100",
    "01001001001111110001111101000011110100100100111111000111110100001111" when "0000100101",
    "01100000011000101100110000000011010110000001100010110011000000001110" when "0000100110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000100111",
    "01111001111000111001000101011111010111100111100011100100010101111101" when "0000101000",
    "01100100100111011111100000000000000110010010011101111110000000000000" when "0000101001",
    "01100001010101010111010001100010000110000101010101011101000110001000" when "0000101010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000101011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000101100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000101101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000101110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000110001",
    "01011111000101111000011011110101100101111100010111100001101111010110" when "0000110010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0000110011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000110100",
    "01101010100100000000000000111001110110101010010000000000000011100111" when "0000110101",
    "01011111111101001000010001101001000101111111110100100001000110100100" when "0000110110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0000110111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000111000",
    "01100010100101110111001111011100000110001010010111011100111101110000" when "0000111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0000111010",
    "01101001000111111100011011000111110110100100011111110001101100011111" when "0000111011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000111100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0000111101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0000111110",
    "01011011100011110110100100001111010101101110001111011010010000111101" when "0000111111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0001000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001000001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001000010",
    "01001110101110100100010110011101110100111010111010010001011001110111" when "0001000011",
    "01001111101111000101010101110111000100111110111100010101010111011100" when "0001000100",
    "01010010101001001100101101101111010101001010100100110010110110111101" when "0001000101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001000110",
    "01110011101111101010000101101111010111001110111110101000010110111101" when "0001000111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001001000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001001001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001001010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001001011",
    "01100110101010111011100110001110000110011010101011101110011000111000" when "0001001100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001001101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001001110",
    "01000011111000111011011000010111110100001111100011101101100001011111" when "0001001111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001010000",
    "01001100010101000100000010110001000100110001010100010000001011000100" when "0001010001",
    "01101010110011010000011011101110100110101011001101000001101110111010" when "0001010010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001010011",
    "01011010111001100100111010100010000101101011100110010011101010001010" when "0001010100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001010101",
    "01100011100110000011111011001101000110001110011000001111101100110100" when "0001010110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001010111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0001011000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001011001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001011011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001011100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001011101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001011110",
    "01011010000111001010111000010000110101101000011100101011100001000011" when "0001011111",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0001100000",
    "01100001001001000001101011001101110110000100100100000110101100110111" when "0001100001",
    "01011010111101011101001100000010110101101011110101110100110000001011" when "0001100010",
    "01000001000110001100010101011100100100000100011000110001010101110010" when "0001100011",
    "01100010011001110100001100000001000110001001100111010000110000000100" when "0001100100",
    "01010000011001011000111011101011010101000001100101100011101110101101" when "0001100101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001100110",
    "01100011000111110011101111001001010110001100011111001110111100100101" when "0001100111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001101000",
    "01001110100111011001010010011000110100111010011101100101001001100011" when "0001101001",
    "01110101000111110000011010101111010111010100011111000001101010111101" when "0001101010",
    "01110001101000110100000110001000010111000110100011010000011000100011" when "0001101011",
    "01101001010111001010110011010100100110100101011100101011001101010010" when "0001101100",
    "01101010001111110111011100111001000110101000111111011101110011100100" when "0001101101",
    "01000100100110010100001000111110010100010010011001010000100011111001" when "0001101110",
    "01101110110010000101000000001101100110111011001000010100000000110110" when "0001101111",
    "01001100000101010101101111110001000100110000010101010110111111000100" when "0001110000",
    "01101110001101101101101100111000110110111000110110110110110011100011" when "0001110001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001110010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001110011",
    "01011010101100011111111001001111110101101010110001111111100100111111" when "0001110100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0001110101",
    "01000110111111110110111011110101100100011011111111011011101111010110" when "0001110110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001110111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0001111000",
    "01101100001001101001100101001010000110110000100110100110010100101000" when "0001111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001111010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0001111011",
    "01001111100111100010000100100110100100111110011110001000010010011010" when "0001111100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0001111101",
    "01111100111010010011101101011010010111110011101001001110110101101001" when "0001111110",
    "01001001000100111001011011100111110100100100010011100101101110011111" when "0001111111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010000000",
    "01111100000001100101101000001001100111110000000110010110100000100110" when "0010000001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010000010",
    "01011001011110001111111101101000010101100101111000111111110110100001" when "0010000011",
    "01111100101010100100010100011001100111110010101010010001010001100110" when "0010000100",
    "01001100001110111111100100110111100100110000111011111110010011011110" when "0010000101",
    "01001011101011101101011111111101000100101110101110110101111111110100" when "0010000110",
    "01101000000111010001001101111010110110100000011101000100110111101011" when "0010000111",
    "01101000110010100000110101001011010110100011001010000011010100101101" when "0010001000",
    "01111110011010010001101000111001100111111001101001000110100011100110" when "0010001001",
    "01100010100101010101000010001011000110001010010101010100001000101100" when "0010001010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0010001011",
    "01000111001100110110010110010101100100011100110011011001011001010110" when "0010001100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0010001101",
    "01111101011001110010111001010110100111110101100111001011100101011010" when "0010001110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010001111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010010000",
    "01100011011010110101010110000111100110001101101011010101011000011110" when "0010010001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010010010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010010011",
    "01101101000100000000011100100100010110110100010000000001110010010001" when "0010010100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0010010101",
    "01000110101100110000000000111010100100011010110011000000000011101010" when "0010010110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010010111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0010011000",
    "01001101010101111111101110000100110100110101010111111110111000010011" when "0010011001",
    "01011010000010001010010101011100000101101000001000101001010101110000" when "0010011010",
    "01101001110100010110110010100001000110100111010001011011001010000100" when "0010011011",
    "01111001100010100111000111110011010111100110001010011100011111001101" when "0010011100",
    "01001100111111111001110011011101110100110011111111100111001101110111" when "0010011101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010011111",
    "01010111111011110101011000000000010101011111101111010101100000000001" when "0010100000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010100001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010100010",
    "01011011011001011000000100111000100101101101100101100000010011100010" when "0010100011",
    "01011111001101111111010001000101100101111100110111111101000100010110" when "0010100100",
    "01100011111000000101001001101011010110001111100000010100100110101101" when "0010100101",
    "01100100001111110111011011110100110110010000111111011101101111010011" when "0010100110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0010100111",
    "01011111110100100000000110010000100101111111010010000000011001000010" when "0010101000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0010101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010101010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010101011",
    "01010101000111001101011001001001000101010100011100110101100100100100" when "0010101100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010101101",
    "01110110010010000001110010011011000111011001001000000111001001101100" when "0010101110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010110001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0010110010",
    "01000000100001010110011101110010110100000010000101011001110111001011" when "0010110011",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0010110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010110110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0010110111",
    "01111010100111101010011001100100100111101010011110101001100110010010" when "0010111000",
    "01111010101000100100000110010101110111101010100010010000011001010111" when "0010111001",
    "01011101010101110100100111110001000101110101010111010010011111000100" when "0010111010",
    "01110011001100010100110011000011110111001100110001010011001100001111" when "0010111011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0010111100",
    "01110110001111100100011001100000000111011000111110010001100110000000" when "0010111101",
    "01111000000001000011111101101111110111100000000100001111110110111111" when "0010111110",
    "01101011011111000100101110100000000110101101111100010010111010000000" when "0010111111",
    "01001001010101111100011100100111000100100101010111110001110010011100" when "0011000000",
    "01101101111001010101011010110110010110110111100101010101101011011001" when "0011000001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011000010",
    "01000011001110001100111111100110000100001100111000110011111110011000" when "0011000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011000100",
    "01100111010010110111001110000110000110011101001011011100111000011000" when "0011000101",
    "01001100110101100010110100111100100100110011010110001011010011110010" when "0011000110",
    "01100110010100000100010101110000000110011001010000010001010111000000" when "0011000111",
    "01011101110011001111111100110111100101110111001100111111110011011110" when "0011001000",
    "01001011000111010001010010111010110100101100011101000101001011101011" when "0011001001",
    "01100011010011110101100100101001010110001101001111010110010010100101" when "0011001010",
    "01100110101000011101010100101011110110011010100001110101010010101111" when "0011001011",
    "01111000111000011100010010110101000111100011100001110001001011010100" when "0011001100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011001101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011001110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011001111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011010000",
    "01001110010101110111100000101001010100111001010111011110000010100101" when "0011010001",
    "01010011001101010101111000110101000101001100110101010111100011010100" when "0011010010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011010011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011010100",
    "01110011101001001011110111100101000111001110100100101111011110010101" when "0011010101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011010110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011010111",
    "01011110100111100100100001010011010101111010011110010010000101001101" when "0011011000",
    "01011001111011001010101010000000010101100111101100101010101000000001" when "0011011001",
    "01001110101000111001111001011101100100111010100011100111100101110110" when "0011011010",
    "01001100100111100001110101001011000100110010011110000111010100101100" when "0011011011",
    "01000111011001000110001101011010010100011101100100011000110101101001" when "0011011100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011011101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011011110",
    "01001101000001110111000001000101010100110100000111011100000100010101" when "0011011111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011100000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011100001",
    "01101101110000010101011111110111110110110111000001010101111111100000" when "0011100010",
    "01111111001100001101101111101100000111111100110000110110111110110000" when "0011100011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011100100",
    "01110000111001001101110001110101010111000011100100110111000111010101" when "0011100101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011100110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011100111",
    "01101100101101111011010001010110000110110010110111101101000101011000" when "0011101000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011101001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011101010",
    "01000101001110010111001110011010000100010100111001011100111001101000" when "0011101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011101100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011101101",
    "01000101000001010010111000110001110100010100000101001011100011000111" when "0011101110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011101111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011110001",
    "01111011101011110010110101100001110111101110101111001011011001000001" when "0011110010",
    "01001001011111111111000001100101000100100101111111111100000110010100" when "0011110011",
    "01110000101100010101111100110010000111000010110001010111110011001000" when "0011110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011110101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011110110",
    "01110100000001101100100000100011000111010000000110110010000010001100" when "0011110111",
    "01100110100110101110101101001000000110011010011010111010110100100000" when "0011111000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0011111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011111010",
    "01001100111000100001110111001101110100110011100010000111011100110111" when "0011111011",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0011111100",
    "01100100110101001000111011010101100110010011010100100011101101010110" when "0011111101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0011111110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0011111111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100000000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100000001",
    "01110100000100101010001000000010110111010000010010101000100000001011" when "0100000010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100000011",
    "01000111111111111000111000000100100100011111111111100011100000010010" when "0100000100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100000101",
    "01100101000011100111100010000011100110010100001110011110001000001110" when "0100000110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100000111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100001000",
    "01100110000001010010111011000001010110011000000101001011101100000101" when "0100001001",
    "01001010001010100011100100010011110100101000101010001110010001001111" when "0100001010",
    "01010111011110111110110111001111110101011101111011111011011101000001" when "0100001011",
    "01110101010001011101101000001011010111010101000101110110100000101101" when "0100001100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100001101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100001110",
    "01110010101010111111110000011111010111001010101011111111000001111101" when "0100001111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100010000",
    "01000010100101010000011100001001010100001010010101000001110000100101" when "0100010001",
    "01100101000000001011011111100111100110010100000000101101111110100100" when "0100010010",
    "01101101001101011010110000101111110110110100110101101011000010111111" when "0100010011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100010100",
    "01001010011110111010000000010001010100101001111011101000000001000101" when "0100010101",
    "01011010010111000100101000100000110101101001011100010010100010000011" when "0100010110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100010111",
    "01101110100101010011100110010111110110111010010101001110011001011111" when "0100011000",
    "01100001010101001100101011000111110110000101010100110010101100011111" when "0100011001",
    "01001011010100001011100101001100110100101101010000101110010100110011" when "0100011010",
    "01010011101010110110110100100011000101001110101011011011010010001101" when "0100011011",
    "01001101011111011111111001011101000100110101111101111111100101110100" when "0100011100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100011101",
    "01110100101001110101111010101011110111010010100111010111101010101111" when "0100011110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100011111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100100000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100100001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100100010",
    "01101000000001000111010010011101000110100000000100011101001001110100" when "0100100011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100100100",
    "01011010101100101101001001111111110101101010110010110100100111111111" when "0100100101",
    "01011110011011011000000100111001010101111001101101100000010011100101" when "0100100110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100100111",
    "01110100001111111010111100000101110111010000111111101011110000010111" when "0100101000",
    "01001111011101100000101011001001100100111101110110000010101100100110" when "0100101001",
    "01101000010010111101100101101110010110100001001011110110010110111001" when "0100101010",
    "01001110110111001110111011011000000100111011011100111011101101100000" when "0100101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100101100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100101101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100101110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100101111",
    "01101001001010010011100111111111100110100100101001001110011111111110" when "0100110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100110001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100110010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0100110011",
    "01101100111110000110101111011110010110110011111000011010111101111001" when "0100110100",
    "01000011000010010010100100111010100100001100001001001010010011101010" when "0100110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0100110110",
    "01010101010101101010010011010001010101010101010110101001001101000101" when "0100110111",
    "01000110011100001010100011101001010100011001110000101010001110100101" when "0100111000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0100111001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0100111010",
    "01011101110101101001010001111111010101110111010110100101000111111101" when "0100111011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0100111100",
    "01000111000011111101001101010110010100011100001111110100110101011001" when "0100111101",
    "01001011010101010010010000011110010100101101010101001001000001111001" when "0100111110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0100111111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101000001",
    "01001010100011111110100000101000110100101010001111111010000010100011" when "0101000010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101000011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101000100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101000101",
    "01001110001101111001011100100000010100111000110111100101110010000001" when "0101000110",
    "01101111000000100100101110101111010110111100000010010010111010111101" when "0101000111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101001000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101001001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0101001010",
    "01101011000101111111110011011000010110101100010111111111001101100001" when "0101001011",
    "01101011000011001100000000101000010110101100001100110000000010100001" when "0101001100",
    "01000111101101101111001100011110110100011110110110111100110001111011" when "0101001101",
    "01001100010110101100100110010001000100110001011010110010011001000100" when "0101001110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101001111",
    "01111000000011111011010011100010100111100000001111101101001110001010" when "0101010000",
    "01101100101110011011110111000000010110110010111001101111011100000001" when "0101010001",
    "01010000111100001010010000101010000101000011110000101001000010101000" when "0101010010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101010011",
    "01001101111001000111001101000111110100110111100100011100110100011111" when "0101010100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101010101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101010110",
    "01000011010110010001100100000110010100001101011001000110010000011001" when "0101010111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101011000",
    "01100000011000100011101111100111110110000001100010001110111110011111" when "0101011001",
    "01001010001100101100010111110000100100101000110010110001011111000010" when "0101011010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0101011011",
    "01000011000110101100011000010001110100001100011010110001100001000111" when "0101011100",
    "01101011111111011011010100100010000110101111111101101101010010001000" when "0101011101",
    "01001011110111110101100100001110110100101111011111010110010000111011" when "0101011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101011111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101100000",
    "01011011000110010100000001010010000101101100011001010000000101001000" when "0101100001",
    "01100100110101101100000111000010000110010011010110110000011100001000" when "0101100010",
    "01101011000100000110010101110111010110101100010000011001010111011101" when "0101100011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101100100",
    "01110111001001110100010101010000100111011100100111010001010101000010" when "0101100101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101100110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101100111",
    "01110100000100010100111110100000000111010000010001010011111010000000" when "0101101000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101101010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101101100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101101101",
    "01100001000000011000011110001010000110000100000001100001111000101000" when "0101101110",
    "01100000000011110010000101001011000110000000001111001000010100101100" when "0101101111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101110001",
    "01100111110101111110000000100110100110011111010111111000000010011010" when "0101110010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101110011",
    "01010010010010100101101110000101100101001001001010010110111000010110" when "0101110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101110101",
    "01100101011000001111110011111111110110010101100000111111001111111111" when "0101110110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101110111",
    "01101111100001000000011111100101010110111110000100000001111110010101" when "0101111000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0101111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101111010",
    "01101011011110110001101001011000100110101101111011000110100101100010" when "0101111011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101111100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0101111101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0101111110",
    "01010111000010000101111000001011110101011100001000010111100000101111" when "0101111111",
    "01111000001111100110010001111100100111100000111110011001000111110010" when "0110000000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110000001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110000010",
    "01111111001011011111000010001011110111111100101101111100001000101111" when "0110000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110000100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110000101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110000110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110000111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110001000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110001001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110001010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110001011",
    "01010011000110011110100001110001010101001100011001111010000111000101" when "0110001100",
    "01101000001011111000111101111000100110100000101111100011110111100010" when "0110001101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110001110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110001111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110010000",
    "01111000101101001101010110000111110111100010110100110101011000011111" when "0110010001",
    "01011011011011110111001100001110000101101101101111011100110000111000" when "0110010010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110010011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110010100",
    "01000110111011111000111110001010100100011011101111100011111000101010" when "0110010101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110010110",
    "01101010010011010101111111101001110110101001001101010111111110100111" when "0110010111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110011000",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0110011001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110011011",
    "01101011111011111111101110000010110110101111101111111110111000001011" when "0110011100",
    "01101110101011011010001111010110100110111010101101101000111101011010" when "0110011101",
    "01100000010110110110011000001001000110000001011011011001100000100100" when "0110011110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110011111",
    "01001111010110001001101101010010000100111101011000100110110101001000" when "0110100000",
    "01010101001000100111001110001001110101010100100010011100111000101000" when "0110100001",
    "01010011111000111001011011101001010101001111100011100101101110100101" when "0110100010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110100011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110100100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110100101",
    "01001100001001111101101100000011000100110000100111110110110000001100" when "0110100110",
    "01101101111110000001100101010010110110110111111000000110010101001011" when "0110100111",
    "01001111011101000101010000110011010100111101110100010101000011001101" when "0110101000",
    "01001000100111110110100111101111010100100010011111011010011110111101" when "0110101001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110101010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110101011",
    "01011110010011111010100010110001110101111001001111101010001011000111" when "0110101100",
    "01101010110011001110010011110101010110101011001100111001001111010110" when "0110101101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0110101110",
    "01111110010100011101011010101110000111111001010001110101101010111000" when "0110101111",
    "01101111100001110100011011100111000110111110000111010001101110011100" when "0110110000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110110001",
    "01101011101100111110011101111110010110101110110011111001110111111001" when "0110110010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110110011",
    "01111111001001101100100101110111110111111100100110110010010111011111" when "0110110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110110101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0110110110",
    "01001011011110011100110011000001110100101101111001110011001100000111" when "0110110111",
    "01100110000001011100000100010101010110011000000101110000010001010101" when "0110111000",
    "01011100111000101101010100100011000101110011100010110101010010001100" when "0110111001",
    "01111100101000010001001011011100000111110010100001000100101101110000" when "0110111010",
    "01000100101010011001110101001110010100010010101001100111010100111001" when "0110111011",
    "01010110010001100010110010110100010101011001000110001011001011010001" when "0110111100",
    "01110111101011000000011011110010000111011110101100000001101111001000" when "0110111101",
    "01110100111010101101001100011000000111010011101010110100110001100000" when "0110111110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0110111111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0111000000",
    "01001111111000101111010110111110010100111111100010111101011011111001" when "0111000001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111000010",
    "01100001110011010111101000011001000110000111001101011110100001100100" when "0111000011",
    "01011100010000100110111010010011100101110001000010011011101001001110" when "0111000100",
    "01000010101000000001010100001011100100001010100000000101010000101110" when "0111000101",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "0111000110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111000111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111001000",
    "01001110100001110100001000110010110100111010000111010000100011001011" when "0111001001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111001010",
    "01110011110111000100110111001010010111001111011100010011011100101001" when "0111001011",
    "01100011101111111101001111000000100110001110111111110100111100000010" when "0111001100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111001101",
    "01110010001000100011011011001001100111001000100010001101101100100111" when "0111001110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111001111",
    "01000001011001101101101101011110000100000101100110110110110101111000" when "0111010000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111010001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111010010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111010011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111010100",
    "01101011001111010110100101000110010110101100111101011010010100011001" when "0111010101",
    "01001010110011011101111110001100010100101011001101110111111000110001" when "0111010110",
    "01011101001010001010011101010000010101110100101000101001110101000001" when "0111010111",
    "01100100111101100001100101110111010110010011110110000110010111011101" when "0111011000",
    "01101001000010011101111010010101010110100100001001110111101001010101" when "0111011001",
    "01001100011000000110100100001001110100110001100000011010010000100111" when "0111011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111011011",
    "01001101101101011001001100011110010100110110110101100100110001111001" when "0111011100",
    "01001100110001110110010000010100000100110011000111011001000001010000" when "0111011101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0111011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111011111",
    "01111000101001110111001101100110100111100010100111011100110110011010" when "0111100000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111100001",
    "01001010111000101101010010110110110100101011100010110101001011011011" when "0111100010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111100011",
    "01110011110111100010101101001111110111001111011110001010110100111111" when "0111100100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111100101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0111100110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "0111100111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111101000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111101001",
    "01000101010111001010101010110101110100010101011100101010101011010111" when "0111101010",
    "01001111110100010011100001000110000100111111010001001110000100011000" when "0111101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0111101100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111101101",
    "01010100111101110000101101010111010101010011110111000010110101011101" when "0111101110",
    "01000000100011110100101110000011100100000010001111010010111000001110" when "0111101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111110000",
    "01001011100111000001000011100000010100101110011100000100001110000001" when "0111110001",
    "01001011001111110111101101010110010100101100111111011110110101011001" when "0111110010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111110011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "0111110101",
    "01010111110011101000001111011100010101011111001110100000111101110001" when "0111110110",
    "01001011000011000100000110001011100100101100001100010000011000101110" when "0111110111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111111000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111111001",
    "01001001000001111001101101010110100100100100000111100110110101011010" when "0111111010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "0111111011",
    "01000011011110000100100001101111110100001101111000010010000110111111" when "0111111100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "0111111101",
    "01011010111000010110011000001011100101101011100001011001100000101110" when "0111111110",
    "01100000001010111110101111001101000110000000101011111010111100110101" when "0111111111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000000000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1000000001",
    "01001010000110100111000101111001100100101000011010011100010111100110" when "1000000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000000011",
    "01101100100101110010011000001011000110110010010111001001100000101100" when "1000000100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000000101",
    "01011001001111001001101110010100010101100100111100100110111001010001" when "1000000110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1000000111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000001000",
    "01000011010100011100101011011100110100001101010001110010101101110011" when "1000001001",
    "01101000001011001111010101000110000110100000101100111101010100011000" when "1000001010",
    "01100001100101011111000000110110110110000110010101111100000011011011" when "1000001011",
    "01001100101001011001011010110010100100110010100101100101101011001010" when "1000001100",
    "01111111101100011100111010101011100111111110110001110011101010110000" when "1000001101",
    "01011000011110001110011100100001110101100001111000111001110010000111" when "1000001110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000001111",
    "01010101010010010011011000100111110101010101001001001101100010011111" when "1000010000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1000010001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000010010",
    "01101011100011111010100111011011000110101110001111101010011101101100" when "1000010011",
    "01100000011110111010001101010001000110000001111011101000110101000100" when "1000010100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1000010101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000010110",
    "01110101010101101011000011101111010111010101010110101100001110111101" when "1000010111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000011000",
    "01000010100010000100010010000011110100001010001000010001001000001111" when "1000011001",
    "01011100001000000110101111110010100101110000100000011010111111001010" when "1000011010",
    "01110110011101101101001000000010010111011001110110110100100000001001" when "1000011011",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1000011100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1000011101",
    "01010101101110100110100010101100010101010110111010011010001010110001" when "1000011110",
    "01111110100001001001000111110100110111111010000100100100011111010011" when "1000011111",
    "01100100000001110000101000111110110110010000000111000010100011111011" when "1000100000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000100001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1000100010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1000100011",
    "01100100100010001001110101001100110110010010001000100111010100110011" when "1000100100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000100101",
    "01011111101101011110111101100000000101111110110101111011110110000000" when "1000100110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000100111",
    "01101101000111101000100110111110110110110100011110100010011011111011" when "1000101000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000101010",
    "01001001101000111010010000101000100100100110100011101001000010100010" when "1000101011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000101100",
    "01101100010000001000000000010110010110110001000000100000000001011001" when "1000101101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000101110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000110000",
    "01100111110010110001110001001000110110011111001011000111000100100011" when "1000110001",
    "01011110100011011001000001101001100101111010001101100100000110100110" when "1000110010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1000110011",
    "01110011110001010100111111011001110111001111000101010011111101100111" when "1000110100",
    "01101100100110101011001011011001100110110010011010101100101101100110" when "1000110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000110110",
    "01011110000101110010001101111000110101111000010111001000110111100011" when "1000110111",
    "01011110100110000110011001101011010101111010011000011001100110101101" when "1000111000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000111001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1000111010",
    "01000110011101010001110000110001100100011001110101000111000011000111" when "1000111011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000111100",
    "01111000011011100101001110111011100111100001101110010100111011101110" when "1000111101",
    "01100010100000110100101111010100000110001010000011010010111101010000" when "1000111110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1000111111",
    "01111001011100000111111000000110110111100101110000011111100000011011" when "1001000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001000001",
    "01011010111011011001111000101101010101101011101101100111100010110101" when "1001000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001000011",
    "01011101111001101010101001101100100101110111100110101010100110110010" when "1001000100",
    "01001011110000110111111010000010010100101111000011011111101000001010" when "1001000101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1001000110",
    "01000000110010110001100111101001100100000011001011000110011110100110" when "1001000111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001001000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001001001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001001010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001001011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001001100",
    "01100010001000110000010000001000000110001000100011000001000000100000" when "1001001101",
    "01101101001001011001001011111100010110110100100101100100101111110001" when "1001001110",
    "01101011100111001001011100100000010110101110011100100101110010000001" when "1001001111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001010000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001010001",
    "01110010000101111001111010010011010111001000010111100111101001001101" when "1001010010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001010011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001010100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001010101",
    "01001100001010111010011001000001110100110000101011101001100100000111" when "1001010110",
    "01110000010110011010110010000110100111000001011001101011001000011010" when "1001010111",
    "01101110010101110010110011000110000110111001010111001011001100011000" when "1001011000",
    "01001110110001011110010011011101100100111011000101111001001101110110" when "1001011001",
    "01110100010110000011101100111010010111010001011000001110110011101001" when "1001011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1001011011",
    "01001100110000001010000110000011000100110011000000101000011000001100" when "1001011100",
    "01000111111110110011010101110001010100011111111011001101010111000101" when "1001011101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001011111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001100000",
    "01011110100001101001000100110010000101111010000110100100010011001000" when "1001100001",
    "01011111111001000000110010111011000101111111100100000011001011110000" when "1001100010",
    "01000100001011111111000001111000100100010000101111111100000111100010" when "1001100011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1001100100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001100101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001100110",
    "01001110100111011001101001111101110100111010011101100110100111110111" when "1001100111",
    "01111011001100110000111101011011100111101100110011000011110101101110" when "1001101000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1001101001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1001101010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001101100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001101101",
    "01010111000110101110010001100101100101011100011010111001000110010110" when "1001101110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001101111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001110000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1001110001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1001110010",
    "01001101000111000111000111001011010100110100011100011100011100101101" when "1001110011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1001110100",
    "01001010111111000100001100000010110100101011111100010000110000001011" when "1001110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001110110",
    "01000011111001111101111010011011110100001111100111110111101001101111" when "1001110111",
    "01010000101101111001110011000100010101000010110111100111001100010001" when "1001111000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001111001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1001111010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001111011",
    "01101101110100110111000111001100010110110111010011011100011100110001" when "1001111100",
    "01010010100011001001101100100100100101001010001100100110110010010010" when "1001111101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001111110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1001111111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010000000",
    "01100101001101001100000000010001110110010100110100110000000001000111" when "1010000001",
    "01111101101010100010101001011100010111110110101010001010100101110001" when "1010000010",
    "01100011000100110011110100000100010110001100010011001111010000010001" when "1010000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010000100",
    "01101001110010101110111101010001110110100111001010111011110101001000" when "1010000101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1010000110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010000111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010001000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010001001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010001010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010001011",
    "01000000001001000000000110000011110100000000100100000000011000010001" when "1010001100",
    "01100000100101011000000111010101000110000010010101100000011101010100" when "1010001101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010001110",
    "01110010000100110111011110101001010111001000010011011101111010100101" when "1010001111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010010000",
    "01000110110101101000111111010111110100011011010110100011111101011111" when "1010010001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010010010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010010011",
    "01001001001000010000110010111111000100100100100001000011001011111100" when "1010010100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010010101",
    "01001000011111011110111100001011110100100001111101111011110000101111" when "1010010110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010010111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1010011000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010011001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1010011011",
    "01100011100100010001001001111100000110001110010001000100100111110000" when "1010011100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010011101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010011111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010100000",
    "01100111001110011100101100100010100110011100111001110010110010001010" when "1010100001",
    "01000110100001010010101110111011100100011010000101001010111011101110" when "1010100010",
    "01000011111010000101011110000000010100001111101000010101111000000001" when "1010100011",
    "01101100110101010100010111001001110110110011010101010001011100100111" when "1010100100",
    "01101010001000010010101010011100010110101000100001001010101001110001" when "1010100101",
    "01001000001111011101111101101101100100100000111101110111110110110110" when "1010100110",
    "01010001111011011010101000001001010101000111101101101010100000100101" when "1010100111",
    "01000001001010010110101011100010010100000100101001011010101110001001" when "1010101000",
    "01111001110111010010110111001101010111100111011101001011011100110101" when "1010101001",
    "01100101111011110010010101001111110110010111101111001001010100111111" when "1010101010",
    "01001110011100100110110010001001000100111001110010011011001000100100" when "1010101011",
    "01001100010110110100110111110100000100110001011011010011011111010000" when "1010101100",
    "01110010111101100010001011011110010111001011110110001000101101111001" when "1010101101",
    "01111001010001111100000111010111100111100101000111110000011101011110" when "1010101110",
    "01011000011001001011110001111111000101100001100100101111000111111100" when "1010101111",
    "01001010001110000000001101011111000100101000111000000000110101111100" when "1010110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010110001",
    "01000110111001101110011010101010000100011011100110111001101010101000" when "1010110010",
    "01000100100110111101000101000110110100010010011011110100010100011011" when "1010110011",
    "01101001100001000110110000011101000110100110000100011011000001110100" when "1010110100",
    "01101011010010010001111000111100100110101101001001000111100011110010" when "1010110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010110110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010110111",
    "01011001111011000010101010011101110101100111101100001010101001110111" when "1010111000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1010111001",
    "01111001010110110101101010101010110111100101011011010110101010101011" when "1010111010",
    "01101000011111101111010101111110110110100001111110111101010111111011" when "1010111011",
    "01111111010001000010011101110111010111111101000100001001110111011101" when "1010111100",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1010111101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1010111110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1010111111",
    "01000101111001001111010010111000010100010111100100111101001011100001" when "1011000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011000001",
    "01111001000000111001011110000110000111100100000011100101111000011000" when "1011000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011000011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1011000100",
    "01000110110101100101101000001101110100011011010110010110100000110111" when "1011000101",
    "01101001110100101011101000101111000110100111010010101110100010111100" when "1011000110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011000111",
    "01001110110011000110010010001101000100111011001100011001001000110100" when "1011001000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1011001001",
    "01000110010111011000011100010111100100011001011101100001110001011110" when "1011001010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011001011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1011001100",
    "01001111100011111010101000010011010100111110001111101010100001001101" when "1011001101",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011001110",
    "01100101110110110100010000001100010110010111011011010001000000110001" when "1011001111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1011010000",
    "01110111010011111000010101111010100111011101001111100001010111101010" when "1011010001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011010010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011010011",
    "01010011010011100110010100101011100101001101001110011001010010101110" when "1011010100",
    "01000101100101000101101011000001110100010110010100010110101100000111" when "1011010101",
    "01111011111010000000101110101100100111101111101000000010111010110010" when "1011010110",
    "01011110011101111001001011111010110101111001110111100100101111101011" when "1011010111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011011000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011011001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1011011010",
    "01100000101100000110110101001100110110000010110000011011010100110011" when "1011011011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011011100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011011101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011011110",
    "01010100000000111111010100011111010101010000000011111101010001111101" when "1011011111",
    "01111000010010001001000011101010110111100001001000100100001110101011" when "1011100000",
    "01011111111010010011110101110010000101111111101001001111010111001000" when "1011100001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011100010",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011100011",
    "01110111100111001000110000100101010111011110011100100011000010010101" when "1011100100",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1011100101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011100110",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1011100111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011101000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1011101001",
    "01100111001010000100111001101011000110011100101000010011100110101100" when "1011101010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011101011",
    "01111111111111101000010100111101100111111111111110100001010101010000" when "1011101100",
    "01010111111010111011011010011111010101011111101011101101101001111101" when "1011101101",
    "01000101100111011110000101010101000100010110011101111000010101010100" when "1011101110",
    "01011101110100111001101110101011100101110111010011100110111010101110" when "1011101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011110000",
    "01101111001001000010010100110110010110111100100100001001010011011001" when "1011110001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011110010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011110011",
    "01011111100101010011000010100011000101111110010101001100001010001100" when "1011110100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1011110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011110110",
    "01111000110011110001011011101101010111100011001111000101101110110101" when "1011110111",
    "01101010100100100100110001011001000110101010010010010011000101100100" when "1011111000",
    "01111000000001000101100111111111010111100000000100010110011111111101" when "1011111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011111010",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1011111011",
    "01000111101110100001110010101101010100011110111010000111001010110101" when "1011111100",
    "01101101000001010111011110010000000110110100000101011101111001000000" when "1011111101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1011111110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1011111111",
    "01000000101111111110101000111011010100000010111111111010100011101101" when "1100000000",
    "01001011100110110100111000100110110100101110011011010011100010011011" when "1100000001",
    "01001101100011100111111010101001100100110110001110011111101010100110" when "1100000010",
    "01111110100100101111101011110011100111111010010010111110101111001110" when "1100000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100000100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100000101",
    "01101011011011010000001111101110000110101101101101000000111110111000" when "1100000110",
    "01010000101101101001011011111111000101000010110110100101101111111100" when "1100000111",
    "01101100001000101110110111111100000110110000100010111011011111110000" when "1100001000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100001001",
    "01101100010101110011101101000110100110110001010111001110110100011010" when "1100001010",
    "01111111011111000101011010110001010111111101111100010101101011000101" when "1100001011",
    "01001110110100101010101110100011110100111011010010101010111010001111" when "1100001100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100001101",
    "01111110111101000110010110001010000111111011110100011001011000101001" when "1100001110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100001111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1100010000",
    "01001010100101110000010110010100000100101010010111000001011001010000" when "1100010001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100010010",
    "01100101011101101110100110101110010110010101110110111010011010111001" when "1100010011",
    "01000000101001110010111111001100000100000010100111001011111100110000" when "1100010100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100010101",
    "01100100010010101100111001110111110110010001001010110011100111011111" when "1100010110",
    "01001000110010101000111100000010110100100011001010100011110000001011" when "1100010111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100011000",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1100011001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100011010",
    "01111110001111111001010000001100110111111000111111100101000000110011" when "1100011011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1100011100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1100011101",
    "01110100111100000010100011001110010111010011110000001010001100111001" when "1100011110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100011111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100100000",
    "01100110110000000110101111011110000110011011000000011010111101111000" when "1100100001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1100100010",
    "01111100001000011010010111001111110111110000100001101001011100111111" when "1100100011",
    "01101100101100100000101001001011100110110010110010000010100100101110" when "1100100100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100100101",
    "01100000010000010000101100111110010110000001000001000010110011111001" when "1100100110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1100100111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100101000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100101001",
    "01011011101001011110001001011100110101101110100101111000100101110011" when "1100101010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100101011",
    "01001110010110001001110101100010000100111001011000100111010110001000" when "1100101100",
    "01110101110000000010010110000011110111010111000000001001011000001111" when "1100101101",
    "01101011100100110010000001011011100110101110010011001000000101101110" when "1100101110",
    "01001101010000000011010100000110110100110101000000001101010000011011" when "1100101111",
    "01101100111110100110110100011010010110110011111010011011010001101001" when "1100110000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100110001",
    "01100101011100001100010000001101000110010101110000110001000000110100" when "1100110010",
    "01111110110000110100111000000000000111111011000011010011100000000000" when "1100110011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100110101",
    "01111001010010000100111010001101000111100101001000010011101000110100" when "1100110110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1100110111",
    "01111111010111110100001001001100110111111101011111010000100100110011" when "1100111000",
    "01110101110101101000000000000011110111010111010110100000000000001111" when "1100111001",
    "01001110101011110010101110010001010100111010101111001010111001000101" when "1100111010",
    "01000110001111010110100010111001110100011000111101011010001011100111" when "1100111011",
    "01111110001010000111001001100111010111111000101000011100100110011101" when "1100111100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100111101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1100111110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1100111111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101000001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101000100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1101000101",
    "01001110000011110111010101101101110100111000001111011101010110110111" when "1101000110",
    "01011100000010000011010010010000010101110000001000001101001001000001" when "1101000111",
    "01000100001001111010001101001100010100010000100111101000110100110001" when "1101001000",
    "01110000111010011010100011001011110111000011101001101010001100101111" when "1101001001",
    "01111011011010101111011100011001010111101101101010111101110001100101" when "1101001010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101001011",
    "01011100100110111011011111110100000101110010011011101101111111010001" when "1101001100",
    "01011010001100111000101011101010010101101000110011100010101110101001" when "1101001101",
    "01000001000110110100011100001000110100000100011011010001110000100011" when "1101001110",
    "01110000001101111110000101100110010111000000110111111000010110011111" when "1101001111",
    "01111100111110000001001100111110110111110011111000000100110011111011" when "1101010000",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1101010001",
    "01001000111100001101111100110110110100100011110000110111110011011011" when "1101010010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101010011",
    "01000011101100110110111111111100000100001110110011011011111111110000" when "1101010100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101010101",
    "01111000000111111111011000010100110111100000011111111101100001010011" when "1101010110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101010111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1101011000",
    "01001001100110001100110110111101010100100110011000110011011011110101" when "1101011001",
    "01011000110001001100100010111000110101100011000100110010001011100100" when "1101011010",
    "01111100000110010101010110110000000111110000011001010101011011000000" when "1101011011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101011100",
    "01101100110100111001011101010010100110110011010011100101110101001010" when "1101011101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1101011110",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1101011111",
    "01101100111000010101011010101001110110110011100001010101101010100111" when "1101100000",
    "01110100011000100001011001101100010111010001100010000101100110110001" when "1101100001",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1101100010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101100011",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1101100100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101100101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1101100110",
    "01111110101101101011001000101100000111111010110110101100100010110000" when "1101100111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101101000",
    "01101110111010010110010110000101110110111011101001011001011000010111" when "1101101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101101010",
    "01000001011010000101000110011011110100000101101000010100011001101111" when "1101101011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101101100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101101101",
    "01001110011000001111110010010001100100111001100000111111001001000110" when "1101101110",
    "01111101001111010100110000100001010111110100111101010011000010000101" when "1101101111",
    "01111001000111100010110011010111110111100100011110001011001101011111" when "1101110000",
    "01000010000101101011101100000010100100001000010110101110110000001010" when "1101110001",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101110010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1101110011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101110101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101110110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101110111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101111000",
    "01011100111010111101010100111101010101110011101011110101010011110101" when "1101111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1101111010",
    "01011101110000110101010000110101110101110111000011010101000011010111" when "1101111011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101111100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1101111101",
    "01111001010111100100100001001011000111100101011110010010000100101100" when "1101111110",
    "01101111111111010010011011011010010110111111111101001001101101101001" when "1101111111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110000000",
    "01010001010011110101010101100101000101000101001111010101010110010100" when "1110000001",
    "01010010010100101110000111010000110101001001010010111000011101000011" when "1110000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110000011",
    "01101111100011001010010111100010000110111110001100101001011110001000" when "1110000100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110000101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110000110",
    "01101010100011011001110110001001100110101010001101100111011000100110" when "1110000111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110001000",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1110001001",
    "01110101001011101011000000001100110111010100101110101100000000110011" when "1110001010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110001011",
    "01101000101100010100111011101000100110100010110001010011101110100010" when "1110001100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110001101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110001110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110001111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110010000",
    "01011011111111000001001000110101010101101111111100000100100011010101" when "1110010001",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110010010",
    "01010010100001001100100110111110100101001010000100110010011011111010" when "1110010011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110010100",
    "01011101101110110100000111010011110101110110111011010000011101001111" when "1110010101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1110010110",
    "01000100111000011001101100001001100100010011100001100110110000100110" when "1110010111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110011000",
    "01101101000101010010011010101001000110110100010101001001101010100100" when "1110011001",
    "01110010001000010101100101110110010111001000100001010110010111011001" when "1110011010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110011011",
    "01101111000010101111110101101100010110111100001010111111010110110001" when "1110011100",
    "01100010100011100010000001110001110110001010001110001000000111001000" when "1110011101",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110011110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110011111",
    "01101010001001101100111110010000110110101000100110110011111001000011" when "1110100000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110100001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110100010",
    "01010100111010011001100111100011000101010011101001100110011110001100" when "1110100011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110100100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110100101",
    "01100100100010111110001111101011100110010010001011111000111110101110" when "1110100110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110100111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110101000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110101010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1110101011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110101100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1110101101",
    "01000110111101110110010110001010110100011011110111011001011000101011" when "1110101110",
    "01001110000000010110100100001110100100111000000001011010010000111010" when "1110101111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110110000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110110001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110110010",
    "01101100110010110011000100100111000110110011001011001100010010011100" when "1110110011",
    "01100011001111111000000100001011110110001100111111100000010000110000" when "1110110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110110110",
    "01001100111100100010110111010001000100110011110010001011011101000100" when "1110110111",
    "01000111110001010011000111111010000100011111000101001100011111101000" when "1110111000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110111001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1110111010",
    "01000001011010011011011110111011110100000101101001101101111011110000" when "1110111011",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1110111100",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1110111101",
    "01110110101110101001000010111001100111011010111010100100001011100110" when "1110111110",
    "01010111010001001001111001111100010101011101000100100111100111110001" when "1110111111",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111000000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111000001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1111000010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111000011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111000100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111000101",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1111000110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111000111",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1111001000",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111001001",
    "01100101011111000010110101110100010110010101111100001011010111010001" when "1111001010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111001011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111001100",
    "01000010101000110110000100110000110100001010100011011000010011000011" when "1111001101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111001110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111001111",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111010000",
    "01000110110010010110011000101011110100011011001001011001100010101111" when "1111010001",
    "01101101101111001010000010111001000110110110111100101000001011100100" when "1111010010",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1111010011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111010100",
    "01010110110100111011011001000000110101011011010011101101100100000011" when "1111010101",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111010110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111010111",
    "01000110010110000101111110100111100100011001011000010111111010011110" when "1111011000",
    "01100111111001100110001101111001010110011111100110011000110111100101" when "1111011001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111011010",
    "01101010101101110101101110010110100110101010110111010110111001011011" when "1111011011",
    "01011111010000110000010010111000100101111101000011000001001011100011" when "1111011100",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1111011101",
    "01111100010001100000001110110111010111110001000110000000111011011101" when "1111011110",
    "01100001101010011001111011110000100110000110101001100111101111000010" when "1111011111",
    "01110011110010110000000000010010010111001111001011000000000001001001" when "1111100000",
    "01001110010010111110000101100100100100111001001011111000010110010010" when "1111100001",
    "00000000000000000000000000000000000000000000000000000000000000000000" when "1111100010",
    "01011001000110111101110010011010100101100100011011110111001001101010" when "1111100011",
    "01101001001101001111010010110011010110100100110100111101001011001101" when "1111100100",
    "01110100100011110110111000100010010111010010001111011011100010001010" when "1111100101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111100110",
    "01001101001001000111000010101000110100110100100100011100001010100011" when "1111100111",
    "01110111000101111001111100010000000111011100010111100111110001000001" when "1111101000",
    "01001111100010110010000100100110000100111110001011001000010010011000" when "1111101001",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111101010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111101011",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111101100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111101101",
    "01101110001111110011100110011101110110111000111111001110011001110111" when "1111101110",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1111101111",
    "00100000000000000000000000000000000010000000000000000000000000000000" when "1111110000",
    "10111111111111111111111111111111111011111111111111111111111111111111" when "1111110001",
    "01110001100000000011000000111111110111000110000000001100000011111111" when "1111110010",
    "10011111111111111111111111111111111001111111111111111111111111111111" when "1111110011",
    "01001000001111100001100001110001010100100000111110000110000111000101" when "1111110100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111110101",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111110110",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111110111",
    "01001000111101101000111111101001000100100011110110100011111110100100" when "1111111000",
    "01100110111101001111101000101000100110011011110100111110100010100010" when "1111111001",
    "01000111101010110111111111111101100100011110101011011111111111110110" when "1111111010",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111111011",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111111100",
    "11011111111111111111111111111111111101111111111111111111111111111111" when "1111111101",
    "01010110101101110011001001101011000101011010110111001100100110101100" when "1111111110",
    "01100101110101111111001000110101110110010111010111111100100011010111" when "1111111111",
    "00000000000000000000000000000000000000000000000000000000000000000000" when others;

end architecture;
